1 0 0 8 0
2 32 1 0
2 1973 1 0
2 1974 1 0
2 1975 1 0
2 1976 1 0
2 1977 1 0
2 1978 1 0
2 1979 1 0
1 1 0 9 0
2 1980 1 1
2 1981 1 1
2 1982 1 1
2 1983 1 1
2 1984 1 1
2 1985 1 1
2 1986 1 1
2 1987 1 1
2 1988 1 1
1 2 0 10 0
2 1989 1 2
2 1990 1 2
2 1991 1 2
2 1992 1 2
2 1993 1 2
2 1994 1 2
2 1995 1 2
2 1996 1 2
2 1997 1 2
2 1998 1 2
1 3 0 11 0
2 1999 1 3
2 2000 1 3
2 2001 1 3
2 2002 1 3
2 2003 1 3
2 2004 1 3
2 2005 1 3
2 2006 1 3
2 2007 1 3
2 2008 1 3
2 2009 1 3
1 4 0 10 0
2 2010 1 4
2 2011 1 4
2 2012 1 4
2 2013 1 4
2 2014 1 4
2 2015 1 4
2 2016 1 4
2 2017 1 4
2 2018 1 4
2 2019 1 4
1 5 0 11 0
2 2020 1 5
2 2021 1 5
2 2022 1 5
2 2023 1 5
2 2024 1 5
2 2025 1 5
2 2026 1 5
2 2027 1 5
2 2028 1 5
2 2029 1 5
2 2030 1 5
1 6 0 10 0
2 2031 1 6
2 2032 1 6
2 2033 1 6
2 2034 1 6
2 2035 1 6
2 2036 1 6
2 2037 1 6
2 2038 1 6
2 2039 1 6
2 2040 1 6
1 7 0 10 0
2 2041 1 7
2 2042 1 7
2 2043 1 7
2 2044 1 7
2 2045 1 7
2 2046 1 7
2 2047 1 7
2 2048 1 7
2 2049 1 7
2 2050 1 7
1 8 0 10 0
2 2051 1 8
2 2052 1 8
2 2053 1 8
2 2054 1 8
2 2055 1 8
2 2056 1 8
2 2057 1 8
2 2058 1 8
2 2059 1 8
2 2060 1 8
1 9 0 10 0
2 2061 1 9
2 2062 1 9
2 2063 1 9
2 2064 1 9
2 2065 1 9
2 2066 1 9
2 2067 1 9
2 2068 1 9
2 2069 1 9
2 2070 1 9
1 10 0 11 0
2 2071 1 10
2 2072 1 10
2 2073 1 10
2 2074 1 10
2 2075 1 10
2 2076 1 10
2 2077 1 10
2 2078 1 10
2 2079 1 10
2 2080 1 10
2 2081 1 10
1 11 0 10 0
2 2082 1 11
2 2083 1 11
2 2084 1 11
2 2085 1 11
2 2086 1 11
2 2087 1 11
2 2088 1 11
2 2089 1 11
2 2090 1 11
2 2091 1 11
1 12 0 10 0
2 2092 1 12
2 2093 1 12
2 2094 1 12
2 2095 1 12
2 2096 1 12
2 2097 1 12
2 2098 1 12
2 2099 1 12
2 2100 1 12
2 2101 1 12
1 13 0 10 0
2 2102 1 13
2 2103 1 13
2 2104 1 13
2 2105 1 13
2 2106 1 13
2 2107 1 13
2 2108 1 13
2 2109 1 13
2 2110 1 13
2 2111 1 13
1 14 0 10 0
2 2112 1 14
2 2113 1 14
2 2114 1 14
2 2115 1 14
2 2116 1 14
2 2117 1 14
2 2118 1 14
2 2119 1 14
2 2120 1 14
2 2121 1 14
1 15 0 10 0
2 2122 1 15
2 2123 1 15
2 2124 1 15
2 2125 1 15
2 2126 1 15
2 2127 1 15
2 2128 1 15
2 2129 1 15
2 2130 1 15
2 2131 1 15
1 16 0 3 0
2 2132 1 16
2 2133 1 16
2 2134 1 16
1 17 0 3 0
2 2135 1 17
2 2136 1 17
2 2137 1 17
1 18 0 3 0
2 2138 1 18
2 2139 1 18
2 2140 1 18
1 19 0 3 0
2 2141 1 19
2 2142 1 19
2 2143 1 19
1 20 0 3 0
2 2144 1 20
2 2145 1 20
2 2146 1 20
1 21 0 3 0
2 2147 1 21
2 2148 1 21
2 2149 1 21
1 22 0 3 0
2 2150 1 22
2 2151 1 22
2 2152 1 22
1 23 0 3 0
2 2153 1 23
2 2154 1 23
2 2155 1 23
1 24 0 3 0
2 2156 1 24
2 2157 1 24
2 2158 1 24
1 25 0 3 0
2 2159 1 25
2 2160 1 25
2 2161 1 25
1 26 0 3 0
2 2162 1 26
2 2163 1 26
2 2164 1 26
1 27 0 3 0
2 2165 1 27
2 2166 1 27
2 2167 1 27
1 28 0 4 0
2 2168 1 28
2 2169 1 28
2 2170 1 28
2 2171 1 28
1 29 0 3 0
2 2172 1 29
2 2173 1 29
2 2174 1 29
1 30 0 4 0
2 2175 1 30
2 2176 1 30
2 2177 1 30
2 2178 1 30
1 31 0 4 0
2 2179 1 31
2 2180 1 31
2 2181 1 31
2 2182 1 31
2 2183 1 34
2 2184 1 34
2 2185 1 35
2 2186 1 35
2 2187 1 36
2 2188 1 36
2 2189 1 37
2 2190 1 37
2 2191 1 38
2 2192 1 38
2 2193 1 39
2 2194 1 39
2 2195 1 40
2 2196 1 40
2 2197 1 41
2 2198 1 41
2 2199 1 42
2 2200 1 42
2 2201 1 43
2 2202 1 43
2 2203 1 44
2 2204 1 44
2 2205 1 45
2 2206 1 45
2 2207 1 46
2 2208 1 46
2 2209 1 47
2 2210 1 47
2 2211 1 48
2 2212 1 48
2 2213 1 48
2 2214 1 49
2 2215 1 49
2 2216 1 49
2 2217 1 50
2 2218 1 50
2 2219 1 50
2 2220 1 51
2 2221 1 51
2 2222 1 51
2 2223 1 52
2 2224 1 52
2 2225 1 52
2 2226 1 53
2 2227 1 53
2 2228 1 53
2 2229 1 54
2 2230 1 54
2 2231 1 54
2 2232 1 55
2 2233 1 55
2 2234 1 55
2 2235 1 56
2 2236 1 56
2 2237 1 56
2 2238 1 57
2 2239 1 57
2 2240 1 57
2 2241 1 58
2 2242 1 58
2 2243 1 58
2 2244 1 59
2 2245 1 59
2 2246 1 59
2 2247 1 60
2 2248 1 60
2 2249 1 60
2 2250 1 60
2 2251 1 61
2 2252 1 61
2 2253 1 61
2 2254 1 62
2 2255 1 62
2 2256 1 63
2 2257 1 63
2 2258 1 64
2 2259 1 64
2 2260 1 66
2 2261 1 66
2 2262 1 66
2 2263 1 68
2 2264 1 68
2 2265 1 74
2 2266 1 74
2 2267 1 76
2 2268 1 76
2 2269 1 81
2 2270 1 81
2 2271 1 84
2 2272 1 84
2 2273 1 87
2 2274 1 87
2 2275 1 89
2 2276 1 89
2 2277 1 90
2 2278 1 90
2 2279 1 95
2 2280 1 95
2 2281 1 98
2 2282 1 98
2 2283 1 103
2 2284 1 103
2 2285 1 104
2 2286 1 104
2 2287 1 105
2 2288 1 105
2 2289 1 108
2 2290 1 108
2 2291 1 111
2 2292 1 111
2 2293 1 113
2 2294 1 113
2 2295 1 114
2 2296 1 114
2 2297 1 119
2 2298 1 119
2 2299 1 122
2 2300 1 122
2 2301 1 127
2 2302 1 127
2 2303 1 127
2 2304 1 129
2 2305 1 129
2 2306 1 132
2 2307 1 132
2 2308 1 135
2 2309 1 135
2 2310 1 137
2 2311 1 137
2 2312 1 138
2 2313 1 138
2 2314 1 143
2 2315 1 143
2 2316 1 146
2 2317 1 146
2 2318 1 151
2 2319 1 151
2 2320 1 151
2 2321 1 153
2 2322 1 153
2 2323 1 156
2 2324 1 156
2 2325 1 159
2 2326 1 159
2 2327 1 161
2 2328 1 161
2 2329 1 162
2 2330 1 162
2 2331 1 167
2 2332 1 167
2 2333 1 170
2 2334 1 170
2 2335 1 175
2 2336 1 175
2 2337 1 175
2 2338 1 177
2 2339 1 177
2 2340 1 180
2 2341 1 180
2 2342 1 183
2 2343 1 183
2 2344 1 185
2 2345 1 185
2 2346 1 186
2 2347 1 186
2 2348 1 191
2 2349 1 191
2 2350 1 194
2 2351 1 194
2 2352 1 199
2 2353 1 199
2 2354 1 199
2 2355 1 201
2 2356 1 201
2 2357 1 204
2 2358 1 204
2 2359 1 207
2 2360 1 207
2 2361 1 209
2 2362 1 209
2 2363 1 210
2 2364 1 210
2 2365 1 215
2 2366 1 215
2 2367 1 218
2 2368 1 218
2 2369 1 223
2 2370 1 223
2 2371 1 223
2 2372 1 225
2 2373 1 225
2 2374 1 228
2 2375 1 228
2 2376 1 231
2 2377 1 231
2 2378 1 233
2 2379 1 233
2 2380 1 234
2 2381 1 234
2 2382 1 239
2 2383 1 239
2 2384 1 242
2 2385 1 242
2 2386 1 247
2 2387 1 247
2 2388 1 247
2 2389 1 249
2 2390 1 249
2 2391 1 252
2 2392 1 252
2 2393 1 255
2 2394 1 255
2 2395 1 257
2 2396 1 257
2 2397 1 258
2 2398 1 258
2 2399 1 263
2 2400 1 263
2 2401 1 266
2 2402 1 266
2 2403 1 271
2 2404 1 271
2 2405 1 271
2 2406 1 273
2 2407 1 273
2 2408 1 276
2 2409 1 276
2 2410 1 279
2 2411 1 279
2 2412 1 281
2 2413 1 281
2 2414 1 282
2 2415 1 282
2 2416 1 287
2 2417 1 287
2 2418 1 290
2 2419 1 290
2 2420 1 295
2 2421 1 295
2 2422 1 295
2 2423 1 297
2 2424 1 297
2 2425 1 300
2 2426 1 300
2 2427 1 303
2 2428 1 303
2 2429 1 305
2 2430 1 305
2 2431 1 306
2 2432 1 306
2 2433 1 311
2 2434 1 311
2 2435 1 314
2 2436 1 314
2 2437 1 319
2 2438 1 319
2 2439 1 319
2 2440 1 321
2 2441 1 321
2 2442 1 324
2 2443 1 324
2 2444 1 327
2 2445 1 327
2 2446 1 329
2 2447 1 329
2 2448 1 330
2 2449 1 330
2 2450 1 335
2 2451 1 335
2 2452 1 338
2 2453 1 338
2 2454 1 343
2 2455 1 343
2 2456 1 343
2 2457 1 345
2 2458 1 345
2 2459 1 348
2 2460 1 348
2 2461 1 351
2 2462 1 351
2 2463 1 353
2 2464 1 353
2 2465 1 354
2 2466 1 354
2 2467 1 359
2 2468 1 359
2 2469 1 362
2 2470 1 362
2 2471 1 367
2 2472 1 367
2 2473 1 367
2 2474 1 369
2 2475 1 369
2 2476 1 372
2 2477 1 372
2 2478 1 375
2 2479 1 375
2 2480 1 377
2 2481 1 377
2 2482 1 378
2 2483 1 378
2 2484 1 383
2 2485 1 383
2 2486 1 386
2 2487 1 386
2 2488 1 391
2 2489 1 391
2 2490 1 391
2 2491 1 393
2 2492 1 393
2 2493 1 396
2 2494 1 396
2 2495 1 399
2 2496 1 399
2 2497 1 401
2 2498 1 401
2 2499 1 402
2 2500 1 402
2 2501 1 407
2 2502 1 407
2 2503 1 410
2 2504 1 410
2 2505 1 415
2 2506 1 415
2 2507 1 415
2 2508 1 417
2 2509 1 417
2 2510 1 420
2 2511 1 420
2 2512 1 423
2 2513 1 423
2 2514 1 425
2 2515 1 425
2 2516 1 426
2 2517 1 426
2 2518 1 431
2 2519 1 431
2 2520 1 434
2 2521 1 434
2 2522 1 439
2 2523 1 439
2 2524 1 439
2 2525 1 441
2 2526 1 441
2 2527 1 444
2 2528 1 444
2 2529 1 447
2 2530 1 447
2 2531 1 449
2 2532 1 449
2 2533 1 450
2 2534 1 450
2 2535 1 455
2 2536 1 455
2 2537 1 458
2 2538 1 458
2 2539 1 463
2 2540 1 463
2 2541 1 463
2 2542 1 465
2 2543 1 465
2 2544 1 468
2 2545 1 468
2 2546 1 471
2 2547 1 471
2 2548 1 473
2 2549 1 473
2 2550 1 474
2 2551 1 474
2 2552 1 479
2 2553 1 479
2 2554 1 482
2 2555 1 482
2 2556 1 487
2 2557 1 487
2 2558 1 487
2 2559 1 489
2 2560 1 489
2 2561 1 492
2 2562 1 492
2 2563 1 495
2 2564 1 495
2 2565 1 497
2 2566 1 497
2 2567 1 498
2 2568 1 498
2 2569 1 503
2 2570 1 503
2 2571 1 506
2 2572 1 506
2 2573 1 511
2 2574 1 511
2 2575 1 511
2 2576 1 513
2 2577 1 513
2 2578 1 516
2 2579 1 516
2 2580 1 519
2 2581 1 519
2 2582 1 521
2 2583 1 521
2 2584 1 522
2 2585 1 522
2 2586 1 527
2 2587 1 527
2 2588 1 530
2 2589 1 530
2 2590 1 535
2 2591 1 535
2 2592 1 535
2 2593 1 537
2 2594 1 537
2 2595 1 540
2 2596 1 540
2 2597 1 543
2 2598 1 543
2 2599 1 545
2 2600 1 545
2 2601 1 546
2 2602 1 546
2 2603 1 551
2 2604 1 551
2 2605 1 554
2 2606 1 554
2 2607 1 559
2 2608 1 559
2 2609 1 559
2 2610 1 561
2 2611 1 561
2 2612 1 564
2 2613 1 564
2 2614 1 567
2 2615 1 567
2 2616 1 569
2 2617 1 569
2 2618 1 570
2 2619 1 570
2 2620 1 575
2 2621 1 575
2 2622 1 578
2 2623 1 578
2 2624 1 583
2 2625 1 583
2 2626 1 583
2 2627 1 585
2 2628 1 585
2 2629 1 588
2 2630 1 588
2 2631 1 591
2 2632 1 591
2 2633 1 593
2 2634 1 593
2 2635 1 594
2 2636 1 594
2 2637 1 599
2 2638 1 599
2 2639 1 602
2 2640 1 602
2 2641 1 607
2 2642 1 607
2 2643 1 607
2 2644 1 609
2 2645 1 609
2 2646 1 612
2 2647 1 612
2 2648 1 615
2 2649 1 615
2 2650 1 617
2 2651 1 617
2 2652 1 618
2 2653 1 618
2 2654 1 623
2 2655 1 623
2 2656 1 626
2 2657 1 626
2 2658 1 631
2 2659 1 631
2 2660 1 631
2 2661 1 633
2 2662 1 633
2 2663 1 636
2 2664 1 636
2 2665 1 639
2 2666 1 639
2 2667 1 641
2 2668 1 641
2 2669 1 642
2 2670 1 642
2 2671 1 647
2 2672 1 647
2 2673 1 650
2 2674 1 650
2 2675 1 655
2 2676 1 655
2 2677 1 655
2 2678 1 657
2 2679 1 657
2 2680 1 660
2 2681 1 660
2 2682 1 663
2 2683 1 663
2 2684 1 665
2 2685 1 665
2 2686 1 666
2 2687 1 666
2 2688 1 671
2 2689 1 671
2 2690 1 674
2 2691 1 674
2 2692 1 679
2 2693 1 679
2 2694 1 679
2 2695 1 681
2 2696 1 681
2 2697 1 686
2 2698 1 686
2 2699 1 687
2 2700 1 687
2 2701 1 687
2 2702 1 689
2 2703 1 689
2 2704 1 694
2 2705 1 694
2 2706 1 697
2 2707 1 697
2 2708 1 702
2 2709 1 702
2 2710 1 708
2 2711 1 708
2 2712 1 711
2 2713 1 711
2 2714 1 713
2 2715 1 713
2 2716 1 722
2 2717 1 722
2 2718 1 728
2 2719 1 728
2 2720 1 730
2 2721 1 730
2 2722 1 732
2 2723 1 732
2 2724 1 735
2 2725 1 735
2 2726 1 736
2 2727 1 736
2 2728 1 740
2 2729 1 740
2 2730 1 743
2 2731 1 743
2 2732 1 744
2 2733 1 744
2 2734 1 746
2 2735 1 746
2 2736 1 747
2 2737 1 747
2 2738 1 748
2 2739 1 748
2 2740 1 750
2 2741 1 750
2 2742 1 755
2 2743 1 755
2 2744 1 756
2 2745 1 756
2 2746 1 759
2 2747 1 759
2 2748 1 762
2 2749 1 762
2 2750 1 765
2 2751 1 765
2 2752 1 766
2 2753 1 766
2 2754 1 770
2 2755 1 770
2 2756 1 773
2 2757 1 773
2 2758 1 774
2 2759 1 774
2 2760 1 776
2 2761 1 776
2 2762 1 779
2 2763 1 779
2 2764 1 780
2 2765 1 780
2 2766 1 784
2 2767 1 784
2 2768 1 787
2 2769 1 787
2 2770 1 788
2 2771 1 788
2 2772 1 792
2 2773 1 792
2 2774 1 795
2 2775 1 795
2 2776 1 796
2 2777 1 796
2 2778 1 800
2 2779 1 800
2 2780 1 803
2 2781 1 803
2 2782 1 804
2 2783 1 804
2 2784 1 806
2 2785 1 806
2 2786 1 808
2 2787 1 808
2 2788 1 810
2 2789 1 810
2 2790 1 816
2 2791 1 816
2 2792 1 819
2 2793 1 819
2 2794 1 819
2 2795 1 822
2 2796 1 822
2 2797 1 825
2 2798 1 825
2 2799 1 826
2 2800 1 826
2 2801 1 830
2 2802 1 830
2 2803 1 833
2 2804 1 833
2 2805 1 834
2 2806 1 834
2 2807 1 838
2 2808 1 838
2 2809 1 841
2 2810 1 841
2 2811 1 842
2 2812 1 842
2 2813 1 846
2 2814 1 846
2 2815 1 849
2 2816 1 849
2 2817 1 850
2 2818 1 850
2 2819 1 852
2 2820 1 852
2 2821 1 854
2 2822 1 854
2 2823 1 855
2 2824 1 855
2 2825 1 856
2 2826 1 856
2 2827 1 857
2 2828 1 857
2 2829 1 858
2 2830 1 858
2 2831 1 861
2 2832 1 861
2 2833 1 862
2 2834 1 862
2 2835 1 866
2 2836 1 866
2 2837 1 869
2 2838 1 869
2 2839 1 870
2 2840 1 870
2 2841 1 874
2 2842 1 874
2 2843 1 877
2 2844 1 877
2 2845 1 878
2 2846 1 878
2 2847 1 882
2 2848 1 882
2 2849 1 885
2 2850 1 885
2 2851 1 886
2 2852 1 886
2 2853 1 890
2 2854 1 890
2 2855 1 893
2 2856 1 893
2 2857 1 894
2 2858 1 894
2 2859 1 898
2 2860 1 898
2 2861 1 901
2 2862 1 901
2 2863 1 902
2 2864 1 902
2 2865 1 906
2 2866 1 906
2 2867 1 909
2 2868 1 909
2 2869 1 910
2 2870 1 910
2 2871 1 914
2 2872 1 914
2 2873 1 917
2 2874 1 917
2 2875 1 918
2 2876 1 918
2 2877 1 920
2 2878 1 920
2 2879 1 923
2 2880 1 923
2 2881 1 926
2 2882 1 926
2 2883 1 930
2 2884 1 930
2 2885 1 933
2 2886 1 933
2 2887 1 934
2 2888 1 934
2 2889 1 938
2 2890 1 938
2 2891 1 941
2 2892 1 941
2 2893 1 942
2 2894 1 942
2 2895 1 944
2 2896 1 944
2 2897 1 947
2 2898 1 947
2 2899 1 948
2 2900 1 948
2 2901 1 950
2 2902 1 950
2 2903 1 956
2 2904 1 956
2 2905 1 959
2 2906 1 959
2 2907 1 962
2 2908 1 962
2 2909 1 965
2 2910 1 965
2 2911 1 968
2 2912 1 968
2 2913 1 972
2 2914 1 972
2 2915 1 975
2 2916 1 975
2 2917 1 976
2 2918 1 976
2 2919 1 980
2 2920 1 980
2 2921 1 983
2 2922 1 983
2 2923 1 984
2 2924 1 984
2 2925 1 986
2 2926 1 986
2 2927 1 989
2 2928 1 989
2 2929 1 992
2 2930 1 992
2 2931 1 996
2 2932 1 996
2 2933 1 999
2 2934 1 999
2 2935 1 1000
2 2936 1 1000
2 2937 1 1004
2 2938 1 1004
2 2939 1 1007
2 2940 1 1007
2 2941 1 1008
2 2942 1 1008
2 2943 1 1012
2 2944 1 1012
2 2945 1 1015
2 2946 1 1015
2 2947 1 1016
2 2948 1 1016
2 2949 1 1020
2 2950 1 1020
2 2951 1 1023
2 2952 1 1023
2 2953 1 1024
2 2954 1 1024
2 2955 1 1028
2 2956 1 1028
2 2957 1 1031
2 2958 1 1031
2 2959 1 1032
2 2960 1 1032
2 2961 1 1034
2 2962 1 1034
2 2963 1 1037
2 2964 1 1037
2 2965 1 1038
2 2966 1 1038
2 2967 1 1042
2 2968 1 1042
2 2969 1 1045
2 2970 1 1045
2 2971 1 1046
2 2972 1 1046
2 2973 1 1048
2 2974 1 1048
2 2975 1 1050
2 2976 1 1050
2 2977 1 1053
2 2978 1 1053
2 2979 1 1054
2 2980 1 1054
2 2981 1 1056
2 2982 1 1056
2 2983 1 1058
2 2984 1 1058
2 2985 1 1060
2 2986 1 1060
2 2987 1 1061
2 2988 1 1061
2 2989 1 1062
2 2990 1 1062
2 2991 1 1063
2 2992 1 1063
2 2993 1 1064
2 2994 1 1064
2 2995 1 1065
2 2996 1 1065
2 2997 1 1066
2 2998 1 1066
2 2999 1 1067
2 3000 1 1067
2 3001 1 1068
2 3002 1 1068
2 3003 1 1071
2 3004 1 1071
2 3005 1 1074
2 3006 1 1074
2 3007 1 1078
2 3008 1 1078
2 3009 1 1081
2 3010 1 1081
2 3011 1 1084
2 3012 1 1084
2 3013 1 1088
2 3014 1 1088
2 3015 1 1091
2 3016 1 1091
2 3017 1 1092
2 3018 1 1092
2 3019 1 1095
2 3020 1 1095
2 3021 1 1096
2 3022 1 1096
2 3023 1 1100
2 3024 1 1100
2 3025 1 1103
2 3026 1 1103
2 3027 1 1104
2 3028 1 1104
2 3029 1 1108
2 3030 1 1108
2 3031 1 1111
2 3032 1 1111
2 3033 1 1112
2 3034 1 1112
2 3035 1 1116
2 3036 1 1116
2 3037 1 1119
2 3038 1 1119
2 3039 1 1122
2 3040 1 1122
2 3041 1 1126
2 3042 1 1126
2 3043 1 1129
2 3044 1 1129
2 3045 1 1132
2 3046 1 1132
2 3047 1 1136
2 3048 1 1136
2 3049 1 1139
2 3050 1 1139
2 3051 1 1140
2 3052 1 1140
2 3053 1 1142
2 3054 1 1142
2 3055 1 1145
2 3056 1 1145
2 3057 1 1146
2 3058 1 1146
2 3059 1 1150
2 3060 1 1150
2 3061 1 1153
2 3062 1 1153
2 3063 1 1154
2 3064 1 1154
2 3065 1 1158
2 3066 1 1158
2 3067 1 1161
2 3068 1 1161
2 3069 1 1162
2 3070 1 1162
2 3071 1 1166
2 3072 1 1166
2 3073 1 1169
2 3074 1 1169
2 3075 1 1170
2 3076 1 1170
2 3077 1 1174
2 3078 1 1174
2 3079 1 1177
2 3080 1 1177
2 3081 1 1178
2 3082 1 1178
2 3083 1 1182
2 3084 1 1182
2 3085 1 1185
2 3086 1 1185
2 3087 1 1186
2 3088 1 1186
2 3089 1 1188
2 3090 1 1188
2 3091 1 1194
2 3092 1 1194
2 3093 1 1197
2 3094 1 1197
2 3095 1 1200
2 3096 1 1200
2 3097 1 1203
2 3098 1 1203
2 3099 1 1206
2 3100 1 1206
2 3101 1 1210
2 3102 1 1210
2 3103 1 1213
2 3104 1 1213
2 3105 1 1214
2 3106 1 1214
2 3107 1 1218
2 3108 1 1218
2 3109 1 1221
2 3110 1 1221
2 3111 1 1222
2 3112 1 1222
2 3113 1 1226
2 3114 1 1226
2 3115 1 1229
2 3116 1 1229
2 3117 1 1230
2 3118 1 1230
2 3119 1 1234
2 3120 1 1234
2 3121 1 1237
2 3122 1 1237
2 3123 1 1238
2 3124 1 1238
2 3125 1 1242
2 3126 1 1242
2 3127 1 1245
2 3128 1 1245
2 3129 1 1246
2 3130 1 1246
2 3131 1 1250
2 3132 1 1250
2 3133 1 1253
2 3134 1 1253
2 3135 1 1254
2 3136 1 1254
2 3137 1 1258
2 3138 1 1258
2 3139 1 1261
2 3140 1 1261
2 3141 1 1262
2 3142 1 1262
2 3143 1 1264
2 3144 1 1264
2 3145 1 1267
2 3146 1 1267
2 3147 1 1270
2 3148 1 1270
2 3149 1 1274
2 3150 1 1274
2 3151 1 1277
2 3152 1 1277
2 3153 1 1278
2 3154 1 1278
2 3155 1 1282
2 3156 1 1282
2 3157 1 1285
2 3158 1 1285
2 3159 1 1286
2 3160 1 1286
2 3161 1 1290
2 3162 1 1290
2 3163 1 1293
2 3164 1 1293
2 3165 1 1294
2 3166 1 1294
2 3167 1 1298
2 3168 1 1298
2 3169 1 1301
2 3170 1 1301
2 3171 1 1302
2 3172 1 1302
2 3173 1 1308
2 3174 1 1308
2 3175 1 1311
2 3176 1 1311
2 3177 1 1312
2 3178 1 1312
2 3179 1 1316
2 3180 1 1316
2 3181 1 1319
2 3182 1 1319
2 3183 1 1320
2 3184 1 1320
2 3185 1 1324
2 3186 1 1324
2 3187 1 1327
2 3188 1 1327
2 3189 1 1328
2 3190 1 1328
2 3191 1 1332
2 3192 1 1332
2 3193 1 1335
2 3194 1 1335
2 3195 1 1336
2 3196 1 1336
2 3197 1 1338
2 3198 1 1338
2 3199 1 1341
2 3200 1 1341
2 3201 1 1344
2 3202 1 1344
2 3203 1 1348
2 3204 1 1348
2 3205 1 1351
2 3206 1 1351
2 3207 1 1352
2 3208 1 1352
2 3209 1 1356
2 3210 1 1356
2 3211 1 1359
2 3212 1 1359
2 3213 1 1362
2 3214 1 1362
2 3215 1 1364
2 3216 1 1364
2 3217 1 1366
2 3218 1 1366
2 3219 1 1368
2 3220 1 1368
2 3221 1 1370
2 3222 1 1370
2 3223 1 1372
2 3224 1 1372
2 3225 1 1374
2 3226 1 1374
2 3227 1 1375
2 3228 1 1375
2 3229 1 1376
2 3230 1 1376
2 3231 1 1376
2 3232 1 1379
2 3233 1 1379
2 3234 1 1382
2 3235 1 1382
2 3236 1 1390
2 3237 1 1390
2 3238 1 1393
2 3239 1 1393
2 3240 1 1394
2 3241 1 1394
2 3242 1 1398
2 3243 1 1398
2 3244 1 1401
2 3245 1 1401
2 3246 1 1404
2 3247 1 1404
2 3248 1 1406
2 3249 1 1406
2 3250 1 1408
2 3251 1 1408
2 3252 1 1410
2 3253 1 1410
2 3254 1 1411
2 3255 1 1411
2 3256 1 1413
2 3257 1 1413
2 3258 1 1414
2 3259 1 1414
2 3260 1 1418
2 3261 1 1418
2 3262 1 1421
2 3263 1 1421
2 3264 1 1422
2 3265 1 1422
2 3266 1 1426
2 3267 1 1426
2 3268 1 1429
2 3269 1 1429
2 3270 1 1430
2 3271 1 1430
2 3272 1 1434
2 3273 1 1434
2 3274 1 1437
2 3275 1 1437
2 3276 1 1438
2 3277 1 1438
2 3278 1 1442
2 3279 1 1442
2 3280 1 1445
2 3281 1 1445
2 3282 1 1446
2 3283 1 1446
2 3284 1 1450
2 3285 1 1450
2 3286 1 1453
2 3287 1 1453
2 3288 1 1454
2 3289 1 1454
2 3290 1 1458
2 3291 1 1458
2 3292 1 1461
2 3293 1 1461
2 3294 1 1462
2 3295 1 1462
2 3296 1 1466
2 3297 1 1466
2 3298 1 1469
2 3299 1 1469
2 3300 1 1470
2 3301 1 1470
2 3302 1 1474
2 3303 1 1474
2 3304 1 1477
2 3305 1 1477
2 3306 1 1478
2 3307 1 1478
2 3308 1 1482
2 3309 1 1482
2 3310 1 1485
2 3311 1 1485
2 3312 1 1486
2 3313 1 1486
2 3314 1 1490
2 3315 1 1490
2 3316 1 1493
2 3317 1 1493
2 3318 1 1494
2 3319 1 1494
2 3320 1 1498
2 3321 1 1498
2 3322 1 1501
2 3323 1 1501
2 3324 1 1502
2 3325 1 1502
2 3326 1 1504
2 3327 1 1504
2 3328 1 1509
2 3329 1 1509
2 3330 1 1512
2 3331 1 1512
2 3332 1 1515
2 3333 1 1515
2 3334 1 1518
2 3335 1 1518
2 3336 1 1521
2 3337 1 1521
2 3338 1 1521
2 3339 1 1522
2 3340 1 1522
2 3341 1 1524
2 3342 1 1524
2 3343 1 1526
2 3344 1 1526
2 3345 1 1528
2 3346 1 1528
2 3347 1 1529
2 3348 1 1529
2 3349 1 1531
2 3350 1 1531
2 3351 1 1534
2 3352 1 1534
2 3353 1 1537
2 3354 1 1537
2 3355 1 1537
2 3356 1 1539
2 3357 1 1539
2 3358 1 1539
2 3359 1 1539
2 3360 1 1542
2 3361 1 1542
2 3362 1 1545
2 3363 1 1545
2 3364 1 1545
2 3365 1 1545
2 3366 1 1545
2 3367 1 1547
2 3368 1 1547
2 3369 1 1550
2 3370 1 1550
2 3371 1 1553
2 3372 1 1553
2 3373 1 1553
2 3374 1 1553
2 3375 1 1554
2 3376 1 1554
2 3377 1 1554
2 3378 1 1556
2 3379 1 1556
2 3380 1 1556
2 3381 1 1556
2 3382 1 1559
2 3383 1 1559
2 3384 1 1562
2 3385 1 1562
2 3386 1 1562
2 3387 1 1562
2 3388 1 1564
2 3389 1 1564
2 3390 1 1564
2 3391 1 1564
2 3392 1 1567
2 3393 1 1567
2 3394 1 1570
2 3395 1 1570
2 3396 1 1570
2 3397 1 1570
2 3398 1 1570
2 3399 1 1572
2 3400 1 1572
2 3401 1 1572
2 3402 1 1572
2 3403 1 1572
2 3404 1 1575
2 3405 1 1575
2 3406 1 1578
2 3407 1 1578
2 3408 1 1578
2 3409 1 1578
2 3410 1 1580
2 3411 1 1580
2 3412 1 1580
2 3413 1 1580
2 3414 1 1583
2 3415 1 1583
2 3416 1 1586
2 3417 1 1586
2 3418 1 1586
2 3419 1 1588
2 3420 1 1588
2 3421 1 1588
2 3422 1 1588
2 3423 1 1591
2 3424 1 1591
2 3425 1 1594
2 3426 1 1594
2 3427 1 1594
2 3428 1 1596
2 3429 1 1596
2 3430 1 1596
2 3431 1 1596
2 3432 1 1599
2 3433 1 1599
2 3434 1 1602
2 3435 1 1602
2 3436 1 1602
2 3437 1 1602
2 3438 1 1604
2 3439 1 1604
2 3440 1 1604
2 3441 1 1604
2 3442 1 1607
2 3443 1 1607
2 3444 1 1610
2 3445 1 1610
2 3446 1 1610
2 3447 1 1610
2 3448 1 1612
2 3449 1 1612
2 3450 1 1612
2 3451 1 1612
2 3452 1 1615
2 3453 1 1615
2 3454 1 1618
2 3455 1 1618
2 3456 1 1618
2 3457 1 1618
2 3458 1 1620
2 3459 1 1620
2 3460 1 1620
2 3461 1 1620
2 3462 1 1623
2 3463 1 1623
2 3464 1 1626
2 3465 1 1626
2 3466 1 1626
2 3467 1 1626
2 3468 1 1628
2 3469 1 1628
2 3470 1 1628
2 3471 1 1628
2 3472 1 1631
2 3473 1 1631
2 3474 1 1634
2 3475 1 1634
2 3476 1 1636
2 3477 1 1636
2 3478 1 1637
2 3479 1 1637
2 3480 1 1641
2 3481 1 1641
2 3482 1 1644
2 3483 1 1644
2 3484 1 1644
2 3485 1 1647
2 3486 1 1647
2 3487 1 1647
2 3488 1 1651
2 3489 1 1651
2 3490 1 1653
2 3491 1 1653
2 3492 1 1655
2 3493 1 1655
2 3494 1 1656
2 3495 1 1656
2 3496 1 1659
2 3497 1 1659
2 3498 1 1660
2 3499 1 1660
2 3500 1 1663
2 3501 1 1663
2 3502 1 1664
2 3503 1 1664
2 3504 1 1667
2 3505 1 1667
2 3506 1 1668
2 3507 1 1668
2 3508 1 1671
2 3509 1 1671
2 3510 1 1677
2 3511 1 1677
2 3512 1 1679
2 3513 1 1679
2 3514 1 1679
2 3515 1 1685
2 3516 1 1685
2 3517 1 1686
2 3518 1 1686
2 3519 1 1689
2 3520 1 1689
2 3521 1 1690
2 3522 1 1690
2 3523 1 1692
2 3524 1 1692
2 3525 1 1692
2 3526 1 1693
2 3527 1 1693
2 3528 1 1693
2 3529 1 1697
2 3530 1 1697
2 3531 1 1701
2 3532 1 1701
2 3533 1 1701
2 3534 1 1702
2 3535 1 1702
2 3536 1 1703
2 3537 1 1703
2 3538 1 1709
2 3539 1 1709
2 3540 1 1711
2 3541 1 1711
2 3542 1 1712
2 3543 1 1712
2 3544 1 1715
2 3545 1 1715
2 3546 1 1717
2 3547 1 1717
2 3548 1 1719
2 3549 1 1719
2 3550 1 1720
2 3551 1 1720
2 3552 1 1723
2 3553 1 1723
2 3554 1 1724
2 3555 1 1724
2 3556 1 1727
2 3557 1 1727
2 3558 1 1729
2 3559 1 1729
2 3560 1 1732
2 3561 1 1732
2 3562 1 1735
2 3563 1 1735
2 3564 1 1739
2 3565 1 1739
2 3566 1 1739
2 3567 1 1740
2 3568 1 1740
2 3569 1 1743
2 3570 1 1743
2 3571 1 1746
2 3572 1 1746
2 3573 1 1749
2 3574 1 1749
2 3575 1 1752
2 3576 1 1752
2 3577 1 1752
2 3578 1 1757
2 3579 1 1757
2 3580 1 1757
2 3581 1 1758
2 3582 1 1758
2 3583 1 1761
2 3584 1 1761
2 3585 1 1762
2 3586 1 1762
2 3587 1 1769
2 3588 1 1769
2 3589 1 1769
2 3590 1 1770
2 3591 1 1770
2 3592 1 1781
2 3593 1 1781
2 3594 1 1782
2 3595 1 1782
2 3596 1 1785
2 3597 1 1785
2 3598 1 1785
2 3599 1 1786
2 3600 1 1786
2 3601 1 1791
2 3602 1 1791
2 3603 1 1791
2 3604 1 1792
2 3605 1 1792
2 3606 1 1797
2 3607 1 1797
2 3608 1 1798
2 3609 1 1798
2 3610 1 1801
2 3611 1 1801
2 3612 1 1802
2 3613 1 1802
2 3614 1 1807
2 3615 1 1807
2 3616 1 1808
2 3617 1 1808
2 3618 1 1811
2 3619 1 1811
2 3620 1 1812
2 3621 1 1812
2 3622 1 1852
2 3623 1 1852
2 3624 1 1854
2 3625 1 1854
0 33 5 1 1 1980
0 34 5 2 1 1989
0 35 5 2 1 1999
0 36 5 2 1 2010
0 37 5 2 1 2020
0 38 5 2 1 2031
0 39 5 2 1 2041
0 40 5 2 1 2051
0 41 5 2 1 2061
0 42 5 2 1 2071
0 43 5 2 1 2082
0 44 5 2 1 2092
0 45 5 2 1 2102
0 46 5 2 1 2112
0 47 5 2 1 2122
0 48 5 3 1 2132
0 49 5 3 1 2135
0 50 5 3 1 2138
0 51 5 3 1 2141
0 52 5 3 1 2144
0 53 5 3 1 2147
0 54 5 3 1 2150
0 55 5 3 1 2153
0 56 5 3 1 2156
0 57 5 3 1 2159
0 58 5 3 1 2162
0 59 5 3 1 2165
0 60 5 4 1 2168
0 61 5 3 1 2172
0 62 5 2 1 2175
0 63 5 2 1 2179
0 64 7 2 2 2251 2254
0 65 5 1 1 2258
0 66 7 3 2 2180 2259
0 67 5 1 1 2260
0 68 7 2 2 2252 2181
0 69 5 1 1 2263
0 70 7 1 2 65 2264
0 71 5 1 1 70
0 72 7 1 2 2173 2256
0 73 5 1 1 72
0 74 7 2 2 71 73
0 75 5 1 1 2265
0 76 7 2 2 2247 2266
0 77 5 1 1 2267
0 78 7 1 2 2176 69
0 79 7 1 2 77 78
0 80 5 1 1 79
0 81 7 2 2 67 80
0 82 5 1 1 2269
0 83 7 1 2 2248 82
0 84 5 2 1 83
0 85 7 1 2 2169 2270
0 86 5 1 1 85
0 87 7 2 2 2271 86
0 88 5 1 1 2273
0 89 7 2 2 2244 2274
0 90 5 2 1 2275
0 91 7 1 2 75 2272
0 92 5 1 1 91
0 93 7 1 2 2249 2261
0 94 5 1 1 93
0 95 7 2 2 92 94
0 96 5 1 1 2279
0 97 7 1 2 2277 96
0 98 5 2 1 97
0 99 7 1 2 2177 2268
0 100 5 1 1 99
0 101 7 1 2 2170 2262
0 102 5 1 1 101
0 103 7 2 2 100 102
0 104 5 2 1 2283
0 105 7 2 2 2281 2284
0 106 5 1 1 2287
0 107 7 1 2 2245 106
0 108 5 2 1 107
0 109 7 1 2 2166 2288
0 110 5 1 1 109
0 111 7 2 2 2289 110
0 112 5 1 1 2291
0 113 7 2 2 2241 2292
0 114 5 2 1 2293
0 115 7 1 2 88 2290
0 116 5 1 1 115
0 117 7 1 2 2276 2285
0 118 5 1 1 117
0 119 7 2 2 116 118
0 120 5 1 1 2297
0 121 7 1 2 2295 120
0 122 5 2 1 121
0 123 7 1 2 2278 2286
0 124 5 1 1 123
0 125 7 1 2 2280 124
0 126 5 1 1 125
0 127 7 3 2 2282 126
0 128 5 1 1 2301
0 129 7 2 2 2299 128
0 130 5 1 1 2304
0 131 7 1 2 2242 130
0 132 5 2 1 131
0 133 7 1 2 2163 2305
0 134 5 1 1 133
0 135 7 2 2 2306 134
0 136 5 1 1 2308
0 137 7 2 2 2238 2309
0 138 5 2 1 2310
0 139 7 1 2 112 2307
0 140 5 1 1 139
0 141 7 1 2 2294 2302
0 142 5 1 1 141
0 143 7 2 2 140 142
0 144 5 1 1 2314
0 145 7 1 2 2312 144
0 146 5 2 1 145
0 147 7 1 2 2296 2303
0 148 5 1 1 147
0 149 7 1 2 2298 148
0 150 5 1 1 149
0 151 7 3 2 2300 150
0 152 5 1 1 2318
0 153 7 2 2 2316 152
0 154 5 1 1 2321
0 155 7 1 2 2239 154
0 156 5 2 1 155
0 157 7 1 2 2160 2322
0 158 5 1 1 157
0 159 7 2 2 2323 158
0 160 5 1 1 2325
0 161 7 2 2 2235 2326
0 162 5 2 1 2327
0 163 7 1 2 136 2324
0 164 5 1 1 163
0 165 7 1 2 2311 2319
0 166 5 1 1 165
0 167 7 2 2 164 166
0 168 5 1 1 2331
0 169 7 1 2 2329 168
0 170 5 2 1 169
0 171 7 1 2 2313 2320
0 172 5 1 1 171
0 173 7 1 2 2315 172
0 174 5 1 1 173
0 175 7 3 2 2317 174
0 176 5 1 1 2335
0 177 7 2 2 2333 176
0 178 5 1 1 2338
0 179 7 1 2 2236 178
0 180 5 2 1 179
0 181 7 1 2 2157 2339
0 182 5 1 1 181
0 183 7 2 2 2340 182
0 184 5 1 1 2342
0 185 7 2 2 2232 2343
0 186 5 2 1 2344
0 187 7 1 2 160 2341
0 188 5 1 1 187
0 189 7 1 2 2328 2336
0 190 5 1 1 189
0 191 7 2 2 188 190
0 192 5 1 1 2348
0 193 7 1 2 2346 192
0 194 5 2 1 193
0 195 7 1 2 2330 2337
0 196 5 1 1 195
0 197 7 1 2 2332 196
0 198 5 1 1 197
0 199 7 3 2 2334 198
0 200 5 1 1 2352
0 201 7 2 2 2350 200
0 202 5 1 1 2355
0 203 7 1 2 2233 202
0 204 5 2 1 203
0 205 7 1 2 2154 2356
0 206 5 1 1 205
0 207 7 2 2 2357 206
0 208 5 1 1 2359
0 209 7 2 2 2229 2360
0 210 5 2 1 2361
0 211 7 1 2 184 2358
0 212 5 1 1 211
0 213 7 1 2 2345 2353
0 214 5 1 1 213
0 215 7 2 2 212 214
0 216 5 1 1 2365
0 217 7 1 2 2363 216
0 218 5 2 1 217
0 219 7 1 2 2347 2354
0 220 5 1 1 219
0 221 7 1 2 2349 220
0 222 5 1 1 221
0 223 7 3 2 2351 222
0 224 5 1 1 2369
0 225 7 2 2 2367 224
0 226 5 1 1 2372
0 227 7 1 2 2230 226
0 228 5 2 1 227
0 229 7 1 2 2151 2373
0 230 5 1 1 229
0 231 7 2 2 2374 230
0 232 5 1 1 2376
0 233 7 2 2 2226 2377
0 234 5 2 1 2378
0 235 7 1 2 208 2375
0 236 5 1 1 235
0 237 7 1 2 2362 2370
0 238 5 1 1 237
0 239 7 2 2 236 238
0 240 5 1 1 2382
0 241 7 1 2 2380 240
0 242 5 2 1 241
0 243 7 1 2 2364 2371
0 244 5 1 1 243
0 245 7 1 2 2366 244
0 246 5 1 1 245
0 247 7 3 2 2368 246
0 248 5 1 1 2386
0 249 7 2 2 2384 248
0 250 5 1 1 2389
0 251 7 1 2 2227 250
0 252 5 2 1 251
0 253 7 1 2 2148 2390
0 254 5 1 1 253
0 255 7 2 2 2391 254
0 256 5 1 1 2393
0 257 7 2 2 2223 2394
0 258 5 2 1 2395
0 259 7 1 2 232 2392
0 260 5 1 1 259
0 261 7 1 2 2379 2387
0 262 5 1 1 261
0 263 7 2 2 260 262
0 264 5 1 1 2399
0 265 7 1 2 2397 264
0 266 5 2 1 265
0 267 7 1 2 2381 2388
0 268 5 1 1 267
0 269 7 1 2 2383 268
0 270 5 1 1 269
0 271 7 3 2 2385 270
0 272 5 1 1 2403
0 273 7 2 2 2401 272
0 274 5 1 1 2406
0 275 7 1 2 2224 274
0 276 5 2 1 275
0 277 7 1 2 2145 2407
0 278 5 1 1 277
0 279 7 2 2 2408 278
0 280 5 1 1 2410
0 281 7 2 2 2220 2411
0 282 5 2 1 2412
0 283 7 1 2 256 2409
0 284 5 1 1 283
0 285 7 1 2 2396 2404
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 2416
0 289 7 1 2 2414 288
0 290 5 2 1 289
0 291 7 1 2 2398 2405
0 292 5 1 1 291
0 293 7 1 2 2400 292
0 294 5 1 1 293
0 295 7 3 2 2402 294
0 296 5 1 1 2420
0 297 7 2 2 2418 296
0 298 5 1 1 2423
0 299 7 1 2 2221 298
0 300 5 2 1 299
0 301 7 1 2 2142 2424
0 302 5 1 1 301
0 303 7 2 2 2425 302
0 304 5 1 1 2427
0 305 7 2 2 2217 2428
0 306 5 2 1 2429
0 307 7 1 2 280 2426
0 308 5 1 1 307
0 309 7 1 2 2413 2421
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 2433
0 313 7 1 2 2431 312
0 314 5 2 1 313
0 315 7 1 2 2415 2422
0 316 5 1 1 315
0 317 7 1 2 2417 316
0 318 5 1 1 317
0 319 7 3 2 2419 318
0 320 5 1 1 2437
0 321 7 2 2 2435 320
0 322 5 1 1 2440
0 323 7 1 2 2218 322
0 324 5 2 1 323
0 325 7 1 2 2139 2441
0 326 5 1 1 325
0 327 7 2 2 2442 326
0 328 5 1 1 2444
0 329 7 2 2 2214 2445
0 330 5 2 1 2446
0 331 7 1 2 304 2443
0 332 5 1 1 331
0 333 7 1 2 2430 2438
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 2450
0 337 7 1 2 2448 336
0 338 5 2 1 337
0 339 7 1 2 2432 2439
0 340 5 1 1 339
0 341 7 1 2 2434 340
0 342 5 1 1 341
0 343 7 3 2 2436 342
0 344 5 1 1 2454
0 345 7 2 2 2452 344
0 346 5 1 1 2457
0 347 7 1 2 2215 346
0 348 5 2 1 347
0 349 7 1 2 2136 2458
0 350 5 1 1 349
0 351 7 2 2 2459 350
0 352 5 1 1 2461
0 353 7 2 2 2211 2462
0 354 5 2 1 2463
0 355 7 1 2 328 2460
0 356 5 1 1 355
0 357 7 1 2 2447 2455
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 2467
0 361 7 1 2 2465 360
0 362 5 2 1 361
0 363 7 1 2 2449 2456
0 364 5 1 1 363
0 365 7 1 2 2451 364
0 366 5 1 1 365
0 367 7 3 2 2453 366
0 368 5 1 1 2471
0 369 7 2 2 2469 368
0 370 5 1 1 2474
0 371 7 1 2 2212 370
0 372 5 2 1 371
0 373 7 1 2 2133 2475
0 374 5 1 1 373
0 375 7 2 2 2476 374
0 376 5 1 1 2478
0 377 7 2 2 2209 2479
0 378 5 2 1 2480
0 379 7 1 2 352 2477
0 380 5 1 1 379
0 381 7 1 2 2464 2472
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 2484
0 385 7 1 2 2482 384
0 386 5 2 1 385
0 387 7 1 2 2466 2473
0 388 5 1 1 387
0 389 7 1 2 2468 388
0 390 5 1 1 389
0 391 7 3 2 2470 390
0 392 5 1 1 2488
0 393 7 2 2 2486 392
0 394 5 1 1 2491
0 395 7 1 2 2210 394
0 396 5 2 1 395
0 397 7 1 2 2123 2492
0 398 5 1 1 397
0 399 7 2 2 2493 398
0 400 5 1 1 2495
0 401 7 2 2 2207 2496
0 402 5 2 1 2497
0 403 7 1 2 376 2494
0 404 5 1 1 403
0 405 7 1 2 2481 2489
0 406 5 1 1 405
0 407 7 2 2 404 406
0 408 5 1 1 2501
0 409 7 1 2 2499 408
0 410 5 2 1 409
0 411 7 1 2 2483 2490
0 412 5 1 1 411
0 413 7 1 2 2485 412
0 414 5 1 1 413
0 415 7 3 2 2487 414
0 416 5 1 1 2505
0 417 7 2 2 2503 416
0 418 5 1 1 2508
0 419 7 1 2 2208 418
0 420 5 2 1 419
0 421 7 1 2 2113 2509
0 422 5 1 1 421
0 423 7 2 2 2510 422
0 424 5 1 1 2512
0 425 7 2 2 2205 2513
0 426 5 2 1 2514
0 427 7 1 2 400 2511
0 428 5 1 1 427
0 429 7 1 2 2498 2506
0 430 5 1 1 429
0 431 7 2 2 428 430
0 432 5 1 1 2518
0 433 7 1 2 2516 432
0 434 5 2 1 433
0 435 7 1 2 2500 2507
0 436 5 1 1 435
0 437 7 1 2 2502 436
0 438 5 1 1 437
0 439 7 3 2 2504 438
0 440 5 1 1 2522
0 441 7 2 2 2520 440
0 442 5 1 1 2525
0 443 7 1 2 2206 442
0 444 5 2 1 443
0 445 7 1 2 2103 2526
0 446 5 1 1 445
0 447 7 2 2 2527 446
0 448 5 1 1 2529
0 449 7 2 2 2203 2530
0 450 5 2 1 2531
0 451 7 1 2 424 2528
0 452 5 1 1 451
0 453 7 1 2 2515 2523
0 454 5 1 1 453
0 455 7 2 2 452 454
0 456 5 1 1 2535
0 457 7 1 2 2533 456
0 458 5 2 1 457
0 459 7 1 2 2517 2524
0 460 5 1 1 459
0 461 7 1 2 2519 460
0 462 5 1 1 461
0 463 7 3 2 2521 462
0 464 5 1 1 2539
0 465 7 2 2 2537 464
0 466 5 1 1 2542
0 467 7 1 2 2204 466
0 468 5 2 1 467
0 469 7 1 2 2093 2543
0 470 5 1 1 469
0 471 7 2 2 2544 470
0 472 5 1 1 2546
0 473 7 2 2 2201 2547
0 474 5 2 1 2548
0 475 7 1 2 448 2545
0 476 5 1 1 475
0 477 7 1 2 2532 2540
0 478 5 1 1 477
0 479 7 2 2 476 478
0 480 5 1 1 2552
0 481 7 1 2 2550 480
0 482 5 2 1 481
0 483 7 1 2 2534 2541
0 484 5 1 1 483
0 485 7 1 2 2536 484
0 486 5 1 1 485
0 487 7 3 2 2538 486
0 488 5 1 1 2556
0 489 7 2 2 2554 488
0 490 5 1 1 2559
0 491 7 1 2 2202 490
0 492 5 2 1 491
0 493 7 1 2 2083 2560
0 494 5 1 1 493
0 495 7 2 2 2561 494
0 496 5 1 1 2563
0 497 7 2 2 2199 2564
0 498 5 2 1 2565
0 499 7 1 2 472 2562
0 500 5 1 1 499
0 501 7 1 2 2549 2557
0 502 5 1 1 501
0 503 7 2 2 500 502
0 504 5 1 1 2569
0 505 7 1 2 2567 504
0 506 5 2 1 505
0 507 7 1 2 2551 2558
0 508 5 1 1 507
0 509 7 1 2 2553 508
0 510 5 1 1 509
0 511 7 3 2 2555 510
0 512 5 1 1 2573
0 513 7 2 2 2571 512
0 514 5 1 1 2576
0 515 7 1 2 2200 514
0 516 5 2 1 515
0 517 7 1 2 2072 2577
0 518 5 1 1 517
0 519 7 2 2 2578 518
0 520 5 1 1 2580
0 521 7 2 2 2197 2581
0 522 5 2 1 2582
0 523 7 1 2 496 2579
0 524 5 1 1 523
0 525 7 1 2 2566 2574
0 526 5 1 1 525
0 527 7 2 2 524 526
0 528 5 1 1 2586
0 529 7 1 2 2584 528
0 530 5 2 1 529
0 531 7 1 2 2568 2575
0 532 5 1 1 531
0 533 7 1 2 2570 532
0 534 5 1 1 533
0 535 7 3 2 2572 534
0 536 5 1 1 2590
0 537 7 2 2 2588 536
0 538 5 1 1 2593
0 539 7 1 2 2198 538
0 540 5 2 1 539
0 541 7 1 2 2062 2594
0 542 5 1 1 541
0 543 7 2 2 2595 542
0 544 5 1 1 2597
0 545 7 2 2 2195 2598
0 546 5 2 1 2599
0 547 7 1 2 520 2596
0 548 5 1 1 547
0 549 7 1 2 2583 2591
0 550 5 1 1 549
0 551 7 2 2 548 550
0 552 5 1 1 2603
0 553 7 1 2 2601 552
0 554 5 2 1 553
0 555 7 1 2 2585 2592
0 556 5 1 1 555
0 557 7 1 2 2587 556
0 558 5 1 1 557
0 559 7 3 2 2589 558
0 560 5 1 1 2607
0 561 7 2 2 2605 560
0 562 5 1 1 2610
0 563 7 1 2 2196 562
0 564 5 2 1 563
0 565 7 1 2 2052 2611
0 566 5 1 1 565
0 567 7 2 2 2612 566
0 568 5 1 1 2614
0 569 7 2 2 2193 2615
0 570 5 2 1 2616
0 571 7 1 2 544 2613
0 572 5 1 1 571
0 573 7 1 2 2600 2608
0 574 5 1 1 573
0 575 7 2 2 572 574
0 576 5 1 1 2620
0 577 7 1 2 2618 576
0 578 5 2 1 577
0 579 7 1 2 2602 2609
0 580 5 1 1 579
0 581 7 1 2 2604 580
0 582 5 1 1 581
0 583 7 3 2 2606 582
0 584 5 1 1 2624
0 585 7 2 2 2622 584
0 586 5 1 1 2627
0 587 7 1 2 2194 586
0 588 5 2 1 587
0 589 7 1 2 2042 2628
0 590 5 1 1 589
0 591 7 2 2 2629 590
0 592 5 1 1 2631
0 593 7 2 2 2191 2632
0 594 5 2 1 2633
0 595 7 1 2 568 2630
0 596 5 1 1 595
0 597 7 1 2 2617 2625
0 598 5 1 1 597
0 599 7 2 2 596 598
0 600 5 1 1 2637
0 601 7 1 2 2635 600
0 602 5 2 1 601
0 603 7 1 2 2619 2626
0 604 5 1 1 603
0 605 7 1 2 2621 604
0 606 5 1 1 605
0 607 7 3 2 2623 606
0 608 5 1 1 2641
0 609 7 2 2 2639 608
0 610 5 1 1 2644
0 611 7 1 2 2192 610
0 612 5 2 1 611
0 613 7 1 2 2032 2645
0 614 5 1 1 613
0 615 7 2 2 2646 614
0 616 5 1 1 2648
0 617 7 2 2 2189 2649
0 618 5 2 1 2650
0 619 7 1 2 592 2647
0 620 5 1 1 619
0 621 7 1 2 2634 2642
0 622 5 1 1 621
0 623 7 2 2 620 622
0 624 5 1 1 2654
0 625 7 1 2 2652 624
0 626 5 2 1 625
0 627 7 1 2 2636 2643
0 628 5 1 1 627
0 629 7 1 2 2638 628
0 630 5 1 1 629
0 631 7 3 2 2640 630
0 632 5 1 1 2658
0 633 7 2 2 2656 632
0 634 5 1 1 2661
0 635 7 1 2 2190 634
0 636 5 2 1 635
0 637 7 1 2 2021 2662
0 638 5 1 1 637
0 639 7 2 2 2663 638
0 640 5 1 1 2665
0 641 7 2 2 2187 2666
0 642 5 2 1 2667
0 643 7 1 2 616 2664
0 644 5 1 1 643
0 645 7 1 2 2651 2659
0 646 5 1 1 645
0 647 7 2 2 644 646
0 648 5 1 1 2671
0 649 7 1 2 2669 648
0 650 5 2 1 649
0 651 7 1 2 2653 2660
0 652 5 1 1 651
0 653 7 1 2 2655 652
0 654 5 1 1 653
0 655 7 3 2 2657 654
0 656 5 1 1 2675
0 657 7 2 2 2673 656
0 658 5 1 1 2678
0 659 7 1 2 2188 658
0 660 5 2 1 659
0 661 7 1 2 2011 2679
0 662 5 1 1 661
0 663 7 2 2 2680 662
0 664 5 1 1 2682
0 665 7 2 2 2185 2683
0 666 5 2 1 2684
0 667 7 1 2 640 2681
0 668 5 1 1 667
0 669 7 1 2 2668 2676
0 670 5 1 1 669
0 671 7 2 2 668 670
0 672 5 1 1 2688
0 673 7 1 2 2686 672
0 674 5 2 1 673
0 675 7 1 2 2670 2677
0 676 5 1 1 675
0 677 7 1 2 2672 676
0 678 5 1 1 677
0 679 7 3 2 2674 678
0 680 5 1 1 2692
0 681 7 2 2 2690 680
0 682 5 1 1 2695
0 683 7 1 2 2000 2696
0 684 5 1 1 683
0 685 7 1 2 2186 682
0 686 5 2 1 685
0 687 7 3 2 684 2697
0 688 7 1 2 2183 2699
0 689 5 2 1 688
0 690 7 1 2 664 2698
0 691 5 1 1 690
0 692 7 1 2 2685 2693
0 693 5 1 1 692
0 694 7 2 2 691 693
0 695 5 1 1 2704
0 696 7 1 2 2702 695
0 697 5 2 1 696
0 698 7 1 2 2687 2694
0 699 5 1 1 698
0 700 7 1 2 2689 699
0 701 5 1 1 700
0 702 7 2 2 2691 701
0 703 5 1 1 2708
0 704 7 1 2 2703 2709
0 705 5 1 1 704
0 706 7 1 2 2705 705
0 707 5 1 1 706
0 708 7 2 2 2706 707
0 709 7 1 2 2700 2710
0 710 5 1 1 709
0 711 7 2 2 2707 703
0 712 5 1 1 2712
0 713 7 2 2 2184 712
0 714 5 1 1 2714
0 715 7 1 2 2711 2715
0 716 5 1 1 715
0 717 7 1 2 1990 2713
0 718 5 1 1 717
0 719 7 1 2 33 714
0 720 7 1 2 718 719
0 721 5 1 1 720
0 722 7 2 2 716 721
0 723 5 1 1 2716
0 724 7 1 2 710 2717
0 725 5 1 1 724
0 726 7 1 2 2701 723
0 727 5 1 1 726
0 728 7 2 2 725 727
0 729 5 1 1 2718
0 730 7 2 2 2012 2124
0 731 5 1 1 2720
0 732 7 2 2 2043 2094
0 733 5 1 1 2722
0 734 7 1 2 2721 2723
0 735 5 2 1 734
0 736 7 2 2 2033 2104
0 737 5 1 1 2726
0 738 7 1 2 731 733
0 739 5 1 1 738
0 740 7 2 2 739 2724
0 741 5 1 1 2728
0 742 7 1 2 2727 2729
0 743 5 2 1 742
0 744 7 2 2 2725 2730
0 745 5 1 1 2732
0 746 7 2 2 2034 2114
0 747 5 2 1 2734
0 748 7 2 2 2044 2105
0 749 5 1 1 2738
0 750 7 2 2 2022 2125
0 751 5 1 1 2740
0 752 7 1 2 749 751
0 753 5 1 1 752
0 754 7 1 2 2739 2741
0 755 5 2 1 754
0 756 7 2 2 753 2742
0 757 5 1 1 2744
0 758 7 1 2 2735 2745
0 759 5 2 1 758
0 760 7 1 2 2736 757
0 761 5 1 1 760
0 762 7 2 2 2746 761
0 763 5 1 1 2748
0 764 7 1 2 745 2749
0 765 5 2 1 764
0 766 7 2 2 2023 2115
0 767 5 1 1 2752
0 768 7 1 2 737 741
0 769 5 1 1 768
0 770 7 2 2 2731 769
0 771 5 1 1 2754
0 772 7 1 2 2753 2755
0 773 5 2 1 772
0 774 7 2 2 2001 2126
0 775 5 1 1 2758
0 776 7 2 2 2045 2084
0 777 5 1 1 2760
0 778 7 1 2 2759 2761
0 779 5 2 1 778
0 780 7 2 2 2035 2095
0 781 5 1 1 2764
0 782 7 1 2 775 777
0 783 5 1 1 782
0 784 7 2 2 783 2762
0 785 5 1 1 2766
0 786 7 1 2 2765 2767
0 787 5 2 1 786
0 788 7 2 2 2763 2768
0 789 5 1 1 2770
0 790 7 1 2 767 771
0 791 5 1 1 790
0 792 7 2 2 2756 791
0 793 5 1 1 2772
0 794 7 1 2 789 2773
0 795 5 2 1 794
0 796 7 2 2 2757 2774
0 797 5 1 1 2776
0 798 7 1 2 2733 763
0 799 5 1 1 798
0 800 7 2 2 2750 799
0 801 5 1 1 2778
0 802 7 1 2 797 2779
0 803 5 2 1 802
0 804 7 2 2 2751 2780
0 805 5 1 1 2782
0 806 7 2 2 2743 2747
0 807 5 1 1 2784
0 808 7 2 2 2036 2127
0 809 5 1 1 2786
0 810 7 2 2 2046 2116
0 811 5 1 1 2788
0 812 7 1 2 809 2789
0 813 5 1 1 812
0 814 7 1 2 2787 811
0 815 5 1 1 814
0 816 7 2 2 813 815
0 817 5 1 1 2790
0 818 7 1 2 807 817
0 819 5 3 1 818
0 820 7 1 2 2785 2791
0 821 5 1 1 820
0 822 7 2 2 2792 821
0 823 5 1 1 2795
0 824 7 1 2 805 2796
0 825 5 2 1 824
0 826 7 2 2 2013 2117
0 827 5 1 1 2799
0 828 7 1 2 781 785
0 829 5 1 1 828
0 830 7 2 2 2769 829
0 831 5 1 1 2801
0 832 7 1 2 2800 2802
0 833 5 2 1 832
0 834 7 2 2 2024 2106
0 835 5 1 1 2805
0 836 7 1 2 827 831
0 837 5 1 1 836
0 838 7 2 2 2803 837
0 839 5 1 1 2807
0 840 7 1 2 2806 2808
0 841 5 2 1 840
0 842 7 2 2 2804 2809
0 843 5 1 1 2811
0 844 7 1 2 2771 793
0 845 5 1 1 844
0 846 7 2 2 2775 845
0 847 5 1 1 2813
0 848 7 1 2 843 2814
0 849 5 2 1 848
0 850 7 2 2 2047 2053
0 851 5 1 1 2817
0 852 7 2 2 2037 2063
0 853 5 1 1 2819
0 854 7 2 2 2818 2820
0 855 5 2 1 2821
0 856 7 2 2 2073 2822
0 857 5 2 1 2825
0 858 7 2 2 1991 2128
0 859 5 1 1 2829
0 860 7 1 2 2826 2830
0 861 5 2 1 860
0 862 7 2 2 2048 2074
0 863 5 1 1 2833
0 864 7 1 2 2827 859
0 865 5 1 1 864
0 866 7 2 2 2831 865
0 867 5 1 1 2835
0 868 7 1 2 2834 2836
0 869 5 2 1 868
0 870 7 2 2 2832 2837
0 871 5 1 1 2839
0 872 7 1 2 835 839
0 873 5 1 1 872
0 874 7 2 2 2810 873
0 875 5 1 1 2841
0 876 7 1 2 871 2842
0 877 5 2 1 876
0 878 7 2 2 2025 2096
0 879 5 1 1 2845
0 880 7 1 2 863 867
0 881 5 1 1 880
0 882 7 2 2 2838 881
0 883 5 1 1 2847
0 884 7 1 2 2846 2848
0 885 5 2 1 884
0 886 7 2 2 2038 2085
0 887 5 1 1 2851
0 888 7 1 2 879 883
0 889 5 1 1 888
0 890 7 2 2 2849 889
0 891 5 1 1 2853
0 892 7 1 2 2852 2854
0 893 5 2 1 892
0 894 7 2 2 2850 2855
0 895 5 1 1 2857
0 896 7 1 2 2840 875
0 897 5 1 1 896
0 898 7 2 2 2843 897
0 899 5 1 1 2859
0 900 7 1 2 895 2860
0 901 5 2 1 900
0 902 7 2 2 2844 2861
0 903 5 1 1 2863
0 904 7 1 2 2812 847
0 905 5 1 1 904
0 906 7 2 2 2815 905
0 907 5 1 1 2865
0 908 7 1 2 903 2866
0 909 5 2 1 908
0 910 7 2 2 2816 2867
0 911 5 1 1 2869
0 912 7 1 2 2777 801
0 913 5 1 1 912
0 914 7 2 2 2781 913
0 915 5 1 1 2871
0 916 7 1 2 911 2872
0 917 5 2 1 916
0 918 7 2 2 2002 2118
0 919 5 1 1 2875
0 920 7 2 2 2014 2107
0 921 5 1 1 2877
0 922 7 1 2 2876 2878
0 923 5 2 1 922
0 924 7 1 2 887 891
0 925 5 1 1 924
0 926 7 2 2 2856 925
0 927 5 1 1 2881
0 928 7 1 2 919 921
0 929 5 1 1 928
0 930 7 2 2 2879 929
0 931 5 1 1 2883
0 932 7 1 2 2882 2884
0 933 5 2 1 932
0 934 7 2 2 2880 2885
0 935 5 1 1 2887
0 936 7 1 2 2858 899
0 937 5 1 1 936
0 938 7 2 2 2862 937
0 939 5 1 1 2889
0 940 7 1 2 935 2890
0 941 5 2 1 940
0 942 7 2 2 2026 2086
0 943 5 1 1 2893
0 944 7 2 2 1992 2119
0 945 5 1 1 2895
0 946 7 1 2 2894 2896
0 947 5 2 1 946
0 948 7 2 2 1981 2129
0 949 5 1 1 2899
0 950 7 2 2 2015 2097
0 951 5 1 1 2901
0 952 7 1 2 2039 2075
0 953 5 1 1 952
0 954 7 1 2 2823 953
0 955 5 1 1 954
0 956 7 2 2 2828 955
0 957 5 1 1 2903
0 958 7 1 2 2902 2904
0 959 5 2 1 958
0 960 7 1 2 951 957
0 961 5 1 1 960
0 962 7 2 2 2905 961
0 963 5 1 1 2907
0 964 7 1 2 2900 2908
0 965 5 2 1 964
0 966 7 1 2 949 963
0 967 5 1 1 966
0 968 7 2 2 2909 967
0 969 5 1 1 2911
0 970 7 1 2 943 945
0 971 5 1 1 970
0 972 7 2 2 2897 971
0 973 5 1 1 2913
0 974 7 1 2 2912 2914
0 975 5 2 1 974
0 976 7 2 2 2898 2915
0 977 5 1 1 2917
0 978 7 1 2 927 931
0 979 5 1 1 978
0 980 7 2 2 2886 979
0 981 5 1 1 2919
0 982 7 1 2 977 2920
0 983 5 2 1 982
0 984 7 2 2 2049 2064
0 985 5 1 1 2923
0 986 7 2 2 2003 2108
0 987 5 1 1 2925
0 988 7 1 2 2924 2926
0 989 5 2 1 988
0 990 7 1 2 969 973
0 991 5 1 1 990
0 992 7 2 2 2916 991
0 993 5 1 1 2929
0 994 7 1 2 985 987
0 995 5 1 1 994
0 996 7 2 2 2927 995
0 997 5 1 1 2931
0 998 7 1 2 2930 2932
0 999 5 2 1 998
0 1000 7 2 2 2928 2933
0 1001 5 1 1 2935
0 1002 7 1 2 2918 981
0 1003 5 1 1 1002
0 1004 7 2 2 2921 1003
0 1005 5 1 1 2937
0 1006 7 1 2 1001 2938
0 1007 5 2 1 1006
0 1008 7 2 2 2922 2939
0 1009 5 1 1 2941
0 1010 7 1 2 2888 939
0 1011 5 1 1 1010
0 1012 7 2 2 2891 1011
0 1013 5 1 1 2943
0 1014 7 1 2 1009 2944
0 1015 5 2 1 1014
0 1016 7 2 2 2892 2945
0 1017 5 1 1 2947
0 1018 7 1 2 2864 907
0 1019 5 1 1 1018
0 1020 7 2 2 2868 1019
0 1021 5 1 1 2949
0 1022 7 1 2 1017 2950
0 1023 5 2 1 1022
0 1024 7 2 2 2906 2910
0 1025 5 1 1 2953
0 1026 7 1 2 2936 1005
0 1027 5 1 1 1026
0 1028 7 2 2 2940 1027
0 1029 5 1 1 2955
0 1030 7 1 2 1025 2956
0 1031 5 2 1 1030
0 1032 7 2 2 2027 2076
0 1033 5 1 1 2959
0 1034 7 2 2 2016 2087
0 1035 5 1 1 2961
0 1036 7 1 2 2960 2962
0 1037 5 2 1 1036
0 1038 7 2 2 1982 2120
0 1039 5 1 1 2965
0 1040 7 1 2 1033 1035
0 1041 5 1 1 1040
0 1042 7 2 2 2963 1041
0 1043 5 1 1 2967
0 1044 7 1 2 2966 2968
0 1045 5 2 1 1044
0 1046 7 2 2 2964 2969
0 1047 5 1 1 2971
0 1048 7 2 2 1993 2109
0 1049 5 1 1 2973
0 1050 7 2 2 32 2130
0 1051 5 1 1 2975
0 1052 7 1 2 2974 2976
0 1053 5 2 1 1052
0 1054 7 2 2 2017 2065
0 1055 5 1 1 2979
0 1056 7 2 2 1973 2088
0 1057 5 1 1 2981
0 1058 7 2 2 1994 2066
0 1059 5 1 1 2983
0 1060 7 2 2 2982 2984
0 1061 5 2 1 2985
0 1062 7 2 2 2004 2986
0 1063 5 2 1 2989
0 1064 7 2 2 2980 2990
0 1065 5 2 1 2993
0 1066 7 2 2 2028 2994
0 1067 5 2 1 2997
0 1068 7 2 2 2005 2098
0 1069 5 1 1 3001
0 1070 7 1 2 2998 3002
0 1071 5 2 1 1070
0 1072 7 1 2 2999 1069
0 1073 5 1 1 1072
0 1074 7 2 2 3003 1073
0 1075 5 1 1 3005
0 1076 7 1 2 851 853
0 1077 5 1 1 1076
0 1078 7 2 2 2824 1077
0 1079 5 1 1 3007
0 1080 7 1 2 3006 3008
0 1081 5 2 1 1080
0 1082 7 1 2 1075 1079
0 1083 5 1 1 1082
0 1084 7 2 2 3009 1083
0 1085 5 1 1 3011
0 1086 7 1 2 1049 1051
0 1087 5 1 1 1086
0 1088 7 2 2 2977 1087
0 1089 5 1 1 3013
0 1090 7 1 2 3012 3014
0 1091 5 2 1 1090
0 1092 7 2 2 2978 3015
0 1093 5 1 1 3017
0 1094 7 1 2 1047 1093
0 1095 5 2 1 1094
0 1096 7 2 2 3004 3010
0 1097 5 1 1 3021
0 1098 7 1 2 2972 3018
0 1099 5 1 1 1098
0 1100 7 2 2 3019 1099
0 1101 5 1 1 3023
0 1102 7 1 2 1097 3024
0 1103 5 2 1 1102
0 1104 7 2 2 3020 3025
0 1105 5 1 1 3027
0 1106 7 1 2 2954 1029
0 1107 5 1 1 1106
0 1108 7 2 2 2957 1107
0 1109 5 1 1 3029
0 1110 7 1 2 1105 3030
0 1111 5 2 1 1110
0 1112 7 2 2 2958 3031
0 1113 5 1 1 3033
0 1114 7 1 2 2942 1013
0 1115 5 1 1 1114
0 1116 7 2 2 2946 1115
0 1117 5 1 1 3035
0 1118 7 1 2 1113 3036
0 1119 5 2 1 1118
0 1120 7 1 2 993 997
0 1121 5 1 1 1120
0 1122 7 2 2 2934 1121
0 1123 5 1 1 3039
0 1124 7 1 2 3022 1101
0 1125 5 1 1 1124
0 1126 7 2 2 3026 1125
0 1127 5 1 1 3041
0 1128 7 1 2 3040 3042
0 1129 5 2 1 1128
0 1130 7 1 2 1039 1043
0 1131 5 1 1 1130
0 1132 7 2 2 2970 1131
0 1133 5 1 1 3045
0 1134 7 1 2 1085 1089
0 1135 5 1 1 1134
0 1136 7 2 2 3016 1135
0 1137 5 1 1 3047
0 1138 7 1 2 3046 3048
0 1139 5 2 1 1138
0 1140 7 2 2 2006 2089
0 1141 5 1 1 3051
0 1142 7 2 2 1995 2099
0 1143 5 1 1 3053
0 1144 7 1 2 3052 3054
0 1145 5 2 1 1144
0 1146 7 2 2 1983 2110
0 1147 5 1 1 3057
0 1148 7 1 2 1141 1143
0 1149 5 1 1 1148
0 1150 7 2 2 3055 1149
0 1151 5 1 1 3059
0 1152 7 1 2 3058 3060
0 1153 5 2 1 1152
0 1154 7 2 2 3056 3061
0 1155 5 1 1 3063
0 1156 7 1 2 1133 1137
0 1157 5 1 1 1156
0 1158 7 2 2 3049 1157
0 1159 5 1 1 3065
0 1160 7 1 2 1155 3066
0 1161 5 2 1 1160
0 1162 7 2 2 3050 3067
0 1163 5 1 1 3069
0 1164 7 1 2 1123 1127
0 1165 5 1 1 1164
0 1166 7 2 2 3043 1165
0 1167 5 1 1 3071
0 1168 7 1 2 1163 3072
0 1169 5 2 1 1168
0 1170 7 2 2 3044 3073
0 1171 5 1 1 3075
0 1172 7 1 2 3028 1109
0 1173 5 1 1 1172
0 1174 7 2 2 3032 1173
0 1175 5 1 1 3077
0 1176 7 1 2 1171 3078
0 1177 5 2 1 1176
0 1178 7 2 2 1974 2121
0 1179 5 1 1 3081
0 1180 7 1 2 1147 1151
0 1181 5 1 1 1180
0 1182 7 2 2 3062 1181
0 1183 5 1 1 3083
0 1184 7 1 2 3082 3084
0 1185 5 2 1 1184
0 1186 7 2 2 2040 2054
0 1187 5 1 1 3087
0 1188 7 2 2 2018 2077
0 1189 5 1 1 3089
0 1190 7 1 2 2029 2067
0 1191 5 1 1 1190
0 1192 7 1 2 2995 1191
0 1193 5 1 1 1192
0 1194 7 2 2 3000 1193
0 1195 5 1 1 3091
0 1196 7 1 2 3090 3092
0 1197 5 2 1 1196
0 1198 7 1 2 1189 1195
0 1199 5 1 1 1198
0 1200 7 2 2 3093 1199
0 1201 5 1 1 3095
0 1202 7 1 2 3088 3096
0 1203 5 2 1 1202
0 1204 7 1 2 1187 1201
0 1205 5 1 1 1204
0 1206 7 2 2 3097 1205
0 1207 5 1 1 3099
0 1208 7 1 2 1179 1183
0 1209 5 1 1 1208
0 1210 7 2 2 3085 1209
0 1211 5 1 1 3101
0 1212 7 1 2 3100 3102
0 1213 5 2 1 1212
0 1214 7 2 2 3086 3103
0 1215 5 1 1 3105
0 1216 7 1 2 3064 1159
0 1217 5 1 1 1216
0 1218 7 2 2 3068 1217
0 1219 5 1 1 3107
0 1220 7 1 2 1215 3108
0 1221 5 2 1 1220
0 1222 7 2 2 3094 3098
0 1223 5 1 1 3111
0 1224 7 1 2 3106 1219
0 1225 5 1 1 1224
0 1226 7 2 2 3109 1225
0 1227 5 1 1 3113
0 1228 7 1 2 1223 3114
0 1229 5 2 1 1228
0 1230 7 2 2 3110 3115
0 1231 5 1 1 3117
0 1232 7 1 2 3070 1167
0 1233 5 1 1 1232
0 1234 7 2 2 3074 1233
0 1235 5 1 1 3119
0 1236 7 1 2 1231 3120
0 1237 5 2 1 1236
0 1238 7 2 2 2007 2078
0 1239 5 1 1 3123
0 1240 7 1 2 1055 2991
0 1241 5 1 1 1240
0 1242 7 2 2 2996 1241
0 1243 5 1 1 3125
0 1244 7 1 2 3124 3126
0 1245 5 2 1 1244
0 1246 7 2 2 2030 2055
0 1247 5 1 1 3129
0 1248 7 1 2 1239 1243
0 1249 5 1 1 1248
0 1250 7 2 2 3127 1249
0 1251 5 1 1 3131
0 1252 7 1 2 3130 3132
0 1253 5 2 1 1252
0 1254 7 2 2 3128 3133
0 1255 5 1 1 3135
0 1256 7 1 2 1207 1211
0 1257 5 1 1 1256
0 1258 7 2 2 3104 1257
0 1259 5 1 1 3137
0 1260 7 1 2 1255 3138
0 1261 5 2 1 1260
0 1262 7 2 2 1996 2090
0 1263 5 1 1 3141
0 1264 7 2 2 1975 2111
0 1265 5 1 1 3143
0 1266 7 1 2 3142 3144
0 1267 5 2 1 1266
0 1268 7 1 2 1247 1251
0 1269 5 1 1 1268
0 1270 7 2 2 3134 1269
0 1271 5 1 1 3147
0 1272 7 1 2 1263 1265
0 1273 5 1 1 1272
0 1274 7 2 2 3145 1273
0 1275 5 1 1 3149
0 1276 7 1 2 3148 3150
0 1277 5 2 1 1276
0 1278 7 2 2 3146 3151
0 1279 5 1 1 3153
0 1280 7 1 2 3136 1259
0 1281 5 1 1 1280
0 1282 7 2 2 3139 1281
0 1283 5 1 1 3155
0 1284 7 1 2 1279 3156
0 1285 5 2 1 1284
0 1286 7 2 2 3140 3157
0 1287 5 1 1 3159
0 1288 7 1 2 3112 1227
0 1289 5 1 1 1288
0 1290 7 2 2 3116 1289
0 1291 5 1 1 3161
0 1292 7 1 2 1287 3162
0 1293 5 2 1 1292
0 1294 7 2 2 1984 2100
0 1295 5 1 1 3165
0 1296 7 1 2 1271 1275
0 1297 5 1 1 1296
0 1298 7 2 2 3152 1297
0 1299 5 1 1 3167
0 1300 7 1 2 3166 3168
0 1301 5 2 1 1300
0 1302 7 2 2 1997 2079
0 1303 5 1 1 3171
0 1304 7 1 2 2008 2068
0 1305 5 1 1 1304
0 1306 7 1 2 2987 1305
0 1307 5 1 1 1306
0 1308 7 2 2 2992 1307
0 1309 5 1 1 3173
0 1310 7 1 2 3172 3174
0 1311 5 2 1 1310
0 1312 7 2 2 2019 2056
0 1313 5 1 1 3177
0 1314 7 1 2 1303 1309
0 1315 5 1 1 1314
0 1316 7 2 2 3175 1315
0 1317 5 1 1 3179
0 1318 7 1 2 3178 3180
0 1319 5 2 1 1318
0 1320 7 2 2 3176 3181
0 1321 5 1 1 3183
0 1322 7 1 2 1295 1299
0 1323 5 1 1 1322
0 1324 7 2 2 3169 1323
0 1325 5 1 1 3185
0 1326 7 1 2 1321 3186
0 1327 5 2 1 1326
0 1328 7 2 2 3170 3187
0 1329 5 1 1 3189
0 1330 7 1 2 3154 1283
0 1331 5 1 1 1330
0 1332 7 2 2 3158 1331
0 1333 5 1 1 3191
0 1334 7 1 2 1329 3192
0 1335 5 2 1 1334
0 1336 7 2 2 1976 2101
0 1337 5 1 1 3195
0 1338 7 2 2 1985 2091
0 1339 5 1 1 3197
0 1340 7 1 2 3196 3198
0 1341 5 2 1 1340
0 1342 7 1 2 1313 1317
0 1343 5 1 1 1342
0 1344 7 2 2 3182 1343
0 1345 5 1 1 3201
0 1346 7 1 2 1337 1339
0 1347 5 1 1 1346
0 1348 7 2 2 3199 1347
0 1349 5 1 1 3203
0 1350 7 1 2 3202 3204
0 1351 5 2 1 1350
0 1352 7 2 2 3200 3205
0 1353 5 1 1 3207
0 1354 7 1 2 3184 1325
0 1355 5 1 1 1354
0 1356 7 2 2 3188 1355
0 1357 5 1 1 3209
0 1358 7 1 2 1353 3210
0 1359 5 2 1 1358
0 1360 7 1 2 1345 1349
0 1361 5 1 1 1360
0 1362 7 2 2 3206 1361
0 1363 5 1 1 3213
0 1364 7 2 2 1986 2080
0 1365 5 1 1 3215
0 1366 7 2 2 2009 2057
0 1367 5 1 1 3217
0 1368 7 2 2 3216 3218
0 1369 5 1 1 3219
0 1370 7 2 2 1987 2069
0 1371 5 1 1 3221
0 1372 7 2 2 1977 2081
0 1373 5 1 1 3223
0 1374 7 2 2 3222 3224
0 1375 5 2 1 3225
0 1376 7 3 2 1369 3227
0 1377 5 1 1 3229
0 1378 7 1 2 3214 1377
0 1379 5 2 1 1378
0 1380 7 1 2 1057 1059
0 1381 5 1 1 1380
0 1382 7 2 2 2988 1381
0 1383 5 1 1 3234
0 1384 7 1 2 1365 1367
0 1385 5 1 1 1384
0 1386 7 1 2 3230 1385
0 1387 5 1 1 1386
0 1388 7 1 2 3220 3226
0 1389 5 1 1 1388
0 1390 7 2 2 1387 1389
0 1391 5 1 1 3236
0 1392 7 1 2 3235 1391
0 1393 5 2 1 1392
0 1394 7 2 2 1998 2058
0 1395 5 1 1 3240
0 1396 7 1 2 1371 1373
0 1397 5 1 1 1396
0 1398 7 2 2 3228 1397
0 1399 5 1 1 3242
0 1400 7 1 2 3241 3243
0 1401 5 2 1 1400
0 1402 7 1 2 1395 1399
0 1403 5 1 1 1402
0 1404 7 2 2 3244 1403
0 1405 5 1 1 3246
0 1406 7 2 2 1978 2070
0 1407 5 1 1 3248
0 1408 7 2 2 1988 2059
0 1409 5 1 1 3250
0 1410 7 2 2 3249 3251
0 1411 5 2 1 3252
0 1412 7 1 2 3247 3253
0 1413 5 2 1 1412
0 1414 7 2 2 3245 3256
0 1415 5 1 1 3258
0 1416 7 1 2 1383 3237
0 1417 5 1 1 1416
0 1418 7 2 2 3238 1417
0 1419 5 1 1 3260
0 1420 7 1 2 1415 3261
0 1421 5 2 1 1420
0 1422 7 2 2 3239 3262
0 1423 5 1 1 3264
0 1424 7 1 2 1363 3231
0 1425 5 1 1 1424
0 1426 7 2 2 3232 1425
0 1427 5 1 1 3266
0 1428 7 1 2 1423 3267
0 1429 5 2 1 1428
0 1430 7 2 2 3233 3268
0 1431 5 1 1 3270
0 1432 7 1 2 3208 1357
0 1433 5 1 1 1432
0 1434 7 2 2 3211 1433
0 1435 5 1 1 3272
0 1436 7 1 2 1431 3273
0 1437 5 2 1 1436
0 1438 7 2 2 3212 3274
0 1439 5 1 1 3276
0 1440 7 1 2 3190 1333
0 1441 5 1 1 1440
0 1442 7 2 2 3193 1441
0 1443 5 1 1 3278
0 1444 7 1 2 1439 3279
0 1445 5 2 1 1444
0 1446 7 2 2 3194 3280
0 1447 5 1 1 3282
0 1448 7 1 2 3160 1291
0 1449 5 1 1 1448
0 1450 7 2 2 3163 1449
0 1451 5 1 1 3284
0 1452 7 1 2 1447 3285
0 1453 5 2 1 1452
0 1454 7 2 2 3164 3286
0 1455 5 1 1 3288
0 1456 7 1 2 3118 1235
0 1457 5 1 1 1456
0 1458 7 2 2 3121 1457
0 1459 5 1 1 3290
0 1460 7 1 2 1455 3291
0 1461 5 2 1 1460
0 1462 7 2 2 3122 3292
0 1463 5 1 1 3294
0 1464 7 1 2 3076 1175
0 1465 5 1 1 1464
0 1466 7 2 2 3079 1465
0 1467 5 1 1 3296
0 1468 7 1 2 1463 3297
0 1469 5 2 1 1468
0 1470 7 2 2 3080 3298
0 1471 5 1 1 3300
0 1472 7 1 2 3034 1117
0 1473 5 1 1 1472
0 1474 7 2 2 3037 1473
0 1475 5 1 1 3302
0 1476 7 1 2 1471 3303
0 1477 5 2 1 1476
0 1478 7 2 2 3038 3304
0 1479 5 1 1 3306
0 1480 7 1 2 2948 1021
0 1481 5 1 1 1480
0 1482 7 2 2 2951 1481
0 1483 5 1 1 3308
0 1484 7 1 2 1479 3309
0 1485 5 2 1 1484
0 1486 7 2 2 2952 3310
0 1487 5 1 1 3312
0 1488 7 1 2 2870 915
0 1489 5 1 1 1488
0 1490 7 2 2 2873 1489
0 1491 5 1 1 3314
0 1492 7 1 2 1487 3315
0 1493 5 2 1 1492
0 1494 7 2 2 2874 3316
0 1495 5 1 1 3318
0 1496 7 1 2 2783 823
0 1497 5 1 1 1496
0 1498 7 2 2 2797 1497
0 1499 5 1 1 3320
0 1500 7 1 2 1495 3321
0 1501 5 2 1 1500
0 1502 7 2 2 2798 3322
0 1503 5 1 1 3324
0 1504 7 2 2 2050 2131
0 1505 5 1 1 3326
0 1506 7 1 2 2737 2793
0 1507 5 1 1 1506
0 1508 7 1 2 3327 1507
0 1509 5 2 1 1508
0 1510 7 1 2 2794 1505
0 1511 5 1 1 1510
0 1512 7 2 2 3328 1511
0 1513 5 1 1 3330
0 1514 7 1 2 1503 3331
0 1515 5 2 1 1514
0 1516 7 1 2 3325 1513
0 1517 5 1 1 1516
0 1518 7 2 2 3332 1517
0 1519 5 1 1 3334
0 1520 7 1 2 2178 1519
0 1521 5 3 1 1520
0 1522 7 2 2 3329 3333
0 1523 5 1 1 3339
0 1524 7 2 2 2182 3340
0 1525 5 1 1 3341
0 1526 7 2 2 3336 1525
0 1527 5 1 1 3343
0 1528 7 2 2 2257 1523
0 1529 5 2 1 3345
0 1530 7 1 2 1527 3347
0 1531 5 2 1 1530
0 1532 7 1 2 3319 1499
0 1533 5 1 1 1532
0 1534 7 2 2 3323 1533
0 1535 5 1 1 3351
0 1536 7 1 2 2174 1535
0 1537 5 3 1 1536
0 1538 7 1 2 2253 3352
0 1539 5 4 1 1538
0 1540 7 1 2 3313 1491
0 1541 5 1 1 1540
0 1542 7 2 2 3317 1541
0 1543 5 1 1 3360
0 1544 7 1 2 2171 1543
0 1545 5 5 1 1544
0 1546 7 1 2 2250 3361
0 1547 5 2 1 1546
0 1548 7 1 2 3307 1483
0 1549 5 1 1 1548
0 1550 7 2 2 3311 1549
0 1551 5 1 1 3369
0 1552 7 1 2 2246 3370
0 1553 5 4 1 1552
0 1554 7 3 2 3367 3371
0 1555 7 1 2 2167 1551
0 1556 5 4 1 1555
0 1557 7 1 2 3301 1475
0 1558 5 1 1 1557
0 1559 7 2 2 3305 1558
0 1560 5 1 1 3382
0 1561 7 1 2 2164 1560
0 1562 5 4 1 1561
0 1563 7 1 2 2243 3383
0 1564 5 4 1 1563
0 1565 7 1 2 3295 1467
0 1566 5 1 1 1565
0 1567 7 2 2 3299 1566
0 1568 5 1 1 3392
0 1569 7 1 2 2161 1568
0 1570 5 5 1 1569
0 1571 7 1 2 2240 3393
0 1572 5 5 1 1571
0 1573 7 1 2 3289 1459
0 1574 5 1 1 1573
0 1575 7 2 2 3293 1574
0 1576 5 1 1 3404
0 1577 7 1 2 2158 1576
0 1578 5 4 1 1577
0 1579 7 1 2 2237 3405
0 1580 5 4 1 1579
0 1581 7 1 2 3283 1451
0 1582 5 1 1 1581
0 1583 7 2 2 3287 1582
0 1584 5 1 1 3414
0 1585 7 1 2 2155 1584
0 1586 5 3 1 1585
0 1587 7 1 2 2234 3415
0 1588 5 4 1 1587
0 1589 7 1 2 3277 1443
0 1590 5 1 1 1589
0 1591 7 2 2 3281 1590
0 1592 5 1 1 3423
0 1593 7 1 2 2152 1592
0 1594 5 3 1 1593
0 1595 7 1 2 2231 3424
0 1596 5 4 1 1595
0 1597 7 1 2 3271 1435
0 1598 5 1 1 1597
0 1599 7 2 2 3275 1598
0 1600 5 1 1 3432
0 1601 7 1 2 2149 1600
0 1602 5 4 1 1601
0 1603 7 1 2 2228 3433
0 1604 5 4 1 1603
0 1605 7 1 2 3265 1427
0 1606 5 1 1 1605
0 1607 7 2 2 3269 1606
0 1608 5 1 1 3442
0 1609 7 1 2 2146 1608
0 1610 5 4 1 1609
0 1611 7 1 2 2225 3443
0 1612 5 4 1 1611
0 1613 7 1 2 3259 1419
0 1614 5 1 1 1613
0 1615 7 2 2 3263 1614
0 1616 5 1 1 3452
0 1617 7 1 2 2143 1616
0 1618 5 4 1 1617
0 1619 7 1 2 2222 3453
0 1620 5 4 1 1619
0 1621 7 1 2 1405 3254
0 1622 5 1 1 1621
0 1623 7 2 2 3257 1622
0 1624 5 1 1 3462
0 1625 7 1 2 2219 3463
0 1626 5 4 1 1625
0 1627 7 1 2 2140 1624
0 1628 5 4 1 1627
0 1629 7 1 2 1407 1409
0 1630 5 1 1 1629
0 1631 7 2 2 3255 1630
0 1632 5 1 1 3472
0 1633 7 1 2 2216 3473
0 1634 5 2 1 1633
0 1635 7 1 2 2137 1632
0 1636 5 2 1 1635
0 1637 7 2 2 1979 2060
0 1638 5 1 1 3478
0 1639 7 1 2 2134 1638
0 1640 5 1 1 1639
0 1641 7 2 2 3476 1640
0 1642 5 1 1 3480
0 1643 7 1 2 3474 1642
0 1644 5 3 1 1643
0 1645 7 1 2 3468 3482
0 1646 5 1 1 1645
0 1647 7 3 2 3464 1646
0 1648 5 1 1 3485
0 1649 7 1 2 3458 3486
0 1650 5 1 1 1649
0 1651 7 2 2 3454 1650
0 1652 5 1 1 3488
0 1653 7 2 2 3448 1652
0 1654 5 1 1 3490
0 1655 7 2 2 3444 1654
0 1656 5 2 1 3492
0 1657 7 1 2 3438 3494
0 1658 5 1 1 1657
0 1659 7 2 2 3434 1658
0 1660 5 2 1 3496
0 1661 7 1 2 3428 3498
0 1662 5 1 1 1661
0 1663 7 2 2 3425 1662
0 1664 5 2 1 3500
0 1665 7 1 2 3419 3502
0 1666 5 1 1 1665
0 1667 7 2 2 3416 1666
0 1668 5 2 1 3504
0 1669 7 1 2 3410 3506
0 1670 5 1 1 1669
0 1671 7 2 2 3406 1670
0 1672 5 1 1 3508
0 1673 7 1 2 3399 1672
0 1674 5 1 1 1673
0 1675 7 1 2 3394 1674
0 1676 5 1 1 1675
0 1677 7 2 2 3388 1676
0 1678 5 1 1 3510
0 1679 7 3 2 3384 1678
0 1680 5 1 1 3512
0 1681 7 1 2 3378 3513
0 1682 5 1 1 1681
0 1683 7 1 2 3375 1682
0 1684 5 1 1 1683
0 1685 7 2 2 3362 1684
0 1686 5 2 1 3515
0 1687 7 1 2 3356 3517
0 1688 5 1 1 1687
0 1689 7 2 2 3353 1688
0 1690 5 2 1 3519
0 1691 7 1 2 2255 3335
0 1692 5 3 1 1691
0 1693 7 3 2 3523 3348
0 1694 5 1 1 3526
0 1695 7 1 2 3521 3527
0 1696 5 1 1 1695
0 1697 7 2 2 3349 1696
0 1698 5 1 1 3529
0 1699 7 1 2 2213 3479
0 1700 5 1 1 1699
0 1701 7 3 2 3475 1700
0 1702 5 2 1 3531
0 1703 7 2 2 3477 3534
0 1704 5 1 1 3536
0 1705 7 1 2 3465 1704
0 1706 5 1 1 1705
0 1707 7 1 2 3469 1706
0 1708 5 1 1 1707
0 1709 7 2 2 3459 1708
0 1710 5 1 1 3538
0 1711 7 2 2 3455 1710
0 1712 5 2 1 3540
0 1713 7 1 2 3449 3542
0 1714 5 1 1 1713
0 1715 7 2 2 3445 1714
0 1716 5 1 1 3544
0 1717 7 2 2 3439 1716
0 1718 5 1 1 3546
0 1719 7 2 2 3435 1718
0 1720 5 2 1 3548
0 1721 7 1 2 3429 3550
0 1722 5 1 1 1721
0 1723 7 2 2 3426 1722
0 1724 5 2 1 3552
0 1725 7 1 2 3420 3554
0 1726 5 1 1 1725
0 1727 7 2 2 3417 1726
0 1728 5 1 1 3556
0 1729 7 2 2 3411 1728
0 1730 5 1 1 3558
0 1731 7 1 2 3407 1730
0 1732 5 2 1 1731
0 1733 7 1 2 3400 3560
0 1734 5 1 1 1733
0 1735 7 2 2 3395 1734
0 1736 5 1 1 3562
0 1737 7 1 2 3389 1736
0 1738 5 1 1 1737
0 1739 7 3 2 3385 1738
0 1740 5 2 1 3564
0 1741 7 1 2 3379 3565
0 1742 5 1 1 1741
0 1743 7 2 2 3376 1742
0 1744 5 1 1 3569
0 1745 7 1 2 3363 1744
0 1746 5 2 1 1745
0 1747 7 1 2 3357 3571
0 1748 5 1 1 1747
0 1749 7 2 2 3354 1748
0 1750 5 1 1 3573
0 1751 7 1 2 3337 3524
0 1752 5 3 1 1751
0 1753 7 1 2 1750 3575
0 1754 5 1 1 1753
0 1755 7 1 2 3525 3342
0 1756 5 1 1 1755
0 1757 7 3 2 3355 3358
0 1758 5 2 1 3578
0 1759 7 1 2 3572 3581
0 1760 5 1 1 1759
0 1761 7 2 2 3372 3380
0 1762 5 2 1 3583
0 1763 7 1 2 3566 3585
0 1764 5 1 1 1763
0 1765 7 1 2 3567 3584
0 1766 5 1 1 1765
0 1767 7 1 2 1764 1766
0 1768 5 1 1 1767
0 1769 7 3 2 3386 3390
0 1770 5 2 1 3587
0 1771 7 1 2 3396 3588
0 1772 5 1 1 1771
0 1773 7 1 2 3561 1772
0 1774 5 1 1 1773
0 1775 7 1 2 3401 3590
0 1776 5 1 1 1775
0 1777 7 1 2 3563 3589
0 1778 5 1 1 1777
0 1779 7 1 2 3408 3559
0 1780 5 1 1 1779
0 1781 7 2 2 3409 3412
0 1782 5 2 1 3592
0 1783 7 1 2 3557 3594
0 1784 5 1 1 1783
0 1785 7 3 2 3418 3421
0 1786 5 2 1 3596
0 1787 7 1 2 3553 3597
0 1788 5 1 1 1787
0 1789 7 1 2 3555 3599
0 1790 5 1 1 1789
0 1791 7 3 2 3427 3430
0 1792 5 2 1 3601
0 1793 7 1 2 3549 3602
0 1794 5 1 1 1793
0 1795 7 1 2 3436 3547
0 1796 5 1 1 1795
0 1797 7 2 2 3437 3440
0 1798 5 2 1 3606
0 1799 7 1 2 3545 3608
0 1800 5 1 1 1799
0 1801 7 2 2 3446 3450
0 1802 5 2 1 3610
0 1803 7 1 2 3541 3611
0 1804 5 1 1 1803
0 1805 7 1 2 3456 3539
0 1806 5 1 1 1805
0 1807 7 2 2 3457 3460
0 1808 5 2 1 3614
0 1809 7 1 2 3470 3616
0 1810 5 1 1 1809
0 1811 7 2 2 3471 3466
0 1812 5 2 1 3618
0 1813 7 1 2 3537 3620
0 1814 5 1 1 1813
0 1815 7 1 2 3532 3481
0 1816 5 1 1 1815
0 1817 7 1 2 1814 1816
0 1818 7 1 2 1810 1817
0 1819 7 1 2 1806 1818
0 1820 5 1 1 1819
0 1821 7 1 2 3543 3612
0 1822 5 1 1 1821
0 1823 7 1 2 1820 1822
0 1824 7 1 2 1804 1823
0 1825 5 1 1 1824
0 1826 7 1 2 1800 1825
0 1827 7 1 2 1796 1826
0 1828 5 1 1 1827
0 1829 7 1 2 3551 3604
0 1830 5 1 1 1829
0 1831 7 1 2 1828 1830
0 1832 7 1 2 1794 1831
0 1833 7 1 2 1790 1832
0 1834 7 1 2 1788 1833
0 1835 5 1 1 1834
0 1836 7 1 2 1784 1835
0 1837 7 1 2 1780 1836
0 1838 5 1 1 1837
0 1839 7 1 2 1778 1838
0 1840 7 1 2 1776 1839
0 1841 7 1 2 1774 1840
0 1842 7 1 2 1768 1841
0 1843 7 1 2 1760 1842
0 1844 7 1 2 1756 1843
0 1845 7 1 2 1754 1844
0 1846 7 1 2 3574 3344
0 1847 5 1 1 1846
0 1848 7 1 2 3364 3570
0 1849 5 1 1 1848
0 1850 7 1 2 3365 3579
0 1851 5 1 1 1850
0 1852 7 2 2 3366 3368
0 1853 5 1 1 3622
0 1854 7 2 2 3381 1853
0 1855 5 1 1 3624
0 1856 7 1 2 3373 3568
0 1857 5 1 1 1856
0 1858 7 1 2 3625 1857
0 1859 7 1 2 1851 1858
0 1860 5 1 1 1859
0 1861 7 1 2 1849 1860
0 1862 5 1 1 1861
0 1863 7 1 2 1847 1862
0 1864 7 1 2 1845 1863
0 1865 7 1 2 1698 1864
0 1866 5 1 1 1865
0 1867 7 1 2 3576 1694
0 1868 5 1 1 1867
0 1869 7 1 2 3522 1868
0 1870 5 1 1 1869
0 1871 7 1 2 3338 3346
0 1872 5 1 1 1871
0 1873 7 1 2 3582 3516
0 1874 5 1 1 1873
0 1875 7 1 2 3580 3518
0 1876 5 1 1 1875
0 1877 7 1 2 3374 1680
0 1878 7 1 2 3623 1877
0 1879 5 1 1 1878
0 1880 7 1 2 3586 3514
0 1881 5 1 1 1880
0 1882 7 1 2 3387 3511
0 1883 5 1 1 1882
0 1884 7 1 2 3397 3591
0 1885 5 1 1 1884
0 1886 7 1 2 3593 3505
0 1887 5 1 1 1886
0 1888 7 1 2 3600 3501
0 1889 5 1 1 1888
0 1890 7 1 2 3598 3503
0 1891 5 1 1 1890
0 1892 7 1 2 3605 3497
0 1893 5 1 1 1892
0 1894 7 1 2 3447 3491
0 1895 5 1 1 1894
0 1896 7 1 2 3613 3489
0 1897 5 1 1 1896
0 1898 7 1 2 3617 3487
0 1899 5 1 1 1898
0 1900 7 1 2 3615 1648
0 1901 5 1 1 1900
0 1902 7 1 2 3619 3483
0 1903 5 1 1 1902
0 1904 7 1 2 3535 3484
0 1905 5 1 1 1904
0 1906 7 1 2 3621 1905
0 1907 5 1 1 1906
0 1908 7 1 2 1903 1907
0 1909 7 1 2 1901 1908
0 1910 7 1 2 1899 1909
0 1911 5 1 1 1910
0 1912 7 1 2 1897 1911
0 1913 7 1 2 1895 1912
0 1914 5 1 1 1913
0 1915 7 1 2 3607 3495
0 1916 5 1 1 1915
0 1917 7 1 2 3609 3493
0 1918 5 1 1 1917
0 1919 7 1 2 1916 1918
0 1920 5 1 1 1919
0 1921 7 1 2 1914 1920
0 1922 5 1 1 1921
0 1923 7 1 2 3603 3499
0 1924 5 1 1 1923
0 1925 7 1 2 1922 1924
0 1926 7 1 2 1893 1925
0 1927 7 1 2 1891 1926
0 1928 7 1 2 1889 1927
0 1929 5 1 1 1928
0 1930 7 1 2 3595 3507
0 1931 5 1 1 1930
0 1932 7 1 2 1929 1931
0 1933 7 1 2 1887 1932
0 1934 5 1 1 1933
0 1935 7 1 2 3398 3402
0 1936 5 1 1 1935
0 1937 7 1 2 3509 1936
0 1938 5 1 1 1937
0 1939 7 1 2 1934 1938
0 1940 7 1 2 1885 1939
0 1941 7 1 2 1883 1940
0 1942 7 1 2 1881 1941
0 1943 7 1 2 1855 1942
0 1944 7 1 2 1879 1943
0 1945 7 1 2 1876 1944
0 1946 7 1 2 1874 1945
0 1947 7 1 2 1872 1946
0 1948 7 1 2 3577 3520
0 1949 5 1 1 1948
0 1950 7 1 2 3350 1949
0 1951 7 1 2 1947 1950
0 1952 7 1 2 1870 1951
0 1953 5 1 1 1952
0 1954 7 1 2 1866 1953
0 1955 7 1 2 729 1954
0 1956 5 1 1 1955
0 1957 7 1 2 3467 3533
0 1958 7 1 2 3461 1957
0 1959 7 1 2 3451 1958
0 1960 7 1 2 3441 1959
0 1961 7 1 2 3431 1960
0 1962 7 1 2 3422 1961
0 1963 7 1 2 3413 1962
0 1964 7 1 2 3403 1963
0 1965 7 1 2 3391 1964
0 1966 7 1 2 3377 1965
0 1967 7 1 2 3359 1966
0 1968 7 1 2 3528 1967
0 1969 7 1 2 3530 1968
0 1970 5 1 1 1969
0 1971 7 1 2 2719 1970
0 1972 5 1 1 1971
3 4099 7 0 2 1956 1972
