1 0 0 2 0
2 49 1 0
2 1812 1 0
1 1 0 3 0
2 1813 1 1
2 1814 1 1
2 1815 1 1
1 2 0 3 0
2 1816 1 2
2 1817 1 2
2 1818 1 2
1 3 0 3 0
2 1819 1 3
2 1820 1 3
2 1821 1 3
1 4 0 3 0
2 1822 1 4
2 1823 1 4
2 1824 1 4
1 5 0 3 0
2 1825 1 5
2 1826 1 5
2 1827 1 5
1 6 0 3 0
2 1828 1 6
2 1829 1 6
2 1830 1 6
1 7 0 3 0
2 1831 1 7
2 1832 1 7
2 1833 1 7
1 8 0 3 0
2 1834 1 8
2 1835 1 8
2 1836 1 8
1 9 0 3 0
2 1837 1 9
2 1838 1 9
2 1839 1 9
1 10 0 3 0
2 1840 1 10
2 1841 1 10
2 1842 1 10
1 11 0 3 0
2 1843 1 11
2 1844 1 11
2 1845 1 11
1 12 0 3 0
2 1846 1 12
2 1847 1 12
2 1848 1 12
1 13 0 3 0
2 1849 1 13
2 1850 1 13
2 1851 1 13
1 14 0 3 0
2 1852 1 14
2 1853 1 14
2 1854 1 14
1 15 0 3 0
2 1855 1 15
2 1856 1 15
2 1857 1 15
1 16 0 3 0
2 1858 1 16
2 1859 1 16
2 1860 1 16
1 17 0 3 0
2 1861 1 17
2 1862 1 17
2 1863 1 17
1 18 0 3 0
2 1864 1 18
2 1865 1 18
2 1866 1 18
1 19 0 3 0
2 1867 1 19
2 1868 1 19
2 1869 1 19
1 20 0 3 0
2 1870 1 20
2 1871 1 20
2 1872 1 20
1 21 0 3 0
2 1873 1 21
2 1874 1 21
2 1875 1 21
1 22 0 3 0
2 1876 1 22
2 1877 1 22
2 1878 1 22
1 23 0 3 0
2 1879 1 23
2 1880 1 23
2 1881 1 23
1 24 0 3 0
2 1882 1 24
2 1883 1 24
2 1884 1 24
1 25 0 3 0
2 1885 1 25
2 1886 1 25
2 1887 1 25
1 26 0 3 0
2 1888 1 26
2 1889 1 26
2 1890 1 26
1 27 0 3 0
2 1891 1 27
2 1892 1 27
2 1893 1 27
1 28 0 3 0
2 1894 1 28
2 1895 1 28
2 1896 1 28
1 29 0 3 0
2 1897 1 29
2 1898 1 29
2 1899 1 29
1 30 0 3 0
2 1900 1 30
2 1901 1 30
2 1902 1 30
1 31 0 3 0
2 1903 1 31
2 1904 1 31
2 1905 1 31
1 32 0 3 0
2 1906 1 32
2 1907 1 32
2 1908 1 32
1 33 0 3 0
2 1909 1 33
2 1910 1 33
2 1911 1 33
1 34 0 3 0
2 1912 1 34
2 1913 1 34
2 1914 1 34
1 35 0 3 0
2 1915 1 35
2 1916 1 35
2 1917 1 35
1 36 0 3 0
2 1918 1 36
2 1919 1 36
2 1920 1 36
1 37 0 3 0
2 1921 1 37
2 1922 1 37
2 1923 1 37
1 38 0 3 0
2 1924 1 38
2 1925 1 38
2 1926 1 38
1 39 0 3 0
2 1927 1 39
2 1928 1 39
2 1929 1 39
1 40 0 3 0
2 1930 1 40
2 1931 1 40
2 1932 1 40
1 41 0 3 0
2 1933 1 41
2 1934 1 41
2 1935 1 41
1 42 0 3 0
2 1936 1 42
2 1937 1 42
2 1938 1 42
1 43 0 3 0
2 1939 1 43
2 1940 1 43
2 1941 1 43
1 44 0 3 0
2 1942 1 44
2 1943 1 44
2 1944 1 44
1 45 0 4 0
2 1945 1 45
2 1946 1 45
2 1947 1 45
2 1948 1 45
1 46 0 3 0
2 1949 1 46
2 1950 1 46
2 1951 1 46
1 47 0 4 0
2 1952 1 47
2 1953 1 47
2 1954 1 47
2 1955 1 47
1 48 0 4 0
2 1956 1 48
2 1957 1 48
2 1958 1 48
2 1959 1 48
2 1960 1 51
2 1961 1 51
2 1962 1 52
2 1963 1 52
2 1964 1 52
2 1965 1 53
2 1966 1 53
2 1967 1 53
2 1968 1 54
2 1969 1 54
2 1970 1 54
2 1971 1 55
2 1972 1 55
2 1973 1 55
2 1974 1 56
2 1975 1 56
2 1976 1 56
2 1977 1 57
2 1978 1 57
2 1979 1 57
2 1980 1 58
2 1981 1 58
2 1982 1 58
2 1983 1 59
2 1984 1 59
2 1985 1 59
2 1986 1 60
2 1987 1 60
2 1988 1 60
2 1989 1 61
2 1990 1 61
2 1991 1 61
2 1992 1 62
2 1993 1 62
2 1994 1 62
2 1995 1 63
2 1996 1 63
2 1997 1 63
2 1998 1 64
2 1999 1 64
2 2000 1 64
2 2001 1 65
2 2002 1 65
2 2003 1 65
2 2004 1 66
2 2005 1 66
2 2006 1 66
2 2007 1 67
2 2008 1 67
2 2009 1 67
2 2010 1 68
2 2011 1 68
2 2012 1 68
2 2013 1 69
2 2014 1 69
2 2015 1 69
2 2016 1 69
2 2017 1 70
2 2018 1 70
2 2019 1 70
2 2020 1 70
2 2021 1 71
2 2022 1 71
2 2023 1 71
2 2024 1 71
2 2025 1 72
2 2026 1 72
2 2027 1 72
2 2028 1 72
2 2029 1 73
2 2030 1 73
2 2031 1 73
2 2032 1 73
2 2033 1 74
2 2034 1 74
2 2035 1 74
2 2036 1 74
2 2037 1 75
2 2038 1 75
2 2039 1 75
2 2040 1 75
2 2041 1 76
2 2042 1 76
2 2043 1 76
2 2044 1 76
2 2045 1 77
2 2046 1 77
2 2047 1 77
2 2048 1 77
2 2049 1 78
2 2050 1 78
2 2051 1 78
2 2052 1 78
2 2053 1 79
2 2054 1 79
2 2055 1 79
2 2056 1 79
2 2057 1 80
2 2058 1 80
2 2059 1 80
2 2060 1 80
2 2061 1 81
2 2062 1 81
2 2063 1 81
2 2064 1 81
2 2065 1 82
2 2066 1 82
2 2067 1 82
2 2068 1 83
2 2069 1 83
2 2070 1 83
2 2071 1 84
2 2072 1 84
2 2073 1 84
2 2074 1 85
2 2075 1 85
2 2076 1 85
2 2077 1 86
2 2078 1 86
2 2079 1 86
2 2080 1 87
2 2081 1 87
2 2082 1 87
2 2083 1 88
2 2084 1 88
2 2085 1 88
2 2086 1 89
2 2087 1 89
2 2088 1 89
2 2089 1 90
2 2090 1 90
2 2091 1 90
2 2092 1 91
2 2093 1 91
2 2094 1 91
2 2095 1 92
2 2096 1 92
2 2097 1 92
2 2098 1 93
2 2099 1 93
2 2100 1 93
2 2101 1 94
2 2102 1 94
2 2103 1 94
2 2104 1 95
2 2105 1 95
2 2106 1 95
2 2107 1 95
2 2108 1 96
2 2109 1 96
2 2110 1 96
2 2111 1 97
2 2112 1 97
2 2113 1 98
2 2114 1 98
2 2115 1 99
2 2116 1 99
2 2117 1 101
2 2118 1 101
2 2119 1 101
2 2120 1 103
2 2121 1 103
2 2122 1 109
2 2123 1 109
2 2124 1 111
2 2125 1 111
2 2126 1 116
2 2127 1 116
2 2128 1 119
2 2129 1 119
2 2130 1 122
2 2131 1 122
2 2132 1 124
2 2133 1 124
2 2134 1 125
2 2135 1 125
2 2136 1 130
2 2137 1 130
2 2138 1 133
2 2139 1 133
2 2140 1 138
2 2141 1 138
2 2142 1 139
2 2143 1 139
2 2144 1 140
2 2145 1 140
2 2146 1 143
2 2147 1 143
2 2148 1 146
2 2149 1 146
2 2150 1 148
2 2151 1 148
2 2152 1 149
2 2153 1 149
2 2154 1 154
2 2155 1 154
2 2156 1 157
2 2157 1 157
2 2158 1 162
2 2159 1 162
2 2160 1 162
2 2161 1 164
2 2162 1 164
2 2163 1 167
2 2164 1 167
2 2165 1 170
2 2166 1 170
2 2167 1 172
2 2168 1 172
2 2169 1 173
2 2170 1 173
2 2171 1 178
2 2172 1 178
2 2173 1 181
2 2174 1 181
2 2175 1 186
2 2176 1 186
2 2177 1 186
2 2178 1 188
2 2179 1 188
2 2180 1 191
2 2181 1 191
2 2182 1 194
2 2183 1 194
2 2184 1 196
2 2185 1 196
2 2186 1 197
2 2187 1 197
2 2188 1 202
2 2189 1 202
2 2190 1 205
2 2191 1 205
2 2192 1 210
2 2193 1 210
2 2194 1 210
2 2195 1 212
2 2196 1 212
2 2197 1 215
2 2198 1 215
2 2199 1 218
2 2200 1 218
2 2201 1 220
2 2202 1 220
2 2203 1 221
2 2204 1 221
2 2205 1 226
2 2206 1 226
2 2207 1 229
2 2208 1 229
2 2209 1 234
2 2210 1 234
2 2211 1 234
2 2212 1 236
2 2213 1 236
2 2214 1 239
2 2215 1 239
2 2216 1 242
2 2217 1 242
2 2218 1 244
2 2219 1 244
2 2220 1 245
2 2221 1 245
2 2222 1 250
2 2223 1 250
2 2224 1 253
2 2225 1 253
2 2226 1 258
2 2227 1 258
2 2228 1 258
2 2229 1 260
2 2230 1 260
2 2231 1 263
2 2232 1 263
2 2233 1 266
2 2234 1 266
2 2235 1 268
2 2236 1 268
2 2237 1 269
2 2238 1 269
2 2239 1 274
2 2240 1 274
2 2241 1 277
2 2242 1 277
2 2243 1 282
2 2244 1 282
2 2245 1 282
2 2246 1 284
2 2247 1 284
2 2248 1 287
2 2249 1 287
2 2250 1 290
2 2251 1 290
2 2252 1 292
2 2253 1 292
2 2254 1 293
2 2255 1 293
2 2256 1 298
2 2257 1 298
2 2258 1 301
2 2259 1 301
2 2260 1 306
2 2261 1 306
2 2262 1 306
2 2263 1 308
2 2264 1 308
2 2265 1 311
2 2266 1 311
2 2267 1 314
2 2268 1 314
2 2269 1 316
2 2270 1 316
2 2271 1 317
2 2272 1 317
2 2273 1 322
2 2274 1 322
2 2275 1 325
2 2276 1 325
2 2277 1 330
2 2278 1 330
2 2279 1 330
2 2280 1 332
2 2281 1 332
2 2282 1 335
2 2283 1 335
2 2284 1 338
2 2285 1 338
2 2286 1 340
2 2287 1 340
2 2288 1 341
2 2289 1 341
2 2290 1 346
2 2291 1 346
2 2292 1 349
2 2293 1 349
2 2294 1 354
2 2295 1 354
2 2296 1 354
2 2297 1 356
2 2298 1 356
2 2299 1 359
2 2300 1 359
2 2301 1 362
2 2302 1 362
2 2303 1 364
2 2304 1 364
2 2305 1 365
2 2306 1 365
2 2307 1 370
2 2308 1 370
2 2309 1 373
2 2310 1 373
2 2311 1 378
2 2312 1 378
2 2313 1 378
2 2314 1 380
2 2315 1 380
2 2316 1 383
2 2317 1 383
2 2318 1 386
2 2319 1 386
2 2320 1 388
2 2321 1 388
2 2322 1 389
2 2323 1 389
2 2324 1 394
2 2325 1 394
2 2326 1 397
2 2327 1 397
2 2328 1 402
2 2329 1 402
2 2330 1 402
2 2331 1 404
2 2332 1 404
2 2333 1 407
2 2334 1 407
2 2335 1 410
2 2336 1 410
2 2337 1 412
2 2338 1 412
2 2339 1 413
2 2340 1 413
2 2341 1 418
2 2342 1 418
2 2343 1 421
2 2344 1 421
2 2345 1 426
2 2346 1 426
2 2347 1 426
2 2348 1 428
2 2349 1 428
2 2350 1 431
2 2351 1 431
2 2352 1 434
2 2353 1 434
2 2354 1 436
2 2355 1 436
2 2356 1 437
2 2357 1 437
2 2358 1 442
2 2359 1 442
2 2360 1 445
2 2361 1 445
2 2362 1 450
2 2363 1 450
2 2364 1 450
2 2365 1 452
2 2366 1 452
2 2367 1 455
2 2368 1 455
2 2369 1 458
2 2370 1 458
2 2371 1 460
2 2372 1 460
2 2373 1 461
2 2374 1 461
2 2375 1 466
2 2376 1 466
2 2377 1 469
2 2378 1 469
2 2379 1 474
2 2380 1 474
2 2381 1 474
2 2382 1 476
2 2383 1 476
2 2384 1 479
2 2385 1 479
2 2386 1 482
2 2387 1 482
2 2388 1 484
2 2389 1 484
2 2390 1 485
2 2391 1 485
2 2392 1 490
2 2393 1 490
2 2394 1 493
2 2395 1 493
2 2396 1 498
2 2397 1 498
2 2398 1 498
2 2399 1 500
2 2400 1 500
2 2401 1 503
2 2402 1 503
2 2403 1 506
2 2404 1 506
2 2405 1 508
2 2406 1 508
2 2407 1 509
2 2408 1 509
2 2409 1 514
2 2410 1 514
2 2411 1 517
2 2412 1 517
2 2413 1 522
2 2414 1 522
2 2415 1 522
2 2416 1 524
2 2417 1 524
2 2418 1 527
2 2419 1 527
2 2420 1 530
2 2421 1 530
2 2422 1 532
2 2423 1 532
2 2424 1 533
2 2425 1 533
2 2426 1 538
2 2427 1 538
2 2428 1 541
2 2429 1 541
2 2430 1 546
2 2431 1 546
2 2432 1 546
2 2433 1 548
2 2434 1 548
2 2435 1 551
2 2436 1 551
2 2437 1 554
2 2438 1 554
2 2439 1 556
2 2440 1 556
2 2441 1 557
2 2442 1 557
2 2443 1 562
2 2444 1 562
2 2445 1 565
2 2446 1 565
2 2447 1 570
2 2448 1 570
2 2449 1 570
2 2450 1 572
2 2451 1 572
2 2452 1 575
2 2453 1 575
2 2454 1 578
2 2455 1 578
2 2456 1 580
2 2457 1 580
2 2458 1 581
2 2459 1 581
2 2460 1 586
2 2461 1 586
2 2462 1 589
2 2463 1 589
2 2464 1 594
2 2465 1 594
2 2466 1 594
2 2467 1 596
2 2468 1 596
2 2469 1 599
2 2470 1 599
2 2471 1 602
2 2472 1 602
2 2473 1 604
2 2474 1 604
2 2475 1 605
2 2476 1 605
2 2477 1 610
2 2478 1 610
2 2479 1 613
2 2480 1 613
2 2481 1 618
2 2482 1 618
2 2483 1 618
2 2484 1 620
2 2485 1 620
2 2486 1 623
2 2487 1 623
2 2488 1 626
2 2489 1 626
2 2490 1 628
2 2491 1 628
2 2492 1 629
2 2493 1 629
2 2494 1 634
2 2495 1 634
2 2496 1 637
2 2497 1 637
2 2498 1 642
2 2499 1 642
2 2500 1 642
2 2501 1 644
2 2502 1 644
2 2503 1 647
2 2504 1 647
2 2505 1 650
2 2506 1 650
2 2507 1 652
2 2508 1 652
2 2509 1 653
2 2510 1 653
2 2511 1 658
2 2512 1 658
2 2513 1 661
2 2514 1 661
2 2515 1 666
2 2516 1 666
2 2517 1 666
2 2518 1 668
2 2519 1 668
2 2520 1 671
2 2521 1 671
2 2522 1 674
2 2523 1 674
2 2524 1 676
2 2525 1 676
2 2526 1 677
2 2527 1 677
2 2528 1 682
2 2529 1 682
2 2530 1 685
2 2531 1 685
2 2532 1 690
2 2533 1 690
2 2534 1 690
2 2535 1 692
2 2536 1 692
2 2537 1 695
2 2538 1 695
2 2539 1 698
2 2540 1 698
2 2541 1 700
2 2542 1 700
2 2543 1 701
2 2544 1 701
2 2545 1 706
2 2546 1 706
2 2547 1 709
2 2548 1 709
2 2549 1 714
2 2550 1 714
2 2551 1 714
2 2552 1 716
2 2553 1 716
2 2554 1 719
2 2555 1 719
2 2556 1 722
2 2557 1 722
2 2558 1 724
2 2559 1 724
2 2560 1 725
2 2561 1 725
2 2562 1 730
2 2563 1 730
2 2564 1 733
2 2565 1 733
2 2566 1 738
2 2567 1 738
2 2568 1 738
2 2569 1 740
2 2570 1 740
2 2571 1 743
2 2572 1 743
2 2573 1 746
2 2574 1 746
2 2575 1 748
2 2576 1 748
2 2577 1 749
2 2578 1 749
2 2579 1 754
2 2580 1 754
2 2581 1 757
2 2582 1 757
2 2583 1 762
2 2584 1 762
2 2585 1 762
2 2586 1 764
2 2587 1 764
2 2588 1 767
2 2589 1 767
2 2590 1 770
2 2591 1 770
2 2592 1 772
2 2593 1 772
2 2594 1 773
2 2595 1 773
2 2596 1 778
2 2597 1 778
2 2598 1 781
2 2599 1 781
2 2600 1 786
2 2601 1 786
2 2602 1 786
2 2603 1 788
2 2604 1 788
2 2605 1 791
2 2606 1 791
2 2607 1 794
2 2608 1 794
2 2609 1 796
2 2610 1 796
2 2611 1 797
2 2612 1 797
2 2613 1 802
2 2614 1 802
2 2615 1 805
2 2616 1 805
2 2617 1 810
2 2618 1 810
2 2619 1 810
2 2620 1 812
2 2621 1 812
2 2622 1 815
2 2623 1 815
2 2624 1 818
2 2625 1 818
2 2626 1 820
2 2627 1 820
2 2628 1 821
2 2629 1 821
2 2630 1 826
2 2631 1 826
2 2632 1 829
2 2633 1 829
2 2634 1 834
2 2635 1 834
2 2636 1 834
2 2637 1 836
2 2638 1 836
2 2639 1 839
2 2640 1 839
2 2641 1 842
2 2642 1 842
2 2643 1 844
2 2644 1 844
2 2645 1 845
2 2646 1 845
2 2647 1 850
2 2648 1 850
2 2649 1 853
2 2650 1 853
2 2651 1 858
2 2652 1 858
2 2653 1 858
2 2654 1 860
2 2655 1 860
2 2656 1 863
2 2657 1 863
2 2658 1 866
2 2659 1 866
2 2660 1 868
2 2661 1 868
2 2662 1 869
2 2663 1 869
2 2664 1 874
2 2665 1 874
2 2666 1 877
2 2667 1 877
2 2668 1 882
2 2669 1 882
2 2670 1 882
2 2671 1 884
2 2672 1 884
2 2673 1 887
2 2674 1 887
2 2675 1 890
2 2676 1 890
2 2677 1 892
2 2678 1 892
2 2679 1 893
2 2680 1 893
2 2681 1 898
2 2682 1 898
2 2683 1 901
2 2684 1 901
2 2685 1 906
2 2686 1 906
2 2687 1 906
2 2688 1 908
2 2689 1 908
2 2690 1 911
2 2691 1 911
2 2692 1 914
2 2693 1 914
2 2694 1 916
2 2695 1 916
2 2696 1 917
2 2697 1 917
2 2698 1 922
2 2699 1 922
2 2700 1 925
2 2701 1 925
2 2702 1 930
2 2703 1 930
2 2704 1 930
2 2705 1 932
2 2706 1 932
2 2707 1 935
2 2708 1 935
2 2709 1 938
2 2710 1 938
2 2711 1 940
2 2712 1 940
2 2713 1 941
2 2714 1 941
2 2715 1 946
2 2716 1 946
2 2717 1 949
2 2718 1 949
2 2719 1 954
2 2720 1 954
2 2721 1 954
2 2722 1 956
2 2723 1 956
2 2724 1 959
2 2725 1 959
2 2726 1 962
2 2727 1 962
2 2728 1 964
2 2729 1 964
2 2730 1 965
2 2731 1 965
2 2732 1 970
2 2733 1 970
2 2734 1 973
2 2735 1 973
2 2736 1 978
2 2737 1 978
2 2738 1 978
2 2739 1 980
2 2740 1 980
2 2741 1 983
2 2742 1 983
2 2743 1 986
2 2744 1 986
2 2745 1 988
2 2746 1 988
2 2747 1 989
2 2748 1 989
2 2749 1 994
2 2750 1 994
2 2751 1 997
2 2752 1 997
2 2753 1 1002
2 2754 1 1002
2 2755 1 1002
2 2756 1 1004
2 2757 1 1004
2 2758 1 1007
2 2759 1 1007
2 2760 1 1010
2 2761 1 1010
2 2762 1 1012
2 2763 1 1012
2 2764 1 1013
2 2765 1 1013
2 2766 1 1018
2 2767 1 1018
2 2768 1 1021
2 2769 1 1021
2 2770 1 1026
2 2771 1 1026
2 2772 1 1026
2 2773 1 1028
2 2774 1 1028
2 2775 1 1031
2 2776 1 1031
2 2777 1 1034
2 2778 1 1034
2 2779 1 1036
2 2780 1 1036
2 2781 1 1037
2 2782 1 1037
2 2783 1 1042
2 2784 1 1042
2 2785 1 1045
2 2786 1 1045
2 2787 1 1050
2 2788 1 1050
2 2789 1 1050
2 2790 1 1052
2 2791 1 1052
2 2792 1 1055
2 2793 1 1055
2 2794 1 1058
2 2795 1 1058
2 2796 1 1060
2 2797 1 1060
2 2798 1 1061
2 2799 1 1061
2 2800 1 1066
2 2801 1 1066
2 2802 1 1069
2 2803 1 1069
2 2804 1 1074
2 2805 1 1074
2 2806 1 1074
2 2807 1 1076
2 2808 1 1076
2 2809 1 1079
2 2810 1 1079
2 2811 1 1082
2 2812 1 1082
2 2813 1 1084
2 2814 1 1084
2 2815 1 1085
2 2816 1 1085
2 2817 1 1090
2 2818 1 1090
2 2819 1 1093
2 2820 1 1093
2 2821 1 1098
2 2822 1 1098
2 2823 1 1098
2 2824 1 1100
2 2825 1 1100
2 2826 1 1103
2 2827 1 1103
2 2828 1 1106
2 2829 1 1106
2 2830 1 1108
2 2831 1 1108
2 2832 1 1109
2 2833 1 1109
2 2834 1 1114
2 2835 1 1114
2 2836 1 1117
2 2837 1 1117
2 2838 1 1122
2 2839 1 1122
2 2840 1 1122
2 2841 1 1124
2 2842 1 1124
2 2843 1 1129
2 2844 1 1129
2 2845 1 1130
2 2846 1 1130
2 2847 1 1132
2 2848 1 1132
2 2849 1 1133
2 2850 1 1133
2 2851 1 1138
2 2852 1 1138
2 2853 1 1141
2 2854 1 1141
2 2855 1 1146
2 2856 1 1146
2 2857 1 1146
2 2858 1 1154
2 2859 1 1154
2 2860 1 1157
2 2861 1 1157
2 2862 1 1160
2 2863 1 1160
2 2864 1 1170
2 2865 1 1170
2 2866 1 1177
2 2867 1 1177
2 2868 1 1180
2 2869 1 1180
2 2870 1 1182
2 2871 1 1182
2 2872 1 1184
2 2873 1 1184
2 2874 1 1186
2 2875 1 1186
2 2876 1 1187
2 2877 1 1187
2 2878 1 1188
2 2879 1 1188
2 2880 1 1188
2 2881 1 1191
2 2882 1 1191
2 2883 1 1192
2 2884 1 1192
2 2885 1 1195
2 2886 1 1195
2 2887 1 1198
2 2888 1 1198
2 2889 1 1200
2 2890 1 1200
2 2891 1 1203
2 2892 1 1203
2 2893 1 1206
2 2894 1 1206
2 2895 1 1208
2 2896 1 1208
2 2897 1 1211
2 2898 1 1211
2 2899 1 1214
2 2900 1 1214
2 2901 1 1216
2 2902 1 1216
2 2903 1 1219
2 2904 1 1219
2 2905 1 1222
2 2906 1 1222
2 2907 1 1224
2 2908 1 1224
2 2909 1 1227
2 2910 1 1227
2 2911 1 1230
2 2912 1 1230
2 2913 1 1232
2 2914 1 1232
2 2915 1 1235
2 2916 1 1235
2 2917 1 1238
2 2918 1 1238
2 2919 1 1240
2 2920 1 1240
2 2921 1 1243
2 2922 1 1243
2 2923 1 1246
2 2924 1 1246
2 2925 1 1248
2 2926 1 1248
2 2927 1 1251
2 2928 1 1251
2 2929 1 1254
2 2930 1 1254
2 2931 1 1256
2 2932 1 1256
2 2933 1 1259
2 2934 1 1259
2 2935 1 1262
2 2936 1 1262
2 2937 1 1264
2 2938 1 1264
2 2939 1 1267
2 2940 1 1267
2 2941 1 1270
2 2942 1 1270
2 2943 1 1272
2 2944 1 1272
2 2945 1 1275
2 2946 1 1275
2 2947 1 1278
2 2948 1 1278
2 2949 1 1280
2 2950 1 1280
2 2951 1 1283
2 2952 1 1283
2 2953 1 1286
2 2954 1 1286
2 2955 1 1288
2 2956 1 1288
2 2957 1 1291
2 2958 1 1291
2 2959 1 1294
2 2960 1 1294
2 2961 1 1296
2 2962 1 1296
2 2963 1 1299
2 2964 1 1299
2 2965 1 1301
2 2966 1 1301
2 2967 1 1302
2 2968 1 1302
2 2969 1 1304
2 2970 1 1304
2 2971 1 1304
2 2972 1 1305
2 2973 1 1305
2 2974 1 1311
2 2975 1 1311
2 2976 1 1314
2 2977 1 1314
2 2978 1 1314
2 2979 1 1314
2 2980 1 1316
2 2981 1 1316
2 2982 1 1316
2 2983 1 1316
2 2984 1 1316
2 2985 1 1317
2 2986 1 1317
2 2987 1 1323
2 2988 1 1323
2 2989 1 1326
2 2990 1 1326
2 2991 1 1326
2 2992 1 1328
2 2993 1 1328
2 2994 1 1328
2 2995 1 1328
2 2996 1 1329
2 2997 1 1329
2 2998 1 1335
2 2999 1 1335
2 3000 1 1338
2 3001 1 1338
2 3002 1 1338
2 3003 1 1340
2 3004 1 1340
2 3005 1 1340
2 3006 1 1340
2 3007 1 1341
2 3008 1 1341
2 3009 1 1347
2 3010 1 1347
2 3011 1 1350
2 3012 1 1350
2 3013 1 1350
2 3014 1 1352
2 3015 1 1352
2 3016 1 1352
2 3017 1 1352
2 3018 1 1353
2 3019 1 1353
2 3020 1 1359
2 3021 1 1359
2 3022 1 1362
2 3023 1 1362
2 3024 1 1362
2 3025 1 1362
2 3026 1 1364
2 3027 1 1364
2 3028 1 1364
2 3029 1 1364
2 3030 1 1365
2 3031 1 1365
2 3032 1 1371
2 3033 1 1371
2 3034 1 1373
2 3035 1 1373
2 3036 1 1374
2 3037 1 1374
2 3038 1 1374
2 3039 1 1374
2 3040 1 1376
2 3041 1 1376
2 3042 1 1376
2 3043 1 1376
2 3044 1 1377
2 3045 1 1377
2 3046 1 1383
2 3047 1 1383
2 3048 1 1386
2 3049 1 1386
2 3050 1 1386
2 3051 1 1386
2 3052 1 1386
2 3053 1 1388
2 3054 1 1388
2 3055 1 1388
2 3056 1 1388
2 3057 1 1389
2 3058 1 1389
2 3059 1 1395
2 3060 1 1395
2 3061 1 1398
2 3062 1 1398
2 3063 1 1398
2 3064 1 1398
2 3065 1 1398
2 3066 1 1400
2 3067 1 1400
2 3068 1 1400
2 3069 1 1401
2 3070 1 1401
2 3071 1 1407
2 3072 1 1407
2 3073 1 1410
2 3074 1 1410
2 3075 1 1410
2 3076 1 1410
2 3077 1 1410
2 3078 1 1412
2 3079 1 1412
2 3080 1 1412
2 3081 1 1412
2 3082 1 1413
2 3083 1 1413
2 3084 1 1419
2 3085 1 1419
2 3086 1 1422
2 3087 1 1422
2 3088 1 1422
2 3089 1 1422
2 3090 1 1423
2 3091 1 1423
2 3092 1 1429
2 3093 1 1429
2 3094 1 1432
2 3095 1 1432
2 3096 1 1432
2 3097 1 1432
2 3098 1 1434
2 3099 1 1434
2 3100 1 1434
2 3101 1 1435
2 3102 1 1435
2 3103 1 1441
2 3104 1 1441
2 3105 1 1444
2 3106 1 1444
2 3107 1 1444
2 3108 1 1444
2 3109 1 1446
2 3110 1 1446
2 3111 1 1446
2 3112 1 1447
2 3113 1 1447
2 3114 1 1453
2 3115 1 1453
2 3116 1 1456
2 3117 1 1456
2 3118 1 1457
2 3119 1 1457
2 3120 1 1463
2 3121 1 1463
2 3122 1 1467
2 3123 1 1467
2 3124 1 1471
2 3125 1 1471
2 3126 1 1475
2 3127 1 1475
2 3128 1 1477
2 3129 1 1477
2 3130 1 1482
2 3131 1 1482
2 3132 1 1482
2 3133 1 1484
2 3134 1 1484
2 3135 1 1485
2 3136 1 1485
2 3137 1 1488
2 3138 1 1488
2 3139 1 1489
2 3140 1 1489
2 3141 1 1492
2 3142 1 1492
2 3143 1 1495
2 3144 1 1495
2 3145 1 1496
2 3146 1 1496
2 3147 1 1502
2 3148 1 1502
2 3149 1 1505
2 3150 1 1505
2 3151 1 1505
2 3152 1 1505
2 3153 1 1507
2 3154 1 1507
2 3155 1 1507
2 3156 1 1507
2 3157 1 1508
2 3158 1 1508
2 3159 1 1512
2 3160 1 1512
2 3161 1 1512
2 3162 1 1512
2 3163 1 1515
2 3164 1 1515
2 3165 1 1522
2 3166 1 1522
2 3167 1 1525
2 3168 1 1525
2 3169 1 1529
2 3170 1 1529
2 3171 1 1531
2 3172 1 1531
2 3173 1 1532
2 3174 1 1532
2 3175 1 1535
2 3176 1 1535
2 3177 1 1536
2 3178 1 1536
2 3179 1 1539
2 3180 1 1539
2 3181 1 1540
2 3182 1 1540
2 3183 1 1543
2 3184 1 1543
2 3185 1 1546
2 3186 1 1546
2 3187 1 1551
2 3188 1 1551
2 3189 1 1553
2 3190 1 1553
2 3191 1 1558
2 3192 1 1558
2 3193 1 1561
2 3194 1 1561
2 3195 1 1561
2 3196 1 1562
2 3197 1 1562
2 3198 1 1567
2 3199 1 1567
2 3200 1 1567
2 3201 1 1568
2 3202 1 1568
2 3203 1 1573
2 3204 1 1573
2 3205 1 1573
2 3206 1 1574
2 3207 1 1574
2 3208 1 1581
2 3209 1 1581
2 3210 1 1582
2 3211 1 1582
2 3212 1 1586
2 3213 1 1586
2 3214 1 1590
2 3215 1 1590
2 3216 1 1595
2 3217 1 1595
2 3218 1 1595
2 3219 1 1602
2 3220 1 1602
2 3221 1 1605
2 3222 1 1605
2 3223 1 1611
2 3224 1 1611
2 3225 1 1614
2 3226 1 1614
2 3227 1 1614
2 3228 1 1615
2 3229 1 1615
2 3230 1 1618
2 3231 1 1618
2 3232 1 1618
2 3233 1 1619
2 3234 1 1619
2 3235 1 1625
2 3236 1 1625
2 3237 1 1625
2 3238 1 1628
2 3239 1 1628
2 3240 1 1661
2 3241 1 1661
2 3242 1 1662
2 3243 1 1662
2 3244 1 1665
2 3245 1 1665
2 3246 1 1666
2 3247 1 1666
2 3248 1 1669
2 3249 1 1669
2 3250 1 1672
2 3251 1 1672
2 3252 1 1680
2 3253 1 1680
2 3254 1 1683
2 3255 1 1683
2 3256 1 1685
2 3257 1 1685
2 3258 1 1688
2 3259 1 1688
2 3260 1 1692
2 3261 1 1692
2 3262 1 1695
2 3263 1 1695
2 3264 1 1696
2 3265 1 1696
2 3266 1 1699
2 3267 1 1699
2 3268 1 1700
2 3269 1 1700
2 3270 1 1703
2 3271 1 1703
2 3272 1 1704
2 3273 1 1704
2 3274 1 1708
2 3275 1 1708
2 3276 1 1711
2 3277 1 1711
0 50 5 1 1 49
0 51 5 2 1 1813
0 52 5 3 1 1816
0 53 5 3 1 1819
0 54 5 3 1 1822
0 55 5 3 1 1825
0 56 5 3 1 1828
0 57 5 3 1 1831
0 58 5 3 1 1834
0 59 5 3 1 1837
0 60 5 3 1 1840
0 61 5 3 1 1843
0 62 5 3 1 1846
0 63 5 3 1 1849
0 64 5 3 1 1852
0 65 5 3 1 1855
0 66 5 3 1 1858
0 67 5 3 1 1861
0 68 5 3 1 1864
0 69 5 4 1 1867
0 70 5 4 1 1870
0 71 5 4 1 1873
0 72 5 4 1 1876
0 73 5 4 1 1879
0 74 5 4 1 1882
0 75 5 4 1 1885
0 76 5 4 1 1888
0 77 5 4 1 1891
0 78 5 4 1 1894
0 79 5 4 1 1897
0 80 5 4 1 1900
0 81 5 4 1 1903
0 82 5 3 1 1906
0 83 5 3 1 1909
0 84 5 3 1 1912
0 85 5 3 1 1915
0 86 5 3 1 1918
0 87 5 3 1 1921
0 88 5 3 1 1924
0 89 5 3 1 1927
0 90 5 3 1 1930
0 91 5 3 1 1933
0 92 5 3 1 1936
0 93 5 3 1 1939
0 94 5 3 1 1942
0 95 5 4 1 1945
0 96 5 3 1 1949
0 97 5 2 1 1952
0 98 5 2 1 1956
0 99 7 2 2 2108 2111
0 100 5 1 1 2115
0 101 7 3 2 1957 2116
0 102 5 1 1 2117
0 103 7 2 2 2109 1958
0 104 5 1 1 2120
0 105 7 1 2 100 2121
0 106 5 1 1 105
0 107 7 1 2 1950 2113
0 108 5 1 1 107
0 109 7 2 2 106 108
0 110 5 1 1 2122
0 111 7 2 2 2104 2123
0 112 5 1 1 2124
0 113 7 1 2 1953 104
0 114 7 1 2 112 113
0 115 5 1 1 114
0 116 7 2 2 102 115
0 117 5 1 1 2126
0 118 7 1 2 2105 117
0 119 5 2 1 118
0 120 7 1 2 1946 2127
0 121 5 1 1 120
0 122 7 2 2 2128 121
0 123 5 1 1 2130
0 124 7 2 2 2101 2131
0 125 5 2 1 2132
0 126 7 1 2 110 2129
0 127 5 1 1 126
0 128 7 1 2 2106 2118
0 129 5 1 1 128
0 130 7 2 2 127 129
0 131 5 1 1 2136
0 132 7 1 2 2134 131
0 133 5 2 1 132
0 134 7 1 2 1954 2125
0 135 5 1 1 134
0 136 7 1 2 1947 2119
0 137 5 1 1 136
0 138 7 2 2 135 137
0 139 5 2 1 2140
0 140 7 2 2 2138 2141
0 141 5 1 1 2144
0 142 7 1 2 2102 141
0 143 5 2 1 142
0 144 7 1 2 1943 2145
0 145 5 1 1 144
0 146 7 2 2 2146 145
0 147 5 1 1 2148
0 148 7 2 2 2098 2149
0 149 5 2 1 2150
0 150 7 1 2 123 2147
0 151 5 1 1 150
0 152 7 1 2 2133 2142
0 153 5 1 1 152
0 154 7 2 2 151 153
0 155 5 1 1 2154
0 156 7 1 2 2152 155
0 157 5 2 1 156
0 158 7 1 2 2135 2143
0 159 5 1 1 158
0 160 7 1 2 2137 159
0 161 5 1 1 160
0 162 7 3 2 2139 161
0 163 5 1 1 2158
0 164 7 2 2 2156 163
0 165 5 1 1 2161
0 166 7 1 2 2099 165
0 167 5 2 1 166
0 168 7 1 2 1940 2162
0 169 5 1 1 168
0 170 7 2 2 2163 169
0 171 5 1 1 2165
0 172 7 2 2 2095 2166
0 173 5 2 1 2167
0 174 7 1 2 147 2164
0 175 5 1 1 174
0 176 7 1 2 2151 2159
0 177 5 1 1 176
0 178 7 2 2 175 177
0 179 5 1 1 2171
0 180 7 1 2 2169 179
0 181 5 2 1 180
0 182 7 1 2 2153 2160
0 183 5 1 1 182
0 184 7 1 2 2155 183
0 185 5 1 1 184
0 186 7 3 2 2157 185
0 187 5 1 1 2175
0 188 7 2 2 2173 187
0 189 5 1 1 2178
0 190 7 1 2 2096 189
0 191 5 2 1 190
0 192 7 1 2 1937 2179
0 193 5 1 1 192
0 194 7 2 2 2180 193
0 195 5 1 1 2182
0 196 7 2 2 2092 2183
0 197 5 2 1 2184
0 198 7 1 2 171 2181
0 199 5 1 1 198
0 200 7 1 2 2168 2176
0 201 5 1 1 200
0 202 7 2 2 199 201
0 203 5 1 1 2188
0 204 7 1 2 2186 203
0 205 5 2 1 204
0 206 7 1 2 2170 2177
0 207 5 1 1 206
0 208 7 1 2 2172 207
0 209 5 1 1 208
0 210 7 3 2 2174 209
0 211 5 1 1 2192
0 212 7 2 2 2190 211
0 213 5 1 1 2195
0 214 7 1 2 2093 213
0 215 5 2 1 214
0 216 7 1 2 1934 2196
0 217 5 1 1 216
0 218 7 2 2 2197 217
0 219 5 1 1 2199
0 220 7 2 2 2089 2200
0 221 5 2 1 2201
0 222 7 1 2 195 2198
0 223 5 1 1 222
0 224 7 1 2 2185 2193
0 225 5 1 1 224
0 226 7 2 2 223 225
0 227 5 1 1 2205
0 228 7 1 2 2203 227
0 229 5 2 1 228
0 230 7 1 2 2187 2194
0 231 5 1 1 230
0 232 7 1 2 2189 231
0 233 5 1 1 232
0 234 7 3 2 2191 233
0 235 5 1 1 2209
0 236 7 2 2 2207 235
0 237 5 1 1 2212
0 238 7 1 2 2090 237
0 239 5 2 1 238
0 240 7 1 2 1931 2213
0 241 5 1 1 240
0 242 7 2 2 2214 241
0 243 5 1 1 2216
0 244 7 2 2 2086 2217
0 245 5 2 1 2218
0 246 7 1 2 219 2215
0 247 5 1 1 246
0 248 7 1 2 2202 2210
0 249 5 1 1 248
0 250 7 2 2 247 249
0 251 5 1 1 2222
0 252 7 1 2 2220 251
0 253 5 2 1 252
0 254 7 1 2 2204 2211
0 255 5 1 1 254
0 256 7 1 2 2206 255
0 257 5 1 1 256
0 258 7 3 2 2208 257
0 259 5 1 1 2226
0 260 7 2 2 2224 259
0 261 5 1 1 2229
0 262 7 1 2 2087 261
0 263 5 2 1 262
0 264 7 1 2 1928 2230
0 265 5 1 1 264
0 266 7 2 2 2231 265
0 267 5 1 1 2233
0 268 7 2 2 2083 2234
0 269 5 2 1 2235
0 270 7 1 2 243 2232
0 271 5 1 1 270
0 272 7 1 2 2219 2227
0 273 5 1 1 272
0 274 7 2 2 271 273
0 275 5 1 1 2239
0 276 7 1 2 2237 275
0 277 5 2 1 276
0 278 7 1 2 2221 2228
0 279 5 1 1 278
0 280 7 1 2 2223 279
0 281 5 1 1 280
0 282 7 3 2 2225 281
0 283 5 1 1 2243
0 284 7 2 2 2241 283
0 285 5 1 1 2246
0 286 7 1 2 2084 285
0 287 5 2 1 286
0 288 7 1 2 1925 2247
0 289 5 1 1 288
0 290 7 2 2 2248 289
0 291 5 1 1 2250
0 292 7 2 2 2080 2251
0 293 5 2 1 2252
0 294 7 1 2 267 2249
0 295 5 1 1 294
0 296 7 1 2 2236 2244
0 297 5 1 1 296
0 298 7 2 2 295 297
0 299 5 1 1 2256
0 300 7 1 2 2254 299
0 301 5 2 1 300
0 302 7 1 2 2238 2245
0 303 5 1 1 302
0 304 7 1 2 2240 303
0 305 5 1 1 304
0 306 7 3 2 2242 305
0 307 5 1 1 2260
0 308 7 2 2 2258 307
0 309 5 1 1 2263
0 310 7 1 2 2081 309
0 311 5 2 1 310
0 312 7 1 2 1922 2264
0 313 5 1 1 312
0 314 7 2 2 2265 313
0 315 5 1 1 2267
0 316 7 2 2 2077 2268
0 317 5 2 1 2269
0 318 7 1 2 291 2266
0 319 5 1 1 318
0 320 7 1 2 2253 2261
0 321 5 1 1 320
0 322 7 2 2 319 321
0 323 5 1 1 2273
0 324 7 1 2 2271 323
0 325 5 2 1 324
0 326 7 1 2 2255 2262
0 327 5 1 1 326
0 328 7 1 2 2257 327
0 329 5 1 1 328
0 330 7 3 2 2259 329
0 331 5 1 1 2277
0 332 7 2 2 2275 331
0 333 5 1 1 2280
0 334 7 1 2 2078 333
0 335 5 2 1 334
0 336 7 1 2 1919 2281
0 337 5 1 1 336
0 338 7 2 2 2282 337
0 339 5 1 1 2284
0 340 7 2 2 2074 2285
0 341 5 2 1 2286
0 342 7 1 2 315 2283
0 343 5 1 1 342
0 344 7 1 2 2270 2278
0 345 5 1 1 344
0 346 7 2 2 343 345
0 347 5 1 1 2290
0 348 7 1 2 2288 347
0 349 5 2 1 348
0 350 7 1 2 2272 2279
0 351 5 1 1 350
0 352 7 1 2 2274 351
0 353 5 1 1 352
0 354 7 3 2 2276 353
0 355 5 1 1 2294
0 356 7 2 2 2292 355
0 357 5 1 1 2297
0 358 7 1 2 2075 357
0 359 5 2 1 358
0 360 7 1 2 1916 2298
0 361 5 1 1 360
0 362 7 2 2 2299 361
0 363 5 1 1 2301
0 364 7 2 2 2071 2302
0 365 5 2 1 2303
0 366 7 1 2 339 2300
0 367 5 1 1 366
0 368 7 1 2 2287 2295
0 369 5 1 1 368
0 370 7 2 2 367 369
0 371 5 1 1 2307
0 372 7 1 2 2305 371
0 373 5 2 1 372
0 374 7 1 2 2289 2296
0 375 5 1 1 374
0 376 7 1 2 2291 375
0 377 5 1 1 376
0 378 7 3 2 2293 377
0 379 5 1 1 2311
0 380 7 2 2 2309 379
0 381 5 1 1 2314
0 382 7 1 2 2072 381
0 383 5 2 1 382
0 384 7 1 2 1913 2315
0 385 5 1 1 384
0 386 7 2 2 2316 385
0 387 5 1 1 2318
0 388 7 2 2 2068 2319
0 389 5 2 1 2320
0 390 7 1 2 363 2317
0 391 5 1 1 390
0 392 7 1 2 2304 2312
0 393 5 1 1 392
0 394 7 2 2 391 393
0 395 5 1 1 2324
0 396 7 1 2 2322 395
0 397 5 2 1 396
0 398 7 1 2 2306 2313
0 399 5 1 1 398
0 400 7 1 2 2308 399
0 401 5 1 1 400
0 402 7 3 2 2310 401
0 403 5 1 1 2328
0 404 7 2 2 2326 403
0 405 5 1 1 2331
0 406 7 1 2 2069 405
0 407 5 2 1 406
0 408 7 1 2 1910 2332
0 409 5 1 1 408
0 410 7 2 2 2333 409
0 411 5 1 1 2335
0 412 7 2 2 2065 2336
0 413 5 2 1 2337
0 414 7 1 2 387 2334
0 415 5 1 1 414
0 416 7 1 2 2321 2329
0 417 5 1 1 416
0 418 7 2 2 415 417
0 419 5 1 1 2341
0 420 7 1 2 2339 419
0 421 5 2 1 420
0 422 7 1 2 2323 2330
0 423 5 1 1 422
0 424 7 1 2 2325 423
0 425 5 1 1 424
0 426 7 3 2 2327 425
0 427 5 1 1 2345
0 428 7 2 2 2343 427
0 429 5 1 1 2348
0 430 7 1 2 2066 429
0 431 5 2 1 430
0 432 7 1 2 1907 2349
0 433 5 1 1 432
0 434 7 2 2 2350 433
0 435 5 1 1 2352
0 436 7 2 2 2061 2353
0 437 5 2 1 2354
0 438 7 1 2 411 2351
0 439 5 1 1 438
0 440 7 1 2 2338 2346
0 441 5 1 1 440
0 442 7 2 2 439 441
0 443 5 1 1 2358
0 444 7 1 2 2356 443
0 445 5 2 1 444
0 446 7 1 2 2340 2347
0 447 5 1 1 446
0 448 7 1 2 2342 447
0 449 5 1 1 448
0 450 7 3 2 2344 449
0 451 5 1 1 2362
0 452 7 2 2 2360 451
0 453 5 1 1 2365
0 454 7 1 2 2062 453
0 455 5 2 1 454
0 456 7 1 2 1904 2366
0 457 5 1 1 456
0 458 7 2 2 2367 457
0 459 5 1 1 2369
0 460 7 2 2 2057 2370
0 461 5 2 1 2371
0 462 7 1 2 435 2368
0 463 5 1 1 462
0 464 7 1 2 2355 2363
0 465 5 1 1 464
0 466 7 2 2 463 465
0 467 5 1 1 2375
0 468 7 1 2 2373 467
0 469 5 2 1 468
0 470 7 1 2 2357 2364
0 471 5 1 1 470
0 472 7 1 2 2359 471
0 473 5 1 1 472
0 474 7 3 2 2361 473
0 475 5 1 1 2379
0 476 7 2 2 2377 475
0 477 5 1 1 2382
0 478 7 1 2 2058 477
0 479 5 2 1 478
0 480 7 1 2 1901 2383
0 481 5 1 1 480
0 482 7 2 2 2384 481
0 483 5 1 1 2386
0 484 7 2 2 2053 2387
0 485 5 2 1 2388
0 486 7 1 2 459 2385
0 487 5 1 1 486
0 488 7 1 2 2372 2380
0 489 5 1 1 488
0 490 7 2 2 487 489
0 491 5 1 1 2392
0 492 7 1 2 2390 491
0 493 5 2 1 492
0 494 7 1 2 2374 2381
0 495 5 1 1 494
0 496 7 1 2 2376 495
0 497 5 1 1 496
0 498 7 3 2 2378 497
0 499 5 1 1 2396
0 500 7 2 2 2394 499
0 501 5 1 1 2399
0 502 7 1 2 2054 501
0 503 5 2 1 502
0 504 7 1 2 1898 2400
0 505 5 1 1 504
0 506 7 2 2 2401 505
0 507 5 1 1 2403
0 508 7 2 2 2049 2404
0 509 5 2 1 2405
0 510 7 1 2 483 2402
0 511 5 1 1 510
0 512 7 1 2 2389 2397
0 513 5 1 1 512
0 514 7 2 2 511 513
0 515 5 1 1 2409
0 516 7 1 2 2407 515
0 517 5 2 1 516
0 518 7 1 2 2391 2398
0 519 5 1 1 518
0 520 7 1 2 2393 519
0 521 5 1 1 520
0 522 7 3 2 2395 521
0 523 5 1 1 2413
0 524 7 2 2 2411 523
0 525 5 1 1 2416
0 526 7 1 2 2050 525
0 527 5 2 1 526
0 528 7 1 2 1895 2417
0 529 5 1 1 528
0 530 7 2 2 2418 529
0 531 5 1 1 2420
0 532 7 2 2 2045 2421
0 533 5 2 1 2422
0 534 7 1 2 507 2419
0 535 5 1 1 534
0 536 7 1 2 2406 2414
0 537 5 1 1 536
0 538 7 2 2 535 537
0 539 5 1 1 2426
0 540 7 1 2 2424 539
0 541 5 2 1 540
0 542 7 1 2 2408 2415
0 543 5 1 1 542
0 544 7 1 2 2410 543
0 545 5 1 1 544
0 546 7 3 2 2412 545
0 547 5 1 1 2430
0 548 7 2 2 2428 547
0 549 5 1 1 2433
0 550 7 1 2 2046 549
0 551 5 2 1 550
0 552 7 1 2 1892 2434
0 553 5 1 1 552
0 554 7 2 2 2435 553
0 555 5 1 1 2437
0 556 7 2 2 2041 2438
0 557 5 2 1 2439
0 558 7 1 2 531 2436
0 559 5 1 1 558
0 560 7 1 2 2423 2431
0 561 5 1 1 560
0 562 7 2 2 559 561
0 563 5 1 1 2443
0 564 7 1 2 2441 563
0 565 5 2 1 564
0 566 7 1 2 2425 2432
0 567 5 1 1 566
0 568 7 1 2 2427 567
0 569 5 1 1 568
0 570 7 3 2 2429 569
0 571 5 1 1 2447
0 572 7 2 2 2445 571
0 573 5 1 1 2450
0 574 7 1 2 2042 573
0 575 5 2 1 574
0 576 7 1 2 1889 2451
0 577 5 1 1 576
0 578 7 2 2 2452 577
0 579 5 1 1 2454
0 580 7 2 2 2037 2455
0 581 5 2 1 2456
0 582 7 1 2 555 2453
0 583 5 1 1 582
0 584 7 1 2 2440 2448
0 585 5 1 1 584
0 586 7 2 2 583 585
0 587 5 1 1 2460
0 588 7 1 2 2458 587
0 589 5 2 1 588
0 590 7 1 2 2442 2449
0 591 5 1 1 590
0 592 7 1 2 2444 591
0 593 5 1 1 592
0 594 7 3 2 2446 593
0 595 5 1 1 2464
0 596 7 2 2 2462 595
0 597 5 1 1 2467
0 598 7 1 2 2038 597
0 599 5 2 1 598
0 600 7 1 2 1886 2468
0 601 5 1 1 600
0 602 7 2 2 2469 601
0 603 5 1 1 2471
0 604 7 2 2 2033 2472
0 605 5 2 1 2473
0 606 7 1 2 579 2470
0 607 5 1 1 606
0 608 7 1 2 2457 2465
0 609 5 1 1 608
0 610 7 2 2 607 609
0 611 5 1 1 2477
0 612 7 1 2 2475 611
0 613 5 2 1 612
0 614 7 1 2 2459 2466
0 615 5 1 1 614
0 616 7 1 2 2461 615
0 617 5 1 1 616
0 618 7 3 2 2463 617
0 619 5 1 1 2481
0 620 7 2 2 2479 619
0 621 5 1 1 2484
0 622 7 1 2 2034 621
0 623 5 2 1 622
0 624 7 1 2 1883 2485
0 625 5 1 1 624
0 626 7 2 2 2486 625
0 627 5 1 1 2488
0 628 7 2 2 2029 2489
0 629 5 2 1 2490
0 630 7 1 2 603 2487
0 631 5 1 1 630
0 632 7 1 2 2474 2482
0 633 5 1 1 632
0 634 7 2 2 631 633
0 635 5 1 1 2494
0 636 7 1 2 2492 635
0 637 5 2 1 636
0 638 7 1 2 2476 2483
0 639 5 1 1 638
0 640 7 1 2 2478 639
0 641 5 1 1 640
0 642 7 3 2 2480 641
0 643 5 1 1 2498
0 644 7 2 2 2496 643
0 645 5 1 1 2501
0 646 7 1 2 2030 645
0 647 5 2 1 646
0 648 7 1 2 1880 2502
0 649 5 1 1 648
0 650 7 2 2 2503 649
0 651 5 1 1 2505
0 652 7 2 2 2025 2506
0 653 5 2 1 2507
0 654 7 1 2 627 2504
0 655 5 1 1 654
0 656 7 1 2 2491 2499
0 657 5 1 1 656
0 658 7 2 2 655 657
0 659 5 1 1 2511
0 660 7 1 2 2509 659
0 661 5 2 1 660
0 662 7 1 2 2493 2500
0 663 5 1 1 662
0 664 7 1 2 2495 663
0 665 5 1 1 664
0 666 7 3 2 2497 665
0 667 5 1 1 2515
0 668 7 2 2 2513 667
0 669 5 1 1 2518
0 670 7 1 2 2026 669
0 671 5 2 1 670
0 672 7 1 2 1877 2519
0 673 5 1 1 672
0 674 7 2 2 2520 673
0 675 5 1 1 2522
0 676 7 2 2 2021 2523
0 677 5 2 1 2524
0 678 7 1 2 651 2521
0 679 5 1 1 678
0 680 7 1 2 2508 2516
0 681 5 1 1 680
0 682 7 2 2 679 681
0 683 5 1 1 2528
0 684 7 1 2 2526 683
0 685 5 2 1 684
0 686 7 1 2 2510 2517
0 687 5 1 1 686
0 688 7 1 2 2512 687
0 689 5 1 1 688
0 690 7 3 2 2514 689
0 691 5 1 1 2532
0 692 7 2 2 2530 691
0 693 5 1 1 2535
0 694 7 1 2 2022 693
0 695 5 2 1 694
0 696 7 1 2 1874 2536
0 697 5 1 1 696
0 698 7 2 2 2537 697
0 699 5 1 1 2539
0 700 7 2 2 2017 2540
0 701 5 2 1 2541
0 702 7 1 2 675 2538
0 703 5 1 1 702
0 704 7 1 2 2525 2533
0 705 5 1 1 704
0 706 7 2 2 703 705
0 707 5 1 1 2545
0 708 7 1 2 2543 707
0 709 5 2 1 708
0 710 7 1 2 2527 2534
0 711 5 1 1 710
0 712 7 1 2 2529 711
0 713 5 1 1 712
0 714 7 3 2 2531 713
0 715 5 1 1 2549
0 716 7 2 2 2547 715
0 717 5 1 1 2552
0 718 7 1 2 2018 717
0 719 5 2 1 718
0 720 7 1 2 1871 2553
0 721 5 1 1 720
0 722 7 2 2 2554 721
0 723 5 1 1 2556
0 724 7 2 2 2013 2557
0 725 5 2 1 2558
0 726 7 1 2 699 2555
0 727 5 1 1 726
0 728 7 1 2 2542 2550
0 729 5 1 1 728
0 730 7 2 2 727 729
0 731 5 1 1 2562
0 732 7 1 2 2560 731
0 733 5 2 1 732
0 734 7 1 2 2544 2551
0 735 5 1 1 734
0 736 7 1 2 2546 735
0 737 5 1 1 736
0 738 7 3 2 2548 737
0 739 5 1 1 2566
0 740 7 2 2 2564 739
0 741 5 1 1 2569
0 742 7 1 2 2014 741
0 743 5 2 1 742
0 744 7 1 2 1868 2570
0 745 5 1 1 744
0 746 7 2 2 2571 745
0 747 5 1 1 2573
0 748 7 2 2 2010 2574
0 749 5 2 1 2575
0 750 7 1 2 723 2572
0 751 5 1 1 750
0 752 7 1 2 2559 2567
0 753 5 1 1 752
0 754 7 2 2 751 753
0 755 5 1 1 2579
0 756 7 1 2 2577 755
0 757 5 2 1 756
0 758 7 1 2 2561 2568
0 759 5 1 1 758
0 760 7 1 2 2563 759
0 761 5 1 1 760
0 762 7 3 2 2565 761
0 763 5 1 1 2583
0 764 7 2 2 2581 763
0 765 5 1 1 2586
0 766 7 1 2 2011 765
0 767 5 2 1 766
0 768 7 1 2 1865 2587
0 769 5 1 1 768
0 770 7 2 2 2588 769
0 771 5 1 1 2590
0 772 7 2 2 2007 2591
0 773 5 2 1 2592
0 774 7 1 2 747 2589
0 775 5 1 1 774
0 776 7 1 2 2576 2584
0 777 5 1 1 776
0 778 7 2 2 775 777
0 779 5 1 1 2596
0 780 7 1 2 2594 779
0 781 5 2 1 780
0 782 7 1 2 2578 2585
0 783 5 1 1 782
0 784 7 1 2 2580 783
0 785 5 1 1 784
0 786 7 3 2 2582 785
0 787 5 1 1 2600
0 788 7 2 2 2598 787
0 789 5 1 1 2603
0 790 7 1 2 2008 789
0 791 5 2 1 790
0 792 7 1 2 1862 2604
0 793 5 1 1 792
0 794 7 2 2 2605 793
0 795 5 1 1 2607
0 796 7 2 2 2004 2608
0 797 5 2 1 2609
0 798 7 1 2 771 2606
0 799 5 1 1 798
0 800 7 1 2 2593 2601
0 801 5 1 1 800
0 802 7 2 2 799 801
0 803 5 1 1 2613
0 804 7 1 2 2611 803
0 805 5 2 1 804
0 806 7 1 2 2595 2602
0 807 5 1 1 806
0 808 7 1 2 2597 807
0 809 5 1 1 808
0 810 7 3 2 2599 809
0 811 5 1 1 2617
0 812 7 2 2 2615 811
0 813 5 1 1 2620
0 814 7 1 2 2005 813
0 815 5 2 1 814
0 816 7 1 2 1859 2621
0 817 5 1 1 816
0 818 7 2 2 2622 817
0 819 5 1 1 2624
0 820 7 2 2 2001 2625
0 821 5 2 1 2626
0 822 7 1 2 795 2623
0 823 5 1 1 822
0 824 7 1 2 2610 2618
0 825 5 1 1 824
0 826 7 2 2 823 825
0 827 5 1 1 2630
0 828 7 1 2 2628 827
0 829 5 2 1 828
0 830 7 1 2 2612 2619
0 831 5 1 1 830
0 832 7 1 2 2614 831
0 833 5 1 1 832
0 834 7 3 2 2616 833
0 835 5 1 1 2634
0 836 7 2 2 2632 835
0 837 5 1 1 2637
0 838 7 1 2 2002 837
0 839 5 2 1 838
0 840 7 1 2 1856 2638
0 841 5 1 1 840
0 842 7 2 2 2639 841
0 843 5 1 1 2641
0 844 7 2 2 1998 2642
0 845 5 2 1 2643
0 846 7 1 2 819 2640
0 847 5 1 1 846
0 848 7 1 2 2627 2635
0 849 5 1 1 848
0 850 7 2 2 847 849
0 851 5 1 1 2647
0 852 7 1 2 2645 851
0 853 5 2 1 852
0 854 7 1 2 2629 2636
0 855 5 1 1 854
0 856 7 1 2 2631 855
0 857 5 1 1 856
0 858 7 3 2 2633 857
0 859 5 1 1 2651
0 860 7 2 2 2649 859
0 861 5 1 1 2654
0 862 7 1 2 1999 861
0 863 5 2 1 862
0 864 7 1 2 1853 2655
0 865 5 1 1 864
0 866 7 2 2 2656 865
0 867 5 1 1 2658
0 868 7 2 2 1995 2659
0 869 5 2 1 2660
0 870 7 1 2 843 2657
0 871 5 1 1 870
0 872 7 1 2 2644 2652
0 873 5 1 1 872
0 874 7 2 2 871 873
0 875 5 1 1 2664
0 876 7 1 2 2662 875
0 877 5 2 1 876
0 878 7 1 2 2646 2653
0 879 5 1 1 878
0 880 7 1 2 2648 879
0 881 5 1 1 880
0 882 7 3 2 2650 881
0 883 5 1 1 2668
0 884 7 2 2 2666 883
0 885 5 1 1 2671
0 886 7 1 2 1996 885
0 887 5 2 1 886
0 888 7 1 2 1850 2672
0 889 5 1 1 888
0 890 7 2 2 2673 889
0 891 5 1 1 2675
0 892 7 2 2 1992 2676
0 893 5 2 1 2677
0 894 7 1 2 867 2674
0 895 5 1 1 894
0 896 7 1 2 2661 2669
0 897 5 1 1 896
0 898 7 2 2 895 897
0 899 5 1 1 2681
0 900 7 1 2 2679 899
0 901 5 2 1 900
0 902 7 1 2 2663 2670
0 903 5 1 1 902
0 904 7 1 2 2665 903
0 905 5 1 1 904
0 906 7 3 2 2667 905
0 907 5 1 1 2685
0 908 7 2 2 2683 907
0 909 5 1 1 2688
0 910 7 1 2 1993 909
0 911 5 2 1 910
0 912 7 1 2 1847 2689
0 913 5 1 1 912
0 914 7 2 2 2690 913
0 915 5 1 1 2692
0 916 7 2 2 1989 2693
0 917 5 2 1 2694
0 918 7 1 2 891 2691
0 919 5 1 1 918
0 920 7 1 2 2678 2686
0 921 5 1 1 920
0 922 7 2 2 919 921
0 923 5 1 1 2698
0 924 7 1 2 2696 923
0 925 5 2 1 924
0 926 7 1 2 2680 2687
0 927 5 1 1 926
0 928 7 1 2 2682 927
0 929 5 1 1 928
0 930 7 3 2 2684 929
0 931 5 1 1 2702
0 932 7 2 2 2700 931
0 933 5 1 1 2705
0 934 7 1 2 1990 933
0 935 5 2 1 934
0 936 7 1 2 1844 2706
0 937 5 1 1 936
0 938 7 2 2 2707 937
0 939 5 1 1 2709
0 940 7 2 2 1986 2710
0 941 5 2 1 2711
0 942 7 1 2 915 2708
0 943 5 1 1 942
0 944 7 1 2 2695 2703
0 945 5 1 1 944
0 946 7 2 2 943 945
0 947 5 1 1 2715
0 948 7 1 2 2713 947
0 949 5 2 1 948
0 950 7 1 2 2697 2704
0 951 5 1 1 950
0 952 7 1 2 2699 951
0 953 5 1 1 952
0 954 7 3 2 2701 953
0 955 5 1 1 2719
0 956 7 2 2 2717 955
0 957 5 1 1 2722
0 958 7 1 2 1987 957
0 959 5 2 1 958
0 960 7 1 2 1841 2723
0 961 5 1 1 960
0 962 7 2 2 2724 961
0 963 5 1 1 2726
0 964 7 2 2 1983 2727
0 965 5 2 1 2728
0 966 7 1 2 939 2725
0 967 5 1 1 966
0 968 7 1 2 2712 2720
0 969 5 1 1 968
0 970 7 2 2 967 969
0 971 5 1 1 2732
0 972 7 1 2 2730 971
0 973 5 2 1 972
0 974 7 1 2 2714 2721
0 975 5 1 1 974
0 976 7 1 2 2716 975
0 977 5 1 1 976
0 978 7 3 2 2718 977
0 979 5 1 1 2736
0 980 7 2 2 2734 979
0 981 5 1 1 2739
0 982 7 1 2 1984 981
0 983 5 2 1 982
0 984 7 1 2 1838 2740
0 985 5 1 1 984
0 986 7 2 2 2741 985
0 987 5 1 1 2743
0 988 7 2 2 1980 2744
0 989 5 2 1 2745
0 990 7 1 2 963 2742
0 991 5 1 1 990
0 992 7 1 2 2729 2737
0 993 5 1 1 992
0 994 7 2 2 991 993
0 995 5 1 1 2749
0 996 7 1 2 2747 995
0 997 5 2 1 996
0 998 7 1 2 2731 2738
0 999 5 1 1 998
0 1000 7 1 2 2733 999
0 1001 5 1 1 1000
0 1002 7 3 2 2735 1001
0 1003 5 1 1 2753
0 1004 7 2 2 2751 1003
0 1005 5 1 1 2756
0 1006 7 1 2 1981 1005
0 1007 5 2 1 1006
0 1008 7 1 2 1835 2757
0 1009 5 1 1 1008
0 1010 7 2 2 2758 1009
0 1011 5 1 1 2760
0 1012 7 2 2 1977 2761
0 1013 5 2 1 2762
0 1014 7 1 2 987 2759
0 1015 5 1 1 1014
0 1016 7 1 2 2746 2754
0 1017 5 1 1 1016
0 1018 7 2 2 1015 1017
0 1019 5 1 1 2766
0 1020 7 1 2 2764 1019
0 1021 5 2 1 1020
0 1022 7 1 2 2748 2755
0 1023 5 1 1 1022
0 1024 7 1 2 2750 1023
0 1025 5 1 1 1024
0 1026 7 3 2 2752 1025
0 1027 5 1 1 2770
0 1028 7 2 2 2768 1027
0 1029 5 1 1 2773
0 1030 7 1 2 1978 1029
0 1031 5 2 1 1030
0 1032 7 1 2 1832 2774
0 1033 5 1 1 1032
0 1034 7 2 2 2775 1033
0 1035 5 1 1 2777
0 1036 7 2 2 1974 2778
0 1037 5 2 1 2779
0 1038 7 1 2 1011 2776
0 1039 5 1 1 1038
0 1040 7 1 2 2763 2771
0 1041 5 1 1 1040
0 1042 7 2 2 1039 1041
0 1043 5 1 1 2783
0 1044 7 1 2 2781 1043
0 1045 5 2 1 1044
0 1046 7 1 2 2765 2772
0 1047 5 1 1 1046
0 1048 7 1 2 2767 1047
0 1049 5 1 1 1048
0 1050 7 3 2 2769 1049
0 1051 5 1 1 2787
0 1052 7 2 2 2785 1051
0 1053 5 1 1 2790
0 1054 7 1 2 1975 1053
0 1055 5 2 1 1054
0 1056 7 1 2 1829 2791
0 1057 5 1 1 1056
0 1058 7 2 2 2792 1057
0 1059 5 1 1 2794
0 1060 7 2 2 1971 2795
0 1061 5 2 1 2796
0 1062 7 1 2 1035 2793
0 1063 5 1 1 1062
0 1064 7 1 2 2780 2788
0 1065 5 1 1 1064
0 1066 7 2 2 1063 1065
0 1067 5 1 1 2800
0 1068 7 1 2 2798 1067
0 1069 5 2 1 1068
0 1070 7 1 2 2782 2789
0 1071 5 1 1 1070
0 1072 7 1 2 2784 1071
0 1073 5 1 1 1072
0 1074 7 3 2 2786 1073
0 1075 5 1 1 2804
0 1076 7 2 2 2802 1075
0 1077 5 1 1 2807
0 1078 7 1 2 1972 1077
0 1079 5 2 1 1078
0 1080 7 1 2 1826 2808
0 1081 5 1 1 1080
0 1082 7 2 2 2809 1081
0 1083 5 1 1 2811
0 1084 7 2 2 1968 2812
0 1085 5 2 1 2813
0 1086 7 1 2 1059 2810
0 1087 5 1 1 1086
0 1088 7 1 2 2797 2805
0 1089 5 1 1 1088
0 1090 7 2 2 1087 1089
0 1091 5 1 1 2817
0 1092 7 1 2 2815 1091
0 1093 5 2 1 1092
0 1094 7 1 2 2799 2806
0 1095 5 1 1 1094
0 1096 7 1 2 2801 1095
0 1097 5 1 1 1096
0 1098 7 3 2 2803 1097
0 1099 5 1 1 2821
0 1100 7 2 2 2819 1099
0 1101 5 1 1 2824
0 1102 7 1 2 1969 1101
0 1103 5 2 1 1102
0 1104 7 1 2 1823 2825
0 1105 5 1 1 1104
0 1106 7 2 2 2826 1105
0 1107 5 1 1 2828
0 1108 7 2 2 1965 2829
0 1109 5 2 1 2830
0 1110 7 1 2 1083 2827
0 1111 5 1 1 1110
0 1112 7 1 2 2814 2822
0 1113 5 1 1 1112
0 1114 7 2 2 1111 1113
0 1115 5 1 1 2834
0 1116 7 1 2 2832 1115
0 1117 5 2 1 1116
0 1118 7 1 2 2816 2823
0 1119 5 1 1 1118
0 1120 7 1 2 2818 1119
0 1121 5 1 1 1120
0 1122 7 3 2 2820 1121
0 1123 5 1 1 2838
0 1124 7 2 2 2836 1123
0 1125 5 1 1 2841
0 1126 7 1 2 1820 2842
0 1127 5 1 1 1126
0 1128 7 1 2 1966 1125
0 1129 5 2 1 1128
0 1130 7 2 2 1127 2843
0 1131 5 1 1 2845
0 1132 7 2 2 1962 2846
0 1133 5 2 1 2847
0 1134 7 1 2 1107 2844
0 1135 5 1 1 1134
0 1136 7 1 2 2831 2839
0 1137 5 1 1 1136
0 1138 7 2 2 1135 1137
0 1139 5 1 1 2851
0 1140 7 1 2 2849 1139
0 1141 5 2 1 1140
0 1142 7 1 2 2833 2840
0 1143 5 1 1 1142
0 1144 7 1 2 2835 1143
0 1145 5 1 1 1144
0 1146 7 3 2 2837 1145
0 1147 5 1 1 2855
0 1148 7 1 2 2850 2856
0 1149 5 1 1 1148
0 1150 7 1 2 2852 1149
0 1151 5 1 1 1150
0 1152 7 1 2 2853 1151
0 1153 5 1 1 1152
0 1154 7 2 2 2854 1147
0 1155 5 1 1 2858
0 1156 7 1 2 1963 1155
0 1157 5 2 1 1156
0 1158 7 1 2 1817 2859
0 1159 5 1 1 1158
0 1160 7 2 2 2860 1159
0 1161 5 1 1 2862
0 1162 7 1 2 1814 1161
0 1163 5 1 1 1162
0 1164 7 1 2 1153 1163
0 1165 5 1 1 1164
0 1166 7 1 2 1131 2861
0 1167 5 1 1 1166
0 1168 7 1 2 2848 2857
0 1169 5 1 1 1168
0 1170 7 2 2 1167 1169
0 1171 5 1 1 2864
0 1172 7 1 2 1165 2865
0 1173 5 1 1 1172
0 1174 7 1 2 1960 2863
0 1175 7 1 2 1171 1174
0 1176 5 1 1 1175
0 1177 7 2 2 1173 1176
0 1178 5 1 1 2866
0 1179 7 1 2 1964 2012
0 1180 5 2 1 1179
0 1181 7 1 2 1818 1866
0 1182 5 2 1 1181
0 1183 7 1 2 1961 2009
0 1184 5 2 1 1183
0 1185 7 1 2 1815 1863
0 1186 5 2 1 1185
0 1187 7 2 2 1812 1860
0 1188 5 3 1 2876
0 1189 7 1 2 2874 2878
0 1190 5 1 1 1189
0 1191 7 2 2 2872 1190
0 1192 5 2 1 2881
0 1193 7 1 2 2870 2883
0 1194 5 1 1 1193
0 1195 7 2 2 2868 1194
0 1196 5 1 1 2885
0 1197 7 1 2 1967 1196
0 1198 5 2 1 1197
0 1199 7 1 2 1821 2886
0 1200 5 2 1 1199
0 1201 7 1 2 2015 2889
0 1202 5 1 1 1201
0 1203 7 2 2 2887 1202
0 1204 5 1 1 2891
0 1205 7 1 2 1970 1204
0 1206 5 2 1 1205
0 1207 7 1 2 1824 2892
0 1208 5 2 1 1207
0 1209 7 1 2 2019 2895
0 1210 5 1 1 1209
0 1211 7 2 2 2893 1210
0 1212 5 1 1 2897
0 1213 7 1 2 1973 1212
0 1214 5 2 1 1213
0 1215 7 1 2 1827 2898
0 1216 5 2 1 1215
0 1217 7 1 2 2023 2901
0 1218 5 1 1 1217
0 1219 7 2 2 2899 1218
0 1220 5 1 1 2903
0 1221 7 1 2 1976 1220
0 1222 5 2 1 1221
0 1223 7 1 2 1830 2904
0 1224 5 2 1 1223
0 1225 7 1 2 2027 2907
0 1226 5 1 1 1225
0 1227 7 2 2 2905 1226
0 1228 5 1 1 2909
0 1229 7 1 2 1979 1228
0 1230 5 2 1 1229
0 1231 7 1 2 1833 2910
0 1232 5 2 1 1231
0 1233 7 1 2 2031 2913
0 1234 5 1 1 1233
0 1235 7 2 2 2911 1234
0 1236 5 1 1 2915
0 1237 7 1 2 1982 1236
0 1238 5 2 1 1237
0 1239 7 1 2 1836 2916
0 1240 5 2 1 1239
0 1241 7 1 2 2035 2919
0 1242 5 1 1 1241
0 1243 7 2 2 2917 1242
0 1244 5 1 1 2921
0 1245 7 1 2 1985 1244
0 1246 5 2 1 1245
0 1247 7 1 2 1839 2922
0 1248 5 2 1 1247
0 1249 7 1 2 2039 2925
0 1250 5 1 1 1249
0 1251 7 2 2 2923 1250
0 1252 5 1 1 2927
0 1253 7 1 2 1988 1252
0 1254 5 2 1 1253
0 1255 7 1 2 1842 2928
0 1256 5 2 1 1255
0 1257 7 1 2 2043 2931
0 1258 5 1 1 1257
0 1259 7 2 2 2929 1258
0 1260 5 1 1 2933
0 1261 7 1 2 1991 1260
0 1262 5 2 1 1261
0 1263 7 1 2 1845 2934
0 1264 5 2 1 1263
0 1265 7 1 2 2047 2937
0 1266 5 1 1 1265
0 1267 7 2 2 2935 1266
0 1268 5 1 1 2939
0 1269 7 1 2 1994 1268
0 1270 5 2 1 1269
0 1271 7 1 2 1848 2940
0 1272 5 2 1 1271
0 1273 7 1 2 2051 2943
0 1274 5 1 1 1273
0 1275 7 2 2 2941 1274
0 1276 5 1 1 2945
0 1277 7 1 2 1997 1276
0 1278 5 2 1 1277
0 1279 7 1 2 1851 2946
0 1280 5 2 1 1279
0 1281 7 1 2 2055 2949
0 1282 5 1 1 1281
0 1283 7 2 2 2947 1282
0 1284 5 1 1 2951
0 1285 7 1 2 2000 1284
0 1286 5 2 1 1285
0 1287 7 1 2 1854 2952
0 1288 5 2 1 1287
0 1289 7 1 2 2059 2955
0 1290 5 1 1 1289
0 1291 7 2 2 2953 1290
0 1292 5 1 1 2957
0 1293 7 1 2 2003 1292
0 1294 5 2 1 1293
0 1295 7 1 2 1857 2958
0 1296 5 2 1 1295
0 1297 7 1 2 2063 2961
0 1298 5 1 1 1297
0 1299 7 2 2 2959 1298
0 1300 5 1 1 2963
0 1301 7 2 2 1959 1300
0 1302 5 2 1 2965
0 1303 7 1 2 2114 2964
0 1304 5 3 1 1303
0 1305 7 2 2 2960 2962
0 1306 5 1 1 2972
0 1307 7 1 2 1905 2973
0 1308 5 1 1 1307
0 1309 7 1 2 2064 1306
0 1310 5 1 1 1309
0 1311 7 2 2 1308 1310
0 1312 5 1 1 2974
0 1313 7 1 2 1955 1312
0 1314 5 4 1 1313
0 1315 7 1 2 2112 2975
0 1316 5 5 1 1315
0 1317 7 2 2 2954 2956
0 1318 5 1 1 2985
0 1319 7 1 2 1902 2986
0 1320 5 1 1 1319
0 1321 7 1 2 2060 1318
0 1322 5 1 1 1321
0 1323 7 2 2 1320 1322
0 1324 5 1 1 2987
0 1325 7 1 2 1951 1324
0 1326 5 3 1 1325
0 1327 7 1 2 2110 2988
0 1328 5 4 1 1327
0 1329 7 2 2 2948 2950
0 1330 5 1 1 2996
0 1331 7 1 2 1899 2997
0 1332 5 1 1 1331
0 1333 7 1 2 2056 1330
0 1334 5 1 1 1333
0 1335 7 2 2 1332 1334
0 1336 5 1 1 2998
0 1337 7 1 2 1948 1336
0 1338 5 3 1 1337
0 1339 7 1 2 2107 2999
0 1340 5 4 1 1339
0 1341 7 2 2 2942 2944
0 1342 5 1 1 3007
0 1343 7 1 2 1896 3008
0 1344 5 1 1 1343
0 1345 7 1 2 2052 1342
0 1346 5 1 1 1345
0 1347 7 2 2 1344 1346
0 1348 5 1 1 3009
0 1349 7 1 2 1944 1348
0 1350 5 3 1 1349
0 1351 7 1 2 2103 3010
0 1352 5 4 1 1351
0 1353 7 2 2 2936 2938
0 1354 5 1 1 3018
0 1355 7 1 2 1893 3019
0 1356 5 1 1 1355
0 1357 7 1 2 2048 1354
0 1358 5 1 1 1357
0 1359 7 2 2 1356 1358
0 1360 5 1 1 3020
0 1361 7 1 2 1941 1360
0 1362 5 4 1 1361
0 1363 7 1 2 2100 3021
0 1364 5 4 1 1363
0 1365 7 2 2 2930 2932
0 1366 5 1 1 3030
0 1367 7 1 2 1890 3031
0 1368 5 1 1 1367
0 1369 7 1 2 2044 1366
0 1370 5 1 1 1369
0 1371 7 2 2 1368 1370
0 1372 5 1 1 3032
0 1373 7 2 2 2097 3033
0 1374 5 4 1 3034
0 1375 7 1 2 1938 1372
0 1376 5 4 1 1375
0 1377 7 2 2 2924 2926
0 1378 5 1 1 3044
0 1379 7 1 2 1887 3045
0 1380 5 1 1 1379
0 1381 7 1 2 2040 1378
0 1382 5 1 1 1381
0 1383 7 2 2 1380 1382
0 1384 5 1 1 3046
0 1385 7 1 2 2094 3047
0 1386 5 5 1 1385
0 1387 7 1 2 1935 1384
0 1388 5 4 1 1387
0 1389 7 2 2 2918 2920
0 1390 5 1 1 3057
0 1391 7 1 2 1884 3058
0 1392 5 1 1 1391
0 1393 7 1 2 2036 1390
0 1394 5 1 1 1393
0 1395 7 2 2 1392 1394
0 1396 5 1 1 3059
0 1397 7 1 2 2091 3060
0 1398 5 5 1 1397
0 1399 7 1 2 1932 1396
0 1400 5 3 1 1399
0 1401 7 2 2 2912 2914
0 1402 5 1 1 3069
0 1403 7 1 2 1881 3070
0 1404 5 1 1 1403
0 1405 7 1 2 2032 1402
0 1406 5 1 1 1405
0 1407 7 2 2 1404 1406
0 1408 5 1 1 3071
0 1409 7 1 2 2088 3072
0 1410 5 5 1 1409
0 1411 7 1 2 1929 1408
0 1412 5 4 1 1411
0 1413 7 2 2 2900 2902
0 1414 5 1 1 3082
0 1415 7 1 2 1875 3083
0 1416 5 1 1 1415
0 1417 7 1 2 2024 1414
0 1418 5 1 1 1417
0 1419 7 2 2 1416 1418
0 1420 5 1 1 3084
0 1421 7 1 2 1923 1420
0 1422 5 4 1 1421
0 1423 7 2 2 2894 2896
0 1424 5 1 1 3090
0 1425 7 1 2 1872 3091
0 1426 5 1 1 1425
0 1427 7 1 2 2020 1424
0 1428 5 1 1 1427
0 1429 7 2 2 1426 1428
0 1430 5 1 1 3092
0 1431 7 1 2 2079 3093
0 1432 5 4 1 1431
0 1433 7 1 2 1920 1430
0 1434 5 3 1 1433
0 1435 7 2 2 2888 2890
0 1436 5 1 1 3101
0 1437 7 1 2 1869 3102
0 1438 5 1 1 1437
0 1439 7 1 2 2016 1436
0 1440 5 1 1 1439
0 1441 7 2 2 1438 1440
0 1442 5 1 1 3103
0 1443 7 1 2 2076 3104
0 1444 5 4 1 1443
0 1445 7 1 2 1917 1442
0 1446 5 3 1 1445
0 1447 7 2 2 2869 2871
0 1448 5 1 1 3112
0 1449 7 1 2 2882 1448
0 1450 5 1 1 1449
0 1451 7 1 2 2884 3113
0 1452 5 1 1 1451
0 1453 7 2 2 1450 1452
0 1454 5 1 1 3114
0 1455 7 1 2 1914 3115
0 1456 5 2 1 1455
0 1457 7 2 2 2873 2875
0 1458 5 1 1 3118
0 1459 7 1 2 2877 1458
0 1460 5 1 1 1459
0 1461 7 1 2 2879 3119
0 1462 5 1 1 1461
0 1463 7 2 2 1460 1462
0 1464 5 1 1 3120
0 1465 7 1 2 1911 3121
0 1466 5 1 1 1465
0 1467 7 2 2 3116 1466
0 1468 5 1 1 3122
0 1469 7 1 2 50 2006
0 1470 5 1 1 1469
0 1471 7 2 2 2880 1470
0 1472 5 1 1 3124
0 1473 7 1 2 1908 1472
0 1474 5 1 1 1473
0 1475 7 2 2 3123 1474
0 1476 5 1 1 3126
0 1477 7 2 2 2070 1464
0 1478 5 1 1 3128
0 1479 7 1 2 3117 3129
0 1480 5 1 1 1479
0 1481 7 1 2 2073 1454
0 1482 5 3 1 1481
0 1483 7 1 2 1480 3130
0 1484 7 2 2 1476 1483
0 1485 5 2 1 3133
0 1486 7 1 2 3109 3135
0 1487 5 1 1 1486
0 1488 7 2 2 3105 1487
0 1489 5 2 1 3137
0 1490 7 1 2 3098 3139
0 1491 5 1 1 1490
0 1492 7 2 2 3094 1491
0 1493 5 1 1 3141
0 1494 7 1 2 3086 1493
0 1495 5 2 1 1494
0 1496 7 2 2 2906 2908
0 1497 5 1 1 3145
0 1498 7 1 2 1878 3146
0 1499 5 1 1 1498
0 1500 7 1 2 2028 1497
0 1501 5 1 1 1500
0 1502 7 2 2 1499 1501
0 1503 5 1 1 3147
0 1504 7 1 2 2085 3148
0 1505 5 4 1 1504
0 1506 7 1 2 2082 3085
0 1507 5 4 1 1506
0 1508 7 2 2 3149 3153
0 1509 7 1 2 3143 3157
0 1510 5 1 1 1509
0 1511 7 1 2 1926 1503
0 1512 5 4 1 1511
0 1513 7 1 2 1510 3159
0 1514 7 1 2 3078 1513
0 1515 5 2 1 1514
0 1516 7 1 2 3073 3163
0 1517 5 1 1 1516
0 1518 7 1 2 3066 1517
0 1519 5 1 1 1518
0 1520 7 1 2 3061 1519
0 1521 5 1 1 1520
0 1522 7 2 2 3053 1521
0 1523 5 1 1 3165
0 1524 7 1 2 3048 1523
0 1525 5 2 1 1524
0 1526 7 1 2 3040 3167
0 1527 5 1 1 1526
0 1528 7 1 2 3036 1527
0 1529 7 2 2 3026 1528
0 1530 5 1 1 3169
0 1531 7 2 2 3022 1530
0 1532 5 2 1 3171
0 1533 7 1 2 3014 3173
0 1534 5 1 1 1533
0 1535 7 2 2 3011 1534
0 1536 5 2 1 3175
0 1537 7 1 2 3003 3177
0 1538 5 1 1 1537
0 1539 7 2 2 3000 1538
0 1540 5 2 1 3179
0 1541 7 1 2 2992 3181
0 1542 5 1 1 1541
0 1543 7 2 2 2989 1542
0 1544 5 1 1 3183
0 1545 7 1 2 2980 1544
0 1546 5 2 1 1545
0 1547 7 1 2 2976 3185
0 1548 5 1 1 1547
0 1549 7 1 2 2969 1548
0 1550 5 1 1 1549
0 1551 7 2 2 2967 1550
0 1552 5 1 1 3187
0 1553 7 2 2 2970 3186
0 1554 5 1 1 3189
0 1555 7 1 2 2977 1554
0 1556 5 1 1 1555
0 1557 7 1 2 2978 2981
0 1558 5 2 1 1557
0 1559 7 1 2 3184 3191
0 1560 5 1 1 1559
0 1561 7 3 2 2990 2993
0 1562 5 2 1 3193
0 1563 7 1 2 3182 3194
0 1564 5 1 1 1563
0 1565 7 1 2 3180 3196
0 1566 5 1 1 1565
0 1567 7 3 2 3001 3004
0 1568 5 2 1 3198
0 1569 7 1 2 3178 3199
0 1570 5 1 1 1569
0 1571 7 1 2 3176 3201
0 1572 5 1 1 1571
0 1573 7 3 2 3012 3015
0 1574 5 2 1 3203
0 1575 7 1 2 3174 3204
0 1576 5 1 1 1575
0 1577 7 1 2 3172 3206
0 1578 5 1 1 1577
0 1579 7 1 2 3023 3170
0 1580 5 1 1 1579
0 1581 7 2 2 3024 3027
0 1582 5 2 1 3208
0 1583 7 1 2 3041 3210
0 1584 5 1 1 1583
0 1585 7 1 2 3042 3037
0 1586 5 2 1 1585
0 1587 7 1 2 3212 3168
0 1588 5 1 1 1587
0 1589 7 1 2 3049 3054
0 1590 5 2 1 1589
0 1591 7 1 2 3062 3214
0 1592 5 1 1 1591
0 1593 7 1 2 3050 3166
0 1594 5 1 1 1593
0 1595 7 3 2 3063 3067
0 1596 5 1 1 3216
0 1597 7 1 2 3164 3217
0 1598 5 1 1 1597
0 1599 7 1 2 3074 1598
0 1600 5 1 1 1599
0 1601 7 1 2 3075 3079
0 1602 5 2 1 1601
0 1603 7 1 2 3150 3219
0 1604 5 1 1 1603
0 1605 7 2 2 3151 3160
0 1606 7 1 2 3144 3221
0 1607 5 1 1 1606
0 1608 7 1 2 3154 1607
0 1609 5 1 1 1608
0 1610 7 1 2 3087 3155
0 1611 5 2 1 1610
0 1612 7 1 2 3142 3223
0 1613 5 1 1 1612
0 1614 7 3 2 3095 3099
0 1615 5 2 1 3225
0 1616 7 1 2 3138 3226
0 1617 5 1 1 1616
0 1618 7 3 2 3106 3110
0 1619 5 2 1 3230
0 1620 7 1 2 3136 3231
0 1621 5 1 1 1620
0 1622 7 1 2 2067 3125
0 1623 5 1 1 1622
0 1624 7 1 2 1478 1623
0 1625 7 3 2 3131 1624
0 1626 5 1 1 3235
0 1627 7 1 2 3127 3236
0 1628 5 2 1 1627
0 1629 7 1 2 3134 3233
0 1630 5 1 1 1629
0 1631 7 1 2 3238 1630
0 1632 7 1 2 1621 1631
0 1633 5 1 1 1632
0 1634 7 1 2 3140 3228
0 1635 5 1 1 1634
0 1636 7 1 2 1633 1635
0 1637 7 1 2 1617 1636
0 1638 5 1 1 1637
0 1639 7 1 2 1613 1638
0 1640 7 1 2 1609 1639
0 1641 7 1 2 1604 1640
0 1642 7 1 2 1600 1641
0 1643 7 1 2 1594 1642
0 1644 7 1 2 1592 1643
0 1645 5 1 1 1644
0 1646 7 1 2 1588 1645
0 1647 7 1 2 1584 1646
0 1648 7 1 2 1580 1647
0 1649 7 1 2 1578 1648
0 1650 7 1 2 1576 1649
0 1651 7 1 2 1572 1650
0 1652 7 1 2 1570 1651
0 1653 7 1 2 1566 1652
0 1654 7 1 2 1564 1653
0 1655 7 1 2 1560 1654
0 1656 7 1 2 1556 1655
0 1657 7 1 2 3188 1656
0 1658 5 1 1 1657
0 1659 7 1 2 1468 3132
0 1660 5 1 1 1659
0 1661 7 2 2 1626 1660
0 1662 5 2 1 3240
0 1663 7 1 2 3107 3242
0 1664 5 1 1 1663
0 1665 7 2 2 3111 1664
0 1666 5 2 1 3244
0 1667 7 1 2 3096 3246
0 1668 5 1 1 1667
0 1669 7 2 2 3100 1668
0 1670 5 1 1 3248
0 1671 7 1 2 3156 1670
0 1672 5 2 1 1671
0 1673 7 1 2 3088 3250
0 1674 7 1 2 3161 1673
0 1675 5 1 1 1674
0 1676 7 1 2 3152 1675
0 1677 7 1 2 3076 1676
0 1678 5 1 1 1677
0 1679 7 1 2 3080 1678
0 1680 5 2 1 1679
0 1681 7 1 2 3064 3252
0 1682 5 1 1 1681
0 1683 7 2 2 3068 1682
0 1684 5 1 1 3254
0 1685 7 2 2 3051 1684
0 1686 5 1 1 3256
0 1687 7 1 2 3055 1686
0 1688 5 2 1 1687
0 1689 7 1 2 3038 3258
0 1690 5 1 1 1689
0 1691 7 1 2 3043 1690
0 1692 5 2 1 1691
0 1693 7 1 2 3028 3260
0 1694 5 1 1 1693
0 1695 7 2 2 3025 1694
0 1696 5 2 1 3262
0 1697 7 1 2 3016 3264
0 1698 5 1 1 1697
0 1699 7 2 2 3013 1698
0 1700 5 2 1 3266
0 1701 7 1 2 3005 3268
0 1702 5 1 1 1701
0 1703 7 2 2 3002 1702
0 1704 5 2 1 3270
0 1705 7 1 2 2994 3272
0 1706 5 1 1 1705
0 1707 7 1 2 2991 1706
0 1708 5 2 1 1707
0 1709 7 1 2 2982 3274
0 1710 5 1 1 1709
0 1711 7 2 2 2968 2979
0 1712 7 1 2 1710 3276
0 1713 5 1 1 1712
0 1714 7 1 2 3192 3275
0 1715 5 1 1 1714
0 1716 7 1 2 2966 2983
0 1717 5 1 1 1716
0 1718 7 1 2 3195 3273
0 1719 5 1 1 1718
0 1720 7 1 2 3197 3271
0 1721 5 1 1 1720
0 1722 7 1 2 1719 1721
0 1723 5 1 1 1722
0 1724 7 1 2 3200 3267
0 1725 5 1 1 1724
0 1726 7 1 2 3202 3269
0 1727 5 1 1 1726
0 1728 7 1 2 3207 3263
0 1729 5 1 1 1728
0 1730 7 1 2 3205 3265
0 1731 5 1 1 1730
0 1732 7 1 2 1729 1731
0 1733 5 1 1 1732
0 1734 7 1 2 3035 3211
0 1735 5 1 1 1734
0 1736 7 1 2 3209 3261
0 1737 5 1 1 1736
0 1738 7 1 2 1735 1737
0 1739 5 1 1 1738
0 1740 7 1 2 3213 3259
0 1741 5 1 1 1740
0 1742 7 1 2 3215 3255
0 1743 5 1 1 1742
0 1744 7 1 2 3056 3257
0 1745 5 1 1 1744
0 1746 7 1 2 3081 1596
0 1747 5 1 1 1746
0 1748 7 1 2 3218 3253
0 1749 5 1 1 1748
0 1750 7 1 2 3162 3220
0 1751 5 1 1 1750
0 1752 7 1 2 3222 3251
0 1753 5 1 1 1752
0 1754 7 1 2 3089 1753
0 1755 5 1 1 1754
0 1756 7 1 2 3224 3249
0 1757 5 1 1 1756
0 1758 7 1 2 3227 3245
0 1759 5 1 1 1758
0 1760 7 1 2 3232 3243
0 1761 5 1 1 1760
0 1762 7 1 2 3234 3241
0 1763 5 1 1 1762
0 1764 7 1 2 3239 1763
0 1765 7 1 2 1761 1764
0 1766 5 1 1 1765
0 1767 7 1 2 3229 3247
0 1768 5 1 1 1767
0 1769 7 1 2 1766 1768
0 1770 7 1 2 1759 1769
0 1771 5 1 1 1770
0 1772 7 1 2 1757 1771
0 1773 7 1 2 1755 1772
0 1774 7 1 2 1751 1773
0 1775 7 1 2 1749 1774
0 1776 7 1 2 1747 1775
0 1777 7 1 2 1745 1776
0 1778 7 1 2 1743 1777
0 1779 5 1 1 1778
0 1780 7 1 2 1741 1779
0 1781 7 1 2 1739 1780
0 1782 7 1 2 1733 1781
0 1783 7 1 2 1727 1782
0 1784 7 1 2 1725 1783
0 1785 7 1 2 2971 1784
0 1786 7 1 2 1723 1785
0 1787 7 1 2 1717 1786
0 1788 7 1 2 1715 1787
0 1789 7 1 2 1713 1788
0 1790 7 1 2 1552 1789
0 1791 5 1 1 1790
0 1792 7 1 2 1658 1791
0 1793 7 1 2 2867 1792
0 1794 5 1 1 1793
0 1795 7 1 2 3108 3237
0 1796 7 1 2 3097 1795
0 1797 7 1 2 3158 1796
0 1798 7 1 2 3077 1797
0 1799 7 1 2 3065 1798
0 1800 7 1 2 3052 1799
0 1801 7 1 2 3039 1800
0 1802 7 1 2 3029 1801
0 1803 7 1 2 3017 1802
0 1804 7 1 2 3006 1803
0 1805 7 1 2 2995 1804
0 1806 7 1 2 2984 1805
0 1807 7 1 2 3277 1806
0 1808 7 1 2 3190 1807
0 1809 5 1 1 1808
0 1810 7 1 2 1178 1809
0 1811 5 1 1 1810
3 4099 7 0 2 1794 1811
