1 0 0 2 0
2 32 1 0
2 33 1 0
1 1 0 2 0
2 34 1 1
2 35 1 1
1 2 0 2 0
2 36 1 2
2 37 1 2
1 3 0 2 0
2 38 1 3
2 39 1 3
1 4 0 2 0
2 40 1 4
2 41 1 4
1 5 0 2 0
2 42 1 5
2 43 1 5
1 6 0 2 0
2 44 1 6
2 45 1 6
1 7 0 2 0
2 46 1 7
2 47 1 7
1 8 0 2 0
2 48 1 8
2 85 1 8
1 9 0 2 0
2 97 1 9
2 112 1 9
1 10 0 2 0
2 127 1 10
2 142 1 10
1 11 0 2 0
2 157 1 11
2 172 1 11
1 12 0 2 0
2 187 1 12
2 202 1 12
1 13 0 2 0
2 217 1 13
2 232 1 13
1 14 0 2 0
2 247 1 14
2 262 1 14
1 15 0 2 0
2 277 1 15
2 292 1 15
1 16 0 2 0
2 308 1 16
2 311 1 16
1 17 0 2 0
2 312 1 17
2 313 1 17
1 18 0 2 0
2 314 1 18
2 315 1 18
1 19 0 2 0
2 316 1 19
2 317 1 19
1 20 0 2 0
2 318 1 20
2 319 1 20
1 21 0 2 0
2 320 1 21
2 321 1 21
1 22 0 2 0
2 322 1 22
2 323 1 22
1 23 0 2 0
2 324 1 23
2 325 1 23
1 24 0 2 0
2 326 1 24
2 327 1 24
1 25 0 2 0
2 328 1 25
2 329 1 25
1 26 0 2 0
2 330 1 26
2 331 1 26
1 27 0 2 0
2 332 1 27
2 333 1 27
1 28 0 2 0
2 334 1 28
2 335 1 28
1 29 0 2 0
2 336 1 29
2 337 1 29
1 30 0 2 0
2 338 1 30
2 339 1 30
1 31 0 2 0
2 340 1 31
2 341 1 31
2 342 1 67
2 343 1 67
2 344 1 68
2 345 1 68
2 346 1 69
2 347 1 69
2 348 1 70
2 349 1 70
2 350 1 71
2 351 1 71
2 352 1 72
2 353 1 72
2 354 1 73
2 355 1 73
2 356 1 74
2 357 1 74
2 358 1 75
2 359 1 75
2 360 1 76
2 361 1 76
2 362 1 77
2 363 1 77
2 364 1 78
2 365 1 78
2 366 1 79
2 367 1 79
2 368 1 81
2 369 1 81
2 370 1 82
2 371 1 82
2 372 1 82
2 373 1 87
2 374 1 87
2 375 1 89
2 376 1 89
2 377 1 90
2 378 1 90
2 379 1 100
2 380 1 100
2 381 1 103
2 382 1 103
2 383 1 105
2 384 1 105
2 385 1 106
2 386 1 106
2 387 1 115
2 388 1 115
2 389 1 118
2 390 1 118
2 391 1 120
2 392 1 120
2 393 1 121
2 394 1 121
2 395 1 130
2 396 1 130
2 397 1 133
2 398 1 133
2 399 1 135
2 400 1 135
2 401 1 136
2 402 1 136
2 403 1 145
2 404 1 145
2 405 1 148
2 406 1 148
2 407 1 150
2 408 1 150
2 409 1 151
2 410 1 151
2 411 1 160
2 412 1 160
2 413 1 163
2 414 1 163
2 415 1 165
2 416 1 165
2 417 1 166
2 418 1 166
2 419 1 175
2 420 1 175
2 421 1 178
2 422 1 178
2 423 1 180
2 424 1 180
2 425 1 181
2 426 1 181
2 427 1 190
2 428 1 190
2 429 1 193
2 430 1 193
2 431 1 195
2 432 1 195
2 433 1 196
2 434 1 196
2 435 1 205
2 436 1 205
2 437 1 208
2 438 1 208
2 439 1 210
2 440 1 210
2 441 1 211
2 442 1 211
2 443 1 220
2 444 1 220
2 445 1 223
2 446 1 223
2 447 1 225
2 448 1 225
2 449 1 226
2 450 1 226
2 451 1 235
2 452 1 235
2 453 1 238
2 454 1 238
2 455 1 240
2 456 1 240
2 457 1 241
2 458 1 241
2 459 1 250
2 460 1 250
2 461 1 253
2 462 1 253
2 463 1 255
2 464 1 255
2 465 1 256
2 466 1 256
2 467 1 265
2 468 1 265
2 469 1 268
2 470 1 268
2 471 1 270
2 472 1 270
2 473 1 271
2 474 1 271
2 475 1 280
2 476 1 280
2 477 1 283
2 478 1 283
2 479 1 285
2 480 1 285
2 481 1 286
2 482 1 286
2 483 1 295
2 484 1 295
2 485 1 296
2 486 1 296
2 487 1 298
2 488 1 298
2 489 1 300
2 490 1 300
2 491 1 301
2 492 1 301
0 49 5 1 1 32
0 50 5 1 1 34
0 51 5 1 1 36
0 52 5 1 1 38
0 53 5 1 1 40
0 54 5 1 1 42
0 55 5 1 1 44
0 56 5 1 1 46
0 57 5 1 1 48
0 58 5 1 1 97
0 59 5 1 1 127
0 60 5 1 1 157
0 61 5 1 1 187
0 62 5 1 1 217
0 63 5 1 1 247
0 64 5 1 1 277
0 65 5 1 1 308
0 66 5 1 1 312
0 67 5 2 1 314
0 68 5 2 1 316
0 69 5 2 1 318
0 70 5 2 1 320
0 71 5 2 1 322
0 72 5 2 1 324
0 73 5 2 1 326
0 74 5 2 1 328
0 75 5 2 1 330
0 76 5 2 1 332
0 77 5 2 1 334
0 78 5 2 1 336
0 79 5 2 1 338
0 80 5 1 1 340
0 81 7 2 2 33 311
0 82 5 3 1 368
0 83 7 1 2 49 65
0 84 5 1 1 83
3 683 7 0 2 370 84
0 86 7 1 2 35 313
0 87 5 2 1 86
0 88 7 1 2 50 66
0 89 5 2 1 88
0 90 7 2 2 373 375
0 91 5 1 1 377
0 92 7 1 2 369 91
0 93 5 1 1 92
0 94 7 1 2 371 378
0 95 5 1 1 94
0 96 7 1 2 93 95
3 684 5 0 1 96
0 98 7 1 2 372 374
0 99 5 1 1 98
0 100 7 2 2 376 99
0 101 5 1 1 379
0 102 7 1 2 51 101
0 103 5 2 1 102
0 104 7 1 2 37 380
0 105 5 2 1 104
0 106 7 2 2 381 383
0 107 5 1 1 385
0 108 7 1 2 315 386
0 109 5 1 1 108
0 110 7 1 2 342 107
0 111 5 1 1 110
3 685 7 0 2 109 111
0 113 7 1 2 343 384
0 114 5 1 1 113
0 115 7 2 2 382 114
0 116 5 1 1 387
0 117 7 1 2 52 116
0 118 5 2 1 117
0 119 7 1 2 39 388
0 120 5 2 1 119
0 121 7 2 2 389 391
0 122 5 1 1 393
0 123 7 1 2 317 394
0 124 5 1 1 123
0 125 7 1 2 344 122
0 126 5 1 1 125
3 686 7 0 2 124 126
0 128 7 1 2 345 392
0 129 5 1 1 128
0 130 7 2 2 390 129
0 131 5 1 1 395
0 132 7 1 2 53 131
0 133 5 2 1 132
0 134 7 1 2 41 396
0 135 5 2 1 134
0 136 7 2 2 397 399
0 137 5 1 1 401
0 138 7 1 2 319 402
0 139 5 1 1 138
0 140 7 1 2 346 137
0 141 5 1 1 140
3 687 7 0 2 139 141
0 143 7 1 2 347 400
0 144 5 1 1 143
0 145 7 2 2 398 144
0 146 5 1 1 403
0 147 7 1 2 54 146
0 148 5 2 1 147
0 149 7 1 2 43 404
0 150 5 2 1 149
0 151 7 2 2 405 407
0 152 5 1 1 409
0 153 7 1 2 321 410
0 154 5 1 1 153
0 155 7 1 2 348 152
0 156 5 1 1 155
3 688 7 0 2 154 156
0 158 7 1 2 349 408
0 159 5 1 1 158
0 160 7 2 2 406 159
0 161 5 1 1 411
0 162 7 1 2 55 161
0 163 5 2 1 162
0 164 7 1 2 45 412
0 165 5 2 1 164
0 166 7 2 2 413 415
0 167 5 1 1 417
0 168 7 1 2 323 418
0 169 5 1 1 168
0 170 7 1 2 350 167
0 171 5 1 1 170
3 689 7 0 2 169 171
0 173 7 1 2 351 416
0 174 5 1 1 173
0 175 7 2 2 414 174
0 176 5 1 1 419
0 177 7 1 2 47 420
0 178 5 2 1 177
0 179 7 1 2 56 176
0 180 5 2 1 179
0 181 7 2 2 421 423
0 182 5 1 1 425
0 183 7 1 2 325 426
0 184 5 1 1 183
0 185 7 1 2 352 182
0 186 5 1 1 185
3 690 7 0 2 184 186
0 188 7 1 2 353 422
0 189 5 1 1 188
0 190 7 2 2 424 189
0 191 5 1 1 427
0 192 7 1 2 57 191
0 193 5 2 1 192
0 194 7 1 2 85 428
0 195 5 2 1 194
0 196 7 2 2 429 431
0 197 5 1 1 433
0 198 7 1 2 327 434
0 199 5 1 1 198
0 200 7 1 2 354 197
0 201 5 1 1 200
3 691 7 0 2 199 201
0 203 7 1 2 355 432
0 204 5 1 1 203
0 205 7 2 2 430 204
0 206 5 1 1 435
0 207 7 1 2 58 206
0 208 5 2 1 207
0 209 7 1 2 112 436
0 210 5 2 1 209
0 211 7 2 2 437 439
0 212 5 1 1 441
0 213 7 1 2 329 442
0 214 5 1 1 213
0 215 7 1 2 356 212
0 216 5 1 1 215
3 692 7 0 2 214 216
0 218 7 1 2 357 440
0 219 5 1 1 218
0 220 7 2 2 438 219
0 221 5 1 1 443
0 222 7 1 2 59 221
0 223 5 2 1 222
0 224 7 1 2 142 444
0 225 5 2 1 224
0 226 7 2 2 445 447
0 227 5 1 1 449
0 228 7 1 2 331 450
0 229 5 1 1 228
0 230 7 1 2 358 227
0 231 5 1 1 230
3 693 7 0 2 229 231
0 233 7 1 2 359 448
0 234 5 1 1 233
0 235 7 2 2 446 234
0 236 5 1 1 451
0 237 7 1 2 60 236
0 238 5 2 1 237
0 239 7 1 2 172 452
0 240 5 2 1 239
0 241 7 2 2 453 455
0 242 5 1 1 457
0 243 7 1 2 333 458
0 244 5 1 1 243
0 245 7 1 2 360 242
0 246 5 1 1 245
3 694 7 0 2 244 246
0 248 7 1 2 361 456
0 249 5 1 1 248
0 250 7 2 2 454 249
0 251 5 1 1 459
0 252 7 1 2 61 251
0 253 5 2 1 252
0 254 7 1 2 202 460
0 255 5 2 1 254
0 256 7 2 2 461 463
0 257 5 1 1 465
0 258 7 1 2 335 466
0 259 5 1 1 258
0 260 7 1 2 362 257
0 261 5 1 1 260
3 695 7 0 2 259 261
0 263 7 1 2 363 464
0 264 5 1 1 263
0 265 7 2 2 462 264
0 266 5 1 1 467
0 267 7 1 2 62 266
0 268 5 2 1 267
0 269 7 1 2 232 468
0 270 5 2 1 269
0 271 7 2 2 469 471
0 272 5 1 1 473
0 273 7 1 2 337 474
0 274 5 1 1 273
0 275 7 1 2 364 272
0 276 5 1 1 275
3 696 7 0 2 274 276
0 278 7 1 2 365 472
0 279 5 1 1 278
0 280 7 2 2 470 279
0 281 5 1 1 475
0 282 7 1 2 262 476
0 283 5 2 1 282
0 284 7 1 2 63 281
0 285 5 2 1 284
0 286 7 2 2 477 479
0 287 5 1 1 481
0 288 7 1 2 339 482
0 289 5 1 1 288
0 290 7 1 2 366 287
0 291 5 1 1 290
3 697 7 0 2 289 291
0 293 7 1 2 367 478
0 294 5 1 1 293
0 295 7 2 2 480 294
0 296 5 2 1 483
0 297 7 1 2 64 80
0 298 5 2 1 297
0 299 7 1 2 292 341
0 300 5 2 1 299
0 301 7 2 2 487 489
0 302 5 1 1 491
0 303 7 1 2 484 302
0 304 5 1 1 303
0 305 7 1 2 485 492
0 306 5 1 1 305
0 307 7 1 2 304 306
3 698 5 0 1 307
0 309 7 1 2 486 490
0 310 5 1 1 309
3 699 7 0 2 488 310
