1 0 0 8 0
2 32 1 0
2 1240 1 0
2 1241 1 0
2 1242 1 0
2 1243 1 0
2 1244 1 0
2 1245 1 0
2 1246 1 0
1 1 0 8 0
2 1247 1 1
2 1248 1 1
2 1249 1 1
2 1250 1 1
2 1251 1 1
2 1252 1 1
2 1253 1 1
2 1254 1 1
1 2 0 8 0
2 1255 1 2
2 1256 1 2
2 1257 1 2
2 1258 1 2
2 1259 1 2
2 1260 1 2
2 1261 1 2
2 1262 1 2
1 3 0 9 0
2 1263 1 3
2 1264 1 3
2 1265 1 3
2 1266 1 3
2 1267 1 3
2 1268 1 3
2 1269 1 3
2 1270 1 3
2 1271 1 3
1 4 0 8 0
2 1272 1 4
2 1273 1 4
2 1274 1 4
2 1275 1 4
2 1276 1 4
2 1277 1 4
2 1278 1 4
2 1279 1 4
1 5 0 9 0
2 1280 1 5
2 1281 1 5
2 1282 1 5
2 1283 1 5
2 1284 1 5
2 1285 1 5
2 1286 1 5
2 1287 1 5
2 1288 1 5
1 6 0 8 0
2 1289 1 6
2 1290 1 6
2 1291 1 6
2 1292 1 6
2 1293 1 6
2 1294 1 6
2 1295 1 6
2 1296 1 6
1 7 0 8 0
2 1297 1 7
2 1298 1 7
2 1299 1 7
2 1300 1 7
2 1301 1 7
2 1302 1 7
2 1303 1 7
2 1304 1 7
1 8 0 8 0
2 1305 1 8
2 1306 1 8
2 1307 1 8
2 1308 1 8
2 1309 1 8
2 1310 1 8
2 1311 1 8
2 1312 1 8
1 9 0 8 0
2 1313 1 9
2 1314 1 9
2 1315 1 9
2 1316 1 9
2 1317 1 9
2 1318 1 9
2 1319 1 9
2 1320 1 9
1 10 0 9 0
2 1321 1 10
2 1322 1 10
2 1323 1 10
2 1324 1 10
2 1325 1 10
2 1326 1 10
2 1327 1 10
2 1328 1 10
2 1329 1 10
1 11 0 8 0
2 1330 1 11
2 1331 1 11
2 1332 1 11
2 1333 1 11
2 1334 1 11
2 1335 1 11
2 1336 1 11
2 1337 1 11
1 12 0 8 0
2 1338 1 12
2 1339 1 12
2 1340 1 12
2 1341 1 12
2 1342 1 12
2 1343 1 12
2 1344 1 12
2 1345 1 12
1 13 0 8 0
2 1346 1 13
2 1347 1 13
2 1348 1 13
2 1349 1 13
2 1350 1 13
2 1351 1 13
2 1352 1 13
2 1353 1 13
1 14 0 8 0
2 1354 1 14
2 1355 1 14
2 1356 1 14
2 1357 1 14
2 1358 1 14
2 1359 1 14
2 1360 1 14
2 1361 1 14
1 15 0 8 0
2 1362 1 15
2 1363 1 15
2 1364 1 15
2 1365 1 15
2 1366 1 15
2 1367 1 15
2 1368 1 15
2 1369 1 15
1 16 0 2 0
2 1370 1 16
2 1371 1 16
1 17 0 2 0
2 1372 1 17
2 1373 1 17
1 18 0 2 0
2 1374 1 18
2 1375 1 18
1 19 0 2 0
2 1376 1 19
2 1377 1 19
1 20 0 2 0
2 1378 1 20
2 1379 1 20
1 21 0 2 0
2 1380 1 21
2 1381 1 21
1 22 0 2 0
2 1382 1 22
2 1383 1 22
1 23 0 2 0
2 1384 1 23
2 1385 1 23
1 24 0 2 0
2 1386 1 24
2 1387 1 24
1 25 0 2 0
2 1388 1 25
2 1389 1 25
1 26 0 2 0
2 1390 1 26
2 1391 1 26
1 27 0 2 0
2 1392 1 27
2 1393 1 27
1 28 0 2 0
2 1394 1 28
2 1395 1 28
1 29 0 2 0
2 1396 1 29
2 1397 1 29
1 30 0 2 0
2 1398 1 30
2 1399 1 30
1 31 0 2 0
2 1400 1 31
2 1401 1 31
2 1402 1 49
2 1403 1 49
2 1404 1 51
2 1405 1 51
2 1406 1 54
2 1407 1 54
2 1408 1 55
2 1409 1 55
2 1410 1 59
2 1411 1 59
2 1412 1 62
2 1413 1 62
2 1414 1 63
2 1415 1 63
2 1416 1 65
2 1417 1 65
2 1418 1 66
2 1419 1 66
2 1420 1 67
2 1421 1 67
2 1422 1 69
2 1423 1 69
2 1424 1 74
2 1425 1 74
2 1426 1 75
2 1427 1 75
2 1428 1 78
2 1429 1 78
2 1430 1 81
2 1431 1 81
2 1432 1 84
2 1433 1 84
2 1434 1 85
2 1435 1 85
2 1436 1 89
2 1437 1 89
2 1438 1 92
2 1439 1 92
2 1440 1 93
2 1441 1 93
2 1442 1 95
2 1443 1 95
2 1444 1 98
2 1445 1 98
2 1446 1 99
2 1447 1 99
2 1448 1 103
2 1449 1 103
2 1450 1 106
2 1451 1 106
2 1452 1 107
2 1453 1 107
2 1454 1 111
2 1455 1 111
2 1456 1 114
2 1457 1 114
2 1458 1 115
2 1459 1 115
2 1460 1 119
2 1461 1 119
2 1462 1 122
2 1463 1 122
2 1464 1 123
2 1465 1 123
2 1466 1 125
2 1467 1 125
2 1468 1 127
2 1469 1 127
2 1470 1 129
2 1471 1 129
2 1472 1 135
2 1473 1 135
2 1474 1 138
2 1475 1 138
2 1476 1 138
2 1477 1 141
2 1478 1 141
2 1479 1 144
2 1480 1 144
2 1481 1 145
2 1482 1 145
2 1483 1 149
2 1484 1 149
2 1485 1 152
2 1486 1 152
2 1487 1 153
2 1488 1 153
2 1489 1 157
2 1490 1 157
2 1491 1 160
2 1492 1 160
2 1493 1 161
2 1494 1 161
2 1495 1 165
2 1496 1 165
2 1497 1 168
2 1498 1 168
2 1499 1 169
2 1500 1 169
2 1501 1 171
2 1502 1 171
2 1503 1 173
2 1504 1 173
2 1505 1 174
2 1506 1 174
2 1507 1 175
2 1508 1 175
2 1509 1 176
2 1510 1 176
2 1511 1 177
2 1512 1 177
2 1513 1 180
2 1514 1 180
2 1515 1 181
2 1516 1 181
2 1517 1 185
2 1518 1 185
2 1519 1 188
2 1520 1 188
2 1521 1 189
2 1522 1 189
2 1523 1 193
2 1524 1 193
2 1525 1 196
2 1526 1 196
2 1527 1 197
2 1528 1 197
2 1529 1 201
2 1530 1 201
2 1531 1 204
2 1532 1 204
2 1533 1 205
2 1534 1 205
2 1535 1 209
2 1536 1 209
2 1537 1 212
2 1538 1 212
2 1539 1 213
2 1540 1 213
2 1541 1 217
2 1542 1 217
2 1543 1 220
2 1544 1 220
2 1545 1 221
2 1546 1 221
2 1547 1 225
2 1548 1 225
2 1549 1 228
2 1550 1 228
2 1551 1 229
2 1552 1 229
2 1553 1 233
2 1554 1 233
2 1555 1 236
2 1556 1 236
2 1557 1 237
2 1558 1 237
2 1559 1 239
2 1560 1 239
2 1561 1 242
2 1562 1 242
2 1563 1 245
2 1564 1 245
2 1565 1 249
2 1566 1 249
2 1567 1 252
2 1568 1 252
2 1569 1 253
2 1570 1 253
2 1571 1 257
2 1572 1 257
2 1573 1 260
2 1574 1 260
2 1575 1 261
2 1576 1 261
2 1577 1 263
2 1578 1 263
2 1579 1 266
2 1580 1 266
2 1581 1 267
2 1582 1 267
2 1583 1 269
2 1584 1 269
2 1585 1 275
2 1586 1 275
2 1587 1 278
2 1588 1 278
2 1589 1 281
2 1590 1 281
2 1591 1 284
2 1592 1 284
2 1593 1 287
2 1594 1 287
2 1595 1 291
2 1596 1 291
2 1597 1 294
2 1598 1 294
2 1599 1 295
2 1600 1 295
2 1601 1 299
2 1602 1 299
2 1603 1 302
2 1604 1 302
2 1605 1 303
2 1606 1 303
2 1607 1 305
2 1608 1 305
2 1609 1 308
2 1610 1 308
2 1611 1 311
2 1612 1 311
2 1613 1 315
2 1614 1 315
2 1615 1 318
2 1616 1 318
2 1617 1 319
2 1618 1 319
2 1619 1 323
2 1620 1 323
2 1621 1 326
2 1622 1 326
2 1623 1 327
2 1624 1 327
2 1625 1 331
2 1626 1 331
2 1627 1 334
2 1628 1 334
2 1629 1 335
2 1630 1 335
2 1631 1 339
2 1632 1 339
2 1633 1 342
2 1634 1 342
2 1635 1 343
2 1636 1 343
2 1637 1 347
2 1638 1 347
2 1639 1 350
2 1640 1 350
2 1641 1 351
2 1642 1 351
2 1643 1 353
2 1644 1 353
2 1645 1 356
2 1646 1 356
2 1647 1 357
2 1648 1 357
2 1649 1 361
2 1650 1 361
2 1651 1 364
2 1652 1 364
2 1653 1 365
2 1654 1 365
2 1655 1 367
2 1656 1 367
2 1657 1 369
2 1658 1 369
2 1659 1 372
2 1660 1 372
2 1661 1 373
2 1662 1 373
2 1663 1 375
2 1664 1 375
2 1665 1 377
2 1666 1 377
2 1667 1 379
2 1668 1 379
2 1669 1 381
2 1670 1 381
2 1671 1 382
2 1672 1 382
2 1673 1 383
2 1674 1 383
2 1675 1 384
2 1676 1 384
2 1677 1 385
2 1678 1 385
2 1679 1 386
2 1680 1 386
2 1681 1 387
2 1682 1 387
2 1683 1 388
2 1684 1 388
2 1685 1 390
2 1686 1 390
2 1687 1 393
2 1688 1 393
2 1689 1 397
2 1690 1 397
2 1691 1 400
2 1692 1 400
2 1693 1 403
2 1694 1 403
2 1695 1 407
2 1696 1 407
2 1697 1 410
2 1698 1 410
2 1699 1 411
2 1700 1 411
2 1701 1 414
2 1702 1 414
2 1703 1 415
2 1704 1 415
2 1705 1 419
2 1706 1 419
2 1707 1 422
2 1708 1 422
2 1709 1 423
2 1710 1 423
2 1711 1 427
2 1712 1 427
2 1713 1 430
2 1714 1 430
2 1715 1 431
2 1716 1 431
2 1717 1 435
2 1718 1 435
2 1719 1 438
2 1720 1 438
2 1721 1 441
2 1722 1 441
2 1723 1 445
2 1724 1 445
2 1725 1 448
2 1726 1 448
2 1727 1 451
2 1728 1 451
2 1729 1 455
2 1730 1 455
2 1731 1 458
2 1732 1 458
2 1733 1 459
2 1734 1 459
2 1735 1 461
2 1736 1 461
2 1737 1 464
2 1738 1 464
2 1739 1 465
2 1740 1 465
2 1741 1 469
2 1742 1 469
2 1743 1 472
2 1744 1 472
2 1745 1 473
2 1746 1 473
2 1747 1 477
2 1748 1 477
2 1749 1 480
2 1750 1 480
2 1751 1 481
2 1752 1 481
2 1753 1 485
2 1754 1 485
2 1755 1 488
2 1756 1 488
2 1757 1 489
2 1758 1 489
2 1759 1 493
2 1760 1 493
2 1761 1 496
2 1762 1 496
2 1763 1 497
2 1764 1 497
2 1765 1 501
2 1766 1 501
2 1767 1 504
2 1768 1 504
2 1769 1 505
2 1770 1 505
2 1771 1 507
2 1772 1 507
2 1773 1 513
2 1774 1 513
2 1775 1 516
2 1776 1 516
2 1777 1 519
2 1778 1 519
2 1779 1 522
2 1780 1 522
2 1781 1 525
2 1782 1 525
2 1783 1 529
2 1784 1 529
2 1785 1 532
2 1786 1 532
2 1787 1 533
2 1788 1 533
2 1789 1 537
2 1790 1 537
2 1791 1 540
2 1792 1 540
2 1793 1 541
2 1794 1 541
2 1795 1 545
2 1796 1 545
2 1797 1 548
2 1798 1 548
2 1799 1 549
2 1800 1 549
2 1801 1 553
2 1802 1 553
2 1803 1 556
2 1804 1 556
2 1805 1 557
2 1806 1 557
2 1807 1 561
2 1808 1 561
2 1809 1 564
2 1810 1 564
2 1811 1 565
2 1812 1 565
2 1813 1 569
2 1814 1 569
2 1815 1 572
2 1816 1 572
2 1817 1 573
2 1818 1 573
2 1819 1 577
2 1820 1 577
2 1821 1 580
2 1822 1 580
2 1823 1 581
2 1824 1 581
2 1825 1 583
2 1826 1 583
2 1827 1 586
2 1828 1 586
2 1829 1 589
2 1830 1 589
2 1831 1 593
2 1832 1 593
2 1833 1 596
2 1834 1 596
2 1835 1 597
2 1836 1 597
2 1837 1 601
2 1838 1 601
2 1839 1 604
2 1840 1 604
2 1841 1 605
2 1842 1 605
2 1843 1 609
2 1844 1 609
2 1845 1 612
2 1846 1 612
2 1847 1 613
2 1848 1 613
2 1849 1 617
2 1850 1 617
2 1851 1 620
2 1852 1 620
2 1853 1 621
2 1854 1 621
2 1855 1 627
2 1856 1 627
2 1857 1 630
2 1858 1 630
2 1859 1 631
2 1860 1 631
2 1861 1 635
2 1862 1 635
2 1863 1 638
2 1864 1 638
2 1865 1 639
2 1866 1 639
2 1867 1 643
2 1868 1 643
2 1869 1 646
2 1870 1 646
2 1871 1 647
2 1872 1 647
2 1873 1 651
2 1874 1 651
2 1875 1 654
2 1876 1 654
2 1877 1 655
2 1878 1 655
2 1879 1 657
2 1880 1 657
2 1881 1 660
2 1882 1 660
2 1883 1 663
2 1884 1 663
2 1885 1 667
2 1886 1 667
2 1887 1 670
2 1888 1 670
2 1889 1 671
2 1890 1 671
2 1891 1 675
2 1892 1 675
2 1893 1 678
2 1894 1 678
2 1895 1 681
2 1896 1 681
2 1897 1 683
2 1898 1 683
2 1899 1 685
2 1900 1 685
2 1901 1 687
2 1902 1 687
2 1903 1 689
2 1904 1 689
2 1905 1 691
2 1906 1 691
2 1907 1 693
2 1908 1 693
2 1909 1 694
2 1910 1 694
2 1911 1 695
2 1912 1 695
2 1913 1 695
2 1914 1 698
2 1915 1 698
2 1916 1 701
2 1917 1 701
2 1918 1 709
2 1919 1 709
2 1920 1 712
2 1921 1 712
2 1922 1 713
2 1923 1 713
2 1924 1 717
2 1925 1 717
2 1926 1 720
2 1927 1 720
2 1928 1 723
2 1929 1 723
2 1930 1 725
2 1931 1 725
2 1932 1 727
2 1933 1 727
2 1934 1 729
2 1935 1 729
2 1936 1 730
2 1937 1 730
2 1938 1 732
2 1939 1 732
2 1940 1 733
2 1941 1 733
2 1942 1 737
2 1943 1 737
2 1944 1 740
2 1945 1 740
2 1946 1 741
2 1947 1 741
2 1948 1 745
2 1949 1 745
2 1950 1 748
2 1951 1 748
2 1952 1 749
2 1953 1 749
2 1954 1 753
2 1955 1 753
2 1956 1 756
2 1957 1 756
2 1958 1 757
2 1959 1 757
2 1960 1 761
2 1961 1 761
2 1962 1 764
2 1963 1 764
2 1964 1 765
2 1965 1 765
2 1966 1 769
2 1967 1 769
2 1968 1 772
2 1969 1 772
2 1970 1 773
2 1971 1 773
2 1972 1 777
2 1973 1 777
2 1974 1 780
2 1975 1 780
2 1976 1 781
2 1977 1 781
2 1978 1 785
2 1979 1 785
2 1980 1 788
2 1981 1 788
2 1982 1 789
2 1983 1 789
2 1984 1 793
2 1985 1 793
2 1986 1 796
2 1987 1 796
2 1988 1 797
2 1989 1 797
2 1990 1 801
2 1991 1 801
2 1992 1 804
2 1993 1 804
2 1994 1 805
2 1995 1 805
2 1996 1 809
2 1997 1 809
2 1998 1 812
2 1999 1 812
2 2000 1 813
2 2001 1 813
2 2002 1 817
2 2003 1 817
2 2004 1 820
2 2005 1 820
2 2006 1 821
2 2007 1 821
2 2008 1 823
2 2009 1 823
2 2010 1 828
2 2011 1 828
2 2012 1 831
2 2013 1 831
2 2014 1 834
2 2015 1 834
2 2016 1 837
2 2017 1 837
2 2018 1 839
2 2019 1 839
2 2020 1 840
2 2021 1 840
2 2022 1 842
2 2023 1 842
2 2024 1 842
2 2025 1 842
2 2026 1 843
2 2027 1 843
2 2028 1 847
2 2029 1 847
2 2030 1 850
2 2031 1 850
2 2032 1 850
2 2033 1 850
2 2034 1 852
2 2035 1 852
2 2036 1 852
2 2037 1 855
2 2038 1 855
2 2039 1 858
2 2040 1 858
2 2041 1 858
2 2042 1 858
2 2043 1 860
2 2044 1 860
2 2045 1 860
2 2046 1 863
2 2047 1 863
2 2048 1 866
2 2049 1 866
2 2050 1 866
2 2051 1 868
2 2052 1 868
2 2053 1 868
2 2054 1 871
2 2055 1 871
2 2056 1 874
2 2057 1 874
2 2058 1 874
2 2059 1 876
2 2060 1 876
2 2061 1 876
2 2062 1 879
2 2063 1 879
2 2064 1 882
2 2065 1 882
2 2066 1 882
2 2067 1 884
2 2068 1 884
2 2069 1 884
2 2070 1 887
2 2071 1 887
2 2072 1 890
2 2073 1 890
2 2074 1 890
2 2075 1 890
2 2076 1 892
2 2077 1 892
2 2078 1 892
2 2079 1 895
2 2080 1 895
2 2081 1 898
2 2082 1 898
2 2083 1 898
2 2084 1 898
2 2085 1 900
2 2086 1 900
2 2087 1 900
2 2088 1 903
2 2089 1 903
2 2090 1 906
2 2091 1 906
2 2092 1 906
2 2093 1 906
2 2094 1 908
2 2095 1 908
2 2096 1 908
2 2097 1 911
2 2098 1 911
2 2099 1 914
2 2100 1 914
2 2101 1 914
2 2102 1 914
2 2103 1 916
2 2104 1 916
2 2105 1 916
2 2106 1 919
2 2107 1 919
2 2108 1 922
2 2109 1 922
2 2110 1 922
2 2111 1 924
2 2112 1 924
2 2113 1 924
2 2114 1 927
2 2115 1 927
2 2116 1 930
2 2117 1 930
2 2118 1 930
2 2119 1 932
2 2120 1 932
2 2121 1 932
2 2122 1 935
2 2123 1 935
2 2124 1 938
2 2125 1 938
2 2126 1 938
2 2127 1 940
2 2128 1 940
2 2129 1 940
2 2130 1 943
2 2131 1 943
2 2132 1 946
2 2133 1 946
2 2134 1 948
2 2135 1 948
2 2136 1 949
2 2137 1 949
2 2138 1 953
2 2139 1 953
2 2140 1 961
2 2141 1 961
2 2142 1 962
2 2143 1 962
2 2144 1 965
2 2145 1 965
2 2146 1 967
2 2147 1 967
2 2148 1 969
2 2149 1 969
2 2150 1 970
2 2151 1 970
2 2152 1 973
2 2153 1 973
2 2154 1 976
2 2155 1 976
2 2156 1 982
2 2157 1 982
2 2158 1 985
2 2159 1 985
2 2160 1 986
2 2161 1 986
2 2162 1 989
2 2163 1 989
2 2164 1 990
2 2165 1 990
2 2166 1 993
2 2167 1 993
2 2168 1 994
2 2169 1 994
2 2170 1 997
2 2171 1 997
2 2172 1 998
2 2173 1 998
2 2174 1 1001
2 2175 1 1001
2 2176 1 1005
2 2177 1 1005
2 2178 1 1007
2 2179 1 1007
2 2180 1 1008
2 2181 1 1008
2 2182 1 1009
2 2183 1 1009
2 2184 1 1019
2 2185 1 1019
2 2186 1 1020
2 2187 1 1020
2 2188 1 1023
2 2189 1 1023
2 2190 1 1032
2 2191 1 1032
2 2192 1 1036
2 2193 1 1036
2 2194 1 1037
2 2195 1 1037
2 2196 1 1040
2 2197 1 1040
2 2198 1 1042
2 2199 1 1042
2 2200 1 1044
2 2201 1 1044
2 2202 1 1045
2 2203 1 1045
2 2204 1 1048
2 2205 1 1048
2 2206 1 1049
2 2207 1 1049
2 2208 1 1052
2 2209 1 1052
2 2210 1 1053
2 2211 1 1053
2 2212 1 1056
2 2213 1 1056
2 2214 1 1057
2 2215 1 1057
2 2216 1 1060
2 2217 1 1060
2 2218 1 1061
2 2219 1 1061
2 2220 1 1064
2 2221 1 1064
2 2222 1 1067
2 2223 1 1067
2 2224 1 1071
2 2225 1 1071
2 2226 1 1079
2 2227 1 1079
2 2228 1 1081
2 2229 1 1081
2 2230 1 1081
2 2231 1 1089
2 2232 1 1089
2 2233 1 1089
2 2234 1 1090
2 2235 1 1090
2 2236 1 1095
2 2237 1 1095
2 2238 1 1095
2 2239 1 1096
2 2240 1 1096
2 2241 1 1101
2 2242 1 1101
2 2243 1 1101
2 2244 1 1102
2 2245 1 1102
2 2246 1 1107
2 2247 1 1107
2 2248 1 1107
2 2249 1 1113
2 2250 1 1113
2 2251 1 1114
2 2252 1 1114
2 2253 1 1117
2 2254 1 1117
2 2255 1 1118
2 2256 1 1118
2 2257 1 1123
2 2258 1 1123
2 2259 1 1124
2 2260 1 1124
2 2261 1 1127
2 2262 1 1127
2 2263 1 1128
2 2264 1 1128
2 2265 1 1135
2 2266 1 1135
2 2267 1 1158
2 2268 1 1158
2 2269 1 1159
2 2270 1 1159
0 33 5 1 1 1370
0 34 5 1 1 1372
0 35 5 1 1 1374
0 36 5 1 1 1376
0 37 5 1 1 1378
0 38 5 1 1 1380
0 39 5 1 1 1382
0 40 5 1 1 1384
0 41 5 1 1 1386
0 42 5 1 1 1388
0 43 5 1 1 1390
0 44 5 1 1 1392
0 45 5 1 1 1394
0 46 5 1 1 1396
0 47 5 1 1 1398
0 48 5 1 1 1400
0 49 7 2 2 1272 1362
0 50 5 1 1 1402
0 51 7 2 2 1297 1338
0 52 5 1 1 1404
0 53 7 1 2 1403 1405
0 54 5 2 1 53
0 55 7 2 2 1289 1346
0 56 5 1 1 1408
0 57 7 1 2 50 52
0 58 5 1 1 57
0 59 7 2 2 1406 58
0 60 5 1 1 1410
0 61 7 1 2 1409 1411
0 62 5 2 1 61
0 63 7 2 2 1407 1412
0 64 5 1 1 1414
0 65 7 2 2 1290 1354
0 66 5 2 1 1416
0 67 7 2 2 1280 1363
0 68 5 1 1 1420
0 69 7 2 2 1298 1347
0 70 5 1 1 1422
0 71 7 1 2 68 70
0 72 5 1 1 71
0 73 7 1 2 1421 1423
0 74 5 2 1 73
0 75 7 2 2 72 1424
0 76 5 1 1 1426
0 77 7 1 2 1417 1427
0 78 5 2 1 77
0 79 7 1 2 1418 76
0 80 5 1 1 79
0 81 7 2 2 1428 80
0 82 5 1 1 1430
0 83 7 1 2 64 1431
0 84 5 2 1 83
0 85 7 2 2 1281 1355
0 86 5 1 1 1434
0 87 7 1 2 56 60
0 88 5 1 1 87
0 89 7 2 2 1413 88
0 90 5 1 1 1436
0 91 7 1 2 1435 1437
0 92 5 2 1 91
0 93 7 2 2 1263 1364
0 94 5 1 1 1440
0 95 7 2 2 1299 1330
0 96 5 1 1 1442
0 97 7 1 2 1441 1443
0 98 5 2 1 97
0 99 7 2 2 1291 1339
0 100 5 1 1 1446
0 101 7 1 2 94 96
0 102 5 1 1 101
0 103 7 2 2 1444 102
0 104 5 1 1 1448
0 105 7 1 2 1447 1449
0 106 5 2 1 105
0 107 7 2 2 1445 1450
0 108 5 1 1 1452
0 109 7 1 2 86 90
0 110 5 1 1 109
0 111 7 2 2 1438 110
0 112 5 1 1 1454
0 113 7 1 2 108 1455
0 114 5 2 1 113
0 115 7 2 2 1439 1456
0 116 5 1 1 1458
0 117 7 1 2 1415 82
0 118 5 1 1 117
0 119 7 2 2 1432 118
0 120 5 1 1 1460
0 121 7 1 2 116 1461
0 122 5 2 1 121
0 123 7 2 2 1433 1462
0 124 5 1 1 1464
0 125 7 2 2 1425 1429
0 126 5 1 1 1466
0 127 7 2 2 1292 1365
0 128 5 1 1 1468
0 129 7 2 2 1300 1356
0 130 5 1 1 1470
0 131 7 1 2 128 1471
0 132 5 1 1 131
0 133 7 1 2 1469 130
0 134 5 1 1 133
0 135 7 2 2 132 134
0 136 5 1 1 1472
0 137 7 1 2 126 136
0 138 5 3 1 137
0 139 7 1 2 1467 1473
0 140 5 1 1 139
0 141 7 2 2 1474 140
0 142 5 1 1 1477
0 143 7 1 2 124 1478
0 144 5 2 1 143
0 145 7 2 2 1273 1357
0 146 5 1 1 1481
0 147 7 1 2 100 104
0 148 5 1 1 147
0 149 7 2 2 1451 148
0 150 5 1 1 1483
0 151 7 1 2 1482 1484
0 152 5 2 1 151
0 153 7 2 2 1282 1348
0 154 5 1 1 1487
0 155 7 1 2 146 150
0 156 5 1 1 155
0 157 7 2 2 1485 156
0 158 5 1 1 1489
0 159 7 1 2 1488 1490
0 160 5 2 1 159
0 161 7 2 2 1486 1491
0 162 5 1 1 1493
0 163 7 1 2 1453 112
0 164 5 1 1 163
0 165 7 2 2 1457 164
0 166 5 1 1 1495
0 167 7 1 2 162 1496
0 168 5 2 1 167
0 169 7 2 2 1301 1305
0 170 5 1 1 1499
0 171 7 2 2 1293 1313
0 172 5 1 1 1501
0 173 7 2 2 1500 1502
0 174 5 2 1 1503
0 175 7 2 2 1321 1504
0 176 5 2 1 1507
0 177 7 2 2 1255 1366
0 178 5 1 1 1511
0 179 7 1 2 1508 1512
0 180 5 2 1 179
0 181 7 2 2 1302 1322
0 182 5 1 1 1515
0 183 7 1 2 1509 178
0 184 5 1 1 183
0 185 7 2 2 1513 184
0 186 5 1 1 1517
0 187 7 1 2 1516 1518
0 188 5 2 1 187
0 189 7 2 2 1514 1519
0 190 5 1 1 1521
0 191 7 1 2 154 158
0 192 5 1 1 191
0 193 7 2 2 1492 192
0 194 5 1 1 1523
0 195 7 1 2 190 1524
0 196 5 2 1 195
0 197 7 2 2 1283 1340
0 198 5 1 1 1527
0 199 7 1 2 182 186
0 200 5 1 1 199
0 201 7 2 2 1520 200
0 202 5 1 1 1529
0 203 7 1 2 1528 1530
0 204 5 2 1 203
0 205 7 2 2 1294 1331
0 206 5 1 1 1533
0 207 7 1 2 198 202
0 208 5 1 1 207
0 209 7 2 2 1531 208
0 210 5 1 1 1535
0 211 7 1 2 1534 1536
0 212 5 2 1 211
0 213 7 2 2 1532 1537
0 214 5 1 1 1539
0 215 7 1 2 1522 194
0 216 5 1 1 215
0 217 7 2 2 1525 216
0 218 5 1 1 1541
0 219 7 1 2 214 1542
0 220 5 2 1 219
0 221 7 2 2 1526 1543
0 222 5 1 1 1545
0 223 7 1 2 1494 166
0 224 5 1 1 223
0 225 7 2 2 1497 224
0 226 5 1 1 1547
0 227 7 1 2 222 1548
0 228 5 2 1 227
0 229 7 2 2 1498 1549
0 230 5 1 1 1551
0 231 7 1 2 1459 120
0 232 5 1 1 231
0 233 7 2 2 1463 232
0 234 5 1 1 1553
0 235 7 1 2 230 1554
0 236 5 2 1 235
0 237 7 2 2 1264 1358
0 238 5 1 1 1557
0 239 7 2 2 1274 1349
0 240 5 1 1 1559
0 241 7 1 2 1558 1560
0 242 5 2 1 241
0 243 7 1 2 206 210
0 244 5 1 1 243
0 245 7 2 2 1538 244
0 246 5 1 1 1563
0 247 7 1 2 238 240
0 248 5 1 1 247
0 249 7 2 2 1561 248
0 250 5 1 1 1565
0 251 7 1 2 1564 1566
0 252 5 2 1 251
0 253 7 2 2 1562 1567
0 254 5 1 1 1569
0 255 7 1 2 1540 218
0 256 5 1 1 255
0 257 7 2 2 1544 256
0 258 5 1 1 1571
0 259 7 1 2 254 1572
0 260 5 2 1 259
0 261 7 2 2 1284 1332
0 262 5 1 1 1575
0 263 7 2 2 1256 1359
0 264 5 1 1 1577
0 265 7 1 2 1576 1578
0 266 5 2 1 265
0 267 7 2 2 1247 1367
0 268 5 1 1 1581
0 269 7 2 2 1275 1341
0 270 5 1 1 1583
0 271 7 1 2 1295 1323
0 272 5 1 1 271
0 273 7 1 2 1505 272
0 274 5 1 1 273
0 275 7 2 2 1510 274
0 276 5 1 1 1585
0 277 7 1 2 1584 1586
0 278 5 2 1 277
0 279 7 1 2 270 276
0 280 5 1 1 279
0 281 7 2 2 1587 280
0 282 5 1 1 1589
0 283 7 1 2 1582 1590
0 284 5 2 1 283
0 285 7 1 2 268 282
0 286 5 1 1 285
0 287 7 2 2 1591 286
0 288 5 1 1 1593
0 289 7 1 2 262 264
0 290 5 1 1 289
0 291 7 2 2 1579 290
0 292 5 1 1 1595
0 293 7 1 2 1594 1596
0 294 5 2 1 293
0 295 7 2 2 1580 1597
0 296 5 1 1 1599
0 297 7 1 2 246 250
0 298 5 1 1 297
0 299 7 2 2 1568 298
0 300 5 1 1 1601
0 301 7 1 2 296 1602
0 302 5 2 1 301
0 303 7 2 2 1303 1314
0 304 5 1 1 1605
0 305 7 2 2 1265 1350
0 306 5 1 1 1607
0 307 7 1 2 1606 1608
0 308 5 2 1 307
0 309 7 1 2 288 292
0 310 5 1 1 309
0 311 7 2 2 1598 310
0 312 5 1 1 1611
0 313 7 1 2 304 306
0 314 5 1 1 313
0 315 7 2 2 1609 314
0 316 5 1 1 1613
0 317 7 1 2 1612 1614
0 318 5 2 1 317
0 319 7 2 2 1610 1615
0 320 5 1 1 1617
0 321 7 1 2 1600 300
0 322 5 1 1 321
0 323 7 2 2 1603 322
0 324 5 1 1 1619
0 325 7 1 2 320 1620
0 326 5 2 1 325
0 327 7 2 2 1604 1621
0 328 5 1 1 1623
0 329 7 1 2 1570 258
0 330 5 1 1 329
0 331 7 2 2 1573 330
0 332 5 1 1 1625
0 333 7 1 2 328 1626
0 334 5 2 1 333
0 335 7 2 2 1574 1627
0 336 5 1 1 1629
0 337 7 1 2 1546 226
0 338 5 1 1 337
0 339 7 2 2 1550 338
0 340 5 1 1 1631
0 341 7 1 2 336 1632
0 342 5 2 1 341
0 343 7 2 2 1588 1592
0 344 5 1 1 1635
0 345 7 1 2 1618 324
0 346 5 1 1 345
0 347 7 2 2 1622 346
0 348 5 1 1 1637
0 349 7 1 2 344 1638
0 350 5 2 1 349
0 351 7 2 2 1285 1324
0 352 5 1 1 1641
0 353 7 2 2 1276 1333
0 354 5 1 1 1643
0 355 7 1 2 1642 1644
0 356 5 2 1 355
0 357 7 2 2 1248 1360
0 358 5 1 1 1647
0 359 7 1 2 352 354
0 360 5 1 1 359
0 361 7 2 2 1645 360
0 362 5 1 1 1649
0 363 7 1 2 1648 1650
0 364 5 2 1 363
0 365 7 2 2 1646 1651
0 366 5 1 1 1653
0 367 7 2 2 1257 1351
0 368 5 1 1 1655
0 369 7 2 2 32 1368
0 370 5 1 1 1657
0 371 7 1 2 1656 1658
0 372 5 2 1 371
0 373 7 2 2 1266 1342
0 374 5 1 1 1661
0 375 7 2 2 1277 1315
0 376 5 1 1 1663
0 377 7 2 2 1240 1334
0 378 5 1 1 1665
0 379 7 2 2 1258 1316
0 380 5 1 1 1667
0 381 7 2 2 1666 1668
0 382 5 2 1 1669
0 383 7 2 2 1267 1670
0 384 5 2 1 1673
0 385 7 2 2 1664 1674
0 386 5 2 1 1677
0 387 7 2 2 1286 1678
0 388 5 2 1 1681
0 389 7 1 2 1662 1682
0 390 5 2 1 389
0 391 7 1 2 374 1683
0 392 5 1 1 391
0 393 7 2 2 1685 392
0 394 5 1 1 1687
0 395 7 1 2 170 172
0 396 5 1 1 395
0 397 7 2 2 1506 396
0 398 5 1 1 1689
0 399 7 1 2 1688 1690
0 400 5 2 1 399
0 401 7 1 2 394 398
0 402 5 1 1 401
0 403 7 2 2 1691 402
0 404 5 1 1 1693
0 405 7 1 2 368 370
0 406 5 1 1 405
0 407 7 2 2 1659 406
0 408 5 1 1 1695
0 409 7 1 2 1694 1696
0 410 5 2 1 409
0 411 7 2 2 1660 1697
0 412 5 1 1 1699
0 413 7 1 2 366 412
0 414 5 2 1 413
0 415 7 2 2 1686 1692
0 416 5 1 1 1703
0 417 7 1 2 1654 1700
0 418 5 1 1 417
0 419 7 2 2 1701 418
0 420 5 1 1 1705
0 421 7 1 2 416 1706
0 422 5 2 1 421
0 423 7 2 2 1702 1707
0 424 5 1 1 1709
0 425 7 1 2 1636 348
0 426 5 1 1 425
0 427 7 2 2 1639 426
0 428 5 1 1 1711
0 429 7 1 2 424 1712
0 430 5 2 1 429
0 431 7 2 2 1640 1713
0 432 5 1 1 1715
0 433 7 1 2 1624 332
0 434 5 1 1 433
0 435 7 2 2 1628 434
0 436 5 1 1 1717
0 437 7 1 2 432 1718
0 438 5 2 1 437
0 439 7 1 2 312 316
0 440 5 1 1 439
0 441 7 2 2 1616 440
0 442 5 1 1 1721
0 443 7 1 2 1704 420
0 444 5 1 1 443
0 445 7 2 2 1708 444
0 446 5 1 1 1723
0 447 7 1 2 1722 1724
0 448 5 2 1 447
0 449 7 1 2 358 362
0 450 5 1 1 449
0 451 7 2 2 1652 450
0 452 5 1 1 1727
0 453 7 1 2 404 408
0 454 5 1 1 453
0 455 7 2 2 1698 454
0 456 5 1 1 1729
0 457 7 1 2 1728 1730
0 458 5 2 1 457
0 459 7 2 2 1268 1335
0 460 5 1 1 1733
0 461 7 2 2 1259 1343
0 462 5 1 1 1735
0 463 7 1 2 1734 1736
0 464 5 2 1 463
0 465 7 2 2 1249 1352
0 466 5 1 1 1739
0 467 7 1 2 460 462
0 468 5 1 1 467
0 469 7 2 2 1737 468
0 470 5 1 1 1741
0 471 7 1 2 1740 1742
0 472 5 2 1 471
0 473 7 2 2 1738 1743
0 474 5 1 1 1745
0 475 7 1 2 452 456
0 476 5 1 1 475
0 477 7 2 2 1731 476
0 478 5 1 1 1747
0 479 7 1 2 474 1748
0 480 5 2 1 479
0 481 7 2 2 1732 1749
0 482 5 1 1 1751
0 483 7 1 2 442 446
0 484 5 1 1 483
0 485 7 2 2 1725 484
0 486 5 1 1 1753
0 487 7 1 2 482 1754
0 488 5 2 1 487
0 489 7 2 2 1726 1755
0 490 5 1 1 1757
0 491 7 1 2 1710 428
0 492 5 1 1 491
0 493 7 2 2 1714 492
0 494 5 1 1 1759
0 495 7 1 2 490 1760
0 496 5 2 1 495
0 497 7 2 2 1241 1361
0 498 5 1 1 1763
0 499 7 1 2 466 470
0 500 5 1 1 499
0 501 7 2 2 1744 500
0 502 5 1 1 1765
0 503 7 1 2 1764 1766
0 504 5 2 1 503
0 505 7 2 2 1296 1306
0 506 5 1 1 1769
0 507 7 2 2 1278 1325
0 508 5 1 1 1771
0 509 7 1 2 1287 1317
0 510 5 1 1 509
0 511 7 1 2 1679 510
0 512 5 1 1 511
0 513 7 2 2 1684 512
0 514 5 1 1 1773
0 515 7 1 2 1772 1774
0 516 5 2 1 515
0 517 7 1 2 508 514
0 518 5 1 1 517
0 519 7 2 2 1775 518
0 520 5 1 1 1777
0 521 7 1 2 1770 1778
0 522 5 2 1 521
0 523 7 1 2 506 520
0 524 5 1 1 523
0 525 7 2 2 1779 524
0 526 5 1 1 1781
0 527 7 1 2 498 502
0 528 5 1 1 527
0 529 7 2 2 1767 528
0 530 5 1 1 1783
0 531 7 1 2 1782 1784
0 532 5 2 1 531
0 533 7 2 2 1768 1785
0 534 5 1 1 1787
0 535 7 1 2 1746 478
0 536 5 1 1 535
0 537 7 2 2 1750 536
0 538 5 1 1 1789
0 539 7 1 2 534 1790
0 540 5 2 1 539
0 541 7 2 2 1776 1780
0 542 5 1 1 1793
0 543 7 1 2 1788 538
0 544 5 1 1 543
0 545 7 2 2 1791 544
0 546 5 1 1 1795
0 547 7 1 2 542 1796
0 548 5 2 1 547
0 549 7 2 2 1792 1797
0 550 5 1 1 1799
0 551 7 1 2 1752 486
0 552 5 1 1 551
0 553 7 2 2 1756 552
0 554 5 1 1 1801
0 555 7 1 2 550 1802
0 556 5 2 1 555
0 557 7 2 2 1269 1326
0 558 5 1 1 1805
0 559 7 1 2 376 1675
0 560 5 1 1 559
0 561 7 2 2 1680 560
0 562 5 1 1 1807
0 563 7 1 2 1806 1808
0 564 5 2 1 563
0 565 7 2 2 1288 1307
0 566 5 1 1 1811
0 567 7 1 2 558 562
0 568 5 1 1 567
0 569 7 2 2 1809 568
0 570 5 1 1 1813
0 571 7 1 2 1812 1814
0 572 5 2 1 571
0 573 7 2 2 1810 1815
0 574 5 1 1 1817
0 575 7 1 2 526 530
0 576 5 1 1 575
0 577 7 2 2 1786 576
0 578 5 1 1 1819
0 579 7 1 2 574 1820
0 580 5 2 1 579
0 581 7 2 2 1260 1336
0 582 5 1 1 1823
0 583 7 2 2 1242 1353
0 584 5 1 1 1825
0 585 7 1 2 1824 1826
0 586 5 2 1 585
0 587 7 1 2 566 570
0 588 5 1 1 587
0 589 7 2 2 1816 588
0 590 5 1 1 1829
0 591 7 1 2 582 584
0 592 5 1 1 591
0 593 7 2 2 1827 592
0 594 5 1 1 1831
0 595 7 1 2 1830 1832
0 596 5 2 1 595
0 597 7 2 2 1828 1833
0 598 5 1 1 1835
0 599 7 1 2 1818 578
0 600 5 1 1 599
0 601 7 2 2 1821 600
0 602 5 1 1 1837
0 603 7 1 2 598 1838
0 604 5 2 1 603
0 605 7 2 2 1822 1839
0 606 5 1 1 1841
0 607 7 1 2 1794 546
0 608 5 1 1 607
0 609 7 2 2 1798 608
0 610 5 1 1 1843
0 611 7 1 2 606 1844
0 612 5 2 1 611
0 613 7 2 2 1250 1344
0 614 5 1 1 1847
0 615 7 1 2 590 594
0 616 5 1 1 615
0 617 7 2 2 1834 616
0 618 5 1 1 1849
0 619 7 1 2 1848 1850
0 620 5 2 1 619
0 621 7 2 2 1261 1327
0 622 5 1 1 1853
0 623 7 1 2 1270 1318
0 624 5 1 1 623
0 625 7 1 2 1671 624
0 626 5 1 1 625
0 627 7 2 2 1676 626
0 628 5 1 1 1855
0 629 7 1 2 1854 1856
0 630 5 2 1 629
0 631 7 2 2 1279 1308
0 632 5 1 1 1859
0 633 7 1 2 622 628
0 634 5 1 1 633
0 635 7 2 2 1857 634
0 636 5 1 1 1861
0 637 7 1 2 1860 1862
0 638 5 2 1 637
0 639 7 2 2 1858 1863
0 640 5 1 1 1865
0 641 7 1 2 614 618
0 642 5 1 1 641
0 643 7 2 2 1851 642
0 644 5 1 1 1867
0 645 7 1 2 640 1868
0 646 5 2 1 645
0 647 7 2 2 1852 1869
0 648 5 1 1 1871
0 649 7 1 2 1836 602
0 650 5 1 1 649
0 651 7 2 2 1840 650
0 652 5 1 1 1873
0 653 7 1 2 648 1874
0 654 5 2 1 653
0 655 7 2 2 1243 1345
0 656 5 1 1 1877
0 657 7 2 2 1251 1337
0 658 5 1 1 1879
0 659 7 1 2 1878 1880
0 660 5 2 1 659
0 661 7 1 2 632 636
0 662 5 1 1 661
0 663 7 2 2 1864 662
0 664 5 1 1 1883
0 665 7 1 2 656 658
0 666 5 1 1 665
0 667 7 2 2 1881 666
0 668 5 1 1 1885
0 669 7 1 2 1884 1886
0 670 5 2 1 669
0 671 7 2 2 1882 1887
0 672 5 1 1 1889
0 673 7 1 2 1866 644
0 674 5 1 1 673
0 675 7 2 2 1870 674
0 676 5 1 1 1891
0 677 7 1 2 672 1892
0 678 5 2 1 677
0 679 7 1 2 664 668
0 680 5 1 1 679
0 681 7 2 2 1888 680
0 682 5 1 1 1895
0 683 7 2 2 1252 1328
0 684 5 1 1 1897
0 685 7 2 2 1271 1309
0 686 5 1 1 1899
0 687 7 2 2 1898 1900
0 688 5 1 1 1901
0 689 7 2 2 1253 1319
0 690 5 1 1 1903
0 691 7 2 2 1244 1329
0 692 5 1 1 1905
0 693 7 2 2 1904 1906
0 694 5 2 1 1907
0 695 7 3 2 688 1909
0 696 5 1 1 1911
0 697 7 1 2 1896 696
0 698 5 2 1 697
0 699 7 1 2 378 380
0 700 5 1 1 699
0 701 7 2 2 1672 700
0 702 5 1 1 1916
0 703 7 1 2 684 686
0 704 5 1 1 703
0 705 7 1 2 1912 704
0 706 5 1 1 705
0 707 7 1 2 1902 1908
0 708 5 1 1 707
0 709 7 2 2 706 708
0 710 5 1 1 1918
0 711 7 1 2 1917 710
0 712 5 2 1 711
0 713 7 2 2 1262 1310
0 714 5 1 1 1922
0 715 7 1 2 690 692
0 716 5 1 1 715
0 717 7 2 2 1910 716
0 718 5 1 1 1924
0 719 7 1 2 1923 1925
0 720 5 2 1 719
0 721 7 1 2 714 718
0 722 5 1 1 721
0 723 7 2 2 1926 722
0 724 5 1 1 1928
0 725 7 2 2 1245 1320
0 726 5 1 1 1930
0 727 7 2 2 1254 1311
0 728 5 1 1 1932
0 729 7 2 2 1931 1933
0 730 5 2 1 1934
0 731 7 1 2 1929 1935
0 732 5 2 1 731
0 733 7 2 2 1927 1938
0 734 5 1 1 1940
0 735 7 1 2 702 1919
0 736 5 1 1 735
0 737 7 2 2 1920 736
0 738 5 1 1 1942
0 739 7 1 2 734 1943
0 740 5 2 1 739
0 741 7 2 2 1921 1944
0 742 5 1 1 1946
0 743 7 1 2 682 1913
0 744 5 1 1 743
0 745 7 2 2 1914 744
0 746 5 1 1 1948
0 747 7 1 2 742 1949
0 748 5 2 1 747
0 749 7 2 2 1915 1950
0 750 5 1 1 1952
0 751 7 1 2 1890 676
0 752 5 1 1 751
0 753 7 2 2 1893 752
0 754 5 1 1 1954
0 755 7 1 2 750 1955
0 756 5 2 1 755
0 757 7 2 2 1894 1956
0 758 5 1 1 1958
0 759 7 1 2 1872 652
0 760 5 1 1 759
0 761 7 2 2 1875 760
0 762 5 1 1 1960
0 763 7 1 2 758 1961
0 764 5 2 1 763
0 765 7 2 2 1876 1962
0 766 5 1 1 1964
0 767 7 1 2 1842 610
0 768 5 1 1 767
0 769 7 2 2 1845 768
0 770 5 1 1 1966
0 771 7 1 2 766 1967
0 772 5 2 1 771
0 773 7 2 2 1846 1968
0 774 5 1 1 1970
0 775 7 1 2 1800 554
0 776 5 1 1 775
0 777 7 2 2 1803 776
0 778 5 1 1 1972
0 779 7 1 2 774 1973
0 780 5 2 1 779
0 781 7 2 2 1804 1974
0 782 5 1 1 1976
0 783 7 1 2 1758 494
0 784 5 1 1 783
0 785 7 2 2 1761 784
0 786 5 1 1 1978
0 787 7 1 2 782 1979
0 788 5 2 1 787
0 789 7 2 2 1762 1980
0 790 5 1 1 1982
0 791 7 1 2 1716 436
0 792 5 1 1 791
0 793 7 2 2 1719 792
0 794 5 1 1 1984
0 795 7 1 2 790 1985
0 796 5 2 1 795
0 797 7 2 2 1720 1986
0 798 5 1 1 1988
0 799 7 1 2 1630 340
0 800 5 1 1 799
0 801 7 2 2 1633 800
0 802 5 1 1 1990
0 803 7 1 2 798 1991
0 804 5 2 1 803
0 805 7 2 2 1634 1992
0 806 5 1 1 1994
0 807 7 1 2 1552 234
0 808 5 1 1 807
0 809 7 2 2 1555 808
0 810 5 1 1 1996
0 811 7 1 2 806 1997
0 812 5 2 1 811
0 813 7 2 2 1556 1998
0 814 5 1 1 2000
0 815 7 1 2 1465 142
0 816 5 1 1 815
0 817 7 2 2 1479 816
0 818 5 1 1 2002
0 819 7 1 2 814 2003
0 820 5 2 1 819
0 821 7 2 2 1480 2004
0 822 5 1 1 2006
0 823 7 2 2 1304 1369
0 824 5 1 1 2008
0 825 7 1 2 1419 1475
0 826 5 1 1 825
0 827 7 1 2 2009 826
0 828 5 2 1 827
0 829 7 1 2 1476 824
0 830 5 1 1 829
0 831 7 2 2 2010 830
0 832 5 1 1 2012
0 833 7 1 2 822 2013
0 834 5 2 1 833
0 835 7 1 2 2007 832
0 836 5 1 1 835
0 837 7 2 2 2014 836
0 838 5 1 1 2016
0 839 7 2 2 47 2017
0 840 5 2 1 2018
0 841 7 1 2 1399 838
0 842 5 4 1 841
0 843 7 2 2 2020 2022
0 844 5 1 1 2026
0 845 7 1 2 2001 818
0 846 5 1 1 845
0 847 7 2 2 2005 846
0 848 5 1 1 2028
0 849 7 1 2 1397 848
0 850 5 4 1 849
0 851 7 1 2 46 2029
0 852 5 3 1 851
0 853 7 1 2 1995 810
0 854 5 1 1 853
0 855 7 2 2 1999 854
0 856 5 1 1 2037
0 857 7 1 2 1395 856
0 858 5 4 1 857
0 859 7 1 2 45 2038
0 860 5 3 1 859
0 861 7 1 2 1989 802
0 862 5 1 1 861
0 863 7 2 2 1993 862
0 864 5 1 1 2046
0 865 7 1 2 1393 864
0 866 5 3 1 865
0 867 7 1 2 44 2047
0 868 5 3 1 867
0 869 7 1 2 1983 794
0 870 5 1 1 869
0 871 7 2 2 1987 870
0 872 5 1 1 2054
0 873 7 1 2 1391 872
0 874 5 3 1 873
0 875 7 1 2 43 2055
0 876 5 3 1 875
0 877 7 1 2 1977 786
0 878 5 1 1 877
0 879 7 2 2 1981 878
0 880 5 1 1 2062
0 881 7 1 2 1389 880
0 882 5 3 1 881
0 883 7 1 2 42 2063
0 884 5 3 1 883
0 885 7 1 2 1971 778
0 886 5 1 1 885
0 887 7 2 2 1975 886
0 888 5 1 1 2070
0 889 7 1 2 1387 888
0 890 5 4 1 889
0 891 7 1 2 41 2071
0 892 5 3 1 891
0 893 7 1 2 1965 770
0 894 5 1 1 893
0 895 7 2 2 1969 894
0 896 5 1 1 2079
0 897 7 1 2 1385 896
0 898 5 4 1 897
0 899 7 1 2 40 2080
0 900 5 3 1 899
0 901 7 1 2 1959 762
0 902 5 1 1 901
0 903 7 2 2 1963 902
0 904 5 1 1 2088
0 905 7 1 2 1383 904
0 906 5 4 1 905
0 907 7 1 2 39 2089
0 908 5 3 1 907
0 909 7 1 2 1953 754
0 910 5 1 1 909
0 911 7 2 2 1957 910
0 912 5 1 1 2097
0 913 7 1 2 1381 912
0 914 5 4 1 913
0 915 7 1 2 38 2098
0 916 5 3 1 915
0 917 7 1 2 1947 746
0 918 5 1 1 917
0 919 7 2 2 1951 918
0 920 5 1 1 2106
0 921 7 1 2 1379 920
0 922 5 3 1 921
0 923 7 1 2 37 2107
0 924 5 3 1 923
0 925 7 1 2 1941 738
0 926 5 1 1 925
0 927 7 2 2 1945 926
0 928 5 1 1 2114
0 929 7 1 2 1377 928
0 930 5 3 1 929
0 931 7 1 2 36 2115
0 932 5 3 1 931
0 933 7 1 2 724 1936
0 934 5 1 1 933
0 935 7 2 2 1939 934
0 936 5 1 1 2122
0 937 7 1 2 35 2123
0 938 5 3 1 937
0 939 7 1 2 1375 936
0 940 5 3 1 939
0 941 7 1 2 726 728
0 942 5 1 1 941
0 943 7 2 2 1937 942
0 944 5 1 1 2130
0 945 7 1 2 1373 944
0 946 5 2 1 945
0 947 7 1 2 34 2131
0 948 5 2 1 947
0 949 7 2 2 1246 1312
0 950 5 1 1 2136
0 951 7 1 2 33 2137
0 952 5 1 1 951
0 953 7 2 2 2134 952
0 954 5 1 1 2138
0 955 7 1 2 2132 954
0 956 7 1 2 2127 955
0 957 5 1 1 956
0 958 7 1 2 2124 957
0 959 7 1 2 2119 958
0 960 5 1 1 959
0 961 7 2 2 2116 960
0 962 5 2 1 2140
0 963 7 1 2 2111 2142
0 964 5 1 1 963
0 965 7 2 2 2108 964
0 966 5 1 1 2144
0 967 7 2 2 2103 966
0 968 5 1 1 2146
0 969 7 2 2 2099 968
0 970 5 2 1 2148
0 971 7 1 2 2094 2150
0 972 5 1 1 971
0 973 7 2 2 2090 972
0 974 5 1 1 2152
0 975 7 1 2 2085 974
0 976 5 2 1 975
0 977 7 1 2 2081 2154
0 978 5 1 1 977
0 979 7 1 2 2076 978
0 980 5 1 1 979
0 981 7 1 2 2072 980
0 982 5 2 1 981
0 983 7 1 2 2067 2156
0 984 5 1 1 983
0 985 7 2 2 2064 984
0 986 5 2 1 2158
0 987 7 1 2 2059 2160
0 988 5 1 1 987
0 989 7 2 2 2056 988
0 990 5 2 1 2162
0 991 7 1 2 2051 2164
0 992 5 1 1 991
0 993 7 2 2 2048 992
0 994 5 2 1 2166
0 995 7 1 2 2043 2168
0 996 5 1 1 995
0 997 7 2 2 2039 996
0 998 5 2 1 2170
0 999 7 1 2 2034 2172
0 1000 5 1 1 999
0 1001 7 2 2 2030 1000
0 1002 5 1 1 2174
0 1003 7 1 2 844 1002
0 1004 5 1 1 1003
0 1005 7 2 2 2011 2015
0 1006 5 1 1 2176
0 1007 7 2 2 1401 2177
0 1008 5 2 1 2178
0 1009 7 2 2 2023 2175
0 1010 5 1 1 2182
0 1011 7 1 2 2180 1010
0 1012 7 1 2 1004 1011
0 1013 5 1 1 1012
0 1014 7 1 2 2019 2179
0 1015 7 1 2 2183 1014
0 1016 5 1 1 1015
0 1017 7 1 2 1013 1016
0 1018 5 1 1 1017
0 1019 7 2 2 48 1006
0 1020 5 2 1 2184
0 1021 7 1 2 1371 950
0 1022 5 1 1 1021
0 1023 7 2 2 2133 1022
0 1024 5 1 1 2188
0 1025 7 1 2 2135 1024
0 1026 7 1 2 2125 1025
0 1027 5 1 1 1026
0 1028 7 1 2 2128 1027
0 1029 5 1 1 1028
0 1030 7 1 2 2120 1029
0 1031 5 1 1 1030
0 1032 7 2 2 2117 1031
0 1033 5 1 1 2190
0 1034 7 1 2 2112 1033
0 1035 5 1 1 1034
0 1036 7 2 2 2109 1035
0 1037 5 2 1 2192
0 1038 7 1 2 2104 2194
0 1039 5 1 1 1038
0 1040 7 2 2 2100 1039
0 1041 5 1 1 2196
0 1042 7 2 2 2095 1041
0 1043 5 1 1 2198
0 1044 7 2 2 2091 1043
0 1045 5 2 1 2200
0 1046 7 1 2 2086 2202
0 1047 5 1 1 1046
0 1048 7 2 2 2082 1047
0 1049 5 2 1 2204
0 1050 7 1 2 2077 2206
0 1051 5 1 1 1050
0 1052 7 2 2 2073 1051
0 1053 5 2 1 2208
0 1054 7 1 2 2068 2210
0 1055 5 1 1 1054
0 1056 7 2 2 2065 1055
0 1057 5 2 1 2212
0 1058 7 1 2 2060 2214
0 1059 5 1 1 1058
0 1060 7 2 2 2057 1059
0 1061 5 2 1 2216
0 1062 7 1 2 2052 2218
0 1063 5 1 1 1062
0 1064 7 2 2 2049 1063
0 1065 5 1 1 2220
0 1066 7 1 2 2044 1065
0 1067 5 2 1 1066
0 1068 7 1 2 2040 2222
0 1069 5 1 1 1068
0 1070 7 1 2 2035 1069
0 1071 5 2 1 1070
0 1072 7 1 2 2031 2224
0 1073 5 1 1 1072
0 1074 7 1 2 2021 1073
0 1075 5 1 1 1074
0 1076 7 1 2 2024 2181
0 1077 7 1 2 1075 1076
0 1078 5 1 1 1077
0 1079 7 2 2 2186 1078
0 1080 5 1 1 2226
0 1081 7 3 2 2032 2036
0 1082 5 1 1 2228
0 1083 7 1 2 2171 1082
0 1084 5 1 1 1083
0 1085 7 1 2 2173 2229
0 1086 5 1 1 1085
0 1087 7 1 2 1084 1086
0 1088 5 1 1 1087
0 1089 7 3 2 2050 2053
0 1090 5 2 1 2231
0 1091 7 1 2 2163 2234
0 1092 5 1 1 1091
0 1093 7 1 2 2165 2232
0 1094 5 1 1 1093
0 1095 7 3 2 2058 2061
0 1096 5 2 1 2236
0 1097 7 1 2 2159 2239
0 1098 5 1 1 1097
0 1099 7 1 2 2161 2237
0 1100 5 1 1 1099
0 1101 7 3 2 2066 2069
0 1102 5 2 1 2241
0 1103 7 1 2 2074 2244
0 1104 5 1 1 1103
0 1105 7 1 2 2157 2242
0 1106 5 1 1 1105
0 1107 7 3 2 2075 2078
0 1108 5 1 1 2246
0 1109 7 1 2 2155 2247
0 1110 5 1 1 1109
0 1111 7 1 2 2083 1110
0 1112 5 1 1 1111
0 1113 7 2 2 2084 2087
0 1114 5 2 1 2249
0 1115 7 1 2 2153 2251
0 1116 5 1 1 1115
0 1117 7 2 2 2092 2096
0 1118 5 2 1 2253
0 1119 7 1 2 2149 2254
0 1120 5 1 1 1119
0 1121 7 1 2 2101 2147
0 1122 5 1 1 1121
0 1123 7 2 2 2102 2105
0 1124 5 2 1 2257
0 1125 7 1 2 2145 2259
0 1126 5 1 1 1125
0 1127 7 2 2 2110 2113
0 1128 5 2 1 2261
0 1129 7 1 2 2141 2262
0 1130 5 1 1 1129
0 1131 7 1 2 2139 2189
0 1132 7 1 2 2126 1131
0 1133 7 1 2 2129 1132
0 1134 7 1 2 2118 1133
0 1135 7 2 2 2121 1134
0 1136 7 1 2 2143 2263
0 1137 5 1 1 1136
0 1138 7 1 2 2265 1137
0 1139 7 1 2 1130 1138
0 1140 5 1 1 1139
0 1141 7 1 2 1126 1140
0 1142 7 1 2 1122 1141
0 1143 5 1 1 1142
0 1144 7 1 2 2151 2255
0 1145 5 1 1 1144
0 1146 7 1 2 1143 1145
0 1147 7 1 2 1120 1146
0 1148 5 1 1 1147
0 1149 7 1 2 1116 1148
0 1150 7 1 2 1112 1149
0 1151 7 1 2 1106 1150
0 1152 7 1 2 1104 1151
0 1153 7 1 2 1100 1152
0 1154 7 1 2 1098 1153
0 1155 7 1 2 1094 1154
0 1156 7 1 2 1092 1155
0 1157 5 1 1 1156
0 1158 7 2 2 2041 2045
0 1159 5 2 1 2267
0 1160 7 1 2 2167 2269
0 1161 5 1 1 1160
0 1162 7 1 2 2169 2268
0 1163 5 1 1 1162
0 1164 7 1 2 1161 1163
0 1165 5 1 1 1164
0 1166 7 1 2 1157 1165
0 1167 7 1 2 2187 1166
0 1168 7 1 2 1088 1167
0 1169 7 1 2 2227 1168
0 1170 7 1 2 1018 1169
0 1171 5 1 1 1170
0 1172 7 1 2 2027 2225
0 1173 5 1 1 1172
0 1174 7 1 2 2033 1173
0 1175 5 1 1 1174
0 1176 7 1 2 2223 2230
0 1177 5 1 1 1176
0 1178 7 1 2 2042 1177
0 1179 5 1 1 1178
0 1180 7 1 2 2025 2185
0 1181 5 1 1 1180
0 1182 7 1 2 2221 2270
0 1183 5 1 1 1182
0 1184 7 1 2 2217 2233
0 1185 5 1 1 1184
0 1186 7 1 2 2219 2235
0 1187 5 1 1 1186
0 1188 7 1 2 2213 2238
0 1189 5 1 1 1188
0 1190 7 1 2 2215 2240
0 1191 5 1 1 1190
0 1192 7 1 2 2209 2243
0 1193 5 1 1 1192
0 1194 7 1 2 2211 2245
0 1195 5 1 1 1194
0 1196 7 1 2 2205 2248
0 1197 5 1 1 1196
0 1198 7 1 2 2207 1108
0 1199 5 1 1 1198
0 1200 7 1 2 2201 2250
0 1201 5 1 1 1200
0 1202 7 1 2 2093 2199
0 1203 5 1 1 1202
0 1204 7 1 2 2197 2256
0 1205 5 1 1 1204
0 1206 7 1 2 2193 2258
0 1207 5 1 1 1206
0 1208 7 1 2 2191 2264
0 1209 5 1 1 1208
0 1210 7 1 2 2266 1209
0 1211 5 1 1 1210
0 1212 7 1 2 2195 2260
0 1213 5 1 1 1212
0 1214 7 1 2 1211 1213
0 1215 7 1 2 1207 1214
0 1216 5 1 1 1215
0 1217 7 1 2 1205 1216
0 1218 7 1 2 1203 1217
0 1219 5 1 1 1218
0 1220 7 1 2 2203 2252
0 1221 5 1 1 1220
0 1222 7 1 2 1219 1221
0 1223 7 1 2 1201 1222
0 1224 7 1 2 1199 1223
0 1225 7 1 2 1197 1224
0 1226 7 1 2 1195 1225
0 1227 7 1 2 1193 1226
0 1228 7 1 2 1191 1227
0 1229 7 1 2 1189 1228
0 1230 7 1 2 1187 1229
0 1231 7 1 2 1185 1230
0 1232 5 1 1 1231
0 1233 7 1 2 1183 1232
0 1234 7 1 2 1181 1233
0 1235 7 1 2 1179 1234
0 1236 7 1 2 1080 1235
0 1237 7 1 2 1175 1236
0 1238 5 1 1 1237
0 1239 7 1 2 1171 1238
3 4299 5 0 1 1239
