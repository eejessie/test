1 0 0 2 0
2 49 1 0
2 718 1 0
1 1 0 2 0
2 719 1 1
2 720 1 1
1 2 0 2 0
2 721 1 2
2 722 1 2
1 3 0 2 0
2 723 1 3
2 724 1 3
1 4 0 2 0
2 725 1 4
2 726 1 4
1 5 0 2 0
2 727 1 5
2 728 1 5
1 6 0 2 0
2 729 1 6
2 730 1 6
1 7 0 2 0
2 731 1 7
2 732 1 7
1 8 0 2 0
2 733 1 8
2 734 1 8
1 9 0 2 0
2 735 1 9
2 736 1 9
1 10 0 2 0
2 737 1 10
2 738 1 10
1 11 0 2 0
2 739 1 11
2 740 1 11
1 12 0 2 0
2 741 1 12
2 742 1 12
1 13 0 2 0
2 743 1 13
2 744 1 13
1 14 0 2 0
2 745 1 14
2 746 1 14
1 15 0 2 0
2 747 1 15
2 748 1 15
1 16 0 2 0
2 749 1 16
2 750 1 16
1 17 0 2 0
2 751 1 17
2 752 1 17
1 18 0 2 0
2 753 1 18
2 754 1 18
1 19 0 2 0
2 755 1 19
2 756 1 19
1 20 0 2 0
2 757 1 20
2 758 1 20
1 21 0 2 0
2 759 1 21
2 760 1 21
1 22 0 2 0
2 761 1 22
2 762 1 22
1 23 0 2 0
2 763 1 23
2 764 1 23
1 24 0 2 0
2 765 1 24
2 766 1 24
1 25 0 2 0
2 767 1 25
2 768 1 25
1 26 0 2 0
2 769 1 26
2 770 1 26
1 27 0 2 0
2 771 1 27
2 772 1 27
1 28 0 2 0
2 773 1 28
2 774 1 28
1 29 0 2 0
2 775 1 29
2 776 1 29
1 30 0 2 0
2 777 1 30
2 778 1 30
1 31 0 2 0
2 779 1 31
2 780 1 31
1 32 0 2 0
2 781 1 32
2 782 1 32
1 33 0 2 0
2 783 1 33
2 784 1 33
1 34 0 2 0
2 785 1 34
2 786 1 34
1 35 0 2 0
2 787 1 35
2 788 1 35
1 36 0 2 0
2 789 1 36
2 790 1 36
1 37 0 2 0
2 791 1 37
2 792 1 37
1 38 0 2 0
2 793 1 38
2 794 1 38
1 39 0 2 0
2 795 1 39
2 796 1 39
1 40 0 2 0
2 797 1 40
2 798 1 40
1 41 0 2 0
2 799 1 41
2 800 1 41
1 42 0 2 0
2 801 1 42
2 802 1 42
1 43 0 2 0
2 803 1 43
2 804 1 43
1 44 0 2 0
2 805 1 44
2 806 1 44
1 45 0 2 0
2 807 1 45
2 808 1 45
1 46 0 2 0
2 809 1 46
2 810 1 46
1 47 0 2 0
2 811 1 47
2 812 1 47
1 48 0 2 0
2 813 1 48
2 814 1 48
2 815 1 69
2 816 1 69
2 817 1 70
2 818 1 70
2 819 1 71
2 820 1 71
2 821 1 72
2 822 1 72
2 823 1 73
2 824 1 73
2 825 1 74
2 826 1 74
2 827 1 75
2 828 1 75
2 829 1 76
2 830 1 76
2 831 1 77
2 832 1 77
2 833 1 78
2 834 1 78
2 835 1 79
2 836 1 79
2 837 1 80
2 838 1 80
2 839 1 81
2 840 1 81
2 841 1 100
2 842 1 100
2 843 1 102
2 844 1 102
2 845 1 104
2 846 1 104
2 847 1 106
2 848 1 106
2 849 1 107
2 850 1 107
2 851 1 108
2 852 1 108
2 853 1 108
2 854 1 111
2 855 1 111
2 856 1 112
2 857 1 112
2 858 1 115
2 859 1 115
2 860 1 118
2 861 1 118
2 862 1 120
2 863 1 120
2 864 1 123
2 865 1 123
2 866 1 126
2 867 1 126
2 868 1 128
2 869 1 128
2 870 1 131
2 871 1 131
2 872 1 134
2 873 1 134
2 874 1 136
2 875 1 136
2 876 1 139
2 877 1 139
2 878 1 142
2 879 1 142
2 880 1 144
2 881 1 144
2 882 1 147
2 883 1 147
2 884 1 150
2 885 1 150
2 886 1 152
2 887 1 152
2 888 1 155
2 889 1 155
2 890 1 158
2 891 1 158
2 892 1 160
2 893 1 160
2 894 1 163
2 895 1 163
2 896 1 166
2 897 1 166
2 898 1 168
2 899 1 168
2 900 1 171
2 901 1 171
2 902 1 174
2 903 1 174
2 904 1 176
2 905 1 176
2 906 1 179
2 907 1 179
2 908 1 182
2 909 1 182
2 910 1 184
2 911 1 184
2 912 1 187
2 913 1 187
2 914 1 190
2 915 1 190
2 916 1 192
2 917 1 192
2 918 1 195
2 919 1 195
2 920 1 198
2 921 1 198
2 922 1 200
2 923 1 200
2 924 1 203
2 925 1 203
2 926 1 206
2 927 1 206
2 928 1 208
2 929 1 208
2 930 1 211
2 931 1 211
2 932 1 214
2 933 1 214
2 934 1 216
2 935 1 216
2 936 1 219
2 937 1 219
2 938 1 221
2 939 1 221
2 940 1 222
2 941 1 222
2 942 1 223
2 943 1 223
2 944 1 229
2 945 1 229
2 946 1 232
2 947 1 232
2 948 1 232
2 949 1 234
2 950 1 234
2 951 1 234
2 952 1 235
2 953 1 235
2 954 1 241
2 955 1 241
2 956 1 244
2 957 1 244
2 958 1 244
2 959 1 244
2 960 1 246
2 961 1 246
2 962 1 246
2 963 1 247
2 964 1 247
2 965 1 253
2 966 1 253
2 967 1 256
2 968 1 256
2 969 1 256
2 970 1 256
2 971 1 258
2 972 1 258
2 973 1 258
2 974 1 259
2 975 1 259
2 976 1 265
2 977 1 265
2 978 1 268
2 979 1 268
2 980 1 268
2 981 1 268
2 982 1 270
2 983 1 270
2 984 1 270
2 985 1 271
2 986 1 271
2 987 1 277
2 988 1 277
2 989 1 280
2 990 1 280
2 991 1 280
2 992 1 282
2 993 1 282
2 994 1 282
2 995 1 283
2 996 1 283
2 997 1 289
2 998 1 289
2 999 1 292
2 1000 1 292
2 1001 1 292
2 1002 1 292
2 1003 1 294
2 1004 1 294
2 1005 1 294
2 1006 1 295
2 1007 1 295
2 1008 1 301
2 1009 1 301
2 1010 1 304
2 1011 1 304
2 1012 1 304
2 1013 1 304
2 1014 1 306
2 1015 1 306
2 1016 1 306
2 1017 1 306
2 1018 1 307
2 1019 1 307
2 1020 1 313
2 1021 1 313
2 1022 1 315
2 1023 1 315
2 1024 1 316
2 1025 1 316
2 1026 1 316
2 1027 1 317
2 1028 1 317
2 1029 1 323
2 1030 1 323
2 1031 1 325
2 1032 1 325
2 1033 1 326
2 1034 1 326
2 1035 1 326
2 1036 1 326
2 1037 1 327
2 1038 1 327
2 1039 1 328
2 1040 1 328
2 1041 1 328
2 1042 1 329
2 1043 1 329
2 1044 1 330
2 1045 1 330
2 1046 1 330
2 1047 1 331
2 1048 1 331
2 1049 1 337
2 1050 1 337
2 1051 1 340
2 1052 1 340
2 1053 1 340
2 1054 1 342
2 1055 1 342
2 1056 1 342
2 1057 1 343
2 1058 1 343
2 1059 1 349
2 1060 1 349
2 1061 1 352
2 1062 1 352
2 1063 1 352
2 1064 1 352
2 1065 1 354
2 1066 1 354
2 1067 1 354
2 1068 1 355
2 1069 1 355
2 1070 1 361
2 1071 1 361
2 1072 1 364
2 1073 1 364
2 1074 1 364
2 1075 1 366
2 1076 1 366
2 1077 1 366
2 1078 1 367
2 1079 1 367
2 1080 1 373
2 1081 1 373
2 1082 1 376
2 1083 1 376
2 1084 1 376
2 1085 1 378
2 1086 1 378
2 1087 1 378
2 1088 1 379
2 1089 1 379
2 1090 1 385
2 1091 1 385
2 1092 1 388
2 1093 1 388
2 1094 1 388
2 1095 1 390
2 1096 1 390
2 1097 1 390
2 1098 1 391
2 1099 1 391
2 1100 1 397
2 1101 1 397
2 1102 1 400
2 1103 1 400
2 1104 1 401
2 1105 1 401
2 1106 1 405
2 1107 1 405
2 1108 1 409
2 1109 1 409
2 1110 1 415
2 1111 1 415
2 1112 1 416
2 1113 1 416
2 1114 1 419
2 1115 1 419
2 1116 1 420
2 1117 1 420
2 1118 1 423
2 1119 1 423
2 1120 1 425
2 1121 1 425
2 1122 1 427
2 1123 1 427
2 1124 1 428
2 1125 1 428
2 1126 1 431
2 1127 1 431
2 1128 1 435
2 1129 1 435
2 1130 1 443
2 1131 1 443
2 1132 1 445
2 1133 1 445
2 1134 1 446
2 1135 1 446
2 1136 1 449
2 1137 1 449
2 1138 1 450
2 1139 1 450
2 1140 1 453
2 1141 1 453
2 1142 1 454
2 1143 1 454
2 1144 1 457
2 1145 1 457
2 1146 1 458
2 1147 1 458
2 1148 1 461
2 1149 1 461
2 1150 1 461
2 1151 1 465
2 1152 1 465
2 1153 1 473
2 1154 1 473
2 1155 1 474
2 1156 1 474
2 1157 1 478
2 1158 1 478
2 1159 1 489
2 1160 1 489
2 1161 1 489
2 1162 1 493
2 1163 1 493
2 1164 1 494
2 1165 1 494
2 1166 1 497
2 1167 1 497
2 1168 1 498
2 1169 1 498
2 1170 1 506
2 1171 1 506
2 1172 1 508
2 1173 1 508
2 1174 1 509
2 1175 1 509
2 1176 1 512
2 1177 1 512
2 1178 1 513
2 1179 1 513
2 1180 1 516
2 1181 1 516
2 1182 1 519
2 1183 1 519
2 1184 1 523
2 1185 1 523
2 1186 1 526
2 1187 1 526
2 1188 1 528
2 1189 1 528
2 1190 1 529
2 1191 1 529
2 1192 1 532
2 1193 1 532
2 1194 1 536
2 1195 1 536
2 1196 1 538
2 1197 1 538
2 1198 1 538
2 1199 1 539
2 1200 1 539
2 1201 1 546
2 1202 1 546
2 1203 1 546
2 1204 1 552
2 1205 1 552
2 1206 1 553
2 1207 1 553
2 1208 1 558
2 1209 1 558
2 1210 1 558
2 1211 1 559
2 1212 1 559
2 1213 1 564
2 1214 1 564
2 1215 1 565
2 1216 1 565
2 1217 1 571
2 1218 1 571
2 1219 1 582
2 1220 1 582
2 1221 1 582
2 1222 1 583
2 1223 1 583
2 1224 1 588
2 1225 1 588
2 1226 1 589
2 1227 1 589
2 1228 1 592
2 1229 1 592
2 1230 1 592
2 1231 1 598
2 1232 1 598
2 1233 1 598
2 1234 1 603
2 1235 1 603
2 1236 1 632
2 1237 1 632
2 1238 1 632
2 1239 1 670
2 1240 1 670
0 50 5 1 1 49
0 51 5 1 1 719
0 52 5 1 1 721
0 53 5 1 1 723
0 54 5 1 1 725
0 55 5 1 1 727
0 56 5 1 1 729
0 57 5 1 1 731
0 58 5 1 1 733
0 59 5 1 1 735
0 60 5 1 1 737
0 61 5 1 1 739
0 62 5 1 1 741
0 63 5 1 1 743
0 64 5 1 1 745
0 65 5 1 1 747
0 66 5 1 1 749
0 67 5 1 1 751
0 68 5 1 1 753
0 69 5 2 1 755
0 70 5 2 1 757
0 71 5 2 1 759
0 72 5 2 1 761
0 73 5 2 1 763
0 74 5 2 1 765
0 75 5 2 1 767
0 76 5 2 1 769
0 77 5 2 1 771
0 78 5 2 1 773
0 79 5 2 1 775
0 80 5 2 1 777
0 81 5 2 1 779
0 82 5 1 1 781
0 83 5 1 1 783
0 84 5 1 1 785
0 85 5 1 1 787
0 86 5 1 1 789
0 87 5 1 1 791
0 88 5 1 1 793
0 89 5 1 1 795
0 90 5 1 1 797
0 91 5 1 1 799
0 92 5 1 1 801
0 93 5 1 1 803
0 94 5 1 1 805
0 95 5 1 1 807
0 96 5 1 1 809
0 97 5 1 1 811
0 98 5 1 1 813
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 722 754
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 720 752
0 106 5 2 1 105
0 107 7 2 2 718 750
0 108 5 3 1 849
0 109 7 1 2 847 851
0 110 5 1 1 109
0 111 7 2 2 845 110
0 112 5 2 1 854
0 113 7 1 2 843 856
0 114 5 1 1 113
0 115 7 2 2 841 114
0 116 5 1 1 858
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 724 859
0 120 5 2 1 119
0 121 7 1 2 815 862
0 122 5 1 1 121
0 123 7 2 2 860 122
0 124 5 1 1 864
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 726 865
0 128 5 2 1 127
0 129 7 1 2 817 868
0 130 5 1 1 129
0 131 7 2 2 866 130
0 132 5 1 1 870
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 728 871
0 136 5 2 1 135
0 137 7 1 2 819 874
0 138 5 1 1 137
0 139 7 2 2 872 138
0 140 5 1 1 876
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 730 877
0 144 5 2 1 143
0 145 7 1 2 821 880
0 146 5 1 1 145
0 147 7 2 2 878 146
0 148 5 1 1 882
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 732 883
0 152 5 2 1 151
0 153 7 1 2 823 886
0 154 5 1 1 153
0 155 7 2 2 884 154
0 156 5 1 1 888
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 734 889
0 160 5 2 1 159
0 161 7 1 2 825 892
0 162 5 1 1 161
0 163 7 2 2 890 162
0 164 5 1 1 894
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 736 895
0 168 5 2 1 167
0 169 7 1 2 827 898
0 170 5 1 1 169
0 171 7 2 2 896 170
0 172 5 1 1 900
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 738 901
0 176 5 2 1 175
0 177 7 1 2 829 904
0 178 5 1 1 177
0 179 7 2 2 902 178
0 180 5 1 1 906
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 740 907
0 184 5 2 1 183
0 185 7 1 2 831 910
0 186 5 1 1 185
0 187 7 2 2 908 186
0 188 5 1 1 912
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 742 913
0 192 5 2 1 191
0 193 7 1 2 833 916
0 194 5 1 1 193
0 195 7 2 2 914 194
0 196 5 1 1 918
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 744 919
0 200 5 2 1 199
0 201 7 1 2 835 922
0 202 5 1 1 201
0 203 7 2 2 920 202
0 204 5 1 1 924
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 746 925
0 208 5 2 1 207
0 209 7 1 2 837 928
0 210 5 1 1 209
0 211 7 2 2 926 210
0 212 5 1 1 930
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 748 931
0 216 5 2 1 215
0 217 7 1 2 839 934
0 218 5 1 1 217
0 219 7 2 2 932 218
0 220 5 1 1 936
0 221 7 2 2 814 220
0 222 5 2 1 938
0 223 7 2 2 933 935
0 224 5 1 1 942
0 225 7 1 2 780 224
0 226 5 1 1 225
0 227 7 1 2 840 943
0 228 5 1 1 227
0 229 7 2 2 226 228
0 230 5 1 1 944
0 231 7 1 2 97 230
0 232 5 3 1 231
0 233 7 1 2 812 945
0 234 5 3 1 233
0 235 7 2 2 927 929
0 236 5 1 1 952
0 237 7 1 2 778 953
0 238 5 1 1 237
0 239 7 1 2 838 236
0 240 5 1 1 239
0 241 7 2 2 238 240
0 242 5 1 1 954
0 243 7 1 2 810 242
0 244 5 4 1 243
0 245 7 1 2 96 955
0 246 5 3 1 245
0 247 7 2 2 921 923
0 248 5 1 1 963
0 249 7 1 2 776 964
0 250 5 1 1 249
0 251 7 1 2 836 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 965
0 255 7 1 2 808 254
0 256 5 4 1 255
0 257 7 1 2 95 966
0 258 5 3 1 257
0 259 7 2 2 915 917
0 260 5 1 1 974
0 261 7 1 2 774 975
0 262 5 1 1 261
0 263 7 1 2 834 260
0 264 5 1 1 263
0 265 7 2 2 262 264
0 266 5 1 1 976
0 267 7 1 2 806 266
0 268 5 4 1 267
0 269 7 1 2 94 977
0 270 5 3 1 269
0 271 7 2 2 909 911
0 272 5 1 1 985
0 273 7 1 2 772 986
0 274 5 1 1 273
0 275 7 1 2 832 272
0 276 5 1 1 275
0 277 7 2 2 274 276
0 278 5 1 1 987
0 279 7 1 2 804 278
0 280 5 3 1 279
0 281 7 1 2 93 988
0 282 5 3 1 281
0 283 7 2 2 903 905
0 284 5 1 1 995
0 285 7 1 2 770 996
0 286 5 1 1 285
0 287 7 1 2 830 284
0 288 5 1 1 287
0 289 7 2 2 286 288
0 290 5 1 1 997
0 291 7 1 2 802 290
0 292 5 4 1 291
0 293 7 1 2 92 998
0 294 5 3 1 293
0 295 7 2 2 897 899
0 296 5 1 1 1006
0 297 7 1 2 768 1007
0 298 5 1 1 297
0 299 7 1 2 828 296
0 300 5 1 1 299
0 301 7 2 2 298 300
0 302 5 1 1 1008
0 303 7 1 2 91 1009
0 304 5 4 1 303
0 305 7 1 2 800 302
0 306 5 4 1 305
0 307 7 2 2 891 893
0 308 5 1 1 1018
0 309 7 1 2 766 1019
0 310 5 1 1 309
0 311 7 1 2 826 308
0 312 5 1 1 311
0 313 7 2 2 310 312
0 314 5 1 1 1020
0 315 7 2 2 90 1021
0 316 5 3 1 1022
0 317 7 2 2 885 887
0 318 5 1 1 1027
0 319 7 1 2 764 1028
0 320 5 1 1 319
0 321 7 1 2 824 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1029
0 325 7 2 2 796 324
0 326 5 4 1 1031
0 327 7 2 2 798 314
0 328 5 3 1 1037
0 329 7 2 2 89 1030
0 330 5 3 1 1042
0 331 7 2 2 879 881
0 332 5 1 1 1047
0 333 7 1 2 762 1048
0 334 5 1 1 333
0 335 7 1 2 822 332
0 336 5 1 1 335
0 337 7 2 2 334 336
0 338 5 1 1 1049
0 339 7 1 2 794 338
0 340 5 3 1 339
0 341 7 1 2 88 1050
0 342 5 3 1 341
0 343 7 2 2 873 875
0 344 5 1 1 1057
0 345 7 1 2 760 1058
0 346 5 1 1 345
0 347 7 1 2 820 344
0 348 5 1 1 347
0 349 7 2 2 346 348
0 350 5 1 1 1059
0 351 7 1 2 792 350
0 352 5 4 1 351
0 353 7 1 2 87 1060
0 354 5 3 1 353
0 355 7 2 2 867 869
0 356 5 1 1 1068
0 357 7 1 2 758 1069
0 358 5 1 1 357
0 359 7 1 2 818 356
0 360 5 1 1 359
0 361 7 2 2 358 360
0 362 5 1 1 1070
0 363 7 1 2 790 362
0 364 5 3 1 363
0 365 7 1 2 86 1071
0 366 5 3 1 365
0 367 7 2 2 861 863
0 368 5 1 1 1078
0 369 7 1 2 756 1079
0 370 5 1 1 369
0 371 7 1 2 816 368
0 372 5 1 1 371
0 373 7 2 2 370 372
0 374 5 1 1 1080
0 375 7 1 2 788 374
0 376 5 3 1 375
0 377 7 1 2 85 1081
0 378 5 3 1 377
0 379 7 2 2 842 844
0 380 5 1 1 1088
0 381 7 1 2 855 380
0 382 5 1 1 381
0 383 7 1 2 857 1089
0 384 5 1 1 383
0 385 7 2 2 382 384
0 386 5 1 1 1090
0 387 7 1 2 786 1091
0 388 5 3 1 387
0 389 7 1 2 84 386
0 390 5 3 1 389
0 391 7 2 2 846 848
0 392 5 1 1 1098
0 393 7 1 2 850 392
0 394 5 1 1 393
0 395 7 1 2 852 1099
0 396 5 1 1 395
0 397 7 2 2 394 396
0 398 5 1 1 1100
0 399 7 1 2 784 1101
0 400 5 2 1 399
0 401 7 2 2 83 398
0 402 5 1 1 1104
0 403 7 1 2 50 66
0 404 5 1 1 403
0 405 7 2 2 853 404
0 406 5 1 1 1106
0 407 7 1 2 82 1107
0 408 5 1 1 407
0 409 7 2 2 402 408
0 410 5 1 1 1108
0 411 7 1 2 1102 410
0 412 5 1 1 411
0 413 7 1 2 1095 412
0 414 5 1 1 413
0 415 7 2 2 1092 414
0 416 5 2 1 1110
0 417 7 1 2 1085 1112
0 418 5 1 1 417
0 419 7 2 2 1082 418
0 420 5 2 1 1114
0 421 7 1 2 1075 1116
0 422 5 1 1 421
0 423 7 2 2 1072 422
0 424 5 1 1 1118
0 425 7 2 2 1065 424
0 426 5 1 1 1120
0 427 7 2 2 1061 426
0 428 5 2 1 1122
0 429 7 1 2 1054 1124
0 430 5 1 1 429
0 431 7 2 2 1051 430
0 432 5 1 1 1126
0 433 7 1 2 1044 432
0 434 5 1 1 433
0 435 7 2 2 1039 434
0 436 7 1 2 1033 1128
0 437 5 1 1 436
0 438 7 1 2 1024 437
0 439 5 1 1 438
0 440 7 1 2 1014 439
0 441 5 1 1 440
0 442 7 1 2 1010 441
0 443 7 2 2 1003 442
0 444 5 1 1 1130
0 445 7 2 2 999 444
0 446 5 2 1 1132
0 447 7 1 2 992 1134
0 448 5 1 1 447
0 449 7 2 2 989 448
0 450 5 2 1 1136
0 451 7 1 2 982 1138
0 452 5 1 1 451
0 453 7 2 2 978 452
0 454 5 2 1 1140
0 455 7 1 2 971 1142
0 456 5 1 1 455
0 457 7 2 2 967 456
0 458 5 2 1 1144
0 459 7 1 2 960 1146
0 460 5 1 1 459
0 461 7 3 2 956 460
0 462 5 1 1 1148
0 463 7 1 2 949 1149
0 464 5 1 1 463
0 465 7 2 2 946 464
0 466 5 1 1 1151
0 467 7 1 2 940 1152
0 468 5 1 1 467
0 469 7 1 2 939 466
0 470 5 1 1 469
0 471 7 1 2 468 470
0 472 5 1 1 471
0 473 7 2 2 98 937
0 474 5 2 1 1153
0 475 7 1 2 782 406
0 476 5 1 1 475
0 477 7 1 2 476 1103
0 478 7 2 2 1093 477
0 479 5 1 1 1157
0 480 7 1 2 1094 1105
0 481 5 1 1 480
0 482 7 1 2 481 1096
0 483 7 1 2 479 482
0 484 7 1 2 1086 483
0 485 5 1 1 484
0 486 7 1 2 1083 485
0 487 7 1 2 1073 486
0 488 5 1 1 487
0 489 7 3 2 1076 488
0 490 5 1 1 1159
0 491 7 1 2 1066 1160
0 492 5 1 1 491
0 493 7 2 2 1062 492
0 494 5 2 1 1162
0 495 7 1 2 1055 1164
0 496 5 1 1 495
0 497 7 2 2 1052 496
0 498 5 2 1 1166
0 499 7 1 2 1045 1168
0 500 5 1 1 499
0 501 7 1 2 1034 500
0 502 5 1 1 501
0 503 7 1 2 1025 502
0 504 5 1 1 503
0 505 7 1 2 504 1040
0 506 7 2 2 1015 505
0 507 5 1 1 1170
0 508 7 2 2 1011 507
0 509 5 2 1 1172
0 510 7 1 2 1000 1174
0 511 5 1 1 510
0 512 7 2 2 1004 511
0 513 5 2 1 1176
0 514 7 1 2 990 1178
0 515 5 1 1 514
0 516 7 2 2 993 515
0 517 5 1 1 1180
0 518 7 1 2 983 1181
0 519 5 2 1 518
0 520 7 1 2 979 1182
0 521 5 1 1 520
0 522 7 1 2 972 521
0 523 5 2 1 522
0 524 7 1 2 968 1184
0 525 5 1 1 524
0 526 7 2 2 961 525
0 527 5 1 1 1186
0 528 7 2 2 957 527
0 529 5 2 1 1188
0 530 7 1 2 947 1190
0 531 5 1 1 530
0 532 7 2 2 950 531
0 533 5 1 1 1192
0 534 7 1 2 1155 533
0 535 5 1 1 534
0 536 7 2 2 941 535
0 537 5 1 1 1194
0 538 7 3 2 951 948
0 539 5 2 1 1196
0 540 7 1 2 1150 1199
0 541 5 1 1 540
0 542 7 1 2 462 1197
0 543 5 1 1 542
0 544 7 1 2 541 543
0 545 5 1 1 544
0 546 7 3 2 969 973
0 547 5 1 1 1201
0 548 7 1 2 1141 1202
0 549 5 1 1 548
0 550 7 1 2 1143 547
0 551 5 1 1 550
0 552 7 2 2 980 984
0 553 5 2 1 1204
0 554 7 1 2 1139 1206
0 555 5 1 1 554
0 556 7 1 2 1137 1205
0 557 5 1 1 556
0 558 7 3 2 994 991
0 559 5 2 1 1208
0 560 7 1 2 1135 1209
0 561 5 1 1 560
0 562 7 1 2 1133 1211
0 563 5 1 1 562
0 564 7 2 2 1005 1001
0 565 5 2 1 1213
0 566 7 1 2 1016 1215
0 567 5 1 1 566
0 568 7 1 2 1002 1131
0 569 5 1 1 568
0 570 7 1 2 1012 1017
0 571 5 2 1 570
0 572 7 1 2 1041 1217
0 573 5 1 1 572
0 574 7 1 2 1026 1129
0 575 5 1 1 574
0 576 7 1 2 1035 575
0 577 5 1 1 576
0 578 7 1 2 1036 1046
0 579 5 1 1 578
0 580 7 1 2 1127 579
0 581 5 1 1 580
0 582 7 3 2 1053 1056
0 583 5 2 1 1219
0 584 7 1 2 1123 1220
0 585 5 1 1 584
0 586 7 1 2 1063 1121
0 587 5 1 1 586
0 588 7 2 2 1064 1067
0 589 5 2 1 1224
0 590 7 1 2 1119 1226
0 591 5 1 1 590
0 592 7 3 2 1077 1074
0 593 5 1 1 1228
0 594 7 1 2 1115 1229
0 595 5 1 1 594
0 596 7 1 2 1117 593
0 597 5 1 1 596
0 598 7 3 2 1084 1087
0 599 5 1 1 1231
0 600 7 1 2 1111 1232
0 601 5 1 1 600
0 602 7 1 2 1097 1109
0 603 7 2 2 1158 602
0 604 7 1 2 1113 599
0 605 5 1 1 604
0 606 7 1 2 1234 605
0 607 7 1 2 601 606
0 608 7 1 2 597 607
0 609 7 1 2 595 608
0 610 5 1 1 609
0 611 7 1 2 591 610
0 612 7 1 2 587 611
0 613 5 1 1 612
0 614 7 1 2 1125 1222
0 615 5 1 1 614
0 616 7 1 2 613 615
0 617 7 1 2 585 616
0 618 5 1 1 617
0 619 7 1 2 581 618
0 620 7 1 2 577 619
0 621 7 1 2 573 620
0 622 7 1 2 569 621
0 623 7 1 2 567 622
0 624 7 1 2 563 623
0 625 7 1 2 561 624
0 626 5 1 1 625
0 627 7 1 2 557 626
0 628 7 1 2 555 627
0 629 7 1 2 551 628
0 630 7 1 2 549 629
0 631 7 1 2 1156 630
0 632 7 3 2 958 962
0 633 5 1 1 1236
0 634 7 1 2 1145 1237
0 635 5 1 1 634
0 636 7 1 2 1147 633
0 637 5 1 1 636
0 638 7 1 2 635 637
0 639 7 1 2 631 638
0 640 7 1 2 545 639
0 641 7 1 2 537 640
0 642 7 1 2 472 641
0 643 5 1 1 642
0 644 7 1 2 1154 1193
0 645 5 1 1 644
0 646 7 1 2 1189 1200
0 647 5 1 1 646
0 648 7 1 2 1191 1198
0 649 5 1 1 648
0 650 7 1 2 1185 1238
0 651 5 1 1 650
0 652 7 1 2 970 651
0 653 5 1 1 652
0 654 7 1 2 959 1187
0 655 5 1 1 654
0 656 7 1 2 1183 1203
0 657 5 1 1 656
0 658 7 1 2 981 657
0 659 5 1 1 658
0 660 7 1 2 517 1207
0 661 5 1 1 660
0 662 7 1 2 1177 1212
0 663 5 1 1 662
0 664 7 1 2 1179 1210
0 665 5 1 1 664
0 666 7 1 2 1173 1216
0 667 5 1 1 666
0 668 7 1 2 1175 1214
0 669 5 1 1 668
0 670 7 2 2 1043 1167
0 671 5 1 1 1239
0 672 7 1 2 1023 1240
0 673 5 1 1 672
0 674 7 1 2 1218 673
0 675 5 1 1 674
0 676 7 1 2 1013 1171
0 677 5 1 1 676
0 678 7 1 2 1038 671
0 679 5 1 1 678
0 680 7 1 2 1032 1169
0 681 5 1 1 680
0 682 7 1 2 1163 1223
0 683 5 1 1 682
0 684 7 1 2 1165 1221
0 685 5 1 1 684
0 686 7 1 2 1161 1227
0 687 5 1 1 686
0 688 7 1 2 1235 1233
0 689 7 1 2 1230 688
0 690 5 1 1 689
0 691 7 1 2 490 1225
0 692 5 1 1 691
0 693 7 1 2 690 692
0 694 7 1 2 687 693
0 695 5 1 1 694
0 696 7 1 2 685 695
0 697 7 1 2 683 696
0 698 5 1 1 697
0 699 7 1 2 681 698
0 700 7 1 2 679 699
0 701 7 1 2 677 700
0 702 7 1 2 675 701
0 703 7 1 2 669 702
0 704 7 1 2 667 703
0 705 7 1 2 665 704
0 706 7 1 2 663 705
0 707 5 1 1 706
0 708 7 1 2 661 707
0 709 7 1 2 659 708
0 710 7 1 2 655 709
0 711 7 1 2 653 710
0 712 7 1 2 649 711
0 713 7 1 2 647 712
0 714 7 1 2 645 713
0 715 7 1 2 1195 714
0 716 5 1 1 715
0 717 7 1 2 643 716
3 3499 5 0 1 717
