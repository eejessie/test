1 0 0 2 0
2 49 1 0
2 1952 1 0
1 1 0 2 0
2 1953 1 1
2 1954 1 1
1 2 0 2 0
2 1955 1 2
2 1956 1 2
1 3 0 2 0
2 1957 1 3
2 1958 1 3
1 4 0 2 0
2 1959 1 4
2 1960 1 4
1 5 0 2 0
2 1961 1 5
2 1962 1 5
1 6 0 2 0
2 1963 1 6
2 1964 1 6
1 7 0 2 0
2 1965 1 7
2 1966 1 7
1 8 0 2 0
2 1967 1 8
2 1968 1 8
1 9 0 2 0
2 1969 1 9
2 1970 1 9
1 10 0 2 0
2 1971 1 10
2 1972 1 10
1 11 0 2 0
2 1973 1 11
2 1974 1 11
1 12 0 2 0
2 1975 1 12
2 1976 1 12
1 13 0 2 0
2 1977 1 13
2 1978 1 13
1 14 0 2 0
2 1979 1 14
2 1980 1 14
1 15 0 2 0
2 1981 1 15
2 1982 1 15
1 16 0 2 0
2 1983 1 16
2 1984 1 16
1 17 0 2 0
2 1985 1 17
2 1986 1 17
1 18 0 2 0
2 1987 1 18
2 1988 1 18
1 19 0 2 0
2 1989 1 19
2 1990 1 19
1 20 0 2 0
2 1991 1 20
2 1992 1 20
1 21 0 2 0
2 1993 1 21
2 1994 1 21
1 22 0 2 0
2 1995 1 22
2 1996 1 22
1 23 0 2 0
2 1997 1 23
2 1998 1 23
1 24 0 2 0
2 1999 1 24
2 2000 1 24
1 25 0 2 0
2 2001 1 25
2 2002 1 25
1 26 0 2 0
2 2003 1 26
2 2004 1 26
1 27 0 2 0
2 2005 1 27
2 2006 1 27
1 28 0 2 0
2 2007 1 28
2 2008 1 28
1 29 0 2 0
2 2009 1 29
2 2010 1 29
1 30 0 2 0
2 2011 1 30
2 2012 1 30
1 31 0 2 0
2 2013 1 31
2 2014 1 31
1 32 0 2 0
2 2015 1 32
2 2016 1 32
1 33 0 2 0
2 2017 1 33
2 2018 1 33
1 34 0 2 0
2 2019 1 34
2 2020 1 34
1 35 0 2 0
2 2021 1 35
2 2022 1 35
1 36 0 2 0
2 2023 1 36
2 2024 1 36
1 37 0 2 0
2 2025 1 37
2 2026 1 37
1 38 0 2 0
2 2027 1 38
2 2028 1 38
1 39 0 2 0
2 2029 1 39
2 2030 1 39
1 40 0 2 0
2 2031 1 40
2 2032 1 40
1 41 0 2 0
2 2033 1 41
2 2034 1 41
1 42 0 2 0
2 2035 1 42
2 2036 1 42
1 43 0 2 0
2 2037 1 43
2 2038 1 43
1 44 0 2 0
2 2039 1 44
2 2040 1 44
1 45 0 2 0
2 2041 1 45
2 2042 1 45
1 46 0 2 0
2 2043 1 46
2 2044 1 46
1 47 0 2 0
2 2045 1 47
2 2046 1 47
1 48 0 2 0
2 2047 1 48
2 2048 1 48
2 2049 1 69
2 2050 1 69
2 2051 1 70
2 2052 1 70
2 2053 1 71
2 2054 1 71
2 2055 1 72
2 2056 1 72
2 2057 1 73
2 2058 1 73
2 2059 1 74
2 2060 1 74
2 2061 1 75
2 2062 1 75
2 2063 1 76
2 2064 1 76
2 2065 1 77
2 2066 1 77
2 2067 1 78
2 2068 1 78
2 2069 1 79
2 2070 1 79
2 2071 1 80
2 2072 1 80
2 2073 1 100
2 2074 1 100
2 2075 1 102
2 2076 1 102
2 2077 1 104
2 2078 1 104
2 2079 1 106
2 2080 1 106
2 2081 1 107
2 2082 1 107
2 2083 1 108
2 2084 1 108
2 2085 1 108
2 2086 1 111
2 2087 1 111
2 2088 1 112
2 2089 1 112
2 2090 1 115
2 2091 1 115
2 2092 1 118
2 2093 1 118
2 2094 1 120
2 2095 1 120
2 2096 1 123
2 2097 1 123
2 2098 1 126
2 2099 1 126
2 2100 1 128
2 2101 1 128
2 2102 1 131
2 2103 1 131
2 2104 1 134
2 2105 1 134
2 2106 1 136
2 2107 1 136
2 2108 1 139
2 2109 1 139
2 2110 1 142
2 2111 1 142
2 2112 1 144
2 2113 1 144
2 2114 1 147
2 2115 1 147
2 2116 1 150
2 2117 1 150
2 2118 1 152
2 2119 1 152
2 2120 1 155
2 2121 1 155
2 2122 1 158
2 2123 1 158
2 2124 1 160
2 2125 1 160
2 2126 1 163
2 2127 1 163
2 2128 1 166
2 2129 1 166
2 2130 1 168
2 2131 1 168
2 2132 1 171
2 2133 1 171
2 2134 1 174
2 2135 1 174
2 2136 1 176
2 2137 1 176
2 2138 1 179
2 2139 1 179
2 2140 1 182
2 2141 1 182
2 2142 1 184
2 2143 1 184
2 2144 1 187
2 2145 1 187
2 2146 1 190
2 2147 1 190
2 2148 1 192
2 2149 1 192
2 2150 1 195
2 2151 1 195
2 2152 1 198
2 2153 1 198
2 2154 1 200
2 2155 1 200
2 2156 1 203
2 2157 1 203
2 2158 1 206
2 2159 1 206
2 2160 1 208
2 2161 1 208
2 2162 1 211
2 2163 1 211
2 2164 1 211
2 2165 1 212
2 2166 1 212
2 2167 1 212
2 2168 1 213
2 2169 1 213
2 2170 1 214
2 2171 1 214
2 2172 1 216
2 2173 1 216
2 2174 1 217
2 2175 1 217
2 2176 1 223
2 2177 1 223
2 2178 1 223
2 2179 1 223
2 2180 1 224
2 2181 1 224
2 2182 1 224
2 2183 1 225
2 2184 1 225
2 2185 1 226
2 2186 1 226
2 2187 1 227
2 2188 1 227
2 2189 1 233
2 2190 1 233
2 2191 1 233
2 2192 1 234
2 2193 1 234
2 2194 1 236
2 2195 1 236
2 2196 1 237
2 2197 1 237
2 2198 1 243
2 2199 1 243
2 2200 1 243
2 2201 1 243
2 2202 1 244
2 2203 1 244
2 2204 1 244
2 2205 1 246
2 2206 1 246
2 2207 1 247
2 2208 1 247
2 2209 1 253
2 2210 1 253
2 2211 1 253
2 2212 1 253
2 2213 1 254
2 2214 1 254
2 2215 1 254
2 2216 1 256
2 2217 1 256
2 2218 1 257
2 2219 1 257
2 2220 1 263
2 2221 1 263
2 2222 1 263
2 2223 1 263
2 2224 1 264
2 2225 1 264
2 2226 1 264
2 2227 1 266
2 2228 1 266
2 2229 1 267
2 2230 1 267
2 2231 1 273
2 2232 1 273
2 2233 1 273
2 2234 1 273
2 2235 1 274
2 2236 1 274
2 2237 1 274
2 2238 1 276
2 2239 1 276
2 2240 1 277
2 2241 1 277
2 2242 1 283
2 2243 1 283
2 2244 1 283
2 2245 1 283
2 2246 1 284
2 2247 1 284
2 2248 1 284
2 2249 1 286
2 2250 1 286
2 2251 1 287
2 2252 1 287
2 2253 1 293
2 2254 1 293
2 2255 1 293
2 2256 1 293
2 2257 1 294
2 2258 1 294
2 2259 1 294
2 2260 1 296
2 2261 1 296
2 2262 1 297
2 2263 1 297
2 2264 1 303
2 2265 1 303
2 2266 1 303
2 2267 1 303
2 2268 1 304
2 2269 1 304
2 2270 1 304
2 2271 1 306
2 2272 1 306
2 2273 1 307
2 2274 1 307
2 2275 1 313
2 2276 1 313
2 2277 1 313
2 2278 1 313
2 2279 1 314
2 2280 1 314
2 2281 1 314
2 2282 1 316
2 2283 1 316
2 2284 1 317
2 2285 1 317
2 2286 1 323
2 2287 1 323
2 2288 1 323
2 2289 1 323
2 2290 1 324
2 2291 1 324
2 2292 1 324
2 2293 1 326
2 2294 1 326
2 2295 1 327
2 2296 1 327
2 2297 1 333
2 2298 1 333
2 2299 1 333
2 2300 1 333
2 2301 1 334
2 2302 1 334
2 2303 1 334
2 2304 1 336
2 2305 1 336
2 2306 1 337
2 2307 1 337
2 2308 1 343
2 2309 1 343
2 2310 1 343
2 2311 1 343
2 2312 1 344
2 2313 1 344
2 2314 1 344
2 2315 1 346
2 2316 1 346
2 2317 1 347
2 2318 1 347
2 2319 1 353
2 2320 1 353
2 2321 1 353
2 2322 1 353
2 2323 1 354
2 2324 1 354
2 2325 1 356
2 2326 1 356
2 2327 1 359
2 2328 1 359
2 2329 1 360
2 2330 1 360
2 2331 1 363
2 2332 1 363
2 2333 1 369
2 2334 1 369
2 2335 1 370
2 2336 1 370
2 2337 1 371
2 2338 1 371
2 2339 1 375
2 2340 1 375
2 2341 1 378
2 2342 1 378
2 2343 1 379
2 2344 1 379
2 2345 1 383
2 2346 1 383
2 2347 1 386
2 2348 1 386
2 2349 1 387
2 2350 1 387
2 2351 1 391
2 2352 1 391
2 2353 1 394
2 2354 1 394
2 2355 1 395
2 2356 1 395
2 2357 1 399
2 2358 1 399
2 2359 1 402
2 2360 1 402
2 2361 1 403
2 2362 1 403
2 2363 1 407
2 2364 1 407
2 2365 1 410
2 2366 1 410
2 2367 1 411
2 2368 1 411
2 2369 1 415
2 2370 1 415
2 2371 1 418
2 2372 1 418
2 2373 1 419
2 2374 1 419
2 2375 1 423
2 2376 1 423
2 2377 1 426
2 2378 1 426
2 2379 1 427
2 2380 1 427
2 2381 1 431
2 2382 1 431
2 2383 1 434
2 2384 1 434
2 2385 1 435
2 2386 1 435
2 2387 1 439
2 2388 1 439
2 2389 1 442
2 2390 1 442
2 2391 1 443
2 2392 1 443
2 2393 1 447
2 2394 1 447
2 2395 1 450
2 2396 1 450
2 2397 1 451
2 2398 1 451
2 2399 1 455
2 2400 1 455
2 2401 1 458
2 2402 1 458
2 2403 1 459
2 2404 1 459
2 2405 1 463
2 2406 1 463
2 2407 1 466
2 2408 1 466
2 2409 1 467
2 2410 1 467
2 2411 1 471
2 2412 1 471
2 2413 1 474
2 2414 1 474
2 2415 1 475
2 2416 1 475
2 2417 1 479
2 2418 1 479
2 2419 1 481
2 2420 1 481
2 2421 1 482
2 2422 1 482
2 2423 1 485
2 2424 1 485
2 2425 1 485
2 2426 1 486
2 2427 1 486
2 2428 1 489
2 2429 1 489
2 2430 1 489
2 2431 1 489
2 2432 1 490
2 2433 1 490
2 2434 1 492
2 2435 1 492
2 2436 1 492
2 2437 1 494
2 2438 1 494
2 2439 1 494
2 2440 1 496
2 2441 1 496
2 2442 1 496
2 2443 1 498
2 2444 1 498
2 2445 1 498
2 2446 1 500
2 2447 1 500
2 2448 1 500
2 2449 1 502
2 2450 1 502
2 2451 1 502
2 2452 1 504
2 2453 1 504
2 2454 1 504
2 2455 1 506
2 2456 1 506
2 2457 1 506
2 2458 1 508
2 2459 1 508
2 2460 1 508
2 2461 1 510
2 2462 1 510
2 2463 1 510
2 2464 1 512
2 2465 1 512
2 2466 1 512
2 2467 1 514
2 2468 1 514
2 2469 1 514
2 2470 1 516
2 2471 1 516
2 2472 1 516
2 2473 1 518
2 2474 1 518
2 2475 1 518
2 2476 1 520
2 2477 1 520
2 2478 1 520
2 2479 1 522
2 2480 1 522
2 2481 1 522
2 2482 1 523
2 2483 1 523
2 2484 1 523
2 2485 1 524
2 2486 1 524
2 2487 1 527
2 2488 1 527
2 2489 1 528
2 2490 1 528
2 2491 1 531
2 2492 1 531
2 2493 1 532
2 2494 1 532
2 2495 1 535
2 2496 1 535
2 2497 1 536
2 2498 1 536
2 2499 1 539
2 2500 1 539
2 2501 1 540
2 2502 1 540
2 2503 1 543
2 2504 1 543
2 2505 1 544
2 2506 1 544
2 2507 1 547
2 2508 1 547
2 2509 1 548
2 2510 1 548
2 2511 1 551
2 2512 1 551
2 2513 1 552
2 2514 1 552
2 2515 1 555
2 2516 1 555
2 2517 1 556
2 2518 1 556
2 2519 1 558
2 2520 1 558
2 2521 1 558
2 2522 1 560
2 2523 1 560
2 2524 1 560
2 2525 1 561
2 2526 1 561
2 2527 1 561
2 2528 1 562
2 2529 1 562
2 2530 1 567
2 2531 1 567
2 2532 1 567
2 2533 1 567
2 2534 1 568
2 2535 1 568
2 2536 1 568
2 2537 1 570
2 2538 1 570
2 2539 1 570
2 2540 1 572
2 2541 1 572
2 2542 1 572
2 2543 1 573
2 2544 1 573
2 2545 1 573
2 2546 1 574
2 2547 1 574
2 2548 1 576
2 2549 1 576
2 2550 1 576
2 2551 1 578
2 2552 1 578
2 2553 1 578
2 2554 1 580
2 2555 1 580
2 2556 1 580
2 2557 1 582
2 2558 1 582
2 2559 1 582
2 2560 1 584
2 2561 1 584
2 2562 1 584
2 2563 1 586
2 2564 1 586
2 2565 1 586
2 2566 1 589
2 2567 1 589
2 2568 1 590
2 2569 1 590
2 2570 1 593
2 2571 1 593
2 2572 1 594
2 2573 1 594
2 2574 1 597
2 2575 1 597
2 2576 1 598
2 2577 1 598
2 2578 1 601
2 2579 1 601
2 2580 1 602
2 2581 1 602
2 2582 1 607
2 2583 1 607
2 2584 1 607
2 2585 1 607
2 2586 1 608
2 2587 1 608
2 2588 1 608
2 2589 1 608
2 2590 1 610
2 2591 1 610
2 2592 1 613
2 2593 1 613
2 2594 1 615
2 2595 1 615
2 2596 1 615
2 2597 1 616
2 2598 1 616
2 2599 1 621
2 2600 1 621
2 2601 1 621
2 2602 1 621
2 2603 1 622
2 2604 1 622
2 2605 1 622
2 2606 1 624
2 2607 1 624
2 2608 1 625
2 2609 1 625
2 2610 1 627
2 2611 1 627
2 2612 1 627
2 2613 1 628
2 2614 1 628
2 2615 1 633
2 2616 1 633
2 2617 1 633
2 2618 1 633
2 2619 1 634
2 2620 1 634
2 2621 1 634
2 2622 1 636
2 2623 1 636
2 2624 1 636
2 2625 1 638
2 2626 1 638
2 2627 1 638
2 2628 1 639
2 2629 1 639
2 2630 1 639
2 2631 1 640
2 2632 1 640
2 2633 1 643
2 2634 1 643
2 2635 1 644
2 2636 1 644
2 2637 1 649
2 2638 1 649
2 2639 1 649
2 2640 1 649
2 2641 1 650
2 2642 1 650
2 2643 1 650
2 2644 1 652
2 2645 1 652
2 2646 1 655
2 2647 1 655
2 2648 1 658
2 2649 1 658
2 2650 1 661
2 2651 1 661
2 2652 1 664
2 2653 1 664
2 2654 1 665
2 2655 1 665
2 2656 1 665
2 2657 1 666
2 2658 1 666
2 2659 1 671
2 2660 1 671
2 2661 1 671
2 2662 1 671
2 2663 1 672
2 2664 1 672
2 2665 1 672
2 2666 1 673
2 2667 1 673
2 2668 1 673
2 2669 1 674
2 2670 1 674
2 2671 1 679
2 2672 1 679
2 2673 1 679
2 2674 1 679
2 2675 1 680
2 2676 1 680
2 2677 1 680
2 2678 1 682
2 2679 1 682
2 2680 1 685
2 2681 1 685
2 2682 1 688
2 2683 1 688
2 2684 1 689
2 2685 1 689
2 2686 1 693
2 2687 1 693
2 2688 1 696
2 2689 1 696
2 2690 1 697
2 2691 1 697
2 2692 1 697
2 2693 1 698
2 2694 1 698
2 2695 1 703
2 2696 1 703
2 2697 1 703
2 2698 1 703
2 2699 1 704
2 2700 1 704
2 2701 1 704
2 2702 1 706
2 2703 1 706
2 2704 1 709
2 2705 1 709
2 2706 1 712
2 2707 1 712
2 2708 1 713
2 2709 1 713
2 2710 1 717
2 2711 1 717
2 2712 1 720
2 2713 1 720
2 2714 1 721
2 2715 1 721
2 2716 1 721
2 2717 1 722
2 2718 1 722
2 2719 1 727
2 2720 1 727
2 2721 1 727
2 2722 1 727
2 2723 1 728
2 2724 1 728
2 2725 1 728
2 2726 1 730
2 2727 1 730
2 2728 1 733
2 2729 1 733
2 2730 1 736
2 2731 1 736
2 2732 1 737
2 2733 1 737
2 2734 1 741
2 2735 1 741
2 2736 1 744
2 2737 1 744
2 2738 1 745
2 2739 1 745
2 2740 1 745
2 2741 1 746
2 2742 1 746
2 2743 1 751
2 2744 1 751
2 2745 1 751
2 2746 1 751
2 2747 1 752
2 2748 1 752
2 2749 1 752
2 2750 1 754
2 2751 1 754
2 2752 1 757
2 2753 1 757
2 2754 1 760
2 2755 1 760
2 2756 1 761
2 2757 1 761
2 2758 1 765
2 2759 1 765
2 2760 1 768
2 2761 1 768
2 2762 1 769
2 2763 1 769
2 2764 1 769
2 2765 1 770
2 2766 1 770
2 2767 1 775
2 2768 1 775
2 2769 1 775
2 2770 1 775
2 2771 1 776
2 2772 1 776
2 2773 1 776
2 2774 1 778
2 2775 1 778
2 2776 1 781
2 2777 1 781
2 2778 1 784
2 2779 1 784
2 2780 1 785
2 2781 1 785
2 2782 1 789
2 2783 1 789
2 2784 1 792
2 2785 1 792
2 2786 1 793
2 2787 1 793
2 2788 1 793
2 2789 1 794
2 2790 1 794
2 2791 1 799
2 2792 1 799
2 2793 1 799
2 2794 1 799
2 2795 1 799
2 2796 1 800
2 2797 1 800
2 2798 1 800
2 2799 1 802
2 2800 1 802
2 2801 1 805
2 2802 1 805
2 2803 1 808
2 2804 1 808
2 2805 1 809
2 2806 1 809
2 2807 1 813
2 2808 1 813
2 2809 1 816
2 2810 1 816
2 2811 1 817
2 2812 1 817
2 2813 1 817
2 2814 1 818
2 2815 1 818
2 2816 1 823
2 2817 1 823
2 2818 1 823
2 2819 1 823
2 2820 1 824
2 2821 1 824
2 2822 1 826
2 2823 1 826
2 2824 1 829
2 2825 1 829
2 2826 1 832
2 2827 1 832
2 2828 1 833
2 2829 1 833
2 2830 1 837
2 2831 1 837
2 2832 1 840
2 2833 1 840
2 2834 1 841
2 2835 1 841
2 2836 1 841
2 2837 1 842
2 2838 1 842
2 2839 1 847
2 2840 1 847
2 2841 1 847
2 2842 1 847
2 2843 1 848
2 2844 1 848
2 2845 1 850
2 2846 1 850
2 2847 1 853
2 2848 1 853
2 2849 1 856
2 2850 1 856
2 2851 1 857
2 2852 1 857
2 2853 1 861
2 2854 1 861
2 2855 1 864
2 2856 1 864
2 2857 1 865
2 2858 1 865
2 2859 1 866
2 2860 1 866
2 2861 1 869
2 2862 1 869
2 2863 1 872
2 2864 1 872
2 2865 1 875
2 2866 1 875
2 2867 1 877
2 2868 1 877
2 2869 1 878
2 2870 1 878
2 2871 1 878
2 2872 1 879
2 2873 1 879
2 2874 1 879
2 2875 1 880
2 2876 1 880
2 2877 1 880
2 2878 1 880
2 2879 1 880
2 2880 1 883
2 2881 1 883
2 2882 1 884
2 2883 1 884
2 2884 1 887
2 2885 1 887
2 2886 1 890
2 2887 1 890
2 2888 1 891
2 2889 1 891
2 2890 1 895
2 2891 1 895
2 2892 1 898
2 2893 1 898
2 2894 1 899
2 2895 1 899
2 2896 1 903
2 2897 1 903
2 2898 1 906
2 2899 1 906
2 2900 1 907
2 2901 1 907
2 2902 1 911
2 2903 1 911
2 2904 1 914
2 2905 1 914
2 2906 1 915
2 2907 1 915
2 2908 1 919
2 2909 1 919
2 2910 1 922
2 2911 1 922
2 2912 1 923
2 2913 1 923
2 2914 1 927
2 2915 1 927
2 2916 1 930
2 2917 1 930
2 2918 1 931
2 2919 1 931
2 2920 1 935
2 2921 1 935
2 2922 1 938
2 2923 1 938
2 2924 1 939
2 2925 1 939
2 2926 1 943
2 2927 1 943
2 2928 1 946
2 2929 1 946
2 2930 1 947
2 2931 1 947
2 2932 1 951
2 2933 1 951
2 2934 1 954
2 2935 1 954
2 2936 1 955
2 2937 1 955
2 2938 1 959
2 2939 1 959
2 2940 1 962
2 2941 1 962
2 2942 1 963
2 2943 1 963
2 2944 1 965
2 2945 1 965
2 2946 1 968
2 2947 1 968
2 2948 1 968
2 2949 1 970
2 2950 1 970
2 2951 1 970
2 2952 1 971
2 2953 1 971
2 2954 1 971
2 2955 1 972
2 2956 1 972
2 2957 1 975
2 2958 1 975
2 2959 1 976
2 2960 1 976
2 2961 1 981
2 2962 1 981
2 2963 1 981
2 2964 1 981
2 2965 1 982
2 2966 1 982
2 2967 1 982
2 2968 1 982
2 2969 1 984
2 2970 1 984
2 2971 1 987
2 2972 1 987
2 2973 1 990
2 2974 1 990
2 2975 1 993
2 2976 1 993
2 2977 1 996
2 2978 1 996
2 2979 1 999
2 2980 1 999
2 2981 1 1002
2 2982 1 1002
2 2983 1 1005
2 2984 1 1005
2 2985 1 1011
2 2986 1 1011
2 2987 1 1011
2 2988 1 1015
2 2989 1 1015
2 2990 1 1019
2 2991 1 1019
2 2992 1 1023
2 2993 1 1023
2 2994 1 1023
2 2995 1 1024
2 2996 1 1024
2 2997 1 1031
2 2998 1 1031
2 2999 1 1031
2 3000 1 1035
2 3001 1 1035
2 3002 1 1039
2 3003 1 1039
2 3004 1 1043
2 3005 1 1043
2 3006 1 1043
2 3007 1 1044
2 3008 1 1044
2 3009 1 1051
2 3010 1 1051
2 3011 1 1055
2 3012 1 1055
2 3013 1 1059
2 3014 1 1059
2 3015 1 1063
2 3016 1 1063
2 3017 1 1063
2 3018 1 1064
2 3019 1 1064
2 3020 1 1071
2 3021 1 1071
2 3022 1 1075
2 3023 1 1075
2 3024 1 1079
2 3025 1 1079
2 3026 1 1083
2 3027 1 1083
2 3028 1 1083
2 3029 1 1084
2 3030 1 1084
2 3031 1 1091
2 3032 1 1091
2 3033 1 1095
2 3034 1 1095
2 3035 1 1099
2 3036 1 1099
2 3037 1 1099
2 3038 1 1100
2 3039 1 1100
2 3040 1 1103
2 3041 1 1103
2 3042 1 1111
2 3043 1 1111
2 3044 1 1111
2 3045 1 1112
2 3046 1 1112
2 3047 1 1113
2 3048 1 1113
2 3049 1 1114
2 3050 1 1114
2 3051 1 1119
2 3052 1 1119
2 3053 1 1127
2 3054 1 1127
2 3055 1 1127
2 3056 1 1128
2 3057 1 1128
2 3058 1 1131
2 3059 1 1131
2 3060 1 1139
2 3061 1 1139
2 3062 1 1139
2 3063 1 1140
2 3064 1 1140
2 3065 1 1145
2 3066 1 1145
2 3067 1 1149
2 3068 1 1149
2 3069 1 1152
2 3070 1 1152
2 3071 1 1154
2 3072 1 1154
2 3073 1 1157
2 3074 1 1157
2 3075 1 1177
2 3076 1 1177
2 3077 1 1189
2 3078 1 1189
2 3079 1 1201
2 3080 1 1201
2 3081 1 1213
2 3082 1 1213
2 3083 1 1225
2 3084 1 1225
2 3085 1 1238
2 3086 1 1238
2 3087 1 1241
2 3088 1 1241
2 3089 1 1241
2 3090 1 1241
2 3091 1 1241
2 3092 1 1242
2 3093 1 1242
2 3094 1 1243
2 3095 1 1243
2 3096 1 1243
2 3097 1 1243
2 3098 1 1243
2 3099 1 1244
2 3100 1 1244
2 3101 1 1248
2 3102 1 1248
2 3103 1 1248
2 3104 1 1249
2 3105 1 1249
2 3106 1 1249
2 3107 1 1254
2 3108 1 1254
2 3109 1 1255
2 3110 1 1255
2 3111 1 1257
2 3112 1 1257
2 3113 1 1260
2 3114 1 1260
2 3115 1 1263
2 3116 1 1263
2 3117 1 1266
2 3118 1 1266
2 3119 1 1269
2 3120 1 1269
2 3121 1 1272
2 3122 1 1272
2 3123 1 1272
2 3124 1 1273
2 3125 1 1273
2 3126 1 1275
2 3127 1 1275
2 3128 1 1278
2 3129 1 1278
2 3130 1 1281
2 3131 1 1281
2 3132 1 1281
2 3133 1 1284
2 3134 1 1284
2 3135 1 1287
2 3136 1 1287
2 3137 1 1288
2 3138 1 1288
2 3139 1 1290
2 3140 1 1290
2 3141 1 1293
2 3142 1 1293
2 3143 1 1303
2 3144 1 1303
2 3145 1 1309
2 3146 1 1309
2 3147 1 1315
2 3148 1 1315
2 3149 1 1332
2 3150 1 1332
2 3151 1 1333
2 3152 1 1333
2 3153 1 1336
2 3154 1 1336
2 3155 1 1337
2 3156 1 1337
2 3157 1 1340
2 3158 1 1340
2 3159 1 1341
2 3160 1 1341
2 3161 1 1344
2 3162 1 1344
2 3163 1 1345
2 3164 1 1345
2 3165 1 1348
2 3166 1 1348
2 3167 1 1349
2 3168 1 1349
2 3169 1 1352
2 3170 1 1352
2 3171 1 1353
2 3172 1 1353
2 3173 1 1356
2 3174 1 1356
2 3175 1 1357
2 3176 1 1357
2 3177 1 1360
2 3178 1 1360
2 3179 1 1361
2 3180 1 1361
2 3181 1 1364
2 3182 1 1364
2 3183 1 1365
2 3184 1 1365
2 3185 1 1368
2 3186 1 1368
2 3187 1 1369
2 3188 1 1369
2 3189 1 1372
2 3190 1 1372
2 3191 1 1373
2 3192 1 1373
2 3193 1 1376
2 3194 1 1376
2 3195 1 1377
2 3196 1 1377
2 3197 1 1380
2 3198 1 1380
2 3199 1 1381
2 3200 1 1381
2 3201 1 1384
2 3202 1 1384
2 3203 1 1385
2 3204 1 1385
2 3205 1 1388
2 3206 1 1388
2 3207 1 1389
2 3208 1 1389
2 3209 1 1411
2 3210 1 1411
2 3211 1 1411
2 3212 1 1411
2 3213 1 1412
2 3214 1 1412
2 3215 1 1412
2 3216 1 1417
2 3217 1 1417
2 3218 1 1418
2 3219 1 1418
2 3220 1 1420
2 3221 1 1420
2 3222 1 1423
2 3223 1 1423
2 3224 1 1429
2 3225 1 1429
2 3226 1 1429
2 3227 1 1429
2 3228 1 1430
2 3229 1 1430
2 3230 1 1430
2 3231 1 1432
2 3232 1 1432
2 3233 1 1433
2 3234 1 1433
2 3235 1 1439
2 3236 1 1439
2 3237 1 1439
2 3238 1 1439
2 3239 1 1440
2 3240 1 1440
2 3241 1 1440
2 3242 1 1445
2 3243 1 1445
2 3244 1 1446
2 3245 1 1446
2 3246 1 1448
2 3247 1 1448
2 3248 1 1451
2 3249 1 1451
2 3250 1 1453
2 3251 1 1453
2 3252 1 1454
2 3253 1 1454
2 3254 1 1457
2 3255 1 1457
2 3256 1 1460
2 3257 1 1460
2 3258 1 1465
2 3259 1 1465
2 3260 1 1465
2 3261 1 1466
2 3262 1 1466
2 3263 1 1466
2 3264 1 1471
2 3265 1 1471
2 3266 1 1471
2 3267 1 1471
2 3268 1 1472
2 3269 1 1472
2 3270 1 1472
2 3271 1 1474
2 3272 1 1474
2 3273 1 1477
2 3274 1 1477
2 3275 1 1480
2 3276 1 1480
2 3277 1 1481
2 3278 1 1481
2 3279 1 1485
2 3280 1 1485
2 3281 1 1488
2 3282 1 1488
2 3283 1 1493
2 3284 1 1493
2 3285 1 1493
2 3286 1 1493
2 3287 1 1494
2 3288 1 1494
2 3289 1 1494
2 3290 1 1496
2 3291 1 1496
2 3292 1 1499
2 3293 1 1499
2 3294 1 1502
2 3295 1 1502
2 3296 1 1503
2 3297 1 1503
2 3298 1 1507
2 3299 1 1507
2 3300 1 1510
2 3301 1 1510
2 3302 1 1515
2 3303 1 1515
2 3304 1 1515
2 3305 1 1515
2 3306 1 1516
2 3307 1 1516
2 3308 1 1516
2 3309 1 1518
2 3310 1 1518
2 3311 1 1521
2 3312 1 1521
2 3313 1 1524
2 3314 1 1524
2 3315 1 1525
2 3316 1 1525
2 3317 1 1529
2 3318 1 1529
2 3319 1 1532
2 3320 1 1532
2 3321 1 1537
2 3322 1 1537
2 3323 1 1537
2 3324 1 1537
2 3325 1 1538
2 3326 1 1538
2 3327 1 1538
2 3328 1 1540
2 3329 1 1540
2 3330 1 1543
2 3331 1 1543
2 3332 1 1546
2 3333 1 1546
2 3334 1 1547
2 3335 1 1547
2 3336 1 1551
2 3337 1 1551
2 3338 1 1554
2 3339 1 1554
2 3340 1 1559
2 3341 1 1559
2 3342 1 1559
2 3343 1 1559
2 3344 1 1560
2 3345 1 1560
2 3346 1 1560
2 3347 1 1562
2 3348 1 1562
2 3349 1 1565
2 3350 1 1565
2 3351 1 1568
2 3352 1 1568
2 3353 1 1569
2 3354 1 1569
2 3355 1 1573
2 3356 1 1573
2 3357 1 1576
2 3358 1 1576
2 3359 1 1581
2 3360 1 1581
2 3361 1 1581
2 3362 1 1581
2 3363 1 1582
2 3364 1 1582
2 3365 1 1582
2 3366 1 1582
2 3367 1 1584
2 3368 1 1584
2 3369 1 1587
2 3370 1 1587
2 3371 1 1590
2 3372 1 1590
2 3373 1 1591
2 3374 1 1591
2 3375 1 1595
2 3376 1 1595
2 3377 1 1598
2 3378 1 1598
2 3379 1 1603
2 3380 1 1603
2 3381 1 1603
2 3382 1 1603
2 3383 1 1604
2 3384 1 1604
2 3385 1 1604
2 3386 1 1606
2 3387 1 1606
2 3388 1 1609
2 3389 1 1609
2 3390 1 1612
2 3391 1 1612
2 3392 1 1613
2 3393 1 1613
2 3394 1 1617
2 3395 1 1617
2 3396 1 1620
2 3397 1 1620
2 3398 1 1625
2 3399 1 1625
2 3400 1 1625
2 3401 1 1625
2 3402 1 1626
2 3403 1 1626
2 3404 1 1628
2 3405 1 1628
2 3406 1 1631
2 3407 1 1631
2 3408 1 1634
2 3409 1 1634
2 3410 1 1635
2 3411 1 1635
2 3412 1 1639
2 3413 1 1639
2 3414 1 1642
2 3415 1 1642
2 3416 1 1643
2 3417 1 1643
2 3418 1 1644
2 3419 1 1644
2 3420 1 1647
2 3421 1 1647
2 3422 1 1650
2 3423 1 1650
2 3424 1 1653
2 3425 1 1653
2 3426 1 1657
2 3427 1 1657
2 3428 1 1658
2 3429 1 1658
2 3430 1 1661
2 3431 1 1661
2 3432 1 1664
2 3433 1 1664
2 3434 1 1665
2 3435 1 1665
2 3436 1 1669
2 3437 1 1669
2 3438 1 1672
2 3439 1 1672
2 3440 1 1673
2 3441 1 1673
2 3442 1 1677
2 3443 1 1677
2 3444 1 1680
2 3445 1 1680
2 3446 1 1681
2 3447 1 1681
2 3448 1 1685
2 3449 1 1685
2 3450 1 1688
2 3451 1 1688
2 3452 1 1689
2 3453 1 1689
2 3454 1 1693
2 3455 1 1693
2 3456 1 1696
2 3457 1 1696
2 3458 1 1697
2 3459 1 1697
2 3460 1 1701
2 3461 1 1701
2 3462 1 1704
2 3463 1 1704
2 3464 1 1705
2 3465 1 1705
2 3466 1 1709
2 3467 1 1709
2 3468 1 1712
2 3469 1 1712
2 3470 1 1713
2 3471 1 1713
2 3472 1 1717
2 3473 1 1717
2 3474 1 1720
2 3475 1 1720
2 3476 1 1721
2 3477 1 1721
2 3478 1 1725
2 3479 1 1725
2 3480 1 1728
2 3481 1 1728
2 3482 1 1729
2 3483 1 1729
2 3484 1 1733
2 3485 1 1733
2 3486 1 1736
2 3487 1 1736
2 3488 1 1737
2 3489 1 1737
2 3490 1 1739
2 3491 1 1739
2 3492 1 1745
2 3493 1 1745
2 3494 1 1746
2 3495 1 1746
2 3496 1 1751
2 3497 1 1751
2 3498 1 1757
2 3499 1 1757
2 3500 1 1758
2 3501 1 1758
2 3502 1 1763
2 3503 1 1763
2 3504 1 1766
2 3505 1 1766
2 3506 1 1769
2 3507 1 1769
2 3508 1 1775
2 3509 1 1775
2 3510 1 1781
2 3511 1 1781
2 3512 1 1789
2 3513 1 1789
2 3514 1 1797
2 3515 1 1797
2 3516 1 1801
2 3517 1 1801
2 3518 1 1809
2 3519 1 1809
2 3520 1 1813
2 3521 1 1813
2 3522 1 1821
2 3523 1 1821
2 3524 1 1825
2 3525 1 1825
2 3526 1 1831
2 3527 1 1831
2 3528 1 1832
2 3529 1 1832
2 3530 1 1837
2 3531 1 1837
2 3532 1 1845
2 3533 1 1845
2 3534 1 1873
2 3535 1 1873
2 3536 1 1885
2 3537 1 1885
2 3538 1 1897
2 3539 1 1897
2 3540 1 1912
2 3541 1 1912
0 50 5 1 1 49
0 51 5 1 1 1953
0 52 5 1 1 1955
0 53 5 1 1 1957
0 54 5 1 1 1959
0 55 5 1 1 1961
0 56 5 1 1 1963
0 57 5 1 1 1965
0 58 5 1 1 1967
0 59 5 1 1 1969
0 60 5 1 1 1971
0 61 5 1 1 1973
0 62 5 1 1 1975
0 63 5 1 1 1977
0 64 5 1 1 1979
0 65 5 1 1 1981
0 66 5 1 1 1983
0 67 5 1 1 1985
0 68 5 1 1 1987
0 69 5 2 1 1989
0 70 5 2 1 1991
0 71 5 2 1 1993
0 72 5 2 1 1995
0 73 5 2 1 1997
0 74 5 2 1 1999
0 75 5 2 1 2001
0 76 5 2 1 2003
0 77 5 2 1 2005
0 78 5 2 1 2007
0 79 5 2 1 2009
0 80 5 2 1 2011
0 81 5 1 1 2013
0 82 5 1 1 2015
0 83 5 1 1 2017
0 84 5 1 1 2019
0 85 5 1 1 2021
0 86 5 1 1 2023
0 87 5 1 1 2025
0 88 5 1 1 2027
0 89 5 1 1 2029
0 90 5 1 1 2031
0 91 5 1 1 2033
0 92 5 1 1 2035
0 93 5 1 1 2037
0 94 5 1 1 2039
0 95 5 1 1 2041
0 96 5 1 1 2043
0 97 5 1 1 2045
0 98 5 1 1 2047
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 1956 1988
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 1954 1986
0 106 5 2 1 105
0 107 7 2 2 1952 1984
0 108 5 3 1 2081
0 109 7 1 2 2079 2083
0 110 5 1 1 109
0 111 7 2 2 2077 110
0 112 5 2 1 2086
0 113 7 1 2 2075 2088
0 114 5 1 1 113
0 115 7 2 2 2073 114
0 116 5 1 1 2090
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 1958 2091
0 120 5 2 1 119
0 121 7 1 2 2049 2094
0 122 5 1 1 121
0 123 7 2 2 2092 122
0 124 5 1 1 2096
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 1960 2097
0 128 5 2 1 127
0 129 7 1 2 2051 2100
0 130 5 1 1 129
0 131 7 2 2 2098 130
0 132 5 1 1 2102
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 1962 2103
0 136 5 2 1 135
0 137 7 1 2 2053 2106
0 138 5 1 1 137
0 139 7 2 2 2104 138
0 140 5 1 1 2108
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 1964 2109
0 144 5 2 1 143
0 145 7 1 2 2055 2112
0 146 5 1 1 145
0 147 7 2 2 2110 146
0 148 5 1 1 2114
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 1966 2115
0 152 5 2 1 151
0 153 7 1 2 2057 2118
0 154 5 1 1 153
0 155 7 2 2 2116 154
0 156 5 1 1 2120
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 1968 2121
0 160 5 2 1 159
0 161 7 1 2 2059 2124
0 162 5 1 1 161
0 163 7 2 2 2122 162
0 164 5 1 1 2126
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 1970 2127
0 168 5 2 1 167
0 169 7 1 2 2061 2130
0 170 5 1 1 169
0 171 7 2 2 2128 170
0 172 5 1 1 2132
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 1972 2133
0 176 5 2 1 175
0 177 7 1 2 2063 2136
0 178 5 1 1 177
0 179 7 2 2 2134 178
0 180 5 1 1 2138
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 1974 2139
0 184 5 2 1 183
0 185 7 1 2 2065 2142
0 186 5 1 1 185
0 187 7 2 2 2140 186
0 188 5 1 1 2144
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 1976 2145
0 192 5 2 1 191
0 193 7 1 2 2067 2148
0 194 5 1 1 193
0 195 7 2 2 2146 194
0 196 5 1 1 2150
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 1978 2151
0 200 5 2 1 199
0 201 7 1 2 2069 2154
0 202 5 1 1 201
0 203 7 2 2 2152 202
0 204 5 1 1 2156
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 1980 2157
0 208 5 2 1 207
0 209 7 1 2 2071 2160
0 210 5 1 1 209
0 211 7 3 2 2158 210
0 212 5 3 1 2162
0 213 7 2 2 1982 2014
0 214 5 2 1 2168
0 215 7 1 2 2163 2169
0 216 5 2 1 215
0 217 7 2 2 2159 2161
0 218 5 1 1 2174
0 219 7 1 2 2012 2175
0 220 5 1 1 219
0 221 7 1 2 2072 218
0 222 5 1 1 221
0 223 7 4 2 220 222
0 224 5 3 1 2176
0 225 7 2 2 65 81
0 226 5 2 1 2183
0 227 7 2 2 2170 2185
0 228 5 1 1 2187
0 229 7 1 2 2164 228
0 230 5 1 1 229
0 231 7 1 2 2165 2188
0 232 5 1 1 231
0 233 7 3 2 230 232
0 234 5 2 1 2189
0 235 7 1 2 2177 2192
0 236 5 2 1 235
0 237 7 2 2 2153 2155
0 238 5 1 1 2196
0 239 7 1 2 2010 2197
0 240 5 1 1 239
0 241 7 1 2 2070 238
0 242 5 1 1 241
0 243 7 4 2 240 242
0 244 5 3 1 2198
0 245 7 1 2 2178 2199
0 246 5 2 1 245
0 247 7 2 2 2147 2149
0 248 5 1 1 2207
0 249 7 1 2 2008 2208
0 250 5 1 1 249
0 251 7 1 2 2068 248
0 252 5 1 1 251
0 253 7 4 2 250 252
0 254 5 3 1 2209
0 255 7 1 2 2200 2210
0 256 5 2 1 255
0 257 7 2 2 2141 2143
0 258 5 1 1 2218
0 259 7 1 2 2006 2219
0 260 5 1 1 259
0 261 7 1 2 2066 258
0 262 5 1 1 261
0 263 7 4 2 260 262
0 264 5 3 1 2220
0 265 7 1 2 2211 2221
0 266 5 2 1 265
0 267 7 2 2 2135 2137
0 268 5 1 1 2229
0 269 7 1 2 2004 2230
0 270 5 1 1 269
0 271 7 1 2 2064 268
0 272 5 1 1 271
0 273 7 4 2 270 272
0 274 5 3 1 2231
0 275 7 1 2 2222 2232
0 276 5 2 1 275
0 277 7 2 2 2129 2131
0 278 5 1 1 2240
0 279 7 1 2 2002 2241
0 280 5 1 1 279
0 281 7 1 2 2062 278
0 282 5 1 1 281
0 283 7 4 2 280 282
0 284 5 3 1 2242
0 285 7 1 2 2233 2243
0 286 5 2 1 285
0 287 7 2 2 2123 2125
0 288 5 1 1 2251
0 289 7 1 2 2000 2252
0 290 5 1 1 289
0 291 7 1 2 2060 288
0 292 5 1 1 291
0 293 7 4 2 290 292
0 294 5 3 1 2253
0 295 7 1 2 2244 2254
0 296 5 2 1 295
0 297 7 2 2 2117 2119
0 298 5 1 1 2262
0 299 7 1 2 1998 2263
0 300 5 1 1 299
0 301 7 1 2 2058 298
0 302 5 1 1 301
0 303 7 4 2 300 302
0 304 5 3 1 2264
0 305 7 1 2 2255 2265
0 306 5 2 1 305
0 307 7 2 2 2111 2113
0 308 5 1 1 2273
0 309 7 1 2 1996 2274
0 310 5 1 1 309
0 311 7 1 2 2056 308
0 312 5 1 1 311
0 313 7 4 2 310 312
0 314 5 3 1 2275
0 315 7 1 2 2266 2276
0 316 5 2 1 315
0 317 7 2 2 2105 2107
0 318 5 1 1 2284
0 319 7 1 2 1994 2285
0 320 5 1 1 319
0 321 7 1 2 2054 318
0 322 5 1 1 321
0 323 7 4 2 320 322
0 324 5 3 1 2286
0 325 7 1 2 2277 2287
0 326 5 2 1 325
0 327 7 2 2 2099 2101
0 328 5 1 1 2295
0 329 7 1 2 1992 2296
0 330 5 1 1 329
0 331 7 1 2 2052 328
0 332 5 1 1 331
0 333 7 4 2 330 332
0 334 5 3 1 2297
0 335 7 1 2 2288 2298
0 336 5 2 1 335
0 337 7 2 2 2093 2095
0 338 5 1 1 2306
0 339 7 1 2 1990 2307
0 340 5 1 1 339
0 341 7 1 2 2050 338
0 342 5 1 1 341
0 343 7 4 2 340 342
0 344 5 3 1 2308
0 345 7 1 2 2299 2309
0 346 5 2 1 345
0 347 7 2 2 2074 2076
0 348 5 1 1 2317
0 349 7 1 2 2087 348
0 350 5 1 1 349
0 351 7 1 2 2089 2318
0 352 5 1 1 351
0 353 7 4 2 350 352
0 354 5 2 1 2319
0 355 7 1 2 2310 2323
0 356 5 2 1 355
0 357 7 1 2 50 66
0 358 5 1 1 357
0 359 7 2 2 2084 358
0 360 5 2 1 2327
0 361 7 1 2 2320 2329
0 362 5 1 1 361
0 363 7 2 2 2078 2080
0 364 5 1 1 2331
0 365 7 1 2 2082 364
0 366 5 1 1 365
0 367 7 1 2 2085 2332
0 368 5 1 1 367
0 369 7 2 2 366 368
0 370 5 2 1 2333
0 371 7 2 2 362 2335
0 372 5 1 1 2337
0 373 7 1 2 2312 2321
0 374 5 1 1 373
0 375 7 2 2 2325 374
0 376 5 1 1 2339
0 377 7 1 2 2338 2340
0 378 5 2 1 377
0 379 7 2 2 2326 2341
0 380 5 1 1 2343
0 381 7 1 2 2301 2313
0 382 5 1 1 381
0 383 7 2 2 2315 382
0 384 5 1 1 2345
0 385 7 1 2 380 2346
0 386 5 2 1 385
0 387 7 2 2 2316 2347
0 388 5 1 1 2349
0 389 7 1 2 2290 2302
0 390 5 1 1 389
0 391 7 2 2 2304 390
0 392 5 1 1 2351
0 393 7 1 2 388 2352
0 394 5 2 1 393
0 395 7 2 2 2305 2353
0 396 5 1 1 2355
0 397 7 1 2 2279 2291
0 398 5 1 1 397
0 399 7 2 2 2293 398
0 400 5 1 1 2357
0 401 7 1 2 396 2358
0 402 5 2 1 401
0 403 7 2 2 2294 2359
0 404 5 1 1 2361
0 405 7 1 2 2268 2280
0 406 5 1 1 405
0 407 7 2 2 2282 406
0 408 5 1 1 2363
0 409 7 1 2 404 2364
0 410 5 2 1 409
0 411 7 2 2 2283 2365
0 412 5 1 1 2367
0 413 7 1 2 2257 2269
0 414 5 1 1 413
0 415 7 2 2 2271 414
0 416 5 1 1 2369
0 417 7 1 2 412 2370
0 418 5 2 1 417
0 419 7 2 2 2272 2371
0 420 5 1 1 2373
0 421 7 1 2 2246 2258
0 422 5 1 1 421
0 423 7 2 2 2260 422
0 424 5 1 1 2375
0 425 7 1 2 420 2376
0 426 5 2 1 425
0 427 7 2 2 2261 2377
0 428 5 1 1 2379
0 429 7 1 2 2235 2247
0 430 5 1 1 429
0 431 7 2 2 2249 430
0 432 5 1 1 2381
0 433 7 1 2 428 2382
0 434 5 2 1 433
0 435 7 2 2 2250 2383
0 436 5 1 1 2385
0 437 7 1 2 2224 2236
0 438 5 1 1 437
0 439 7 2 2 2238 438
0 440 5 1 1 2387
0 441 7 1 2 436 2388
0 442 5 2 1 441
0 443 7 2 2 2239 2389
0 444 5 1 1 2391
0 445 7 1 2 2213 2225
0 446 5 1 1 445
0 447 7 2 2 2227 446
0 448 5 1 1 2393
0 449 7 1 2 444 2394
0 450 5 2 1 449
0 451 7 2 2 2228 2395
0 452 5 1 1 2397
0 453 7 1 2 2202 2214
0 454 5 1 1 453
0 455 7 2 2 2216 454
0 456 5 1 1 2399
0 457 7 1 2 452 2400
0 458 5 2 1 457
0 459 7 2 2 2217 2401
0 460 5 1 1 2403
0 461 7 1 2 2180 2203
0 462 5 1 1 461
0 463 7 2 2 2205 462
0 464 5 1 1 2405
0 465 7 1 2 460 2406
0 466 5 2 1 465
0 467 7 2 2 2206 2407
0 468 5 1 1 2409
0 469 7 1 2 2181 2190
0 470 5 1 1 469
0 471 7 2 2 2194 470
0 472 5 1 1 2411
0 473 7 1 2 468 2412
0 474 5 2 1 473
0 475 7 2 2 2195 2413
0 476 5 1 1 2415
0 477 7 1 2 2166 2184
0 478 5 1 1 477
0 479 7 2 2 2172 478
0 480 5 1 1 2417
0 481 7 2 2 476 2418
0 482 5 2 1 2419
0 483 7 1 2 2167 2171
0 484 5 1 1 483
0 485 7 3 2 2186 484
0 486 5 2 1 2423
0 487 7 1 2 2420 2424
0 488 5 1 1 487
0 489 7 4 2 2173 488
0 490 5 2 1 2428
0 491 7 1 2 90 2256
0 492 5 3 1 491
0 493 7 1 2 2032 2259
0 494 5 3 1 493
0 495 7 1 2 89 2267
0 496 5 3 1 495
0 497 7 1 2 2030 2270
0 498 5 3 1 497
0 499 7 1 2 88 2278
0 500 5 3 1 499
0 501 7 1 2 2028 2281
0 502 5 3 1 501
0 503 7 1 2 87 2289
0 504 5 3 1 503
0 505 7 1 2 2026 2292
0 506 5 3 1 505
0 507 7 1 2 86 2300
0 508 5 3 1 507
0 509 7 1 2 2024 2303
0 510 5 3 1 509
0 511 7 1 2 85 2311
0 512 5 3 1 511
0 513 7 1 2 2022 2314
0 514 5 3 1 513
0 515 7 1 2 84 2324
0 516 5 3 1 515
0 517 7 1 2 2020 2322
0 518 5 3 1 517
0 519 7 1 2 83 2336
0 520 5 3 1 519
0 521 7 1 2 2018 2334
0 522 5 3 1 521
0 523 7 3 2 82 2328
0 524 5 2 1 2482
0 525 7 1 2 2479 2483
0 526 5 1 1 525
0 527 7 2 2 2476 526
0 528 5 2 1 2487
0 529 7 1 2 2473 2489
0 530 5 1 1 529
0 531 7 2 2 2470 530
0 532 5 2 1 2491
0 533 7 1 2 2467 2493
0 534 5 1 1 533
0 535 7 2 2 2464 534
0 536 5 2 1 2495
0 537 7 1 2 2461 2497
0 538 5 1 1 537
0 539 7 2 2 2458 538
0 540 5 2 1 2499
0 541 7 1 2 2455 2501
0 542 5 1 1 541
0 543 7 2 2 2452 542
0 544 5 2 1 2503
0 545 7 1 2 2449 2505
0 546 5 1 1 545
0 547 7 2 2 2446 546
0 548 5 2 1 2507
0 549 7 1 2 2443 2509
0 550 5 1 1 549
0 551 7 2 2 2440 550
0 552 5 2 1 2511
0 553 7 1 2 2437 2513
0 554 5 1 1 553
0 555 7 2 2 2434 554
0 556 5 2 1 2515
0 557 7 1 2 91 2245
0 558 5 3 1 557
0 559 7 1 2 2034 2248
0 560 5 3 1 559
0 561 7 3 2 2519 2522
0 562 5 2 1 2525
0 563 7 1 2 2517 2526
0 564 5 1 1 563
0 565 7 1 2 2516 2528
0 566 5 1 1 565
0 567 7 4 2 564 566
0 568 5 3 1 2530
0 569 7 1 2 2042 2204
0 570 5 3 1 569
0 571 7 1 2 95 2201
0 572 5 3 1 571
0 573 7 3 2 2537 2540
0 574 5 2 1 2543
0 575 7 1 2 94 2212
0 576 5 3 1 575
0 577 7 1 2 2040 2215
0 578 5 3 1 577
0 579 7 1 2 93 2223
0 580 5 3 1 579
0 581 7 1 2 2038 2226
0 582 5 3 1 581
0 583 7 1 2 92 2234
0 584 5 3 1 583
0 585 7 1 2 2036 2237
0 586 5 3 1 585
0 587 7 1 2 2523 2518
0 588 5 1 1 587
0 589 7 2 2 2520 588
0 590 5 2 1 2566
0 591 7 1 2 2563 2568
0 592 5 1 1 591
0 593 7 2 2 2560 592
0 594 5 2 1 2570
0 595 7 1 2 2557 2572
0 596 5 1 1 595
0 597 7 2 2 2554 596
0 598 5 2 1 2574
0 599 7 1 2 2551 2576
0 600 5 1 1 599
0 601 7 2 2 2548 600
0 602 5 2 1 2578
0 603 7 1 2 2544 2579
0 604 5 1 1 603
0 605 7 1 2 2546 2580
0 606 5 1 1 605
0 607 7 4 2 604 606
0 608 5 4 1 2582
0 609 7 1 2 2534 2583
0 610 5 2 1 609
0 611 7 1 2 2531 2586
0 612 5 1 1 611
0 613 7 2 2 2590 612
0 614 5 1 1 2592
0 615 7 3 2 2561 2564
0 616 5 2 1 2594
0 617 7 1 2 2569 2595
0 618 5 1 1 617
0 619 7 1 2 2567 2597
0 620 5 1 1 619
0 621 7 4 2 618 620
0 622 5 3 1 2599
0 623 7 1 2 2593 2603
0 624 5 2 1 623
0 625 7 2 2 2591 2606
0 626 5 1 1 2608
0 627 7 3 2 2555 2558
0 628 5 2 1 2610
0 629 7 1 2 2571 2613
0 630 5 1 1 629
0 631 7 1 2 2573 2611
0 632 5 1 1 631
0 633 7 4 2 630 632
0 634 5 3 1 2615
0 635 7 1 2 2044 2182
0 636 5 3 1 635
0 637 7 1 2 96 2179
0 638 5 3 1 637
0 639 7 3 2 2622 2625
0 640 5 2 1 2628
0 641 7 1 2 2538 2581
0 642 5 1 1 641
0 643 7 2 2 2541 642
0 644 5 2 1 2633
0 645 7 1 2 2629 2634
0 646 5 1 1 645
0 647 7 1 2 2631 2635
0 648 5 1 1 647
0 649 7 4 2 646 648
0 650 5 3 1 2637
0 651 7 1 2 2604 2638
0 652 5 2 1 651
0 653 7 1 2 2600 2641
0 654 5 1 1 653
0 655 7 2 2 2644 654
0 656 5 1 1 2646
0 657 7 1 2 2619 2647
0 658 5 2 1 657
0 659 7 1 2 2616 656
0 660 5 1 1 659
0 661 7 2 2 2648 660
0 662 5 1 1 2650
0 663 7 1 2 626 2651
0 664 5 2 1 663
0 665 7 3 2 2552 2549
0 666 5 2 1 2654
0 667 7 1 2 2657 2575
0 668 5 1 1 667
0 669 7 1 2 2655 2577
0 670 5 1 1 669
0 671 7 4 2 668 670
0 672 5 3 1 2659
0 673 7 3 2 2435 2438
0 674 5 2 1 2666
0 675 7 1 2 2512 2669
0 676 5 1 1 675
0 677 7 1 2 2514 2667
0 678 5 1 1 677
0 679 7 4 2 676 678
0 680 5 3 1 2671
0 681 7 1 2 2663 2675
0 682 5 2 1 681
0 683 7 1 2 2660 2672
0 684 5 1 1 683
0 685 7 2 2 2678 684
0 686 5 1 1 2680
0 687 7 1 2 2681 2535
0 688 5 2 1 687
0 689 7 2 2 2679 2682
0 690 5 1 1 2684
0 691 7 1 2 614 2601
0 692 5 1 1 691
0 693 7 2 2 2607 692
0 694 5 1 1 2686
0 695 7 1 2 690 2687
0 696 5 2 1 695
0 697 7 3 2 2441 2444
0 698 5 2 1 2690
0 699 7 1 2 2508 2693
0 700 5 1 1 699
0 701 7 1 2 2510 2691
0 702 5 1 1 701
0 703 7 4 2 700 702
0 704 5 3 1 2695
0 705 7 1 2 2620 2699
0 706 5 2 1 705
0 707 7 1 2 2617 2696
0 708 5 1 1 707
0 709 7 2 2 2702 708
0 710 5 1 1 2704
0 711 7 1 2 2676 2705
0 712 5 2 1 711
0 713 7 2 2 2703 2706
0 714 5 1 1 2708
0 715 7 1 2 686 2532
0 716 5 1 1 715
0 717 7 2 2 2683 716
0 718 5 1 1 2710
0 719 7 1 2 714 2711
0 720 5 2 1 719
0 721 7 3 2 2447 2450
0 722 5 2 1 2714
0 723 7 1 2 2504 2717
0 724 5 1 1 723
0 725 7 1 2 2506 2715
0 726 5 1 1 725
0 727 7 4 2 724 726
0 728 5 3 1 2719
0 729 7 1 2 2605 2723
0 730 5 2 1 729
0 731 7 1 2 2602 2720
0 732 5 1 1 731
0 733 7 2 2 2726 732
0 734 5 1 1 2728
0 735 7 1 2 2700 2729
0 736 5 2 1 735
0 737 7 2 2 2727 2730
0 738 5 1 1 2732
0 739 7 1 2 2673 710
0 740 5 1 1 739
0 741 7 2 2 2707 740
0 742 5 1 1 2734
0 743 7 1 2 738 2735
0 744 5 2 1 743
0 745 7 3 2 2453 2456
0 746 5 2 1 2738
0 747 7 1 2 2500 2741
0 748 5 1 1 747
0 749 7 1 2 2502 2739
0 750 5 1 1 749
0 751 7 4 2 748 750
0 752 5 3 1 2743
0 753 7 1 2 2536 2747
0 754 5 2 1 753
0 755 7 1 2 2533 2744
0 756 5 1 1 755
0 757 7 2 2 2750 756
0 758 5 1 1 2752
0 759 7 1 2 2724 2753
0 760 5 2 1 759
0 761 7 2 2 2751 2754
0 762 5 1 1 2756
0 763 7 1 2 2697 734
0 764 5 1 1 763
0 765 7 2 2 2731 764
0 766 5 1 1 2758
0 767 7 1 2 762 2759
0 768 5 2 1 767
0 769 7 3 2 2459 2462
0 770 5 2 1 2762
0 771 7 1 2 2496 2765
0 772 5 1 1 771
0 773 7 1 2 2498 2763
0 774 5 1 1 773
0 775 7 4 2 772 774
0 776 5 3 1 2767
0 777 7 1 2 2677 2771
0 778 5 2 1 777
0 779 7 1 2 2674 2768
0 780 5 1 1 779
0 781 7 2 2 2774 780
0 782 5 1 1 2776
0 783 7 1 2 2748 2777
0 784 5 2 1 783
0 785 7 2 2 2775 2778
0 786 5 1 1 2780
0 787 7 1 2 2721 758
0 788 5 1 1 787
0 789 7 2 2 2755 788
0 790 5 1 1 2782
0 791 7 1 2 786 2783
0 792 5 2 1 791
0 793 7 3 2 2465 2468
0 794 5 2 1 2786
0 795 7 1 2 2492 2789
0 796 5 1 1 795
0 797 7 1 2 2494 2787
0 798 5 1 1 797
0 799 7 5 2 796 798
0 800 5 3 1 2791
0 801 7 1 2 2701 2796
0 802 5 2 1 801
0 803 7 1 2 2698 2792
0 804 5 1 1 803
0 805 7 2 2 2799 804
0 806 5 1 1 2801
0 807 7 1 2 2772 2802
0 808 5 2 1 807
0 809 7 2 2 2800 2803
0 810 5 1 1 2805
0 811 7 1 2 2745 782
0 812 5 1 1 811
0 813 7 2 2 2779 812
0 814 5 1 1 2807
0 815 7 1 2 810 2808
0 816 5 2 1 815
0 817 7 3 2 2471 2474
0 818 5 2 1 2811
0 819 7 1 2 2488 2814
0 820 5 1 1 819
0 821 7 1 2 2490 2812
0 822 5 1 1 821
0 823 7 4 2 820 822
0 824 5 2 1 2816
0 825 7 1 2 2725 2820
0 826 5 2 1 825
0 827 7 1 2 2722 2817
0 828 5 1 1 827
0 829 7 2 2 2822 828
0 830 5 1 1 2824
0 831 7 1 2 2797 2825
0 832 5 2 1 831
0 833 7 2 2 2823 2826
0 834 5 1 1 2828
0 835 7 1 2 2769 806
0 836 5 1 1 835
0 837 7 2 2 2804 836
0 838 5 1 1 2830
0 839 7 1 2 834 2831
0 840 5 2 1 839
0 841 7 3 2 2477 2480
0 842 5 2 1 2834
0 843 7 1 2 2485 2835
0 844 5 1 1 843
0 845 7 1 2 2484 2837
0 846 5 1 1 845
0 847 7 4 2 844 846
0 848 5 2 1 2839
0 849 7 1 2 2749 2840
0 850 5 2 1 849
0 851 7 1 2 2746 2843
0 852 5 1 1 851
0 853 7 2 2 2845 852
0 854 5 1 1 2847
0 855 7 1 2 2821 2848
0 856 5 2 1 855
0 857 7 2 2 2846 2849
0 858 5 1 1 2851
0 859 7 1 2 2793 830
0 860 5 1 1 859
0 861 7 2 2 2827 860
0 862 5 1 1 2853
0 863 7 1 2 858 2854
0 864 5 2 1 863
0 865 7 2 2 2773 2841
0 866 5 2 1 2857
0 867 7 1 2 2818 854
0 868 5 1 1 867
0 869 7 2 2 2850 868
0 870 5 1 1 2861
0 871 7 1 2 2858 2862
0 872 5 2 1 871
0 873 7 1 2 2859 870
0 874 5 1 1 873
0 875 7 2 2 2863 874
0 876 5 1 1 2865
0 877 7 2 2 2016 2330
0 878 5 3 1 2867
0 879 7 3 2 2486 2869
0 880 5 5 1 2872
0 881 7 1 2 2770 2844
0 882 5 1 1 881
0 883 7 2 2 2860 882
0 884 5 2 1 2880
0 885 7 1 2 2794 2882
0 886 5 1 1 885
0 887 7 2 2 2875 886
0 888 5 1 1 2884
0 889 7 1 2 2866 2885
0 890 5 2 1 889
0 891 7 2 2 2864 2886
0 892 5 1 1 2888
0 893 7 1 2 2852 862
0 894 5 1 1 893
0 895 7 2 2 2855 894
0 896 5 1 1 2890
0 897 7 1 2 892 2891
0 898 5 2 1 897
0 899 7 2 2 2856 2892
0 900 5 1 1 2894
0 901 7 1 2 2829 838
0 902 5 1 1 901
0 903 7 2 2 2832 902
0 904 5 1 1 2896
0 905 7 1 2 900 2897
0 906 5 2 1 905
0 907 7 2 2 2833 2898
0 908 5 1 1 2900
0 909 7 1 2 2806 814
0 910 5 1 1 909
0 911 7 2 2 2809 910
0 912 5 1 1 2902
0 913 7 1 2 908 2903
0 914 5 2 1 913
0 915 7 2 2 2810 2904
0 916 5 1 1 2906
0 917 7 1 2 2781 790
0 918 5 1 1 917
0 919 7 2 2 2784 918
0 920 5 1 1 2908
0 921 7 1 2 916 2909
0 922 5 2 1 921
0 923 7 2 2 2785 2910
0 924 5 1 1 2912
0 925 7 1 2 2757 766
0 926 5 1 1 925
0 927 7 2 2 2760 926
0 928 5 1 1 2914
0 929 7 1 2 924 2915
0 930 5 2 1 929
0 931 7 2 2 2761 2916
0 932 5 1 1 2918
0 933 7 1 2 2733 742
0 934 5 1 1 933
0 935 7 2 2 2736 934
0 936 5 1 1 2920
0 937 7 1 2 932 2921
0 938 5 2 1 937
0 939 7 2 2 2737 2922
0 940 5 1 1 2924
0 941 7 1 2 2709 718
0 942 5 1 1 941
0 943 7 2 2 2712 942
0 944 5 1 1 2926
0 945 7 1 2 940 2927
0 946 5 2 1 945
0 947 7 2 2 2713 2928
0 948 5 1 1 2930
0 949 7 1 2 2685 694
0 950 5 1 1 949
0 951 7 2 2 2688 950
0 952 5 1 1 2932
0 953 7 1 2 948 2933
0 954 5 2 1 953
0 955 7 2 2 2689 2934
0 956 5 1 1 2936
0 957 7 1 2 2609 662
0 958 5 1 1 957
0 959 7 2 2 2652 958
0 960 5 1 1 2938
0 961 7 1 2 956 2939
0 962 5 2 1 961
0 963 7 2 2 2653 2940
0 964 5 1 1 2942
0 965 7 2 2 2645 2649
0 966 5 1 1 2944
0 967 7 1 2 2046 2191
0 968 5 3 1 967
0 969 7 1 2 97 2193
0 970 5 3 1 969
0 971 7 3 2 2946 2949
0 972 5 2 1 2952
0 973 7 1 2 2623 2636
0 974 5 1 1 973
0 975 7 2 2 2626 974
0 976 5 2 1 2957
0 977 7 1 2 2953 2959
0 978 5 1 1 977
0 979 7 1 2 2955 2958
0 980 5 1 1 979
0 981 7 4 2 978 980
0 982 5 4 1 2961
0 983 7 1 2 2621 2965
0 984 5 2 1 983
0 985 7 1 2 2618 2962
0 986 5 1 1 985
0 987 7 2 2 2969 986
0 988 5 1 1 2971
0 989 7 1 2 2664 2972
0 990 5 2 1 989
0 991 7 1 2 2661 988
0 992 5 1 1 991
0 993 7 2 2 2973 992
0 994 5 1 1 2975
0 995 7 1 2 966 2976
0 996 5 2 1 995
0 997 7 1 2 2945 994
0 998 5 1 1 997
0 999 7 2 2 2977 998
0 1000 5 1 1 2979
0 1001 7 1 2 964 2980
0 1002 5 2 1 1001
0 1003 7 1 2 2943 1000
0 1004 5 1 1 1003
0 1005 7 2 2 2981 1004
0 1006 5 1 1 2983
0 1007 7 1 2 2432 1006
0 1008 5 1 1 1007
0 1009 7 1 2 2421 2426
0 1010 5 1 1 1009
0 1011 7 3 2 2429 1010
0 1012 5 1 1 2985
0 1013 7 1 2 2937 960
0 1014 5 1 1 1013
0 1015 7 2 2 2941 1014
0 1016 5 1 1 2988
0 1017 7 1 2 2931 952
0 1018 5 1 1 1017
0 1019 7 2 2 2935 1018
0 1020 5 1 1 2990
0 1021 7 1 2 2416 480
0 1022 5 1 1 1021
0 1023 7 3 2 2422 1022
0 1024 5 2 1 2992
0 1025 7 1 2 1020 2993
0 1026 5 1 1 1025
0 1027 7 1 2 2991 2995
0 1028 5 1 1 1027
0 1029 7 1 2 2410 472
0 1030 5 1 1 1029
0 1031 7 3 2 2414 1030
0 1032 5 1 1 2997
0 1033 7 1 2 2925 944
0 1034 5 1 1 1033
0 1035 7 2 2 2929 1034
0 1036 5 1 1 3000
0 1037 7 1 2 2919 936
0 1038 5 1 1 1037
0 1039 7 2 2 2923 1038
0 1040 5 1 1 3002
0 1041 7 1 2 2404 464
0 1042 5 1 1 1041
0 1043 7 3 2 2408 1042
0 1044 5 2 1 3004
0 1045 7 1 2 1040 3005
0 1046 5 1 1 1045
0 1047 7 1 2 3003 3007
0 1048 5 1 1 1047
0 1049 7 1 2 2398 456
0 1050 5 1 1 1049
0 1051 7 2 2 2402 1050
0 1052 5 1 1 3009
0 1053 7 1 2 2913 928
0 1054 5 1 1 1053
0 1055 7 2 2 2917 1054
0 1056 5 1 1 3011
0 1057 7 1 2 2907 920
0 1058 5 1 1 1057
0 1059 7 2 2 2911 1058
0 1060 5 1 1 3013
0 1061 7 1 2 2392 448
0 1062 5 1 1 1061
0 1063 7 3 2 2396 1062
0 1064 5 2 1 3015
0 1065 7 1 2 1060 3016
0 1066 5 1 1 1065
0 1067 7 1 2 3014 3018
0 1068 5 1 1 1067
0 1069 7 1 2 2386 440
0 1070 5 1 1 1069
0 1071 7 2 2 2390 1070
0 1072 5 1 1 3020
0 1073 7 1 2 2901 912
0 1074 5 1 1 1073
0 1075 7 2 2 2905 1074
0 1076 5 1 1 3022
0 1077 7 1 2 2895 904
0 1078 5 1 1 1077
0 1079 7 2 2 2899 1078
0 1080 5 1 1 3024
0 1081 7 1 2 2380 432
0 1082 5 1 1 1081
0 1083 7 3 2 2384 1082
0 1084 5 2 1 3026
0 1085 7 1 2 1080 3027
0 1086 5 1 1 1085
0 1087 7 1 2 3025 3029
0 1088 5 1 1 1087
0 1089 7 1 2 2374 424
0 1090 5 1 1 1089
0 1091 7 2 2 2378 1090
0 1092 5 1 1 3031
0 1093 7 1 2 2889 896
0 1094 5 1 1 1093
0 1095 7 2 2 2893 1094
0 1096 5 1 1 3033
0 1097 7 1 2 2368 416
0 1098 5 1 1 1097
0 1099 7 3 2 2372 1098
0 1100 5 2 1 3035
0 1101 7 1 2 876 888
0 1102 5 1 1 1101
0 1103 7 2 2 2887 1102
0 1104 5 1 1 3040
0 1105 7 1 2 3036 1104
0 1106 5 1 1 1105
0 1107 7 1 2 3038 3041
0 1108 5 1 1 1107
0 1109 7 1 2 2362 408
0 1110 5 1 1 1109
0 1111 7 3 2 2366 1110
0 1112 5 2 1 3042
0 1113 7 2 2 2795 2876
0 1114 5 2 1 3047
0 1115 7 1 2 2881 3049
0 1116 5 1 1 1115
0 1117 7 1 2 2883 3048
0 1118 5 1 1 1117
0 1119 7 2 2 1116 1118
0 1120 5 1 1 3051
0 1121 7 1 2 3043 3052
0 1122 5 1 1 1121
0 1123 7 1 2 3045 1120
0 1124 5 1 1 1123
0 1125 7 1 2 2356 400
0 1126 5 1 1 1125
0 1127 7 3 2 2360 1126
0 1128 5 2 1 3053
0 1129 7 1 2 2798 2873
0 1130 5 1 1 1129
0 1131 7 2 2 3050 1130
0 1132 5 1 1 3058
0 1133 7 1 2 3054 3059
0 1134 5 1 1 1133
0 1135 7 1 2 3056 1132
0 1136 5 1 1 1135
0 1137 7 1 2 2350 392
0 1138 5 1 1 1137
0 1139 7 3 2 2354 1138
0 1140 5 2 1 3060
0 1141 7 1 2 372 376
0 1142 5 1 1 1141
0 1143 7 1 2 2342 1142
0 1144 5 1 1 1143
0 1145 7 2 2 2877 1144
0 1146 5 1 1 3065
0 1147 7 1 2 2344 384
0 1148 5 1 1 1147
0 1149 7 2 2 2348 1148
0 1150 5 1 1 3067
0 1151 7 1 2 3066 1150
0 1152 5 2 1 1151
0 1153 7 1 2 1146 3068
0 1154 5 2 1 1153
0 1155 7 1 2 2842 3071
0 1156 5 1 1 1155
0 1157 7 2 2 3069 1156
0 1158 5 1 1 3073
0 1159 7 1 2 3063 1158
0 1160 5 1 1 1159
0 1161 7 1 2 2819 1160
0 1162 5 1 1 1161
0 1163 7 1 2 3061 3074
0 1164 5 1 1 1163
0 1165 7 1 2 1162 1164
0 1166 5 1 1 1165
0 1167 7 1 2 1136 1166
0 1168 5 1 1 1167
0 1169 7 1 2 1134 1168
0 1170 5 1 1 1169
0 1171 7 1 2 1124 1170
0 1172 5 1 1 1171
0 1173 7 1 2 1122 1172
0 1174 5 1 1 1173
0 1175 7 1 2 1108 1174
0 1176 5 1 1 1175
0 1177 7 2 2 1106 1176
0 1178 5 1 1 3075
0 1179 7 1 2 3034 3076
0 1180 5 1 1 1179
0 1181 7 1 2 3032 1180
0 1182 5 1 1 1181
0 1183 7 1 2 1096 1178
0 1184 5 1 1 1183
0 1185 7 1 2 1182 1184
0 1186 5 1 1 1185
0 1187 7 1 2 1088 1186
0 1188 5 1 1 1187
0 1189 7 2 2 1086 1188
0 1190 5 1 1 3077
0 1191 7 1 2 3023 3078
0 1192 5 1 1 1191
0 1193 7 1 2 3021 1192
0 1194 5 1 1 1193
0 1195 7 1 2 1076 1190
0 1196 5 1 1 1195
0 1197 7 1 2 1194 1196
0 1198 5 1 1 1197
0 1199 7 1 2 1068 1198
0 1200 5 1 1 1199
0 1201 7 2 2 1066 1200
0 1202 5 1 1 3079
0 1203 7 1 2 3012 3080
0 1204 5 1 1 1203
0 1205 7 1 2 3010 1204
0 1206 5 1 1 1205
0 1207 7 1 2 1056 1202
0 1208 5 1 1 1207
0 1209 7 1 2 1206 1208
0 1210 5 1 1 1209
0 1211 7 1 2 1048 1210
0 1212 5 1 1 1211
0 1213 7 2 2 1046 1212
0 1214 5 1 1 3081
0 1215 7 1 2 3001 3082
0 1216 5 1 1 1215
0 1217 7 1 2 2998 1216
0 1218 5 1 1 1217
0 1219 7 1 2 1036 1214
0 1220 5 1 1 1219
0 1221 7 1 2 1218 1220
0 1222 5 1 1 1221
0 1223 7 1 2 1028 1222
0 1224 5 1 1 1223
0 1225 7 2 2 1026 1224
0 1226 5 1 1 3083
0 1227 7 1 2 2989 3084
0 1228 5 1 1 1227
0 1229 7 1 2 2986 1228
0 1230 5 1 1 1229
0 1231 7 1 2 1016 1226
0 1232 5 1 1 1231
0 1233 7 1 2 1230 1232
0 1234 7 1 2 1008 1233
0 1235 5 1 1 1234
0 1236 7 1 2 2430 2984
0 1237 5 1 1 1236
0 1238 7 2 2 2970 2974
0 1239 5 1 1 3085
0 1240 7 1 2 2048 2427
0 1241 5 5 1 1240
0 1242 7 2 2 98 2425
0 1243 5 5 1 3092
0 1244 7 2 2 3087 3094
0 1245 5 1 1 3099
0 1246 7 1 2 2947 2960
0 1247 5 1 1 1246
0 1248 7 3 2 2950 1247
0 1249 5 3 1 3101
0 1250 7 1 2 3100 3104
0 1251 5 1 1 1250
0 1252 7 1 2 1245 3102
0 1253 5 1 1 1252
0 1254 7 2 2 1251 1253
0 1255 5 2 1 3107
0 1256 7 1 2 2665 3109
0 1257 5 2 1 1256
0 1258 7 1 2 2662 3108
0 1259 5 1 1 1258
0 1260 7 2 2 3111 1259
0 1261 5 1 1 3113
0 1262 7 1 2 2584 3114
0 1263 5 2 1 1262
0 1264 7 1 2 2587 1261
0 1265 5 1 1 1264
0 1266 7 2 2 3115 1265
0 1267 5 1 1 3117
0 1268 7 1 2 1239 3118
0 1269 5 2 1 1268
0 1270 7 1 2 3088 3105
0 1271 5 1 1 1270
0 1272 7 3 2 3095 1271
0 1273 5 2 1 3121
0 1274 7 1 2 2966 3124
0 1275 5 2 1 1274
0 1276 7 1 2 2963 3122
0 1277 5 1 1 1276
0 1278 7 2 2 3126 1277
0 1279 5 1 1 3128
0 1280 7 1 2 2639 3129
0 1281 5 3 1 1280
0 1282 7 1 2 2642 1279
0 1283 5 1 1 1282
0 1284 7 2 2 3130 1283
0 1285 5 1 1 3133
0 1286 7 1 2 2640 3125
0 1287 5 2 1 1286
0 1288 7 2 2 2643 3123
0 1289 5 1 1 3137
0 1290 7 2 2 1289 3135
0 1291 5 1 1 3139
0 1292 7 1 2 2585 3140
0 1293 5 2 1 1292
0 1294 7 1 2 3136 3141
0 1295 5 1 1 1294
0 1296 7 1 2 3134 1295
0 1297 5 1 1 1296
0 1298 7 1 2 3119 1297
0 1299 7 1 2 3089 3103
0 1300 5 1 1 1299
0 1301 7 1 2 3096 3106
0 1302 5 1 1 1301
0 1303 7 2 2 1300 1302
0 1304 5 1 1 3143
0 1305 7 1 2 2964 3144
0 1306 5 1 1 1305
0 1307 7 1 2 2967 1304
0 1308 5 1 1 1307
0 1309 7 2 2 1306 1308
0 1310 5 1 1 3145
0 1311 7 1 2 3127 3131
0 1312 5 1 1 1311
0 1313 7 1 2 1310 1312
0 1314 5 1 1 1313
0 1315 7 2 2 3112 3116
0 1316 5 1 1 3147
0 1317 7 1 2 2588 1291
0 1318 5 1 1 1317
0 1319 7 1 2 3142 1318
0 1320 7 1 2 1316 1319
0 1321 5 1 1 1320
0 1322 7 1 2 1314 1321
0 1323 7 1 2 1298 1322
0 1324 7 1 2 3086 1267
0 1325 5 1 1 1324
0 1326 7 1 2 3120 1325
0 1327 5 1 1 1326
0 1328 7 1 2 2968 3110
0 1329 5 1 1 1328
0 1330 7 1 2 2481 2870
0 1331 5 1 1 1330
0 1332 7 2 2 2478 1331
0 1333 5 2 1 3149
0 1334 7 1 2 2475 3151
0 1335 5 1 1 1334
0 1336 7 2 2 2472 1335
0 1337 5 2 1 3153
0 1338 7 1 2 2469 3155
0 1339 5 1 1 1338
0 1340 7 2 2 2466 1339
0 1341 5 2 1 3157
0 1342 7 1 2 2463 3159
0 1343 5 1 1 1342
0 1344 7 2 2 2460 1343
0 1345 5 2 1 3161
0 1346 7 1 2 2457 3163
0 1347 5 1 1 1346
0 1348 7 2 2 2454 1347
0 1349 5 2 1 3165
0 1350 7 1 2 2451 3167
0 1351 5 1 1 1350
0 1352 7 2 2 2448 1351
0 1353 5 2 1 3169
0 1354 7 1 2 2445 3171
0 1355 5 1 1 1354
0 1356 7 2 2 2442 1355
0 1357 5 2 1 3173
0 1358 7 1 2 2439 3175
0 1359 5 1 1 1358
0 1360 7 2 2 2436 1359
0 1361 5 2 1 3177
0 1362 7 1 2 2524 3179
0 1363 5 1 1 1362
0 1364 7 2 2 2521 1363
0 1365 5 2 1 3181
0 1366 7 1 2 2565 3183
0 1367 5 1 1 1366
0 1368 7 2 2 2562 1367
0 1369 5 2 1 3185
0 1370 7 1 2 2559 3187
0 1371 5 1 1 1370
0 1372 7 2 2 2556 1371
0 1373 5 2 1 3189
0 1374 7 1 2 2553 3191
0 1375 5 1 1 1374
0 1376 7 2 2 2550 1375
0 1377 5 2 1 3193
0 1378 7 1 2 2539 3195
0 1379 5 1 1 1378
0 1380 7 2 2 2542 1379
0 1381 5 2 1 3197
0 1382 7 1 2 2624 3199
0 1383 5 1 1 1382
0 1384 7 2 2 2627 1383
0 1385 5 2 1 3201
0 1386 7 1 2 2948 3203
0 1387 5 1 1 1386
0 1388 7 2 2 2951 1387
0 1389 5 2 1 3205
0 1390 7 1 2 3090 3207
0 1391 5 1 1 1390
0 1392 7 1 2 2589 3097
0 1393 7 1 2 1391 1392
0 1394 7 1 2 3138 1393
0 1395 7 1 2 1329 1394
0 1396 7 1 2 3146 1395
0 1397 7 1 2 2978 3132
0 1398 7 1 2 1396 1397
0 1399 7 1 2 1285 3148
0 1400 7 1 2 1398 1399
0 1401 7 1 2 2982 1400
0 1402 7 1 2 1327 1401
0 1403 7 1 2 1323 1402
0 1404 7 1 2 1237 1403
0 1405 7 1 2 1235 1404
0 1406 5 1 1 1405
0 1407 7 1 2 2527 3180
0 1408 5 1 1 1407
0 1409 7 1 2 2529 3178
0 1410 5 1 1 1409
0 1411 7 4 2 1408 1410
0 1412 5 3 1 3209
0 1413 7 1 2 2547 3194
0 1414 5 1 1 1413
0 1415 7 1 2 2545 3196
0 1416 5 1 1 1415
0 1417 7 2 2 1414 1416
0 1418 5 2 1 3216
0 1419 7 1 2 3210 3217
0 1420 5 2 1 1419
0 1421 7 1 2 3213 3218
0 1422 5 1 1 1421
0 1423 7 2 2 3220 1422
0 1424 5 1 1 3222
0 1425 7 1 2 2596 3184
0 1426 5 1 1 1425
0 1427 7 1 2 2598 3182
0 1428 5 1 1 1427
0 1429 7 4 2 1426 1428
0 1430 5 3 1 3224
0 1431 7 1 2 3223 3225
0 1432 5 2 1 1431
0 1433 7 2 2 3221 3231
0 1434 5 1 1 3233
0 1435 7 1 2 2614 3186
0 1436 5 1 1 1435
0 1437 7 1 2 2612 3188
0 1438 5 1 1 1437
0 1439 7 4 2 1436 1438
0 1440 5 3 1 3235
0 1441 7 1 2 2630 3200
0 1442 5 1 1 1441
0 1443 7 1 2 2632 3198
0 1444 5 1 1 1443
0 1445 7 2 2 1442 1444
0 1446 5 2 1 3242
0 1447 7 1 2 3226 3243
0 1448 5 2 1 1447
0 1449 7 1 2 3228 3244
0 1450 5 1 1 1449
0 1451 7 2 2 3246 1450
0 1452 5 1 1 3248
0 1453 7 2 2 3236 3249
0 1454 5 2 1 3250
0 1455 7 1 2 3239 1452
0 1456 5 1 1 1455
0 1457 7 2 2 3252 1456
0 1458 5 1 1 3254
0 1459 7 1 2 1434 3255
0 1460 5 2 1 1459
0 1461 7 1 2 2658 3190
0 1462 5 1 1 1461
0 1463 7 1 2 2656 3192
0 1464 5 1 1 1463
0 1465 7 3 2 1462 1464
0 1466 5 3 1 3258
0 1467 7 1 2 2670 3174
0 1468 5 1 1 1467
0 1469 7 1 2 2668 3176
0 1470 5 1 1 1469
0 1471 7 4 2 1468 1470
0 1472 5 3 1 3264
0 1473 7 1 2 3259 3265
0 1474 5 2 1 1473
0 1475 7 1 2 3261 3268
0 1476 5 1 1 1475
0 1477 7 2 2 3271 1476
0 1478 5 1 1 3273
0 1479 7 1 2 3274 3211
0 1480 5 2 1 1479
0 1481 7 2 2 3272 3275
0 1482 5 1 1 3277
0 1483 7 1 2 1424 3229
0 1484 5 1 1 1483
0 1485 7 2 2 3232 1484
0 1486 5 1 1 3279
0 1487 7 1 2 1482 3280
0 1488 5 2 1 1487
0 1489 7 1 2 2694 3170
0 1490 5 1 1 1489
0 1491 7 1 2 2692 3172
0 1492 5 1 1 1491
0 1493 7 4 2 1490 1492
0 1494 5 3 1 3283
0 1495 7 1 2 3237 3284
0 1496 5 2 1 1495
0 1497 7 1 2 3240 3287
0 1498 5 1 1 1497
0 1499 7 2 2 3290 1498
0 1500 5 1 1 3292
0 1501 7 1 2 3266 3293
0 1502 5 2 1 1501
0 1503 7 2 2 3291 3294
0 1504 5 1 1 3296
0 1505 7 1 2 1478 3214
0 1506 5 1 1 1505
0 1507 7 2 2 3276 1506
0 1508 5 1 1 3298
0 1509 7 1 2 1504 3299
0 1510 5 2 1 1509
0 1511 7 1 2 2718 3166
0 1512 5 1 1 1511
0 1513 7 1 2 2716 3168
0 1514 5 1 1 1513
0 1515 7 4 2 1512 1514
0 1516 5 3 1 3302
0 1517 7 1 2 3227 3303
0 1518 5 2 1 1517
0 1519 7 1 2 3230 3306
0 1520 5 1 1 1519
0 1521 7 2 2 3309 1520
0 1522 5 1 1 3311
0 1523 7 1 2 3285 3312
0 1524 5 2 1 1523
0 1525 7 2 2 3310 3313
0 1526 5 1 1 3315
0 1527 7 1 2 3269 1500
0 1528 5 1 1 1527
0 1529 7 2 2 3295 1528
0 1530 5 1 1 3317
0 1531 7 1 2 1526 3318
0 1532 5 2 1 1531
0 1533 7 1 2 2742 3162
0 1534 5 1 1 1533
0 1535 7 1 2 2740 3164
0 1536 5 1 1 1535
0 1537 7 4 2 1534 1536
0 1538 5 3 1 3321
0 1539 7 1 2 3212 3322
0 1540 5 2 1 1539
0 1541 7 1 2 3215 3325
0 1542 5 1 1 1541
0 1543 7 2 2 3328 1542
0 1544 5 1 1 3330
0 1545 7 1 2 3304 3331
0 1546 5 2 1 1545
0 1547 7 2 2 3329 3332
0 1548 5 1 1 3334
0 1549 7 1 2 3288 1522
0 1550 5 1 1 1549
0 1551 7 2 2 3314 1550
0 1552 5 1 1 3336
0 1553 7 1 2 1548 3337
0 1554 5 2 1 1553
0 1555 7 1 2 2766 3158
0 1556 5 1 1 1555
0 1557 7 1 2 2764 3160
0 1558 5 1 1 1557
0 1559 7 4 2 1556 1558
0 1560 5 3 1 3340
0 1561 7 1 2 3267 3341
0 1562 5 2 1 1561
0 1563 7 1 2 3270 3344
0 1564 5 1 1 1563
0 1565 7 2 2 3347 1564
0 1566 5 1 1 3349
0 1567 7 1 2 3323 3350
0 1568 5 2 1 1567
0 1569 7 2 2 3348 3351
0 1570 5 1 1 3353
0 1571 7 1 2 3307 1544
0 1572 5 1 1 1571
0 1573 7 2 2 3333 1572
0 1574 5 1 1 3355
0 1575 7 1 2 1570 3356
0 1576 5 2 1 1575
0 1577 7 1 2 2790 3154
0 1578 5 1 1 1577
0 1579 7 1 2 2788 3156
0 1580 5 1 1 1579
0 1581 7 4 2 1578 1580
0 1582 5 4 1 3359
0 1583 7 1 2 3286 3360
0 1584 5 2 1 1583
0 1585 7 1 2 3289 3363
0 1586 5 1 1 1585
0 1587 7 2 2 3367 1586
0 1588 5 1 1 3369
0 1589 7 1 2 3342 3370
0 1590 5 2 1 1589
0 1591 7 2 2 3368 3371
0 1592 5 1 1 3373
0 1593 7 1 2 3326 1566
0 1594 5 1 1 1593
0 1595 7 2 2 3352 1594
0 1596 5 1 1 3375
0 1597 7 1 2 1592 3376
0 1598 5 2 1 1597
0 1599 7 1 2 2813 3152
0 1600 5 1 1 1599
0 1601 7 1 2 2815 3150
0 1602 5 1 1 1601
0 1603 7 4 2 1600 1602
0 1604 5 3 1 3379
0 1605 7 1 2 3305 3380
0 1606 5 2 1 1605
0 1607 7 1 2 3308 3383
0 1608 5 1 1 1607
0 1609 7 2 2 3386 1608
0 1610 5 1 1 3388
0 1611 7 1 2 3361 3389
0 1612 5 2 1 1611
0 1613 7 2 2 3387 3390
0 1614 5 1 1 3392
0 1615 7 1 2 3345 1588
0 1616 5 1 1 1615
0 1617 7 2 2 3372 1616
0 1618 5 1 1 3394
0 1619 7 1 2 1614 3395
0 1620 5 2 1 1619
0 1621 7 1 2 2836 2871
0 1622 5 1 1 1621
0 1623 7 1 2 2838 2868
0 1624 5 1 1 1623
0 1625 7 4 2 1622 1624
0 1626 5 2 1 3398
0 1627 7 1 2 3324 3399
0 1628 5 2 1 1627
0 1629 7 1 2 3327 3402
0 1630 5 1 1 1629
0 1631 7 2 2 3404 1630
0 1632 5 1 1 3406
0 1633 7 1 2 3381 3407
0 1634 5 2 1 1633
0 1635 7 2 2 3405 3408
0 1636 5 1 1 3410
0 1637 7 1 2 3364 1610
0 1638 5 1 1 1637
0 1639 7 2 2 3391 1638
0 1640 5 1 1 3412
0 1641 7 1 2 1636 3413
0 1642 5 2 1 1641
0 1643 7 2 2 3343 3400
0 1644 5 2 1 3416
0 1645 7 1 2 3384 1632
0 1646 5 1 1 1645
0 1647 7 2 2 3409 1646
0 1648 5 1 1 3420
0 1649 7 1 2 3417 3421
0 1650 5 2 1 1649
0 1651 7 1 2 3418 1648
0 1652 5 1 1 1651
0 1653 7 2 2 3422 1652
0 1654 5 1 1 3424
0 1655 7 1 2 3346 3403
0 1656 5 1 1 1655
0 1657 7 2 2 3419 1656
0 1658 5 2 1 3426
0 1659 7 1 2 3365 3428
0 1660 5 1 1 1659
0 1661 7 2 2 2878 1660
0 1662 5 1 1 3430
0 1663 7 1 2 3425 3431
0 1664 5 2 1 1663
0 1665 7 2 2 3423 3432
0 1666 5 1 1 3434
0 1667 7 1 2 3411 1640
0 1668 5 1 1 1667
0 1669 7 2 2 3414 1668
0 1670 5 1 1 3436
0 1671 7 1 2 1666 3437
0 1672 5 2 1 1671
0 1673 7 2 2 3415 3438
0 1674 5 1 1 3440
0 1675 7 1 2 3393 1618
0 1676 5 1 1 1675
0 1677 7 2 2 3396 1676
0 1678 5 1 1 3442
0 1679 7 1 2 1674 3443
0 1680 5 2 1 1679
0 1681 7 2 2 3397 3444
0 1682 5 1 1 3446
0 1683 7 1 2 3374 1596
0 1684 5 1 1 1683
0 1685 7 2 2 3377 1684
0 1686 5 1 1 3448
0 1687 7 1 2 1682 3449
0 1688 5 2 1 1687
0 1689 7 2 2 3378 3450
0 1690 5 1 1 3452
0 1691 7 1 2 3354 1574
0 1692 5 1 1 1691
0 1693 7 2 2 3357 1692
0 1694 5 1 1 3454
0 1695 7 1 2 1690 3455
0 1696 5 2 1 1695
0 1697 7 2 2 3358 3456
0 1698 5 1 1 3458
0 1699 7 1 2 3335 1552
0 1700 5 1 1 1699
0 1701 7 2 2 3338 1700
0 1702 5 1 1 3460
0 1703 7 1 2 1698 3461
0 1704 5 2 1 1703
0 1705 7 2 2 3339 3462
0 1706 5 1 1 3464
0 1707 7 1 2 3316 1530
0 1708 5 1 1 1707
0 1709 7 2 2 3319 1708
0 1710 5 1 1 3466
0 1711 7 1 2 1706 3467
0 1712 5 2 1 1711
0 1713 7 2 2 3320 3468
0 1714 5 1 1 3470
0 1715 7 1 2 3297 1508
0 1716 5 1 1 1715
0 1717 7 2 2 3300 1716
0 1718 5 1 1 3472
0 1719 7 1 2 1714 3473
0 1720 5 2 1 1719
0 1721 7 2 2 3301 3474
0 1722 5 1 1 3476
0 1723 7 1 2 3278 1486
0 1724 5 1 1 1723
0 1725 7 2 2 3281 1724
0 1726 5 1 1 3478
0 1727 7 1 2 1722 3479
0 1728 5 2 1 1727
0 1729 7 2 2 3282 3480
0 1730 5 1 1 3482
0 1731 7 1 2 3234 1458
0 1732 5 1 1 1731
0 1733 7 2 2 3256 1732
0 1734 5 1 1 3484
0 1735 7 1 2 1730 3485
0 1736 5 2 1 1735
0 1737 7 2 2 3257 3486
0 1738 5 1 1 3488
0 1739 7 2 2 3247 3253
0 1740 5 1 1 3490
0 1741 7 1 2 2954 3204
0 1742 5 1 1 1741
0 1743 7 1 2 2956 3202
0 1744 5 1 1 1743
0 1745 7 2 2 1742 1744
0 1746 5 2 1 3492
0 1747 7 1 2 3262 3238
0 1748 5 1 1 1747
0 1749 7 1 2 3260 3241
0 1750 5 1 1 1749
0 1751 7 2 2 1748 1750
0 1752 5 1 1 3496
0 1753 7 1 2 3493 3497
0 1754 5 1 1 1753
0 1755 7 1 2 3494 1752
0 1756 5 1 1 1755
0 1757 7 2 2 1754 1756
0 1758 5 2 1 3498
0 1759 7 1 2 3491 3500
0 1760 5 1 1 1759
0 1761 7 1 2 1740 3499
0 1762 5 1 1 1761
0 1763 7 2 2 1760 1762
0 1764 5 1 1 3502
0 1765 7 1 2 1738 1764
0 1766 5 2 1 1765
0 1767 7 1 2 3489 3503
0 1768 5 1 1 1767
0 1769 7 2 2 3504 1768
0 1770 5 1 1 3506
0 1771 7 1 2 2433 1770
0 1772 5 1 1 1771
0 1773 7 1 2 3483 1734
0 1774 5 1 1 1773
0 1775 7 2 2 3487 1774
0 1776 5 1 1 3508
0 1777 7 1 2 1012 3509
0 1778 5 1 1 1777
0 1779 7 1 2 3471 1718
0 1780 5 1 1 1779
0 1781 7 2 2 3475 1780
0 1782 5 1 1 3510
0 1783 7 1 2 2999 1782
0 1784 5 1 1 1783
0 1785 7 1 2 1032 3511
0 1786 5 1 1 1785
0 1787 7 1 2 3465 1710
0 1788 5 1 1 1787
0 1789 7 2 2 3469 1788
0 1790 5 1 1 3512
0 1791 7 1 2 3006 1790
0 1792 5 1 1 1791
0 1793 7 1 2 3008 3513
0 1794 5 1 1 1793
0 1795 7 1 2 3459 1702
0 1796 5 1 1 1795
0 1797 7 2 2 3463 1796
0 1798 5 1 1 3514
0 1799 7 1 2 3453 1694
0 1800 5 1 1 1799
0 1801 7 2 2 3457 1800
0 1802 5 1 1 3516
0 1803 7 1 2 3019 3517
0 1804 5 1 1 1803
0 1805 7 1 2 3017 1802
0 1806 5 1 1 1805
0 1807 7 1 2 3447 1686
0 1808 5 1 1 1807
0 1809 7 2 2 3451 1808
0 1810 5 1 1 3518
0 1811 7 1 2 3441 1678
0 1812 5 1 1 1811
0 1813 7 2 2 3445 1812
0 1814 5 1 1 3520
0 1815 7 1 2 3030 3521
0 1816 5 1 1 1815
0 1817 7 1 2 3028 1814
0 1818 5 1 1 1817
0 1819 7 1 2 3435 1670
0 1820 5 1 1 1819
0 1821 7 2 2 3439 1820
0 1822 5 1 1 3522
0 1823 7 1 2 1654 1662
0 1824 5 1 1 1823
0 1825 7 2 2 3433 1824
0 1826 5 1 1 3524
0 1827 7 1 2 3039 3525
0 1828 5 1 1 1827
0 1829 7 1 2 3037 1826
0 1830 5 1 1 1829
0 1831 7 2 2 2879 3366
0 1832 5 2 1 3526
0 1833 7 1 2 3427 3528
0 1834 5 1 1 1833
0 1835 7 1 2 3429 3527
0 1836 5 1 1 1835
0 1837 7 2 2 1834 1836
0 1838 5 1 1 3530
0 1839 7 1 2 3046 1838
0 1840 5 1 1 1839
0 1841 7 1 2 3044 3531
0 1842 5 1 1 1841
0 1843 7 1 2 2874 3362
0 1844 5 1 1 1843
0 1845 7 2 2 3529 1844
0 1846 5 1 1 3532
0 1847 7 1 2 3057 1846
0 1848 5 1 1 1847
0 1849 7 1 2 3055 3533
0 1850 5 1 1 1849
0 1851 7 1 2 3064 3382
0 1852 5 1 1 1851
0 1853 7 1 2 3062 3385
0 1854 5 1 1 1853
0 1855 7 1 2 3072 3401
0 1856 5 1 1 1855
0 1857 7 1 2 3070 1856
0 1858 5 1 1 1857
0 1859 7 1 2 1854 1858
0 1860 5 1 1 1859
0 1861 7 1 2 1852 1860
0 1862 5 1 1 1861
0 1863 7 1 2 1850 1862
0 1864 5 1 1 1863
0 1865 7 1 2 1848 1864
0 1866 5 1 1 1865
0 1867 7 1 2 1842 1866
0 1868 5 1 1 1867
0 1869 7 1 2 1840 1868
0 1870 5 1 1 1869
0 1871 7 1 2 1830 1870
0 1872 5 1 1 1871
0 1873 7 2 2 1828 1872
0 1874 5 1 1 3534
0 1875 7 1 2 3523 1874
0 1876 5 1 1 1875
0 1877 7 1 2 1822 3535
0 1878 5 1 1 1877
0 1879 7 1 2 1092 1878
0 1880 5 1 1 1879
0 1881 7 1 2 1876 1880
0 1882 5 1 1 1881
0 1883 7 1 2 1818 1882
0 1884 5 1 1 1883
0 1885 7 2 2 1816 1884
0 1886 5 1 1 3536
0 1887 7 1 2 3519 1886
0 1888 5 1 1 1887
0 1889 7 1 2 1810 3537
0 1890 5 1 1 1889
0 1891 7 1 2 1072 1890
0 1892 5 1 1 1891
0 1893 7 1 2 1888 1892
0 1894 5 1 1 1893
0 1895 7 1 2 1806 1894
0 1896 5 1 1 1895
0 1897 7 2 2 1804 1896
0 1898 5 1 1 3538
0 1899 7 1 2 3515 1898
0 1900 5 1 1 1899
0 1901 7 1 2 1798 3539
0 1902 5 1 1 1901
0 1903 7 1 2 1052 1902
0 1904 5 1 1 1903
0 1905 7 1 2 1900 1904
0 1906 7 1 2 1794 1905
0 1907 5 1 1 1906
0 1908 7 1 2 1792 1907
0 1909 5 1 1 1908
0 1910 7 1 2 1786 1909
0 1911 5 1 1 1910
0 1912 7 2 2 1784 1911
0 1913 5 1 1 3540
0 1914 7 1 2 2996 3541
0 1915 5 1 1 1914
0 1916 7 1 2 2994 1913
0 1917 5 1 1 1916
0 1918 7 1 2 3477 1726
0 1919 5 1 1 1918
0 1920 7 1 2 3481 1919
0 1921 7 1 2 1917 1920
0 1922 5 1 1 1921
0 1923 7 1 2 1915 1922
0 1924 7 1 2 1778 1923
0 1925 5 1 1 1924
0 1926 7 1 2 2987 1776
0 1927 5 1 1 1926
0 1928 7 1 2 1925 1927
0 1929 7 1 2 1772 1928
0 1930 5 1 1 1929
0 1931 7 1 2 2431 3507
0 1932 5 1 1 1931
0 1933 7 1 2 3251 3501
0 1934 5 1 1 1933
0 1935 7 1 2 3098 3208
0 1936 5 1 1 1935
0 1937 7 1 2 3093 3206
0 1938 5 1 1 1937
0 1939 7 1 2 1936 1938
0 1940 5 1 1 1939
0 1941 7 1 2 3263 3219
0 1942 7 1 2 3091 1941
0 1943 7 1 2 3245 1942
0 1944 7 1 2 3495 1943
0 1945 7 1 2 1940 1944
0 1946 7 1 2 1934 1945
0 1947 7 1 2 3505 1946
0 1948 7 1 2 1932 1947
0 1949 7 1 2 1930 1948
0 1950 5 1 1 1949
0 1951 7 1 2 1406 1950
3 3999 5 0 1 1951
