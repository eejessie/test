1 0 0 2 0
2 97 1 0
2 1479 1 0
1 1 0 2 0
2 1480 1 1
2 1481 1 1
1 2 0 2 0
2 1482 1 2
2 1483 1 2
1 3 0 2 0
2 1484 1 3
2 1485 1 3
1 4 0 2 0
2 1486 1 4
2 1487 1 4
1 5 0 2 0
2 1488 1 5
2 1489 1 5
1 6 0 2 0
2 1490 1 6
2 1491 1 6
1 7 0 2 0
2 1492 1 7
2 1493 1 7
1 8 0 2 0
2 1494 1 8
2 1495 1 8
1 9 0 2 0
2 1496 1 9
2 1497 1 9
1 10 0 2 0
2 1498 1 10
2 1499 1 10
1 11 0 2 0
2 1500 1 11
2 1501 1 11
1 12 0 2 0
2 1502 1 12
2 1503 1 12
1 13 0 2 0
2 1504 1 13
2 1505 1 13
1 14 0 2 0
2 1506 1 14
2 1507 1 14
1 15 0 2 0
2 1508 1 15
2 1509 1 15
1 16 0 2 0
2 1510 1 16
2 1511 1 16
1 17 0 2 0
2 1512 1 17
2 1513 1 17
1 18 0 2 0
2 1514 1 18
2 1515 1 18
1 19 0 2 0
2 1516 1 19
2 1517 1 19
1 20 0 2 0
2 1518 1 20
2 1519 1 20
1 21 0 2 0
2 1520 1 21
2 1521 1 21
1 22 0 2 0
2 1522 1 22
2 1523 1 22
1 23 0 2 0
2 1524 1 23
2 1525 1 23
1 24 0 2 0
2 1526 1 24
2 1527 1 24
1 25 0 2 0
2 1528 1 25
2 1529 1 25
1 26 0 2 0
2 1530 1 26
2 1531 1 26
1 27 0 2 0
2 1532 1 27
2 1533 1 27
1 28 0 2 0
2 1534 1 28
2 1535 1 28
1 29 0 2 0
2 1536 1 29
2 1537 1 29
1 30 0 2 0
2 1538 1 30
2 1539 1 30
1 31 0 2 0
2 1540 1 31
2 1541 1 31
1 32 0 2 0
2 1542 1 32
2 1543 1 32
1 33 0 2 0
2 1544 1 33
2 1545 1 33
1 34 0 2 0
2 1546 1 34
2 1547 1 34
1 35 0 2 0
2 1548 1 35
2 1549 1 35
1 36 0 2 0
2 1550 1 36
2 1551 1 36
1 37 0 2 0
2 1552 1 37
2 1553 1 37
1 38 0 2 0
2 1554 1 38
2 1555 1 38
1 39 0 2 0
2 1556 1 39
2 1557 1 39
1 40 0 2 0
2 1558 1 40
2 1559 1 40
1 41 0 2 0
2 1560 1 41
2 1561 1 41
1 42 0 2 0
2 1562 1 42
2 1563 1 42
1 43 0 2 0
2 1564 1 43
2 1565 1 43
1 44 0 2 0
2 1566 1 44
2 1567 1 44
1 45 0 2 0
2 1568 1 45
2 1569 1 45
1 46 0 2 0
2 1570 1 46
2 1571 1 46
1 47 0 2 0
2 1572 1 47
2 1573 1 47
1 48 0 2 0
2 1574 1 48
2 1575 1 48
1 49 0 2 0
2 1576 1 49
2 1577 1 49
1 50 0 2 0
2 1578 1 50
2 1579 1 50
1 51 0 2 0
2 1580 1 51
2 1581 1 51
1 52 0 2 0
2 1582 1 52
2 1583 1 52
1 53 0 2 0
2 1584 1 53
2 1585 1 53
1 54 0 2 0
2 1586 1 54
2 1587 1 54
1 55 0 2 0
2 1588 1 55
2 1589 1 55
1 56 0 2 0
2 1590 1 56
2 1591 1 56
1 57 0 2 0
2 1592 1 57
2 1593 1 57
1 58 0 2 0
2 1594 1 58
2 1595 1 58
1 59 0 2 0
2 1596 1 59
2 1597 1 59
1 60 0 2 0
2 1598 1 60
2 1599 1 60
1 61 0 2 0
2 1600 1 61
2 1601 1 61
1 62 0 2 0
2 1602 1 62
2 1603 1 62
1 63 0 2 0
2 1604 1 63
2 1605 1 63
1 64 0 2 0
2 1606 1 64
2 1607 1 64
1 65 0 2 0
2 1608 1 65
2 1609 1 65
1 66 0 2 0
2 1610 1 66
2 1611 1 66
1 67 0 2 0
2 1612 1 67
2 1613 1 67
1 68 0 2 0
2 1614 1 68
2 1615 1 68
1 69 0 2 0
2 1616 1 69
2 1617 1 69
1 70 0 2 0
2 1618 1 70
2 1619 1 70
1 71 0 2 0
2 1620 1 71
2 1621 1 71
1 72 0 2 0
2 1622 1 72
2 1623 1 72
1 73 0 2 0
2 1624 1 73
2 1625 1 73
1 74 0 2 0
2 1626 1 74
2 1627 1 74
1 75 0 2 0
2 1628 1 75
2 1629 1 75
1 76 0 2 0
2 1630 1 76
2 1631 1 76
1 77 0 2 0
2 1632 1 77
2 1633 1 77
1 78 0 2 0
2 1634 1 78
2 1635 1 78
1 79 0 2 0
2 1636 1 79
2 1637 1 79
1 80 0 2 0
2 1638 1 80
2 1639 1 80
1 81 0 2 0
2 1640 1 81
2 1641 1 81
1 82 0 2 0
2 1642 1 82
2 1643 1 82
1 83 0 2 0
2 1644 1 83
2 1645 1 83
1 84 0 2 0
2 1646 1 84
2 1647 1 84
1 85 0 2 0
2 1648 1 85
2 1649 1 85
1 86 0 2 0
2 1650 1 86
2 1651 1 86
1 87 0 2 0
2 1652 1 87
2 1653 1 87
1 88 0 2 0
2 1654 1 88
2 1655 1 88
1 89 0 2 0
2 1656 1 89
2 1657 1 89
1 90 0 2 0
2 1658 1 90
2 1659 1 90
1 91 0 2 0
2 1660 1 91
2 1661 1 91
1 92 0 2 0
2 1662 1 92
2 1663 1 92
1 93 0 2 0
2 1664 1 93
2 1665 1 93
1 94 0 2 0
2 1666 1 94
2 1667 1 94
1 95 0 2 0
2 1668 1 95
2 1669 1 95
1 96 0 2 0
2 1670 1 96
2 1671 1 96
2 1672 1 133
2 1673 1 133
2 1674 1 134
2 1675 1 134
2 1676 1 135
2 1677 1 135
2 1678 1 136
2 1679 1 136
2 1680 1 137
2 1681 1 137
2 1682 1 138
2 1683 1 138
2 1684 1 139
2 1685 1 139
2 1686 1 140
2 1687 1 140
2 1688 1 141
2 1689 1 141
2 1690 1 142
2 1691 1 142
2 1692 1 143
2 1693 1 143
2 1694 1 144
2 1695 1 144
2 1696 1 145
2 1697 1 145
2 1698 1 146
2 1699 1 146
2 1700 1 147
2 1701 1 147
2 1702 1 148
2 1703 1 148
2 1704 1 149
2 1705 1 149
2 1706 1 150
2 1707 1 150
2 1708 1 151
2 1709 1 151
2 1710 1 152
2 1711 1 152
2 1712 1 153
2 1713 1 153
2 1714 1 154
2 1715 1 154
2 1716 1 155
2 1717 1 155
2 1718 1 156
2 1719 1 156
2 1720 1 157
2 1721 1 157
2 1722 1 158
2 1723 1 158
2 1724 1 159
2 1725 1 159
2 1726 1 160
2 1727 1 160
2 1728 1 196
2 1729 1 196
2 1730 1 196
2 1731 1 198
2 1732 1 198
2 1733 1 200
2 1734 1 200
2 1735 1 202
2 1736 1 202
2 1737 1 204
2 1738 1 204
2 1739 1 206
2 1740 1 206
2 1741 1 207
2 1742 1 207
2 1743 1 208
2 1744 1 208
2 1745 1 208
2 1746 1 211
2 1747 1 211
2 1748 1 212
2 1749 1 212
2 1750 1 215
2 1751 1 215
2 1752 1 218
2 1753 1 218
2 1754 1 220
2 1755 1 220
2 1756 1 223
2 1757 1 223
2 1758 1 226
2 1759 1 226
2 1760 1 228
2 1761 1 228
2 1762 1 231
2 1763 1 231
2 1764 1 234
2 1765 1 234
2 1766 1 236
2 1767 1 236
2 1768 1 239
2 1769 1 239
2 1770 1 242
2 1771 1 242
2 1772 1 244
2 1773 1 244
2 1774 1 247
2 1775 1 247
2 1776 1 250
2 1777 1 250
2 1778 1 252
2 1779 1 252
2 1780 1 255
2 1781 1 255
2 1782 1 258
2 1783 1 258
2 1784 1 260
2 1785 1 260
2 1786 1 263
2 1787 1 263
2 1788 1 266
2 1789 1 266
2 1790 1 268
2 1791 1 268
2 1792 1 271
2 1793 1 271
2 1794 1 274
2 1795 1 274
2 1796 1 276
2 1797 1 276
2 1798 1 279
2 1799 1 279
2 1800 1 282
2 1801 1 282
2 1802 1 284
2 1803 1 284
2 1804 1 287
2 1805 1 287
2 1806 1 290
2 1807 1 290
2 1808 1 292
2 1809 1 292
2 1810 1 295
2 1811 1 295
2 1812 1 298
2 1813 1 298
2 1814 1 300
2 1815 1 300
2 1816 1 303
2 1817 1 303
2 1818 1 306
2 1819 1 306
2 1820 1 308
2 1821 1 308
2 1822 1 311
2 1823 1 311
2 1824 1 314
2 1825 1 314
2 1826 1 316
2 1827 1 316
2 1828 1 319
2 1829 1 319
2 1830 1 322
2 1831 1 322
2 1832 1 324
2 1833 1 324
2 1834 1 327
2 1835 1 327
2 1836 1 330
2 1837 1 330
2 1838 1 332
2 1839 1 332
2 1840 1 335
2 1841 1 335
2 1842 1 338
2 1843 1 338
2 1844 1 340
2 1845 1 340
2 1846 1 343
2 1847 1 343
2 1848 1 346
2 1849 1 346
2 1850 1 348
2 1851 1 348
2 1852 1 351
2 1853 1 351
2 1854 1 354
2 1855 1 354
2 1856 1 356
2 1857 1 356
2 1858 1 359
2 1859 1 359
2 1860 1 362
2 1861 1 362
2 1862 1 364
2 1863 1 364
2 1864 1 367
2 1865 1 367
2 1866 1 370
2 1867 1 370
2 1868 1 372
2 1869 1 372
2 1870 1 375
2 1871 1 375
2 1872 1 378
2 1873 1 378
2 1874 1 380
2 1875 1 380
2 1876 1 383
2 1877 1 383
2 1878 1 386
2 1879 1 386
2 1880 1 388
2 1881 1 388
2 1882 1 391
2 1883 1 391
2 1884 1 394
2 1885 1 394
2 1886 1 396
2 1887 1 396
2 1888 1 399
2 1889 1 399
2 1890 1 402
2 1891 1 402
2 1892 1 404
2 1893 1 404
2 1894 1 407
2 1895 1 407
2 1896 1 410
2 1897 1 410
2 1898 1 412
2 1899 1 412
2 1900 1 415
2 1901 1 415
2 1902 1 418
2 1903 1 418
2 1904 1 420
2 1905 1 420
2 1906 1 423
2 1907 1 423
2 1908 1 426
2 1909 1 426
2 1910 1 428
2 1911 1 428
2 1912 1 431
2 1913 1 431
2 1914 1 434
2 1915 1 434
2 1916 1 436
2 1917 1 436
2 1918 1 439
2 1919 1 439
2 1920 1 441
2 1921 1 441
2 1922 1 443
2 1923 1 443
2 1924 1 445
2 1925 1 445
2 1926 1 446
2 1927 1 446
2 1928 1 448
2 1929 1 448
2 1930 1 455
2 1931 1 455
2 1932 1 457
2 1933 1 457
2 1934 1 458
2 1935 1 458
2 1936 1 458
2 1937 1 459
2 1938 1 459
2 1939 1 460
2 1940 1 460
2 1941 1 460
2 1942 1 461
2 1943 1 461
2 1944 1 467
2 1945 1 467
2 1946 1 470
2 1947 1 470
2 1948 1 470
2 1949 1 470
2 1950 1 472
2 1951 1 472
2 1952 1 472
2 1953 1 473
2 1954 1 473
2 1955 1 479
2 1956 1 479
2 1957 1 482
2 1958 1 482
2 1959 1 482
2 1960 1 482
2 1961 1 484
2 1962 1 484
2 1963 1 484
2 1964 1 484
2 1965 1 485
2 1966 1 485
2 1967 1 491
2 1968 1 491
2 1969 1 494
2 1970 1 494
2 1971 1 494
2 1972 1 494
2 1973 1 495
2 1974 1 495
2 1975 1 501
2 1976 1 501
2 1977 1 504
2 1978 1 504
2 1979 1 504
2 1980 1 504
2 1981 1 505
2 1982 1 505
2 1983 1 511
2 1984 1 511
2 1985 1 514
2 1986 1 514
2 1987 1 514
2 1988 1 514
2 1989 1 516
2 1990 1 516
2 1991 1 516
2 1992 1 516
2 1993 1 517
2 1994 1 517
2 1995 1 523
2 1996 1 523
2 1997 1 526
2 1998 1 526
2 1999 1 526
2 2000 1 526
2 2001 1 528
2 2002 1 528
2 2003 1 528
2 2004 1 528
2 2005 1 529
2 2006 1 529
2 2007 1 535
2 2008 1 535
2 2009 1 538
2 2010 1 538
2 2011 1 538
2 2012 1 540
2 2013 1 540
2 2014 1 540
2 2015 1 540
2 2016 1 541
2 2017 1 541
2 2018 1 547
2 2019 1 547
2 2020 1 550
2 2021 1 550
2 2022 1 550
2 2023 1 552
2 2024 1 552
2 2025 1 552
2 2026 1 552
2 2027 1 553
2 2028 1 553
2 2029 1 559
2 2030 1 559
2 2031 1 562
2 2032 1 562
2 2033 1 562
2 2034 1 562
2 2035 1 564
2 2036 1 564
2 2037 1 564
2 2038 1 565
2 2039 1 565
2 2040 1 571
2 2041 1 571
2 2042 1 574
2 2043 1 574
2 2044 1 574
2 2045 1 576
2 2046 1 576
2 2047 1 576
2 2048 1 577
2 2049 1 577
2 2050 1 583
2 2051 1 583
2 2052 1 586
2 2053 1 586
2 2054 1 586
2 2055 1 588
2 2056 1 588
2 2057 1 588
2 2058 1 589
2 2059 1 589
2 2060 1 595
2 2061 1 595
2 2062 1 598
2 2063 1 598
2 2064 1 598
2 2065 1 598
2 2066 1 600
2 2067 1 600
2 2068 1 600
2 2069 1 601
2 2070 1 601
2 2071 1 607
2 2072 1 607
2 2073 1 610
2 2074 1 610
2 2075 1 610
2 2076 1 612
2 2077 1 612
2 2078 1 612
2 2079 1 613
2 2080 1 613
2 2081 1 619
2 2082 1 619
2 2083 1 622
2 2084 1 622
2 2085 1 622
2 2086 1 622
2 2087 1 624
2 2088 1 624
2 2089 1 624
2 2090 1 625
2 2091 1 625
2 2092 1 631
2 2093 1 631
2 2094 1 634
2 2095 1 634
2 2096 1 634
2 2097 1 634
2 2098 1 636
2 2099 1 636
2 2100 1 636
2 2101 1 637
2 2102 1 637
2 2103 1 643
2 2104 1 643
2 2105 1 646
2 2106 1 646
2 2107 1 646
2 2108 1 648
2 2109 1 648
2 2110 1 648
2 2111 1 649
2 2112 1 649
2 2113 1 655
2 2114 1 655
2 2115 1 658
2 2116 1 658
2 2117 1 658
2 2118 1 660
2 2119 1 660
2 2120 1 660
2 2121 1 661
2 2122 1 661
2 2123 1 667
2 2124 1 667
2 2125 1 670
2 2126 1 670
2 2127 1 670
2 2128 1 672
2 2129 1 672
2 2130 1 672
2 2131 1 673
2 2132 1 673
2 2133 1 679
2 2134 1 679
2 2135 1 681
2 2136 1 681
2 2137 1 682
2 2138 1 682
2 2139 1 682
2 2140 1 684
2 2141 1 684
2 2142 1 684
2 2143 1 684
2 2144 1 685
2 2145 1 685
2 2146 1 691
2 2147 1 691
2 2148 1 694
2 2149 1 694
2 2150 1 694
2 2151 1 696
2 2152 1 696
2 2153 1 696
2 2154 1 696
2 2155 1 697
2 2156 1 697
2 2157 1 703
2 2158 1 703
2 2159 1 705
2 2160 1 705
2 2161 1 706
2 2162 1 706
2 2163 1 706
2 2164 1 707
2 2165 1 707
2 2166 1 708
2 2167 1 708
2 2168 1 708
2 2169 1 708
2 2170 1 709
2 2171 1 709
2 2172 1 715
2 2173 1 715
2 2174 1 717
2 2175 1 717
2 2176 1 718
2 2177 1 718
2 2178 1 718
2 2179 1 719
2 2180 1 719
2 2181 1 719
2 2182 1 720
2 2183 1 720
2 2184 1 720
2 2185 1 720
2 2186 1 721
2 2187 1 721
2 2188 1 727
2 2189 1 727
2 2190 1 730
2 2191 1 730
2 2192 1 730
2 2193 1 732
2 2194 1 732
2 2195 1 732
2 2196 1 733
2 2197 1 733
2 2198 1 739
2 2199 1 739
2 2200 1 742
2 2201 1 742
2 2202 1 742
2 2203 1 742
2 2204 1 744
2 2205 1 744
2 2206 1 744
2 2207 1 745
2 2208 1 745
2 2209 1 751
2 2210 1 751
2 2211 1 754
2 2212 1 754
2 2213 1 754
2 2214 1 754
2 2215 1 755
2 2216 1 755
2 2217 1 761
2 2218 1 761
2 2219 1 764
2 2220 1 764
2 2221 1 764
2 2222 1 764
2 2223 1 766
2 2224 1 766
2 2225 1 766
2 2226 1 767
2 2227 1 767
2 2228 1 773
2 2229 1 773
2 2230 1 776
2 2231 1 776
2 2232 1 776
2 2233 1 776
2 2234 1 778
2 2235 1 778
2 2236 1 778
2 2237 1 778
2 2238 1 779
2 2239 1 779
2 2240 1 785
2 2241 1 785
2 2242 1 788
2 2243 1 788
2 2244 1 788
2 2245 1 790
2 2246 1 790
2 2247 1 790
2 2248 1 791
2 2249 1 791
2 2250 1 797
2 2251 1 797
2 2252 1 800
2 2253 1 800
2 2254 1 800
2 2255 1 802
2 2256 1 802
2 2257 1 802
2 2258 1 803
2 2259 1 803
2 2260 1 809
2 2261 1 809
2 2262 1 812
2 2263 1 812
2 2264 1 815
2 2265 1 815
2 2266 1 820
2 2267 1 820
2 2268 1 823
2 2269 1 823
2 2270 1 824
2 2271 1 824
2 2272 1 827
2 2273 1 827
2 2274 1 828
2 2275 1 828
2 2276 1 831
2 2277 1 831
2 2278 1 833
2 2279 1 833
2 2280 1 835
2 2281 1 835
2 2282 1 837
2 2283 1 837
2 2284 1 840
2 2285 1 840
2 2286 1 844
2 2287 1 844
2 2288 1 844
2 2289 1 844
2 2290 1 846
2 2291 1 846
2 2292 1 848
2 2293 1 848
2 2294 1 849
2 2295 1 849
2 2296 1 852
2 2297 1 852
2 2298 1 859
2 2299 1 859
2 2300 1 862
2 2301 1 862
2 2302 1 866
2 2303 1 866
2 2304 1 867
2 2305 1 867
2 2306 1 870
2 2307 1 870
2 2308 1 871
2 2309 1 871
2 2310 1 874
2 2311 1 874
2 2312 1 875
2 2313 1 875
2 2314 1 878
2 2315 1 878
2 2316 1 880
2 2317 1 880
2 2318 1 882
2 2319 1 882
2 2320 1 884
2 2321 1 884
2 2322 1 886
2 2323 1 886
2 2324 1 887
2 2325 1 887
2 2326 1 890
2 2327 1 890
2 2328 1 892
2 2329 1 892
2 2330 1 894
2 2331 1 894
2 2332 1 895
2 2333 1 895
2 2334 1 898
2 2335 1 898
2 2336 1 899
2 2337 1 899
2 2338 1 902
2 2339 1 902
2 2340 1 904
2 2341 1 904
2 2342 1 906
2 2343 1 906
2 2344 1 907
2 2345 1 907
2 2346 1 910
2 2347 1 910
2 2348 1 911
2 2349 1 911
2 2350 1 914
2 2351 1 914
2 2352 1 916
2 2353 1 916
2 2354 1 918
2 2355 1 918
2 2356 1 921
2 2357 1 921
2 2358 1 926
2 2359 1 926
2 2360 1 926
2 2361 1 928
2 2362 1 928
2 2363 1 928
2 2364 1 929
2 2365 1 929
2 2366 1 931
2 2367 1 931
2 2368 1 935
2 2369 1 935
2 2370 1 940
2 2371 1 940
2 2372 1 945
2 2373 1 945
2 2374 1 948
2 2375 1 948
2 2376 1 952
2 2377 1 952
2 2378 1 958
2 2379 1 958
2 2380 1 958
2 2381 1 964
2 2382 1 964
2 2383 1 970
2 2384 1 970
2 2385 1 974
2 2386 1 974
2 2387 1 979
2 2388 1 979
2 2389 1 985
2 2390 1 985
2 2391 1 989
2 2392 1 989
2 2393 1 989
2 2394 1 995
2 2395 1 995
2 2396 1 996
2 2397 1 996
2 2398 1 1003
2 2399 1 1003
2 2400 1 1004
2 2401 1 1004
2 2402 1 1007
2 2403 1 1007
2 2404 1 1007
2 2405 1 1008
2 2406 1 1008
2 2407 1 1013
2 2408 1 1013
2 2409 1 1013
2 2410 1 1014
2 2411 1 1014
2 2412 1 1021
2 2413 1 1021
2 2414 1 1022
2 2415 1 1022
2 2416 1 1025
2 2417 1 1025
2 2418 1 1025
2 2419 1 1026
2 2420 1 1026
2 2421 1 1033
2 2422 1 1033
2 2423 1 1034
2 2424 1 1034
2 2425 1 1039
2 2426 1 1039
2 2427 1 1040
2 2428 1 1040
2 2429 1 1043
2 2430 1 1043
2 2431 1 1043
2 2432 1 1044
2 2433 1 1044
2 2434 1 1049
2 2435 1 1049
2 2436 1 1049
2 2437 1 1050
2 2438 1 1050
2 2439 1 1055
2 2440 1 1055
2 2441 1 1056
2 2442 1 1056
2 2443 1 1056
2 2444 1 1064
2 2445 1 1064
2 2446 1 1067
2 2447 1 1067
2 2448 1 1068
2 2449 1 1068
2 2450 1 1077
2 2451 1 1077
2 2452 1 1077
2 2453 1 1078
2 2454 1 1078
2 2455 1 1081
2 2456 1 1081
2 2457 1 1082
2 2458 1 1082
2 2459 1 1088
2 2460 1 1088
2 2461 1 1093
2 2462 1 1093
2 2463 1 1094
2 2464 1 1094
2 2465 1 1100
2 2466 1 1100
2 2467 1 1103
2 2468 1 1103
2 2469 1 1103
2 2470 1 1104
2 2471 1 1104
2 2472 1 1109
2 2473 1 1109
2 2474 1 1109
2 2475 1 1110
2 2476 1 1110
2 2477 1 1179
2 2478 1 1179
2 2479 1 1184
2 2480 1 1184
2 2481 1 1185
2 2482 1 1185
2 2483 1 1188
2 2484 1 1188
2 2485 1 1188
2 2486 1 1192
2 2487 1 1192
2 2488 1 1194
2 2489 1 1194
2 2490 1 1196
2 2491 1 1196
2 2492 1 1197
2 2493 1 1197
2 2494 1 1200
2 2495 1 1200
2 2496 1 1204
2 2497 1 1204
2 2498 1 1208
2 2499 1 1208
2 2500 1 1209
2 2501 1 1209
2 2502 1 1212
2 2503 1 1212
2 2504 1 1213
2 2505 1 1213
2 2506 1 1225
2 2507 1 1225
2 2508 1 1227
2 2509 1 1227
2 2510 1 1228
2 2511 1 1228
2 2512 1 1231
2 2513 1 1231
2 2514 1 1232
2 2515 1 1232
2 2516 1 1235
2 2517 1 1235
2 2518 1 1236
2 2519 1 1236
2 2520 1 1239
2 2521 1 1239
2 2522 1 1240
2 2523 1 1240
2 2524 1 1243
2 2525 1 1243
2 2526 1 1244
2 2527 1 1244
2 2528 1 1247
2 2529 1 1247
2 2530 1 1248
2 2531 1 1248
2 2532 1 1251
2 2533 1 1251
2 2534 1 1252
2 2535 1 1252
2 2536 1 1255
2 2537 1 1255
2 2538 1 1256
2 2539 1 1256
2 2540 1 1259
2 2541 1 1259
2 2542 1 1260
2 2543 1 1260
2 2544 1 1263
2 2545 1 1263
2 2546 1 1264
2 2547 1 1264
2 2548 1 1267
2 2549 1 1267
2 2550 1 1270
2 2551 1 1270
2 2552 1 1274
2 2553 1 1274
2 2554 1 1278
2 2555 1 1278
2 2556 1 1282
2 2557 1 1282
2 2558 1 1286
2 2559 1 1286
2 2560 1 1293
2 2561 1 1293
2 2562 1 1296
2 2563 1 1296
2 2564 1 1297
2 2565 1 1297
0 98 5 1 1 97
0 99 5 1 1 1480
0 100 5 1 1 1482
0 101 5 1 1 1484
0 102 5 1 1 1486
0 103 5 1 1 1488
0 104 5 1 1 1490
0 105 5 1 1 1492
0 106 5 1 1 1494
0 107 5 1 1 1496
0 108 5 1 1 1498
0 109 5 1 1 1500
0 110 5 1 1 1502
0 111 5 1 1 1504
0 112 5 1 1 1506
0 113 5 1 1 1508
0 114 5 1 1 1510
0 115 5 1 1 1512
0 116 5 1 1 1514
0 117 5 1 1 1516
0 118 5 1 1 1518
0 119 5 1 1 1520
0 120 5 1 1 1522
0 121 5 1 1 1524
0 122 5 1 1 1526
0 123 5 1 1 1528
0 124 5 1 1 1530
0 125 5 1 1 1532
0 126 5 1 1 1534
0 127 5 1 1 1536
0 128 5 1 1 1538
0 129 5 1 1 1540
0 130 5 1 1 1542
0 131 5 1 1 1544
0 132 5 1 1 1546
0 133 5 2 1 1548
0 134 5 2 1 1550
0 135 5 2 1 1552
0 136 5 2 1 1554
0 137 5 2 1 1556
0 138 5 2 1 1558
0 139 5 2 1 1560
0 140 5 2 1 1562
0 141 5 2 1 1564
0 142 5 2 1 1566
0 143 5 2 1 1568
0 144 5 2 1 1570
0 145 5 2 1 1572
0 146 5 2 1 1574
0 147 5 2 1 1576
0 148 5 2 1 1578
0 149 5 2 1 1580
0 150 5 2 1 1582
0 151 5 2 1 1584
0 152 5 2 1 1586
0 153 5 2 1 1588
0 154 5 2 1 1590
0 155 5 2 1 1592
0 156 5 2 1 1594
0 157 5 2 1 1596
0 158 5 2 1 1598
0 159 5 2 1 1600
0 160 5 2 1 1602
0 161 5 1 1 1604
0 162 5 1 1 1606
0 163 5 1 1 1608
0 164 5 1 1 1610
0 165 5 1 1 1612
0 166 5 1 1 1614
0 167 5 1 1 1616
0 168 5 1 1 1618
0 169 5 1 1 1620
0 170 5 1 1 1622
0 171 5 1 1 1624
0 172 5 1 1 1626
0 173 5 1 1 1628
0 174 5 1 1 1630
0 175 5 1 1 1632
0 176 5 1 1 1634
0 177 5 1 1 1636
0 178 5 1 1 1638
0 179 5 1 1 1640
0 180 5 1 1 1642
0 181 5 1 1 1644
0 182 5 1 1 1646
0 183 5 1 1 1648
0 184 5 1 1 1650
0 185 5 1 1 1652
0 186 5 1 1 1654
0 187 5 1 1 1656
0 188 5 1 1 1658
0 189 5 1 1 1660
0 190 5 1 1 1662
0 191 5 1 1 1664
0 192 5 1 1 1666
0 193 5 1 1 1668
0 194 5 1 1 1670
0 195 7 1 2 129 161
0 196 5 3 1 195
0 197 7 1 2 1541 1605
0 198 5 2 1 197
0 199 7 1 2 100 132
0 200 5 2 1 199
0 201 7 1 2 1483 1547
0 202 5 2 1 201
0 203 7 1 2 99 131
0 204 5 2 1 203
0 205 7 1 2 1481 1545
0 206 5 2 1 205
0 207 7 2 2 1479 1543
0 208 5 3 1 1741
0 209 7 1 2 1739 1743
0 210 5 1 1 209
0 211 7 2 2 1737 210
0 212 5 2 1 1746
0 213 7 1 2 1735 1748
0 214 5 1 1 213
0 215 7 2 2 1733 214
0 216 5 1 1 1750
0 217 7 1 2 101 216
0 218 5 2 1 217
0 219 7 1 2 1485 1751
0 220 5 2 1 219
0 221 7 1 2 1672 1754
0 222 5 1 1 221
0 223 7 2 2 1752 222
0 224 5 1 1 1756
0 225 7 1 2 102 224
0 226 5 2 1 225
0 227 7 1 2 1487 1757
0 228 5 2 1 227
0 229 7 1 2 1674 1760
0 230 5 1 1 229
0 231 7 2 2 1758 230
0 232 5 1 1 1762
0 233 7 1 2 103 232
0 234 5 2 1 233
0 235 7 1 2 1489 1763
0 236 5 2 1 235
0 237 7 1 2 1676 1766
0 238 5 1 1 237
0 239 7 2 2 1764 238
0 240 5 1 1 1768
0 241 7 1 2 104 240
0 242 5 2 1 241
0 243 7 1 2 1491 1769
0 244 5 2 1 243
0 245 7 1 2 1678 1772
0 246 5 1 1 245
0 247 7 2 2 1770 246
0 248 5 1 1 1774
0 249 7 1 2 105 248
0 250 5 2 1 249
0 251 7 1 2 1493 1775
0 252 5 2 1 251
0 253 7 1 2 1680 1778
0 254 5 1 1 253
0 255 7 2 2 1776 254
0 256 5 1 1 1780
0 257 7 1 2 106 256
0 258 5 2 1 257
0 259 7 1 2 1495 1781
0 260 5 2 1 259
0 261 7 1 2 1682 1784
0 262 5 1 1 261
0 263 7 2 2 1782 262
0 264 5 1 1 1786
0 265 7 1 2 107 264
0 266 5 2 1 265
0 267 7 1 2 1497 1787
0 268 5 2 1 267
0 269 7 1 2 1684 1790
0 270 5 1 1 269
0 271 7 2 2 1788 270
0 272 5 1 1 1792
0 273 7 1 2 108 272
0 274 5 2 1 273
0 275 7 1 2 1499 1793
0 276 5 2 1 275
0 277 7 1 2 1686 1796
0 278 5 1 1 277
0 279 7 2 2 1794 278
0 280 5 1 1 1798
0 281 7 1 2 109 280
0 282 5 2 1 281
0 283 7 1 2 1501 1799
0 284 5 2 1 283
0 285 7 1 2 1688 1802
0 286 5 1 1 285
0 287 7 2 2 1800 286
0 288 5 1 1 1804
0 289 7 1 2 110 288
0 290 5 2 1 289
0 291 7 1 2 1503 1805
0 292 5 2 1 291
0 293 7 1 2 1690 1808
0 294 5 1 1 293
0 295 7 2 2 1806 294
0 296 5 1 1 1810
0 297 7 1 2 111 296
0 298 5 2 1 297
0 299 7 1 2 1505 1811
0 300 5 2 1 299
0 301 7 1 2 1692 1814
0 302 5 1 1 301
0 303 7 2 2 1812 302
0 304 5 1 1 1816
0 305 7 1 2 112 304
0 306 5 2 1 305
0 307 7 1 2 1507 1817
0 308 5 2 1 307
0 309 7 1 2 1694 1820
0 310 5 1 1 309
0 311 7 2 2 1818 310
0 312 5 1 1 1822
0 313 7 1 2 113 312
0 314 5 2 1 313
0 315 7 1 2 1509 1823
0 316 5 2 1 315
0 317 7 1 2 1696 1826
0 318 5 1 1 317
0 319 7 2 2 1824 318
0 320 5 1 1 1828
0 321 7 1 2 114 320
0 322 5 2 1 321
0 323 7 1 2 1511 1829
0 324 5 2 1 323
0 325 7 1 2 1698 1832
0 326 5 1 1 325
0 327 7 2 2 1830 326
0 328 5 1 1 1834
0 329 7 1 2 115 328
0 330 5 2 1 329
0 331 7 1 2 1513 1835
0 332 5 2 1 331
0 333 7 1 2 1700 1838
0 334 5 1 1 333
0 335 7 2 2 1836 334
0 336 5 1 1 1840
0 337 7 1 2 116 336
0 338 5 2 1 337
0 339 7 1 2 1515 1841
0 340 5 2 1 339
0 341 7 1 2 1702 1844
0 342 5 1 1 341
0 343 7 2 2 1842 342
0 344 5 1 1 1846
0 345 7 1 2 117 344
0 346 5 2 1 345
0 347 7 1 2 1517 1847
0 348 5 2 1 347
0 349 7 1 2 1704 1850
0 350 5 1 1 349
0 351 7 2 2 1848 350
0 352 5 1 1 1852
0 353 7 1 2 118 352
0 354 5 2 1 353
0 355 7 1 2 1519 1853
0 356 5 2 1 355
0 357 7 1 2 1706 1856
0 358 5 1 1 357
0 359 7 2 2 1854 358
0 360 5 1 1 1858
0 361 7 1 2 119 360
0 362 5 2 1 361
0 363 7 1 2 1521 1859
0 364 5 2 1 363
0 365 7 1 2 1708 1862
0 366 5 1 1 365
0 367 7 2 2 1860 366
0 368 5 1 1 1864
0 369 7 1 2 120 368
0 370 5 2 1 369
0 371 7 1 2 1523 1865
0 372 5 2 1 371
0 373 7 1 2 1710 1868
0 374 5 1 1 373
0 375 7 2 2 1866 374
0 376 5 1 1 1870
0 377 7 1 2 121 376
0 378 5 2 1 377
0 379 7 1 2 1525 1871
0 380 5 2 1 379
0 381 7 1 2 1712 1874
0 382 5 1 1 381
0 383 7 2 2 1872 382
0 384 5 1 1 1876
0 385 7 1 2 122 384
0 386 5 2 1 385
0 387 7 1 2 1527 1877
0 388 5 2 1 387
0 389 7 1 2 1714 1880
0 390 5 1 1 389
0 391 7 2 2 1878 390
0 392 5 1 1 1882
0 393 7 1 2 123 392
0 394 5 2 1 393
0 395 7 1 2 1529 1883
0 396 5 2 1 395
0 397 7 1 2 1716 1886
0 398 5 1 1 397
0 399 7 2 2 1884 398
0 400 5 1 1 1888
0 401 7 1 2 124 400
0 402 5 2 1 401
0 403 7 1 2 1531 1889
0 404 5 2 1 403
0 405 7 1 2 1718 1892
0 406 5 1 1 405
0 407 7 2 2 1890 406
0 408 5 1 1 1894
0 409 7 1 2 125 408
0 410 5 2 1 409
0 411 7 1 2 1533 1895
0 412 5 2 1 411
0 413 7 1 2 1720 1898
0 414 5 1 1 413
0 415 7 2 2 1896 414
0 416 5 1 1 1900
0 417 7 1 2 126 416
0 418 5 2 1 417
0 419 7 1 2 1535 1901
0 420 5 2 1 419
0 421 7 1 2 1722 1904
0 422 5 1 1 421
0 423 7 2 2 1902 422
0 424 5 1 1 1906
0 425 7 1 2 127 424
0 426 5 2 1 425
0 427 7 1 2 1537 1907
0 428 5 2 1 427
0 429 7 1 2 1724 1910
0 430 5 1 1 429
0 431 7 2 2 1908 430
0 432 5 1 1 1912
0 433 7 1 2 128 432
0 434 5 2 1 433
0 435 7 1 2 1539 1913
0 436 5 2 1 435
0 437 7 1 2 1726 1916
0 438 5 1 1 437
0 439 7 2 2 1914 438
0 440 5 1 1 1918
0 441 7 2 2 1731 440
0 442 5 1 1 1920
0 443 7 2 2 1728 442
0 444 5 1 1 1922
0 445 7 2 2 194 1923
0 446 5 2 1 1924
0 447 7 1 2 1671 444
0 448 5 2 1 447
0 449 7 1 2 1729 1732
0 450 5 1 1 449
0 451 7 1 2 1919 450
0 452 5 1 1 451
0 453 7 1 2 1730 1921
0 454 5 1 1 453
0 455 7 2 2 452 454
0 456 5 1 1 1930
0 457 7 2 2 193 456
0 458 5 3 1 1932
0 459 7 2 2 1669 1931
0 460 5 3 1 1937
0 461 7 2 2 1915 1917
0 462 5 1 1 1942
0 463 7 1 2 1603 1943
0 464 5 1 1 463
0 465 7 1 2 1727 462
0 466 5 1 1 465
0 467 7 2 2 464 466
0 468 5 1 1 1944
0 469 7 1 2 1667 468
0 470 5 4 1 469
0 471 7 1 2 192 1945
0 472 5 3 1 471
0 473 7 2 2 1909 1911
0 474 5 1 1 1953
0 475 7 1 2 1601 1954
0 476 5 1 1 475
0 477 7 1 2 1725 474
0 478 5 1 1 477
0 479 7 2 2 476 478
0 480 5 1 1 1955
0 481 7 1 2 1665 480
0 482 5 4 1 481
0 483 7 1 2 191 1956
0 484 5 4 1 483
0 485 7 2 2 1903 1905
0 486 5 1 1 1965
0 487 7 1 2 1599 1966
0 488 5 1 1 487
0 489 7 1 2 1723 486
0 490 5 1 1 489
0 491 7 2 2 488 490
0 492 5 1 1 1967
0 493 7 1 2 1663 492
0 494 5 4 1 493
0 495 7 2 2 1897 1899
0 496 5 1 1 1973
0 497 7 1 2 1597 1974
0 498 5 1 1 497
0 499 7 1 2 1721 496
0 500 5 1 1 499
0 501 7 2 2 498 500
0 502 5 1 1 1975
0 503 7 1 2 1661 502
0 504 5 4 1 503
0 505 7 2 2 1891 1893
0 506 5 1 1 1981
0 507 7 1 2 1595 1982
0 508 5 1 1 507
0 509 7 1 2 1719 506
0 510 5 1 1 509
0 511 7 2 2 508 510
0 512 5 1 1 1983
0 513 7 1 2 1659 512
0 514 5 4 1 513
0 515 7 1 2 188 1984
0 516 5 4 1 515
0 517 7 2 2 1885 1887
0 518 5 1 1 1993
0 519 7 1 2 1593 1994
0 520 5 1 1 519
0 521 7 1 2 1717 518
0 522 5 1 1 521
0 523 7 2 2 520 522
0 524 5 1 1 1995
0 525 7 1 2 1657 524
0 526 5 4 1 525
0 527 7 1 2 187 1996
0 528 5 4 1 527
0 529 7 2 2 1879 1881
0 530 5 1 1 2005
0 531 7 1 2 1591 2006
0 532 5 1 1 531
0 533 7 1 2 1715 530
0 534 5 1 1 533
0 535 7 2 2 532 534
0 536 5 1 1 2007
0 537 7 1 2 1655 536
0 538 5 3 1 537
0 539 7 1 2 186 2008
0 540 5 4 1 539
0 541 7 2 2 1873 1875
0 542 5 1 1 2016
0 543 7 1 2 1589 2017
0 544 5 1 1 543
0 545 7 1 2 1713 542
0 546 5 1 1 545
0 547 7 2 2 544 546
0 548 5 1 1 2018
0 549 7 1 2 1653 548
0 550 5 3 1 549
0 551 7 1 2 185 2019
0 552 5 4 1 551
0 553 7 2 2 1867 1869
0 554 5 1 1 2027
0 555 7 1 2 1587 2028
0 556 5 1 1 555
0 557 7 1 2 1711 554
0 558 5 1 1 557
0 559 7 2 2 556 558
0 560 5 1 1 2029
0 561 7 1 2 1651 560
0 562 5 4 1 561
0 563 7 1 2 184 2030
0 564 5 3 1 563
0 565 7 2 2 1861 1863
0 566 5 1 1 2038
0 567 7 1 2 1585 2039
0 568 5 1 1 567
0 569 7 1 2 1709 566
0 570 5 1 1 569
0 571 7 2 2 568 570
0 572 5 1 1 2040
0 573 7 1 2 1649 572
0 574 5 3 1 573
0 575 7 1 2 183 2041
0 576 5 3 1 575
0 577 7 2 2 1855 1857
0 578 5 1 1 2048
0 579 7 1 2 1583 2049
0 580 5 1 1 579
0 581 7 1 2 1707 578
0 582 5 1 1 581
0 583 7 2 2 580 582
0 584 5 1 1 2050
0 585 7 1 2 1647 584
0 586 5 3 1 585
0 587 7 1 2 182 2051
0 588 5 3 1 587
0 589 7 2 2 1849 1851
0 590 5 1 1 2058
0 591 7 1 2 1581 2059
0 592 5 1 1 591
0 593 7 1 2 1705 590
0 594 5 1 1 593
0 595 7 2 2 592 594
0 596 5 1 1 2060
0 597 7 1 2 1645 596
0 598 5 4 1 597
0 599 7 1 2 181 2061
0 600 5 3 1 599
0 601 7 2 2 1843 1845
0 602 5 1 1 2069
0 603 7 1 2 1579 2070
0 604 5 1 1 603
0 605 7 1 2 1703 602
0 606 5 1 1 605
0 607 7 2 2 604 606
0 608 5 1 1 2071
0 609 7 1 2 1643 608
0 610 5 3 1 609
0 611 7 1 2 180 2072
0 612 5 3 1 611
0 613 7 2 2 1837 1839
0 614 5 1 1 2079
0 615 7 1 2 1577 2080
0 616 5 1 1 615
0 617 7 1 2 1701 614
0 618 5 1 1 617
0 619 7 2 2 616 618
0 620 5 1 1 2081
0 621 7 1 2 1641 620
0 622 5 4 1 621
0 623 7 1 2 179 2082
0 624 5 3 1 623
0 625 7 2 2 1831 1833
0 626 5 1 1 2090
0 627 7 1 2 1575 2091
0 628 5 1 1 627
0 629 7 1 2 1699 626
0 630 5 1 1 629
0 631 7 2 2 628 630
0 632 5 1 1 2092
0 633 7 1 2 1639 632
0 634 5 4 1 633
0 635 7 1 2 178 2093
0 636 5 3 1 635
0 637 7 2 2 1825 1827
0 638 5 1 1 2101
0 639 7 1 2 1573 2102
0 640 5 1 1 639
0 641 7 1 2 1697 638
0 642 5 1 1 641
0 643 7 2 2 640 642
0 644 5 1 1 2103
0 645 7 1 2 1637 644
0 646 5 3 1 645
0 647 7 1 2 177 2104
0 648 5 3 1 647
0 649 7 2 2 1819 1821
0 650 5 1 1 2111
0 651 7 1 2 1571 2112
0 652 5 1 1 651
0 653 7 1 2 1695 650
0 654 5 1 1 653
0 655 7 2 2 652 654
0 656 5 1 1 2113
0 657 7 1 2 1635 656
0 658 5 3 1 657
0 659 7 1 2 176 2114
0 660 5 3 1 659
0 661 7 2 2 1813 1815
0 662 5 1 1 2121
0 663 7 1 2 1569 2122
0 664 5 1 1 663
0 665 7 1 2 1693 662
0 666 5 1 1 665
0 667 7 2 2 664 666
0 668 5 1 1 2123
0 669 7 1 2 1633 668
0 670 5 3 1 669
0 671 7 1 2 175 2124
0 672 5 3 1 671
0 673 7 2 2 1807 1809
0 674 5 1 1 2131
0 675 7 1 2 1567 2132
0 676 5 1 1 675
0 677 7 1 2 1691 674
0 678 5 1 1 677
0 679 7 2 2 676 678
0 680 5 1 1 2133
0 681 7 2 2 1631 680
0 682 5 3 1 2135
0 683 7 1 2 174 2134
0 684 5 4 1 683
0 685 7 2 2 1801 1803
0 686 5 1 1 2144
0 687 7 1 2 1565 2145
0 688 5 1 1 687
0 689 7 1 2 1689 686
0 690 5 1 1 689
0 691 7 2 2 688 690
0 692 5 1 1 2146
0 693 7 1 2 1629 692
0 694 5 3 1 693
0 695 7 1 2 173 2147
0 696 5 4 1 695
0 697 7 2 2 1795 1797
0 698 5 1 1 2155
0 699 7 1 2 1563 2156
0 700 5 1 1 699
0 701 7 1 2 1687 698
0 702 5 1 1 701
0 703 7 2 2 700 702
0 704 5 1 1 2157
0 705 7 2 2 1627 704
0 706 5 3 1 2159
0 707 7 2 2 172 2158
0 708 5 4 1 2164
0 709 7 2 2 1789 1791
0 710 5 1 1 2170
0 711 7 1 2 1561 2171
0 712 5 1 1 711
0 713 7 1 2 1685 710
0 714 5 1 1 713
0 715 7 2 2 712 714
0 716 5 1 1 2172
0 717 7 2 2 171 2173
0 718 5 3 1 2174
0 719 7 3 2 1625 716
0 720 5 4 1 2179
0 721 7 2 2 1783 1785
0 722 5 1 1 2186
0 723 7 1 2 1559 2187
0 724 5 1 1 723
0 725 7 1 2 1683 722
0 726 5 1 1 725
0 727 7 2 2 724 726
0 728 5 1 1 2188
0 729 7 1 2 1623 728
0 730 5 3 1 729
0 731 7 1 2 170 2189
0 732 5 3 1 731
0 733 7 2 2 1777 1779
0 734 5 1 1 2196
0 735 7 1 2 1557 2197
0 736 5 1 1 735
0 737 7 1 2 1681 734
0 738 5 1 1 737
0 739 7 2 2 736 738
0 740 5 1 1 2198
0 741 7 1 2 1621 740
0 742 5 4 1 741
0 743 7 1 2 169 2199
0 744 5 3 1 743
0 745 7 2 2 1771 1773
0 746 5 1 1 2207
0 747 7 1 2 1555 2208
0 748 5 1 1 747
0 749 7 1 2 1679 746
0 750 5 1 1 749
0 751 7 2 2 748 750
0 752 5 1 1 2209
0 753 7 1 2 1619 752
0 754 5 4 1 753
0 755 7 2 2 1765 1767
0 756 5 1 1 2215
0 757 7 1 2 1553 2216
0 758 5 1 1 757
0 759 7 1 2 1677 756
0 760 5 1 1 759
0 761 7 2 2 758 760
0 762 5 1 1 2217
0 763 7 1 2 167 2218
0 764 5 4 1 763
0 765 7 1 2 1617 762
0 766 5 3 1 765
0 767 7 2 2 1759 1761
0 768 5 1 1 2226
0 769 7 1 2 1551 2227
0 770 5 1 1 769
0 771 7 1 2 1675 768
0 772 5 1 1 771
0 773 7 2 2 770 772
0 774 5 1 1 2228
0 775 7 1 2 1615 774
0 776 5 4 1 775
0 777 7 1 2 166 2229
0 778 5 4 1 777
0 779 7 2 2 1753 1755
0 780 5 1 1 2238
0 781 7 1 2 1549 2239
0 782 5 1 1 781
0 783 7 1 2 1673 780
0 784 5 1 1 783
0 785 7 2 2 782 784
0 786 5 1 1 2240
0 787 7 1 2 165 2241
0 788 5 3 1 787
0 789 7 1 2 1613 786
0 790 5 3 1 789
0 791 7 2 2 1734 1736
0 792 5 1 1 2248
0 793 7 1 2 1747 792
0 794 5 1 1 793
0 795 7 1 2 1749 2249
0 796 5 1 1 795
0 797 7 2 2 794 796
0 798 5 1 1 2250
0 799 7 1 2 164 798
0 800 5 3 1 799
0 801 7 1 2 1611 2251
0 802 5 3 1 801
0 803 7 2 2 1738 1740
0 804 5 1 1 2258
0 805 7 1 2 1742 804
0 806 5 1 1 805
0 807 7 1 2 1744 2259
0 808 5 1 1 807
0 809 7 2 2 806 808
0 810 5 1 1 2260
0 811 7 1 2 163 810
0 812 5 2 1 811
0 813 7 1 2 98 130
0 814 5 1 1 813
0 815 7 2 2 1745 814
0 816 5 1 1 2264
0 817 7 1 2 1607 816
0 818 5 1 1 817
0 819 7 1 2 1609 2261
0 820 5 2 1 819
0 821 7 1 2 818 2266
0 822 5 1 1 821
0 823 7 2 2 2262 822
0 824 5 2 1 2268
0 825 7 1 2 2255 2270
0 826 5 1 1 825
0 827 7 2 2 2252 826
0 828 5 2 1 2272
0 829 7 1 2 2245 2274
0 830 5 1 1 829
0 831 7 2 2 2242 830
0 832 5 1 1 2276
0 833 7 2 2 2234 2277
0 834 5 1 1 2278
0 835 7 2 2 2230 834
0 836 5 1 1 2280
0 837 7 2 2 2223 2281
0 838 5 1 1 2282
0 839 7 1 2 2219 838
0 840 5 2 1 839
0 841 7 1 2 2211 2284
0 842 5 1 1 841
0 843 7 1 2 168 2210
0 844 5 4 1 843
0 845 7 1 2 842 2286
0 846 7 2 2 2204 845
0 847 5 1 1 2290
0 848 7 2 2 2200 847
0 849 5 2 1 2292
0 850 7 1 2 2193 2294
0 851 5 1 1 850
0 852 7 2 2 2190 851
0 853 7 1 2 2182 2296
0 854 5 1 1 853
0 855 7 1 2 2176 854
0 856 7 1 2 2166 855
0 857 5 1 1 856
0 858 7 1 2 2161 857
0 859 5 2 1 858
0 860 7 1 2 2151 2298
0 861 5 1 1 860
0 862 7 2 2 2148 861
0 863 5 1 1 2300
0 864 7 1 2 2140 863
0 865 5 1 1 864
0 866 7 2 2 2137 865
0 867 5 2 1 2302
0 868 7 1 2 2128 2304
0 869 5 1 1 868
0 870 7 2 2 2125 869
0 871 5 2 1 2306
0 872 7 1 2 2118 2308
0 873 5 1 1 872
0 874 7 2 2 2115 873
0 875 5 2 1 2310
0 876 7 1 2 2108 2312
0 877 5 1 1 876
0 878 7 2 2 2105 877
0 879 5 1 1 2314
0 880 7 2 2 2098 879
0 881 5 1 1 2316
0 882 7 2 2 2094 881
0 883 5 1 1 2318
0 884 7 2 2 2087 883
0 885 5 1 1 2320
0 886 7 2 2 2083 885
0 887 5 2 1 2322
0 888 7 1 2 2076 2324
0 889 5 1 1 888
0 890 7 2 2 2073 889
0 891 5 1 1 2326
0 892 7 2 2 2066 891
0 893 5 1 1 2328
0 894 7 2 2 2062 893
0 895 5 2 1 2330
0 896 7 1 2 2055 2332
0 897 5 1 1 896
0 898 7 2 2 2052 897
0 899 5 2 1 2334
0 900 7 1 2 2045 2336
0 901 5 1 1 900
0 902 7 2 2 2042 901
0 903 5 1 1 2338
0 904 7 2 2 2035 903
0 905 5 1 1 2340
0 906 7 2 2 2031 905
0 907 5 2 1 2342
0 908 7 1 2 2023 2344
0 909 5 1 1 908
0 910 7 2 2 2020 909
0 911 5 2 1 2346
0 912 7 1 2 2012 2348
0 913 5 1 1 912
0 914 7 2 2 2009 913
0 915 5 1 1 2350
0 916 7 2 2 2001 915
0 917 5 1 1 2352
0 918 7 2 2 1997 917
0 919 5 1 1 2354
0 920 7 1 2 1989 919
0 921 5 2 1 920
0 922 7 1 2 1985 2356
0 923 7 1 2 1977 922
0 924 5 1 1 923
0 925 7 1 2 190 1968
0 926 5 3 1 925
0 927 7 1 2 189 1976
0 928 5 3 1 927
0 929 7 2 2 2358 2361
0 930 7 1 2 924 2364
0 931 5 2 1 930
0 932 7 1 2 1969 2366
0 933 5 1 1 932
0 934 7 1 2 1961 933
0 935 5 2 1 934
0 936 7 1 2 1957 2368
0 937 5 1 1 936
0 938 7 1 2 1950 937
0 939 5 1 1 938
0 940 7 2 2 1946 939
0 941 5 1 1 2370
0 942 7 1 2 1939 2371
0 943 5 1 1 942
0 944 7 1 2 1934 943
0 945 5 2 1 944
0 946 7 1 2 1928 2372
0 947 5 1 1 946
0 948 7 2 2 1926 947
0 949 5 1 1 2374
0 950 7 1 2 1925 2373
0 951 5 1 1 950
0 952 7 2 2 1935 1940
0 953 5 1 1 2376
0 954 7 1 2 941 2377
0 955 5 1 1 954
0 956 7 1 2 1947 953
0 957 5 1 1 956
0 958 7 3 2 1948 1951
0 959 5 1 1 2378
0 960 7 1 2 2369 2379
0 961 5 1 1 960
0 962 7 1 2 1958 961
0 963 5 1 1 962
0 964 7 2 2 1959 1962
0 965 5 1 1 2381
0 966 7 1 2 2367 2382
0 967 5 1 1 966
0 968 7 1 2 1970 967
0 969 5 1 1 968
0 970 7 2 2 1971 2359
0 971 5 1 1 2383
0 972 7 1 2 1978 971
0 973 5 1 1 972
0 974 7 2 2 1979 2362
0 975 7 1 2 2357 2385
0 976 5 1 1 975
0 977 7 1 2 1986 976
0 978 5 1 1 977
0 979 7 2 2 1987 1990
0 980 5 1 1 2387
0 981 7 1 2 2355 980
0 982 5 1 1 981
0 983 7 1 2 1998 2353
0 984 5 1 1 983
0 985 7 2 2 1999 2002
0 986 5 1 1 2389
0 987 7 1 2 2351 986
0 988 5 1 1 987
0 989 7 3 2 2010 2013
0 990 5 1 1 2391
0 991 7 1 2 2347 990
0 992 5 1 1 991
0 993 7 1 2 2349 2392
0 994 5 1 1 993
0 995 7 2 2 2021 2024
0 996 5 2 1 2394
0 997 7 1 2 2343 2396
0 998 5 1 1 997
0 999 7 1 2 2345 2395
0 1000 5 1 1 999
0 1001 7 1 2 2032 2341
0 1002 5 1 1 1001
0 1003 7 2 2 2033 2036
0 1004 5 2 1 2398
0 1005 7 1 2 2339 2400
0 1006 5 1 1 1005
0 1007 7 3 2 2043 2046
0 1008 5 2 1 2402
0 1009 7 1 2 2335 2405
0 1010 5 1 1 1009
0 1011 7 1 2 2337 2403
0 1012 5 1 1 1011
0 1013 7 3 2 2053 2056
0 1014 5 2 1 2407
0 1015 7 1 2 2331 2410
0 1016 5 1 1 1015
0 1017 7 1 2 2333 2408
0 1018 5 1 1 1017
0 1019 7 1 2 2063 2329
0 1020 5 1 1 1019
0 1021 7 2 2 2064 2067
0 1022 5 2 1 2412
0 1023 7 1 2 2327 2414
0 1024 5 1 1 1023
0 1025 7 3 2 2074 2077
0 1026 5 2 1 2416
0 1027 7 1 2 2323 2419
0 1028 5 1 1 1027
0 1029 7 1 2 2325 2417
0 1030 5 1 1 1029
0 1031 7 1 2 2084 2321
0 1032 5 1 1 1031
0 1033 7 2 2 2085 2088
0 1034 5 2 1 2421
0 1035 7 1 2 2319 2423
0 1036 5 1 1 1035
0 1037 7 1 2 2095 2317
0 1038 5 1 1 1037
0 1039 7 2 2 2096 2099
0 1040 5 2 1 2425
0 1041 7 1 2 2315 2427
0 1042 5 1 1 1041
0 1043 7 3 2 2106 2109
0 1044 5 2 1 2429
0 1045 7 1 2 2311 2432
0 1046 5 1 1 1045
0 1047 7 1 2 2313 2430
0 1048 5 1 1 1047
0 1049 7 3 2 2116 2119
0 1050 5 2 1 2434
0 1051 7 1 2 2309 2435
0 1052 5 1 1 1051
0 1053 7 1 2 2307 2437
0 1054 5 1 1 1053
0 1055 7 2 2 2126 2129
0 1056 5 3 1 2439
0 1057 7 1 2 2136 2441
0 1058 5 1 1 1057
0 1059 7 1 2 2305 1058
0 1060 5 1 1 1059
0 1061 7 1 2 2303 2442
0 1062 5 1 1 1061
0 1063 7 1 2 2138 2141
0 1064 5 2 1 1063
0 1065 7 1 2 2301 2444
0 1066 5 1 1 1065
0 1067 7 2 2 2149 2152
0 1068 5 2 1 2446
0 1069 7 1 2 2160 2180
0 1070 5 1 1 1069
0 1071 7 1 2 2448 1070
0 1072 5 1 1 1071
0 1073 7 1 2 2299 2447
0 1074 5 1 1 1073
0 1075 7 1 2 2165 2183
0 1076 5 1 1 1075
0 1077 7 3 2 2191 2194
0 1078 5 2 1 2450
0 1079 7 1 2 2293 2451
0 1080 5 1 1 1079
0 1081 7 2 2 2201 2205
0 1082 5 2 1 2455
0 1083 7 1 2 2212 2457
0 1084 5 1 1 1083
0 1085 7 1 2 2202 2291
0 1086 5 1 1 1085
0 1087 7 1 2 2213 2287
0 1088 5 2 1 1087
0 1089 7 1 2 2285 2459
0 1090 5 1 1 1089
0 1091 7 1 2 2220 2283
0 1092 5 1 1 1091
0 1093 7 2 2 2221 2224
0 1094 5 2 1 2461
0 1095 7 1 2 836 2463
0 1096 5 1 1 1095
0 1097 7 1 2 2231 2279
0 1098 5 1 1 1097
0 1099 7 1 2 2232 2235
0 1100 5 2 1 1099
0 1101 7 1 2 832 2465
0 1102 5 1 1 1101
0 1103 7 3 2 2243 2246
0 1104 5 2 1 2467
0 1105 7 1 2 2275 2468
0 1106 5 1 1 1105
0 1107 7 1 2 2273 2470
0 1108 5 1 1 1107
0 1109 7 3 2 2253 2256
0 1110 5 2 1 2472
0 1111 7 1 2 2271 2473
0 1112 5 1 1 1111
0 1113 7 1 2 2269 2475
0 1114 5 1 1 1113
0 1115 7 1 2 1112 1114
0 1116 7 1 2 1108 1115
0 1117 7 1 2 1106 1116
0 1118 5 1 1 1117
0 1119 7 1 2 1102 1118
0 1120 7 1 2 1098 1119
0 1121 5 1 1 1120
0 1122 7 1 2 1096 1121
0 1123 7 1 2 1092 1122
0 1124 5 1 1 1123
0 1125 7 1 2 1090 1124
0 1126 7 1 2 1086 1125
0 1127 7 1 2 1084 1126
0 1128 5 1 1 1127
0 1129 7 1 2 2295 2453
0 1130 5 1 1 1129
0 1131 7 1 2 1128 1130
0 1132 7 1 2 1080 1131
0 1133 5 1 1 1132
0 1134 7 1 2 2177 2184
0 1135 5 1 1 1134
0 1136 7 1 2 2297 1135
0 1137 5 1 1 1136
0 1138 7 1 2 1133 1137
0 1139 7 1 2 1076 1138
0 1140 7 1 2 1074 1139
0 1141 7 1 2 1072 1140
0 1142 7 1 2 1066 1141
0 1143 7 1 2 1062 1142
0 1144 7 1 2 1060 1143
0 1145 7 1 2 1054 1144
0 1146 7 1 2 1052 1145
0 1147 7 1 2 1048 1146
0 1148 7 1 2 1046 1147
0 1149 7 1 2 1042 1148
0 1150 7 1 2 1038 1149
0 1151 7 1 2 1036 1150
0 1152 7 1 2 1032 1151
0 1153 7 1 2 1030 1152
0 1154 7 1 2 1028 1153
0 1155 7 1 2 1024 1154
0 1156 7 1 2 1020 1155
0 1157 7 1 2 1018 1156
0 1158 7 1 2 1016 1157
0 1159 7 1 2 1012 1158
0 1160 7 1 2 1010 1159
0 1161 7 1 2 1006 1160
0 1162 7 1 2 1002 1161
0 1163 7 1 2 1000 1162
0 1164 7 1 2 998 1163
0 1165 7 1 2 994 1164
0 1166 7 1 2 992 1165
0 1167 7 1 2 988 1166
0 1168 7 1 2 984 1167
0 1169 7 1 2 982 1168
0 1170 7 1 2 978 1169
0 1171 7 1 2 973 1170
0 1172 7 1 2 969 1171
0 1173 7 1 2 963 1172
0 1174 7 1 2 957 1173
0 1175 7 1 2 955 1174
0 1176 7 1 2 951 1175
0 1177 7 1 2 949 1176
0 1178 5 1 1 1177
0 1179 7 2 2 1927 1929
0 1180 5 1 1 2477
0 1181 7 1 2 162 2265
0 1182 7 1 2 2267 1181
0 1183 5 1 1 1182
0 1184 7 2 2 2263 1183
0 1185 5 2 1 2479
0 1186 7 1 2 2257 2481
0 1187 5 1 1 1186
0 1188 7 3 2 2254 1187
0 1189 5 1 1 2483
0 1190 7 1 2 2244 2484
0 1191 5 1 1 1190
0 1192 7 2 2 2247 1191
0 1193 5 1 1 2486
0 1194 7 2 2 2233 2487
0 1195 5 1 1 2488
0 1196 7 2 2 2236 1195
0 1197 5 2 1 2490
0 1198 7 1 2 2225 2492
0 1199 5 1 1 1198
0 1200 7 2 2 2222 1199
0 1201 5 1 1 2494
0 1202 7 1 2 2214 1201
0 1203 5 1 1 1202
0 1204 7 2 2 2288 1203
0 1205 5 1 1 2496
0 1206 7 1 2 2206 2497
0 1207 5 1 1 1206
0 1208 7 2 2 2203 1207
0 1209 5 2 1 2498
0 1210 7 1 2 2195 2500
0 1211 5 1 1 1210
0 1212 7 2 2 2192 1211
0 1213 5 2 1 2502
0 1214 7 1 2 2178 2504
0 1215 5 1 1 1214
0 1216 7 1 2 2185 1215
0 1217 7 1 2 2162 1216
0 1218 5 1 1 1217
0 1219 7 1 2 2167 1218
0 1220 5 1 1 1219
0 1221 7 1 2 2150 1220
0 1222 5 1 1 1221
0 1223 7 1 2 2153 1222
0 1224 5 1 1 1223
0 1225 7 2 2 2139 1224
0 1226 5 1 1 2506
0 1227 7 2 2 2142 1226
0 1228 5 2 1 2508
0 1229 7 1 2 2127 2510
0 1230 5 1 1 1229
0 1231 7 2 2 2130 1230
0 1232 5 2 1 2512
0 1233 7 1 2 2117 2514
0 1234 5 1 1 1233
0 1235 7 2 2 2120 1234
0 1236 5 2 1 2516
0 1237 7 1 2 2107 2518
0 1238 5 1 1 1237
0 1239 7 2 2 2110 1238
0 1240 5 2 1 2520
0 1241 7 1 2 2097 2522
0 1242 5 1 1 1241
0 1243 7 2 2 2100 1242
0 1244 5 2 1 2524
0 1245 7 1 2 2086 2526
0 1246 5 1 1 1245
0 1247 7 2 2 2089 1246
0 1248 5 2 1 2528
0 1249 7 1 2 2075 2530
0 1250 5 1 1 1249
0 1251 7 2 2 2078 1250
0 1252 5 2 1 2532
0 1253 7 1 2 2065 2534
0 1254 5 1 1 1253
0 1255 7 2 2 2068 1254
0 1256 5 2 1 2536
0 1257 7 1 2 2054 2538
0 1258 5 1 1 1257
0 1259 7 2 2 2057 1258
0 1260 5 2 1 2540
0 1261 7 1 2 2044 2542
0 1262 5 1 1 1261
0 1263 7 2 2 2047 1262
0 1264 5 2 1 2544
0 1265 7 1 2 2034 2546
0 1266 5 1 1 1265
0 1267 7 2 2 2037 1266
0 1268 5 1 1 2548
0 1269 7 1 2 2022 1268
0 1270 5 2 1 1269
0 1271 7 1 2 2025 2550
0 1272 5 1 1 1271
0 1273 7 1 2 2011 1272
0 1274 5 2 1 1273
0 1275 7 1 2 2014 2552
0 1276 5 1 1 1275
0 1277 7 1 2 2000 1276
0 1278 5 2 1 1277
0 1279 7 1 2 2003 2554
0 1280 5 1 1 1279
0 1281 7 1 2 1988 1280
0 1282 5 2 1 1281
0 1283 7 1 2 1991 2556
0 1284 5 1 1 1283
0 1285 7 1 2 1980 1284
0 1286 5 2 1 1285
0 1287 7 1 2 2365 2558
0 1288 5 1 1 1287
0 1289 7 1 2 1972 1288
0 1290 7 1 2 1960 1289
0 1291 5 1 1 1290
0 1292 7 1 2 1963 1291
0 1293 5 2 1 1292
0 1294 7 1 2 1949 2560
0 1295 5 1 1 1294
0 1296 7 2 2 1952 1295
0 1297 5 2 1 2562
0 1298 7 1 2 1941 2564
0 1299 5 1 1 1298
0 1300 7 1 2 2478 1299
0 1301 5 1 1 1300
0 1302 7 1 2 1936 1301
0 1303 5 1 1 1302
0 1304 7 1 2 1180 2565
0 1305 5 1 1 1304
0 1306 7 1 2 1933 1305
0 1307 5 1 1 1306
0 1308 7 1 2 1938 2563
0 1309 5 1 1 1308
0 1310 7 1 2 1964 959
0 1311 5 1 1 1310
0 1312 7 1 2 2380 2561
0 1313 5 1 1 1312
0 1314 7 1 2 2360 965
0 1315 5 1 1 1314
0 1316 7 1 2 2384 2559
0 1317 5 1 1 1316
0 1318 7 1 2 2363 1317
0 1319 5 1 1 1318
0 1320 7 1 2 2386 2557
0 1321 5 1 1 1320
0 1322 7 1 2 1992 1321
0 1323 5 1 1 1322
0 1324 7 1 2 2388 2555
0 1325 5 1 1 1324
0 1326 7 1 2 2004 1325
0 1327 5 1 1 1326
0 1328 7 1 2 2390 2553
0 1329 5 1 1 1328
0 1330 7 1 2 2015 1329
0 1331 5 1 1 1330
0 1332 7 1 2 2393 2551
0 1333 5 1 1 1332
0 1334 7 1 2 2026 1333
0 1335 5 1 1 1334
0 1336 7 1 2 2397 2549
0 1337 5 1 1 1336
0 1338 7 1 2 2399 2547
0 1339 5 1 1 1338
0 1340 7 1 2 2401 2545
0 1341 5 1 1 1340
0 1342 7 1 2 2406 2541
0 1343 5 1 1 1342
0 1344 7 1 2 2404 2543
0 1345 5 1 1 1344
0 1346 7 1 2 2411 2537
0 1347 5 1 1 1346
0 1348 7 1 2 2409 2539
0 1349 5 1 1 1348
0 1350 7 1 2 2415 2533
0 1351 5 1 1 1350
0 1352 7 1 2 2413 2535
0 1353 5 1 1 1352
0 1354 7 1 2 2420 2531
0 1355 5 1 1 1354
0 1356 7 1 2 2418 2529
0 1357 5 1 1 1356
0 1358 7 1 2 1355 1357
0 1359 5 1 1 1358
0 1360 7 1 2 2424 2525
0 1361 5 1 1 1360
0 1362 7 1 2 2422 2527
0 1363 5 1 1 1362
0 1364 7 1 2 2426 2523
0 1365 5 1 1 1364
0 1366 7 1 2 2428 2521
0 1367 5 1 1 1366
0 1368 7 1 2 2433 2519
0 1369 5 1 1 1368
0 1370 7 1 2 2431 2517
0 1371 5 1 1 1370
0 1372 7 1 2 1369 1371
0 1373 5 1 1 1372
0 1374 7 1 2 2438 2513
0 1375 5 1 1 1374
0 1376 7 1 2 2436 2515
0 1377 5 1 1 1376
0 1378 7 1 2 2443 2511
0 1379 5 1 1 1378
0 1380 7 1 2 2440 2509
0 1381 5 1 1 1380
0 1382 7 1 2 1379 1381
0 1383 5 1 1 1382
0 1384 7 1 2 2143 2507
0 1385 5 1 1 1384
0 1386 7 1 2 2154 2445
0 1387 5 1 1 1386
0 1388 7 1 2 2168 2449
0 1389 5 1 1 1388
0 1390 7 1 2 2175 2503
0 1391 5 1 1 1390
0 1392 7 1 2 2163 2169
0 1393 5 1 1 1392
0 1394 7 1 2 1391 1393
0 1395 5 1 1 1394
0 1396 7 1 2 2181 2505
0 1397 5 1 1 1396
0 1398 7 1 2 2454 2499
0 1399 5 1 1 1398
0 1400 7 1 2 2289 2458
0 1401 5 1 1 1400
0 1402 7 1 2 2456 1205
0 1403 5 1 1 1402
0 1404 7 1 2 2460 2495
0 1405 5 1 1 1404
0 1406 7 1 2 2462 2491
0 1407 5 1 1 1406
0 1408 7 1 2 2237 2489
0 1409 5 1 1 1408
0 1410 7 1 2 2466 1193
0 1411 5 1 1 1410
0 1412 7 1 2 2469 2485
0 1413 5 1 1 1412
0 1414 7 1 2 2476 2480
0 1415 5 1 1 1414
0 1416 7 1 2 2474 2482
0 1417 5 1 1 1416
0 1418 7 1 2 1415 1417
0 1419 5 1 1 1418
0 1420 7 1 2 2471 1189
0 1421 5 1 1 1420
0 1422 7 1 2 1419 1421
0 1423 7 1 2 1413 1422
0 1424 5 1 1 1423
0 1425 7 1 2 1411 1424
0 1426 7 1 2 1409 1425
0 1427 5 1 1 1426
0 1428 7 1 2 2464 2493
0 1429 5 1 1 1428
0 1430 7 1 2 1427 1429
0 1431 7 1 2 1407 1430
0 1432 5 1 1 1431
0 1433 7 1 2 1405 1432
0 1434 7 1 2 1403 1433
0 1435 7 1 2 1401 1434
0 1436 5 1 1 1435
0 1437 7 1 2 2452 2501
0 1438 5 1 1 1437
0 1439 7 1 2 1436 1438
0 1440 7 1 2 1399 1439
0 1441 5 1 1 1440
0 1442 7 1 2 1397 1441
0 1443 7 1 2 1395 1442
0 1444 7 1 2 1389 1443
0 1445 7 1 2 1387 1444
0 1446 7 1 2 1385 1445
0 1447 7 1 2 1383 1446
0 1448 7 1 2 1377 1447
0 1449 7 1 2 1375 1448
0 1450 7 1 2 1373 1449
0 1451 7 1 2 1367 1450
0 1452 7 1 2 1365 1451
0 1453 7 1 2 1363 1452
0 1454 7 1 2 1361 1453
0 1455 7 1 2 1359 1454
0 1456 7 1 2 1353 1455
0 1457 7 1 2 1351 1456
0 1458 7 1 2 1349 1457
0 1459 7 1 2 1347 1458
0 1460 7 1 2 1345 1459
0 1461 7 1 2 1343 1460
0 1462 7 1 2 1341 1461
0 1463 7 1 2 1339 1462
0 1464 7 1 2 1337 1463
0 1465 7 1 2 1335 1464
0 1466 7 1 2 1331 1465
0 1467 7 1 2 1327 1466
0 1468 7 1 2 1323 1467
0 1469 7 1 2 1319 1468
0 1470 7 1 2 1315 1469
0 1471 7 1 2 1313 1470
0 1472 7 1 2 1311 1471
0 1473 7 1 2 1309 1472
0 1474 7 1 2 1307 1473
0 1475 7 1 2 1303 1474
0 1476 7 1 2 2375 1475
0 1477 5 1 1 1476
0 1478 7 1 2 1178 1477
3 2999 5 0 1 1478
