1 0 0 100 0
2 25 1 0
2 26 1 0
2 21756 1 0
2 21757 1 0
2 21758 1 0
2 21759 1 0
2 21760 1 0
2 21761 1 0
2 21762 1 0
2 21763 1 0
2 21764 1 0
2 21765 1 0
2 21766 1 0
2 21767 1 0
2 21768 1 0
2 21769 1 0
2 21770 1 0
2 21771 1 0
2 21772 1 0
2 21773 1 0
2 21774 1 0
2 21775 1 0
2 21776 1 0
2 21777 1 0
2 21778 1 0
2 21779 1 0
2 21780 1 0
2 21781 1 0
2 21782 1 0
2 21783 1 0
2 21784 1 0
2 21785 1 0
2 21786 1 0
2 21787 1 0
2 21788 1 0
2 21789 1 0
2 21790 1 0
2 21791 1 0
2 21792 1 0
2 21793 1 0
2 21794 1 0
2 21795 1 0
2 21796 1 0
2 21797 1 0
2 21798 1 0
2 21799 1 0
2 21800 1 0
2 21801 1 0
2 21802 1 0
2 21803 1 0
2 21804 1 0
2 21805 1 0
2 21806 1 0
2 21807 1 0
2 21808 1 0
2 21809 1 0
2 21810 1 0
2 21811 1 0
2 21812 1 0
2 21813 1 0
2 21814 1 0
2 21815 1 0
2 21816 1 0
2 21817 1 0
2 21818 1 0
2 21819 1 0
2 21820 1 0
2 21821 1 0
2 21822 1 0
2 21823 1 0
2 21824 1 0
2 21825 1 0
2 21826 1 0
2 21827 1 0
2 21828 1 0
2 21829 1 0
2 21830 1 0
2 21831 1 0
2 21832 1 0
2 21833 1 0
2 21834 1 0
2 21835 1 0
2 21836 1 0
2 21837 1 0
2 21838 1 0
2 21839 1 0
2 21840 1 0
2 21841 1 0
2 21842 1 0
2 21843 1 0
2 21844 1 0
2 21845 1 0
2 21846 1 0
2 21847 1 0
2 21848 1 0
2 21849 1 0
2 21850 1 0
2 21851 1 0
2 21852 1 0
2 21853 1 0
1 1 0 118 0
2 21854 1 1
2 21855 1 1
2 21856 1 1
2 21857 1 1
2 21858 1 1
2 21859 1 1
2 21860 1 1
2 21861 1 1
2 21862 1 1
2 21863 1 1
2 21864 1 1
2 21865 1 1
2 21866 1 1
2 21867 1 1
2 21868 1 1
2 21869 1 1
2 21870 1 1
2 21871 1 1
2 21872 1 1
2 21873 1 1
2 21874 1 1
2 21875 1 1
2 21876 1 1
2 21877 1 1
2 21878 1 1
2 21879 1 1
2 21880 1 1
2 21881 1 1
2 21882 1 1
2 21883 1 1
2 21884 1 1
2 21885 1 1
2 21886 1 1
2 21887 1 1
2 21888 1 1
2 21889 1 1
2 21890 1 1
2 21891 1 1
2 21892 1 1
2 21893 1 1
2 21894 1 1
2 21895 1 1
2 21896 1 1
2 21897 1 1
2 21898 1 1
2 21899 1 1
2 21900 1 1
2 21901 1 1
2 21902 1 1
2 21903 1 1
2 21904 1 1
2 21905 1 1
2 21906 1 1
2 21907 1 1
2 21908 1 1
2 21909 1 1
2 21910 1 1
2 21911 1 1
2 21912 1 1
2 21913 1 1
2 21914 1 1
2 21915 1 1
2 21916 1 1
2 21917 1 1
2 21918 1 1
2 21919 1 1
2 21920 1 1
2 21921 1 1
2 21922 1 1
2 21923 1 1
2 21924 1 1
2 21925 1 1
2 21926 1 1
2 21927 1 1
2 21928 1 1
2 21929 1 1
2 21930 1 1
2 21931 1 1
2 21932 1 1
2 21933 1 1
2 21934 1 1
2 21935 1 1
2 21936 1 1
2 21937 1 1
2 21938 1 1
2 21939 1 1
2 21940 1 1
2 21941 1 1
2 21942 1 1
2 21943 1 1
2 21944 1 1
2 21945 1 1
2 21946 1 1
2 21947 1 1
2 21948 1 1
2 21949 1 1
2 21950 1 1
2 21951 1 1
2 21952 1 1
2 21953 1 1
2 21954 1 1
2 21955 1 1
2 21956 1 1
2 21957 1 1
2 21958 1 1
2 21959 1 1
2 21960 1 1
2 21961 1 1
2 21962 1 1
2 21963 1 1
2 21964 1 1
2 21965 1 1
2 21966 1 1
2 21967 1 1
2 21968 1 1
2 21969 1 1
2 21970 1 1
2 21971 1 1
1 2 0 143 0
2 21972 1 2
2 21973 1 2
2 21974 1 2
2 21975 1 2
2 21976 1 2
2 21977 1 2
2 21978 1 2
2 21979 1 2
2 21980 1 2
2 21981 1 2
2 21982 1 2
2 21983 1 2
2 21984 1 2
2 21985 1 2
2 21986 1 2
2 21987 1 2
2 21988 1 2
2 21989 1 2
2 21990 1 2
2 21991 1 2
2 21992 1 2
2 21993 1 2
2 21994 1 2
2 21995 1 2
2 21996 1 2
2 21997 1 2
2 21998 1 2
2 21999 1 2
2 22000 1 2
2 22001 1 2
2 22002 1 2
2 22003 1 2
2 22004 1 2
2 22005 1 2
2 22006 1 2
2 22007 1 2
2 22008 1 2
2 22009 1 2
2 22010 1 2
2 22011 1 2
2 22012 1 2
2 22013 1 2
2 22014 1 2
2 22015 1 2
2 22016 1 2
2 22017 1 2
2 22018 1 2
2 22019 1 2
2 22020 1 2
2 22021 1 2
2 22022 1 2
2 22023 1 2
2 22024 1 2
2 22025 1 2
2 22026 1 2
2 22027 1 2
2 22028 1 2
2 22029 1 2
2 22030 1 2
2 22031 1 2
2 22032 1 2
2 22033 1 2
2 22034 1 2
2 22035 1 2
2 22036 1 2
2 22037 1 2
2 22038 1 2
2 22039 1 2
2 22040 1 2
2 22041 1 2
2 22042 1 2
2 22043 1 2
2 22044 1 2
2 22045 1 2
2 22046 1 2
2 22047 1 2
2 22048 1 2
2 22049 1 2
2 22050 1 2
2 22051 1 2
2 22052 1 2
2 22053 1 2
2 22054 1 2
2 22055 1 2
2 22056 1 2
2 22057 1 2
2 22058 1 2
2 22059 1 2
2 22060 1 2
2 22061 1 2
2 22062 1 2
2 22063 1 2
2 22064 1 2
2 22065 1 2
2 22066 1 2
2 22067 1 2
2 22068 1 2
2 22069 1 2
2 22070 1 2
2 22071 1 2
2 22072 1 2
2 22073 1 2
2 22074 1 2
2 22075 1 2
2 22076 1 2
2 22077 1 2
2 22078 1 2
2 22079 1 2
2 22080 1 2
2 22081 1 2
2 22082 1 2
2 22083 1 2
2 22084 1 2
2 22085 1 2
2 22086 1 2
2 22087 1 2
2 22088 1 2
2 22089 1 2
2 22090 1 2
2 22091 1 2
2 22092 1 2
2 22093 1 2
2 22094 1 2
2 22095 1 2
2 22096 1 2
2 22097 1 2
2 22098 1 2
2 22099 1 2
2 22100 1 2
2 22101 1 2
2 22102 1 2
2 22103 1 2
2 22104 1 2
2 22105 1 2
2 22106 1 2
2 22107 1 2
2 22108 1 2
2 22109 1 2
2 22110 1 2
2 22111 1 2
2 22112 1 2
2 22113 1 2
2 22114 1 2
1 3 0 51 0
2 22115 1 3
2 22116 1 3
2 22117 1 3
2 22118 1 3
2 22119 1 3
2 22120 1 3
2 22121 1 3
2 22122 1 3
2 22123 1 3
2 22124 1 3
2 22125 1 3
2 22126 1 3
2 22127 1 3
2 22128 1 3
2 22129 1 3
2 22130 1 3
2 22131 1 3
2 22132 1 3
2 22133 1 3
2 22134 1 3
2 22135 1 3
2 22136 1 3
2 22137 1 3
2 22138 1 3
2 22139 1 3
2 22140 1 3
2 22141 1 3
2 22142 1 3
2 22143 1 3
2 22144 1 3
2 22145 1 3
2 22146 1 3
2 22147 1 3
2 22148 1 3
2 22149 1 3
2 22150 1 3
2 22151 1 3
2 22152 1 3
2 22153 1 3
2 22154 1 3
2 22155 1 3
2 22156 1 3
2 22157 1 3
2 22158 1 3
2 22159 1 3
2 22160 1 3
2 22161 1 3
2 22162 1 3
2 22163 1 3
2 22164 1 3
2 22165 1 3
1 4 0 75 0
2 22166 1 4
2 22167 1 4
2 22168 1 4
2 22169 1 4
2 22170 1 4
2 22171 1 4
2 22172 1 4
2 22173 1 4
2 22174 1 4
2 22175 1 4
2 22176 1 4
2 22177 1 4
2 22178 1 4
2 22179 1 4
2 22180 1 4
2 22181 1 4
2 22182 1 4
2 22183 1 4
2 22184 1 4
2 22185 1 4
2 22186 1 4
2 22187 1 4
2 22188 1 4
2 22189 1 4
2 22190 1 4
2 22191 1 4
2 22192 1 4
2 22193 1 4
2 22194 1 4
2 22195 1 4
2 22196 1 4
2 22197 1 4
2 22198 1 4
2 22199 1 4
2 22200 1 4
2 22201 1 4
2 22202 1 4
2 22203 1 4
2 22204 1 4
2 22205 1 4
2 22206 1 4
2 22207 1 4
2 22208 1 4
2 22209 1 4
2 22210 1 4
2 22211 1 4
2 22212 1 4
2 22213 1 4
2 22214 1 4
2 22215 1 4
2 22216 1 4
2 22217 1 4
2 22218 1 4
2 22219 1 4
2 22220 1 4
2 22221 1 4
2 22222 1 4
2 22223 1 4
2 22224 1 4
2 22225 1 4
2 22226 1 4
2 22227 1 4
2 22228 1 4
2 22229 1 4
2 22230 1 4
2 22231 1 4
2 22232 1 4
2 22233 1 4
2 22234 1 4
2 22235 1 4
2 22236 1 4
2 22237 1 4
2 22238 1 4
2 22239 1 4
2 22240 1 4
1 5 0 40 0
2 22241 1 5
2 22242 1 5
2 22243 1 5
2 22244 1 5
2 22245 1 5
2 22246 1 5
2 22247 1 5
2 22248 1 5
2 22249 1 5
2 22250 1 5
2 22251 1 5
2 22252 1 5
2 22253 1 5
2 22254 1 5
2 22255 1 5
2 22256 1 5
2 22257 1 5
2 22258 1 5
2 22259 1 5
2 22260 1 5
2 22261 1 5
2 22262 1 5
2 22263 1 5
2 22264 1 5
2 22265 1 5
2 22266 1 5
2 22267 1 5
2 22268 1 5
2 22269 1 5
2 22270 1 5
2 22271 1 5
2 22272 1 5
2 22273 1 5
2 22274 1 5
2 22275 1 5
2 22276 1 5
2 22277 1 5
2 22278 1 5
2 22279 1 5
2 22280 1 5
1 6 0 68 0
2 22281 1 6
2 22282 1 6
2 22283 1 6
2 22284 1 6
2 22285 1 6
2 22286 1 6
2 22287 1 6
2 22288 1 6
2 22289 1 6
2 22290 1 6
2 22291 1 6
2 22292 1 6
2 22293 1 6
2 22294 1 6
2 22295 1 6
2 22296 1 6
2 22297 1 6
2 22298 1 6
2 22299 1 6
2 22300 1 6
2 22301 1 6
2 22302 1 6
2 22303 1 6
2 22304 1 6
2 22305 1 6
2 22306 1 6
2 22307 1 6
2 22308 1 6
2 22309 1 6
2 22310 1 6
2 22311 1 6
2 22312 1 6
2 22313 1 6
2 22314 1 6
2 22315 1 6
2 22316 1 6
2 22317 1 6
2 22318 1 6
2 22319 1 6
2 22320 1 6
2 22321 1 6
2 22322 1 6
2 22323 1 6
2 22324 1 6
2 22325 1 6
2 22326 1 6
2 22327 1 6
2 22328 1 6
2 22329 1 6
2 22330 1 6
2 22331 1 6
2 22332 1 6
2 22333 1 6
2 22334 1 6
2 22335 1 6
2 22336 1 6
2 22337 1 6
2 22338 1 6
2 22339 1 6
2 22340 1 6
2 22341 1 6
2 22342 1 6
2 22343 1 6
2 22344 1 6
2 22345 1 6
2 22346 1 6
2 22347 1 6
2 22348 1 6
1 7 0 79 0
2 22349 1 7
2 22350 1 7
2 22351 1 7
2 22352 1 7
2 22353 1 7
2 22354 1 7
2 22355 1 7
2 22356 1 7
2 22357 1 7
2 22358 1 7
2 22359 1 7
2 22360 1 7
2 22361 1 7
2 22362 1 7
2 22363 1 7
2 22364 1 7
2 22365 1 7
2 22366 1 7
2 22367 1 7
2 22368 1 7
2 22369 1 7
2 22370 1 7
2 22371 1 7
2 22372 1 7
2 22373 1 7
2 22374 1 7
2 22375 1 7
2 22376 1 7
2 22377 1 7
2 22378 1 7
2 22379 1 7
2 22380 1 7
2 22381 1 7
2 22382 1 7
2 22383 1 7
2 22384 1 7
2 22385 1 7
2 22386 1 7
2 22387 1 7
2 22388 1 7
2 22389 1 7
2 22390 1 7
2 22391 1 7
2 22392 1 7
2 22393 1 7
2 22394 1 7
2 22395 1 7
2 22396 1 7
2 22397 1 7
2 22398 1 7
2 22399 1 7
2 22400 1 7
2 22401 1 7
2 22402 1 7
2 22403 1 7
2 22404 1 7
2 22405 1 7
2 22406 1 7
2 22407 1 7
2 22408 1 7
2 22409 1 7
2 22410 1 7
2 22411 1 7
2 22412 1 7
2 22413 1 7
2 22414 1 7
2 22415 1 7
2 22416 1 7
2 22417 1 7
2 22418 1 7
2 22419 1 7
2 22420 1 7
2 22421 1 7
2 22422 1 7
2 22423 1 7
2 22424 1 7
2 22425 1 7
2 22426 1 7
2 22427 1 7
1 8 0 65 0
2 22428 1 8
2 22429 1 8
2 22430 1 8
2 22431 1 8
2 22432 1 8
2 22433 1 8
2 22434 1 8
2 22435 1 8
2 22436 1 8
2 22437 1 8
2 22438 1 8
2 22439 1 8
2 22440 1 8
2 22441 1 8
2 22442 1 8
2 22443 1 8
2 22444 1 8
2 22445 1 8
2 22446 1 8
2 22447 1 8
2 22448 1 8
2 22449 1 8
2 22450 1 8
2 22451 1 8
2 22452 1 8
2 22453 1 8
2 22454 1 8
2 22455 1 8
2 22456 1 8
2 22457 1 8
2 22458 1 8
2 22459 1 8
2 22460 1 8
2 22461 1 8
2 22462 1 8
2 22463 1 8
2 22464 1 8
2 22465 1 8
2 22466 1 8
2 22467 1 8
2 22468 1 8
2 22469 1 8
2 22470 1 8
2 22471 1 8
2 22472 1 8
2 22473 1 8
2 22474 1 8
2 22475 1 8
2 22476 1 8
2 22477 1 8
2 22478 1 8
2 22479 1 8
2 22480 1 8
2 22481 1 8
2 22482 1 8
2 22483 1 8
2 22484 1 8
2 22485 1 8
2 22486 1 8
2 22487 1 8
2 22488 1 8
2 22489 1 8
2 22490 1 8
2 22491 1 8
2 22492 1 8
1 9 0 93 0
2 22493 1 9
2 22494 1 9
2 22495 1 9
2 22496 1 9
2 22497 1 9
2 22498 1 9
2 22499 1 9
2 22500 1 9
2 22501 1 9
2 22502 1 9
2 22503 1 9
2 22504 1 9
2 22505 1 9
2 22506 1 9
2 22507 1 9
2 22508 1 9
2 22509 1 9
2 22510 1 9
2 22511 1 9
2 22512 1 9
2 22513 1 9
2 22514 1 9
2 22515 1 9
2 22516 1 9
2 22517 1 9
2 22518 1 9
2 22519 1 9
2 22520 1 9
2 22521 1 9
2 22522 1 9
2 22523 1 9
2 22524 1 9
2 22525 1 9
2 22526 1 9
2 22527 1 9
2 22528 1 9
2 22529 1 9
2 22530 1 9
2 22531 1 9
2 22532 1 9
2 22533 1 9
2 22534 1 9
2 22535 1 9
2 22536 1 9
2 22537 1 9
2 22538 1 9
2 22539 1 9
2 22540 1 9
2 22541 1 9
2 22542 1 9
2 22543 1 9
2 22544 1 9
2 22545 1 9
2 22546 1 9
2 22547 1 9
2 22548 1 9
2 22549 1 9
2 22550 1 9
2 22551 1 9
2 22552 1 9
2 22553 1 9
2 22554 1 9
2 22555 1 9
2 22556 1 9
2 22557 1 9
2 22558 1 9
2 22559 1 9
2 22560 1 9
2 22561 1 9
2 22562 1 9
2 22563 1 9
2 22564 1 9
2 22565 1 9
2 22566 1 9
2 22567 1 9
2 22568 1 9
2 22569 1 9
2 22570 1 9
2 22571 1 9
2 22572 1 9
2 22573 1 9
2 22574 1 9
2 22575 1 9
2 22576 1 9
2 22577 1 9
2 22578 1 9
2 22579 1 9
2 22580 1 9
2 22581 1 9
2 22582 1 9
2 22583 1 9
2 22584 1 9
2 22585 1 9
1 10 0 101 0
2 22586 1 10
2 22587 1 10
2 22588 1 10
2 22589 1 10
2 22590 1 10
2 22591 1 10
2 22592 1 10
2 22593 1 10
2 22594 1 10
2 22595 1 10
2 22596 1 10
2 22597 1 10
2 22598 1 10
2 22599 1 10
2 22600 1 10
2 22601 1 10
2 22602 1 10
2 22603 1 10
2 22604 1 10
2 22605 1 10
2 22606 1 10
2 22607 1 10
2 22608 1 10
2 22609 1 10
2 22610 1 10
2 22611 1 10
2 22612 1 10
2 22613 1 10
2 22614 1 10
2 22615 1 10
2 22616 1 10
2 22617 1 10
2 22618 1 10
2 22619 1 10
2 22620 1 10
2 22621 1 10
2 22622 1 10
2 22623 1 10
2 22624 1 10
2 22625 1 10
2 22626 1 10
2 22627 1 10
2 22628 1 10
2 22629 1 10
2 22630 1 10
2 22631 1 10
2 22632 1 10
2 22633 1 10
2 22634 1 10
2 22635 1 10
2 22636 1 10
2 22637 1 10
2 22638 1 10
2 22639 1 10
2 22640 1 10
2 22641 1 10
2 22642 1 10
2 22643 1 10
2 22644 1 10
2 22645 1 10
2 22646 1 10
2 22647 1 10
2 22648 1 10
2 22649 1 10
2 22650 1 10
2 22651 1 10
2 22652 1 10
2 22653 1 10
2 22654 1 10
2 22655 1 10
2 22656 1 10
2 22657 1 10
2 22658 1 10
2 22659 1 10
2 22660 1 10
2 22661 1 10
2 22662 1 10
2 22663 1 10
2 22664 1 10
2 22665 1 10
2 22666 1 10
2 22667 1 10
2 22668 1 10
2 22669 1 10
2 22670 1 10
2 22671 1 10
2 22672 1 10
2 22673 1 10
2 22674 1 10
2 22675 1 10
2 22676 1 10
2 22677 1 10
2 22678 1 10
2 22679 1 10
2 22680 1 10
2 22681 1 10
2 22682 1 10
2 22683 1 10
2 22684 1 10
2 22685 1 10
2 22686 1 10
1 11 0 39 0
2 22687 1 11
2 22688 1 11
2 22689 1 11
2 22690 1 11
2 22691 1 11
2 22692 1 11
2 22693 1 11
2 22694 1 11
2 22695 1 11
2 22696 1 11
2 22697 1 11
2 22698 1 11
2 22699 1 11
2 22700 1 11
2 22701 1 11
2 22702 1 11
2 22703 1 11
2 22704 1 11
2 22705 1 11
2 22706 1 11
2 22707 1 11
2 22708 1 11
2 22709 1 11
2 22710 1 11
2 22711 1 11
2 22712 1 11
2 22713 1 11
2 22714 1 11
2 22715 1 11
2 22716 1 11
2 22717 1 11
2 22718 1 11
2 22719 1 11
2 22720 1 11
2 22721 1 11
2 22722 1 11
2 22723 1 11
2 22724 1 11
2 22725 1 11
1 12 0 59 0
2 22726 1 12
2 22727 1 12
2 22728 1 12
2 22729 1 12
2 22730 1 12
2 22731 1 12
2 22732 1 12
2 22733 1 12
2 22734 1 12
2 22735 1 12
2 22736 1 12
2 22737 1 12
2 22738 1 12
2 22739 1 12
2 22740 1 12
2 22741 1 12
2 22742 1 12
2 22743 1 12
2 22744 1 12
2 22745 1 12
2 22746 1 12
2 22747 1 12
2 22748 1 12
2 22749 1 12
2 22750 1 12
2 22751 1 12
2 22752 1 12
2 22753 1 12
2 22754 1 12
2 22755 1 12
2 22756 1 12
2 22757 1 12
2 22758 1 12
2 22759 1 12
2 22760 1 12
2 22761 1 12
2 22762 1 12
2 22763 1 12
2 22764 1 12
2 22765 1 12
2 22766 1 12
2 22767 1 12
2 22768 1 12
2 22769 1 12
2 22770 1 12
2 22771 1 12
2 22772 1 12
2 22773 1 12
2 22774 1 12
2 22775 1 12
2 22776 1 12
2 22777 1 12
2 22778 1 12
2 22779 1 12
2 22780 1 12
2 22781 1 12
2 22782 1 12
2 22783 1 12
2 22784 1 12
1 13 0 37 0
2 22785 1 13
2 22786 1 13
2 22787 1 13
2 22788 1 13
2 22789 1 13
2 22790 1 13
2 22791 1 13
2 22792 1 13
2 22793 1 13
2 22794 1 13
2 22795 1 13
2 22796 1 13
2 22797 1 13
2 22798 1 13
2 22799 1 13
2 22800 1 13
2 22801 1 13
2 22802 1 13
2 22803 1 13
2 22804 1 13
2 22805 1 13
2 22806 1 13
2 22807 1 13
2 22808 1 13
2 22809 1 13
2 22810 1 13
2 22811 1 13
2 22812 1 13
2 22813 1 13
2 22814 1 13
2 22815 1 13
2 22816 1 13
2 22817 1 13
2 22818 1 13
2 22819 1 13
2 22820 1 13
2 22821 1 13
1 14 0 63 0
2 22822 1 14
2 22823 1 14
2 22824 1 14
2 22825 1 14
2 22826 1 14
2 22827 1 14
2 22828 1 14
2 22829 1 14
2 22830 1 14
2 22831 1 14
2 22832 1 14
2 22833 1 14
2 22834 1 14
2 22835 1 14
2 22836 1 14
2 22837 1 14
2 22838 1 14
2 22839 1 14
2 22840 1 14
2 22841 1 14
2 22842 1 14
2 22843 1 14
2 22844 1 14
2 22845 1 14
2 22846 1 14
2 22847 1 14
2 22848 1 14
2 22849 1 14
2 22850 1 14
2 22851 1 14
2 22852 1 14
2 22853 1 14
2 22854 1 14
2 22855 1 14
2 22856 1 14
2 22857 1 14
2 22858 1 14
2 22859 1 14
2 22860 1 14
2 22861 1 14
2 22862 1 14
2 22863 1 14
2 22864 1 14
2 22865 1 14
2 22866 1 14
2 22867 1 14
2 22868 1 14
2 22869 1 14
2 22870 1 14
2 22871 1 14
2 22872 1 14
2 22873 1 14
2 22874 1 14
2 22875 1 14
2 22876 1 14
2 22877 1 14
2 22878 1 14
2 22879 1 14
2 22880 1 14
2 22881 1 14
2 22882 1 14
2 22883 1 14
2 22884 1 14
1 15 0 70 0
2 22885 1 15
2 22886 1 15
2 22887 1 15
2 22888 1 15
2 22889 1 15
2 22890 1 15
2 22891 1 15
2 22892 1 15
2 22893 1 15
2 22894 1 15
2 22895 1 15
2 22896 1 15
2 22897 1 15
2 22898 1 15
2 22899 1 15
2 22900 1 15
2 22901 1 15
2 22902 1 15
2 22903 1 15
2 22904 1 15
2 22905 1 15
2 22906 1 15
2 22907 1 15
2 22908 1 15
2 22909 1 15
2 22910 1 15
2 22911 1 15
2 22912 1 15
2 22913 1 15
2 22914 1 15
2 22915 1 15
2 22916 1 15
2 22917 1 15
2 22918 1 15
2 22919 1 15
2 22920 1 15
2 22921 1 15
2 22922 1 15
2 22923 1 15
2 22924 1 15
2 22925 1 15
2 22926 1 15
2 22927 1 15
2 22928 1 15
2 22929 1 15
2 22930 1 15
2 22931 1 15
2 22932 1 15
2 22933 1 15
2 22934 1 15
2 22935 1 15
2 22936 1 15
2 22937 1 15
2 22938 1 15
2 22939 1 15
2 22940 1 15
2 22941 1 15
2 22942 1 15
2 22943 1 15
2 22944 1 15
2 22945 1 15
2 22946 1 15
2 22947 1 15
2 22948 1 15
2 22949 1 15
2 22950 1 15
2 22951 1 15
2 22952 1 15
2 22953 1 15
2 22954 1 15
1 16 0 78 0
2 22955 1 16
2 22956 1 16
2 22957 1 16
2 22958 1 16
2 22959 1 16
2 22960 1 16
2 22961 1 16
2 22962 1 16
2 22963 1 16
2 22964 1 16
2 22965 1 16
2 22966 1 16
2 22967 1 16
2 22968 1 16
2 22969 1 16
2 22970 1 16
2 22971 1 16
2 22972 1 16
2 22973 1 16
2 22974 1 16
2 22975 1 16
2 22976 1 16
2 22977 1 16
2 22978 1 16
2 22979 1 16
2 22980 1 16
2 22981 1 16
2 22982 1 16
2 22983 1 16
2 22984 1 16
2 22985 1 16
2 22986 1 16
2 22987 1 16
2 22988 1 16
2 22989 1 16
2 22990 1 16
2 22991 1 16
2 22992 1 16
2 22993 1 16
2 22994 1 16
2 22995 1 16
2 22996 1 16
2 22997 1 16
2 22998 1 16
2 22999 1 16
2 23000 1 16
2 23001 1 16
2 23002 1 16
2 23003 1 16
2 23004 1 16
2 23005 1 16
2 23006 1 16
2 23007 1 16
2 23008 1 16
2 23009 1 16
2 23010 1 16
2 23011 1 16
2 23012 1 16
2 23013 1 16
2 23014 1 16
2 23015 1 16
2 23016 1 16
2 23017 1 16
2 23018 1 16
2 23019 1 16
2 23020 1 16
2 23021 1 16
2 23022 1 16
2 23023 1 16
2 23024 1 16
2 23025 1 16
2 23026 1 16
2 23027 1 16
2 23028 1 16
2 23029 1 16
2 23030 1 16
2 23031 1 16
2 23032 1 16
1 17 0 123 0
2 23033 1 17
2 23034 1 17
2 23035 1 17
2 23036 1 17
2 23037 1 17
2 23038 1 17
2 23039 1 17
2 23040 1 17
2 23041 1 17
2 23042 1 17
2 23043 1 17
2 23044 1 17
2 23045 1 17
2 23046 1 17
2 23047 1 17
2 23048 1 17
2 23049 1 17
2 23050 1 17
2 23051 1 17
2 23052 1 17
2 23053 1 17
2 23054 1 17
2 23055 1 17
2 23056 1 17
2 23057 1 17
2 23058 1 17
2 23059 1 17
2 23060 1 17
2 23061 1 17
2 23062 1 17
2 23063 1 17
2 23064 1 17
2 23065 1 17
2 23066 1 17
2 23067 1 17
2 23068 1 17
2 23069 1 17
2 23070 1 17
2 23071 1 17
2 23072 1 17
2 23073 1 17
2 23074 1 17
2 23075 1 17
2 23076 1 17
2 23077 1 17
2 23078 1 17
2 23079 1 17
2 23080 1 17
2 23081 1 17
2 23082 1 17
2 23083 1 17
2 23084 1 17
2 23085 1 17
2 23086 1 17
2 23087 1 17
2 23088 1 17
2 23089 1 17
2 23090 1 17
2 23091 1 17
2 23092 1 17
2 23093 1 17
2 23094 1 17
2 23095 1 17
2 23096 1 17
2 23097 1 17
2 23098 1 17
2 23099 1 17
2 23100 1 17
2 23101 1 17
2 23102 1 17
2 23103 1 17
2 23104 1 17
2 23105 1 17
2 23106 1 17
2 23107 1 17
2 23108 1 17
2 23109 1 17
2 23110 1 17
2 23111 1 17
2 23112 1 17
2 23113 1 17
2 23114 1 17
2 23115 1 17
2 23116 1 17
2 23117 1 17
2 23118 1 17
2 23119 1 17
2 23120 1 17
2 23121 1 17
2 23122 1 17
2 23123 1 17
2 23124 1 17
2 23125 1 17
2 23126 1 17
2 23127 1 17
2 23128 1 17
2 23129 1 17
2 23130 1 17
2 23131 1 17
2 23132 1 17
2 23133 1 17
2 23134 1 17
2 23135 1 17
2 23136 1 17
2 23137 1 17
2 23138 1 17
2 23139 1 17
2 23140 1 17
2 23141 1 17
2 23142 1 17
2 23143 1 17
2 23144 1 17
2 23145 1 17
2 23146 1 17
2 23147 1 17
2 23148 1 17
2 23149 1 17
2 23150 1 17
2 23151 1 17
2 23152 1 17
2 23153 1 17
2 23154 1 17
2 23155 1 17
1 18 0 85 0
2 23156 1 18
2 23157 1 18
2 23158 1 18
2 23159 1 18
2 23160 1 18
2 23161 1 18
2 23162 1 18
2 23163 1 18
2 23164 1 18
2 23165 1 18
2 23166 1 18
2 23167 1 18
2 23168 1 18
2 23169 1 18
2 23170 1 18
2 23171 1 18
2 23172 1 18
2 23173 1 18
2 23174 1 18
2 23175 1 18
2 23176 1 18
2 23177 1 18
2 23178 1 18
2 23179 1 18
2 23180 1 18
2 23181 1 18
2 23182 1 18
2 23183 1 18
2 23184 1 18
2 23185 1 18
2 23186 1 18
2 23187 1 18
2 23188 1 18
2 23189 1 18
2 23190 1 18
2 23191 1 18
2 23192 1 18
2 23193 1 18
2 23194 1 18
2 23195 1 18
2 23196 1 18
2 23197 1 18
2 23198 1 18
2 23199 1 18
2 23200 1 18
2 23201 1 18
2 23202 1 18
2 23203 1 18
2 23204 1 18
2 23205 1 18
2 23206 1 18
2 23207 1 18
2 23208 1 18
2 23209 1 18
2 23210 1 18
2 23211 1 18
2 23212 1 18
2 23213 1 18
2 23214 1 18
2 23215 1 18
2 23216 1 18
2 23217 1 18
2 23218 1 18
2 23219 1 18
2 23220 1 18
2 23221 1 18
2 23222 1 18
2 23223 1 18
2 23224 1 18
2 23225 1 18
2 23226 1 18
2 23227 1 18
2 23228 1 18
2 23229 1 18
2 23230 1 18
2 23231 1 18
2 23232 1 18
2 23233 1 18
2 23234 1 18
2 23235 1 18
2 23236 1 18
2 23237 1 18
2 23238 1 18
2 23239 1 18
2 23240 1 18
1 19 0 90 0
2 23241 1 19
2 23242 1 19
2 23243 1 19
2 23244 1 19
2 23245 1 19
2 23246 1 19
2 23247 1 19
2 23248 1 19
2 23249 1 19
2 23250 1 19
2 23251 1 19
2 23252 1 19
2 23253 1 19
2 23254 1 19
2 23255 1 19
2 23256 1 19
2 23257 1 19
2 23258 1 19
2 23259 1 19
2 23260 1 19
2 23261 1 19
2 23262 1 19
2 23263 1 19
2 23264 1 19
2 23265 1 19
2 23266 1 19
2 23267 1 19
2 23268 1 19
2 23269 1 19
2 23270 1 19
2 23271 1 19
2 23272 1 19
2 23273 1 19
2 23274 1 19
2 23275 1 19
2 23276 1 19
2 23277 1 19
2 23278 1 19
2 23279 1 19
2 23280 1 19
2 23281 1 19
2 23282 1 19
2 23283 1 19
2 23284 1 19
2 23285 1 19
2 23286 1 19
2 23287 1 19
2 23288 1 19
2 23289 1 19
2 23290 1 19
2 23291 1 19
2 23292 1 19
2 23293 1 19
2 23294 1 19
2 23295 1 19
2 23296 1 19
2 23297 1 19
2 23298 1 19
2 23299 1 19
2 23300 1 19
2 23301 1 19
2 23302 1 19
2 23303 1 19
2 23304 1 19
2 23305 1 19
2 23306 1 19
2 23307 1 19
2 23308 1 19
2 23309 1 19
2 23310 1 19
2 23311 1 19
2 23312 1 19
2 23313 1 19
2 23314 1 19
2 23315 1 19
2 23316 1 19
2 23317 1 19
2 23318 1 19
2 23319 1 19
2 23320 1 19
2 23321 1 19
2 23322 1 19
2 23323 1 19
2 23324 1 19
2 23325 1 19
2 23326 1 19
2 23327 1 19
2 23328 1 19
2 23329 1 19
2 23330 1 19
1 20 0 63 0
2 23331 1 20
2 23332 1 20
2 23333 1 20
2 23334 1 20
2 23335 1 20
2 23336 1 20
2 23337 1 20
2 23338 1 20
2 23339 1 20
2 23340 1 20
2 23341 1 20
2 23342 1 20
2 23343 1 20
2 23344 1 20
2 23345 1 20
2 23346 1 20
2 23347 1 20
2 23348 1 20
2 23349 1 20
2 23350 1 20
2 23351 1 20
2 23352 1 20
2 23353 1 20
2 23354 1 20
2 23355 1 20
2 23356 1 20
2 23357 1 20
2 23358 1 20
2 23359 1 20
2 23360 1 20
2 23361 1 20
2 23362 1 20
2 23363 1 20
2 23364 1 20
2 23365 1 20
2 23366 1 20
2 23367 1 20
2 23368 1 20
2 23369 1 20
2 23370 1 20
2 23371 1 20
2 23372 1 20
2 23373 1 20
2 23374 1 20
2 23375 1 20
2 23376 1 20
2 23377 1 20
2 23378 1 20
2 23379 1 20
2 23380 1 20
2 23381 1 20
2 23382 1 20
2 23383 1 20
2 23384 1 20
2 23385 1 20
2 23386 1 20
2 23387 1 20
2 23388 1 20
2 23389 1 20
2 23390 1 20
2 23391 1 20
2 23392 1 20
2 23393 1 20
1 21 0 88 0
2 23394 1 21
2 23395 1 21
2 23396 1 21
2 23397 1 21
2 23398 1 21
2 23399 1 21
2 23400 1 21
2 23401 1 21
2 23402 1 21
2 23403 1 21
2 23404 1 21
2 23405 1 21
2 23406 1 21
2 23407 1 21
2 23408 1 21
2 23409 1 21
2 23410 1 21
2 23411 1 21
2 23412 1 21
2 23413 1 21
2 23414 1 21
2 23415 1 21
2 23416 1 21
2 23417 1 21
2 23418 1 21
2 23419 1 21
2 23420 1 21
2 23421 1 21
2 23422 1 21
2 23423 1 21
2 23424 1 21
2 23425 1 21
2 23426 1 21
2 23427 1 21
2 23428 1 21
2 23429 1 21
2 23430 1 21
2 23431 1 21
2 23432 1 21
2 23433 1 21
2 23434 1 21
2 23435 1 21
2 23436 1 21
2 23437 1 21
2 23438 1 21
2 23439 1 21
2 23440 1 21
2 23441 1 21
2 23442 1 21
2 23443 1 21
2 23444 1 21
2 23445 1 21
2 23446 1 21
2 23447 1 21
2 23448 1 21
2 23449 1 21
2 23450 1 21
2 23451 1 21
2 23452 1 21
2 23453 1 21
2 23454 1 21
2 23455 1 21
2 23456 1 21
2 23457 1 21
2 23458 1 21
2 23459 1 21
2 23460 1 21
2 23461 1 21
2 23462 1 21
2 23463 1 21
2 23464 1 21
2 23465 1 21
2 23466 1 21
2 23467 1 21
2 23468 1 21
2 23469 1 21
2 23470 1 21
2 23471 1 21
2 23472 1 21
2 23473 1 21
2 23474 1 21
2 23475 1 21
2 23476 1 21
2 23477 1 21
2 23478 1 21
2 23479 1 21
2 23480 1 21
2 23481 1 21
1 22 0 109 0
2 23482 1 22
2 23483 1 22
2 23484 1 22
2 23485 1 22
2 23486 1 22
2 23487 1 22
2 23488 1 22
2 23489 1 22
2 23490 1 22
2 23491 1 22
2 23492 1 22
2 23493 1 22
2 23494 1 22
2 23495 1 22
2 23496 1 22
2 23497 1 22
2 23498 1 22
2 23499 1 22
2 23500 1 22
2 23501 1 22
2 23502 1 22
2 23503 1 22
2 23504 1 22
2 23505 1 22
2 23506 1 22
2 23507 1 22
2 23508 1 22
2 23509 1 22
2 23510 1 22
2 23511 1 22
2 23512 1 22
2 23513 1 22
2 23514 1 22
2 23515 1 22
2 23516 1 22
2 23517 1 22
2 23518 1 22
2 23519 1 22
2 23520 1 22
2 23521 1 22
2 23522 1 22
2 23523 1 22
2 23524 1 22
2 23525 1 22
2 23526 1 22
2 23527 1 22
2 23528 1 22
2 23529 1 22
2 23530 1 22
2 23531 1 22
2 23532 1 22
2 23533 1 22
2 23534 1 22
2 23535 1 22
2 23536 1 22
2 23537 1 22
2 23538 1 22
2 23539 1 22
2 23540 1 22
2 23541 1 22
2 23542 1 22
2 23543 1 22
2 23544 1 22
2 23545 1 22
2 23546 1 22
2 23547 1 22
2 23548 1 22
2 23549 1 22
2 23550 1 22
2 23551 1 22
2 23552 1 22
2 23553 1 22
2 23554 1 22
2 23555 1 22
2 23556 1 22
2 23557 1 22
2 23558 1 22
2 23559 1 22
2 23560 1 22
2 23561 1 22
2 23562 1 22
2 23563 1 22
2 23564 1 22
2 23565 1 22
2 23566 1 22
2 23567 1 22
2 23568 1 22
2 23569 1 22
2 23570 1 22
2 23571 1 22
2 23572 1 22
2 23573 1 22
2 23574 1 22
2 23575 1 22
2 23576 1 22
2 23577 1 22
2 23578 1 22
2 23579 1 22
2 23580 1 22
2 23581 1 22
2 23582 1 22
2 23583 1 22
2 23584 1 22
2 23585 1 22
2 23586 1 22
2 23587 1 22
2 23588 1 22
2 23589 1 22
2 23590 1 22
1 23 0 110 0
2 23591 1 23
2 23592 1 23
2 23593 1 23
2 23594 1 23
2 23595 1 23
2 23596 1 23
2 23597 1 23
2 23598 1 23
2 23599 1 23
2 23600 1 23
2 23601 1 23
2 23602 1 23
2 23603 1 23
2 23604 1 23
2 23605 1 23
2 23606 1 23
2 23607 1 23
2 23608 1 23
2 23609 1 23
2 23610 1 23
2 23611 1 23
2 23612 1 23
2 23613 1 23
2 23614 1 23
2 23615 1 23
2 23616 1 23
2 23617 1 23
2 23618 1 23
2 23619 1 23
2 23620 1 23
2 23621 1 23
2 23622 1 23
2 23623 1 23
2 23624 1 23
2 23625 1 23
2 23626 1 23
2 23627 1 23
2 23628 1 23
2 23629 1 23
2 23630 1 23
2 23631 1 23
2 23632 1 23
2 23633 1 23
2 23634 1 23
2 23635 1 23
2 23636 1 23
2 23637 1 23
2 23638 1 23
2 23639 1 23
2 23640 1 23
2 23641 1 23
2 23642 1 23
2 23643 1 23
2 23644 1 23
2 23645 1 23
2 23646 1 23
2 23647 1 23
2 23648 1 23
2 23649 1 23
2 23650 1 23
2 23651 1 23
2 23652 1 23
2 23653 1 23
2 23654 1 23
2 23655 1 23
2 23656 1 23
2 23657 1 23
2 23658 1 23
2 23659 1 23
2 23660 1 23
2 23661 1 23
2 23662 1 23
2 23663 1 23
2 23664 1 23
2 23665 1 23
2 23666 1 23
2 23667 1 23
2 23668 1 23
2 23669 1 23
2 23670 1 23
2 23671 1 23
2 23672 1 23
2 23673 1 23
2 23674 1 23
2 23675 1 23
2 23676 1 23
2 23677 1 23
2 23678 1 23
2 23679 1 23
2 23680 1 23
2 23681 1 23
2 23682 1 23
2 23683 1 23
2 23684 1 23
2 23685 1 23
2 23686 1 23
2 23687 1 23
2 23688 1 23
2 23689 1 23
2 23690 1 23
2 23691 1 23
2 23692 1 23
2 23693 1 23
2 23694 1 23
2 23695 1 23
2 23696 1 23
2 23697 1 23
2 23698 1 23
2 23699 1 23
2 23700 1 23
1 24 0 71 0
2 23701 1 24
2 23702 1 24
2 23703 1 24
2 23704 1 24
2 23705 1 24
2 23706 1 24
2 23707 1 24
2 23708 1 24
2 23709 1 24
2 23710 1 24
2 23711 1 24
2 23712 1 24
2 23713 1 24
2 23714 1 24
2 23715 1 24
2 23716 1 24
2 23717 1 24
2 23718 1 24
2 23719 1 24
2 23720 1 24
2 23721 1 24
2 23722 1 24
2 23723 1 24
2 23724 1 24
2 23725 1 24
2 23726 1 24
2 23727 1 24
2 23728 1 24
2 23729 1 24
2 23730 1 24
2 23731 1 24
2 23732 1 24
2 23733 1 24
2 23734 1 24
2 23735 1 24
2 23736 1 24
2 23737 1 24
2 23738 1 24
2 23739 1 24
2 23740 1 24
2 23741 1 24
2 23742 1 24
2 23743 1 24
2 23744 1 24
2 23745 1 24
2 23746 1 24
2 23747 1 24
2 23748 1 24
2 23749 1 24
2 23750 1 24
2 23751 1 24
2 23752 1 24
2 23753 1 24
2 23754 1 24
2 23755 1 24
2 23756 1 24
2 23757 1 24
2 23758 1 24
2 23759 1 24
2 23760 1 24
2 23761 1 24
2 23762 1 24
2 23763 1 24
2 23764 1 24
2 23765 1 24
2 23766 1 24
2 23767 1 24
2 23768 1 24
2 23769 1 24
2 23770 1 24
2 23771 1 24
2 23772 1 27
2 23773 1 27
2 23774 1 27
2 23775 1 27
2 23776 1 27
2 23777 1 27
2 23778 1 27
2 23779 1 27
2 23780 1 27
2 23781 1 27
2 23782 1 27
2 23783 1 27
2 23784 1 27
2 23785 1 27
2 23786 1 27
2 23787 1 27
2 23788 1 27
2 23789 1 27
2 23790 1 27
2 23791 1 27
2 23792 1 27
2 23793 1 27
2 23794 1 27
2 23795 1 27
2 23796 1 27
2 23797 1 27
2 23798 1 27
2 23799 1 27
2 23800 1 27
2 23801 1 27
2 23802 1 27
2 23803 1 27
2 23804 1 27
2 23805 1 27
2 23806 1 27
2 23807 1 27
2 23808 1 27
2 23809 1 27
2 23810 1 27
2 23811 1 27
2 23812 1 27
2 23813 1 27
2 23814 1 27
2 23815 1 27
2 23816 1 27
2 23817 1 27
2 23818 1 27
2 23819 1 27
2 23820 1 27
2 23821 1 27
2 23822 1 27
2 23823 1 27
2 23824 1 27
2 23825 1 27
2 23826 1 27
2 23827 1 27
2 23828 1 27
2 23829 1 27
2 23830 1 27
2 23831 1 27
2 23832 1 27
2 23833 1 27
2 23834 1 27
2 23835 1 27
2 23836 1 27
2 23837 1 27
2 23838 1 27
2 23839 1 27
2 23840 1 27
2 23841 1 27
2 23842 1 27
2 23843 1 27
2 23844 1 27
2 23845 1 27
2 23846 1 27
2 23847 1 27
2 23848 1 27
2 23849 1 27
2 23850 1 27
2 23851 1 27
2 23852 1 27
2 23853 1 27
2 23854 1 27
2 23855 1 27
2 23856 1 27
2 23857 1 27
2 23858 1 27
2 23859 1 27
2 23860 1 27
2 23861 1 27
2 23862 1 27
2 23863 1 27
2 23864 1 27
2 23865 1 27
2 23866 1 27
2 23867 1 27
2 23868 1 27
2 23869 1 27
2 23870 1 27
2 23871 1 27
2 23872 1 27
2 23873 1 27
2 23874 1 27
2 23875 1 27
2 23876 1 27
2 23877 1 27
2 23878 1 27
2 23879 1 27
2 23880 1 27
2 23881 1 27
2 23882 1 27
2 23883 1 27
2 23884 1 27
2 23885 1 27
2 23886 1 27
2 23887 1 27
2 23888 1 27
2 23889 1 27
2 23890 1 27
2 23891 1 27
2 23892 1 28
2 23893 1 28
2 23894 1 28
2 23895 1 28
2 23896 1 28
2 23897 1 28
2 23898 1 28
2 23899 1 28
2 23900 1 28
2 23901 1 28
2 23902 1 28
2 23903 1 28
2 23904 1 28
2 23905 1 28
2 23906 1 28
2 23907 1 28
2 23908 1 28
2 23909 1 28
2 23910 1 28
2 23911 1 28
2 23912 1 28
2 23913 1 28
2 23914 1 28
2 23915 1 28
2 23916 1 28
2 23917 1 28
2 23918 1 28
2 23919 1 28
2 23920 1 28
2 23921 1 28
2 23922 1 28
2 23923 1 28
2 23924 1 28
2 23925 1 28
2 23926 1 28
2 23927 1 28
2 23928 1 28
2 23929 1 28
2 23930 1 28
2 23931 1 28
2 23932 1 28
2 23933 1 28
2 23934 1 28
2 23935 1 28
2 23936 1 28
2 23937 1 28
2 23938 1 28
2 23939 1 28
2 23940 1 28
2 23941 1 28
2 23942 1 28
2 23943 1 28
2 23944 1 28
2 23945 1 28
2 23946 1 28
2 23947 1 28
2 23948 1 28
2 23949 1 28
2 23950 1 28
2 23951 1 28
2 23952 1 28
2 23953 1 28
2 23954 1 28
2 23955 1 28
2 23956 1 28
2 23957 1 28
2 23958 1 28
2 23959 1 28
2 23960 1 28
2 23961 1 28
2 23962 1 28
2 23963 1 28
2 23964 1 28
2 23965 1 28
2 23966 1 28
2 23967 1 28
2 23968 1 28
2 23969 1 28
2 23970 1 28
2 23971 1 28
2 23972 1 28
2 23973 1 28
2 23974 1 28
2 23975 1 28
2 23976 1 28
2 23977 1 28
2 23978 1 28
2 23979 1 28
2 23980 1 28
2 23981 1 28
2 23982 1 28
2 23983 1 28
2 23984 1 28
2 23985 1 28
2 23986 1 28
2 23987 1 28
2 23988 1 28
2 23989 1 28
2 23990 1 28
2 23991 1 28
2 23992 1 28
2 23993 1 28
2 23994 1 28
2 23995 1 28
2 23996 1 28
2 23997 1 28
2 23998 1 28
2 23999 1 28
2 24000 1 28
2 24001 1 28
2 24002 1 28
2 24003 1 28
2 24004 1 28
2 24005 1 28
2 24006 1 28
2 24007 1 29
2 24008 1 29
2 24009 1 29
2 24010 1 29
2 24011 1 29
2 24012 1 29
2 24013 1 29
2 24014 1 29
2 24015 1 29
2 24016 1 29
2 24017 1 29
2 24018 1 29
2 24019 1 29
2 24020 1 29
2 24021 1 29
2 24022 1 29
2 24023 1 29
2 24024 1 29
2 24025 1 29
2 24026 1 29
2 24027 1 29
2 24028 1 29
2 24029 1 29
2 24030 1 29
2 24031 1 29
2 24032 1 29
2 24033 1 29
2 24034 1 29
2 24035 1 29
2 24036 1 29
2 24037 1 29
2 24038 1 29
2 24039 1 29
2 24040 1 29
2 24041 1 29
2 24042 1 29
2 24043 1 29
2 24044 1 29
2 24045 1 29
2 24046 1 29
2 24047 1 29
2 24048 1 29
2 24049 1 29
2 24050 1 29
2 24051 1 29
2 24052 1 29
2 24053 1 29
2 24054 1 29
2 24055 1 29
2 24056 1 29
2 24057 1 29
2 24058 1 29
2 24059 1 29
2 24060 1 29
2 24061 1 29
2 24062 1 29
2 24063 1 29
2 24064 1 29
2 24065 1 29
2 24066 1 29
2 24067 1 29
2 24068 1 29
2 24069 1 29
2 24070 1 29
2 24071 1 29
2 24072 1 29
2 24073 1 29
2 24074 1 29
2 24075 1 29
2 24076 1 29
2 24077 1 29
2 24078 1 29
2 24079 1 29
2 24080 1 29
2 24081 1 29
2 24082 1 29
2 24083 1 29
2 24084 1 29
2 24085 1 29
2 24086 1 29
2 24087 1 29
2 24088 1 29
2 24089 1 29
2 24090 1 29
2 24091 1 29
2 24092 1 29
2 24093 1 29
2 24094 1 29
2 24095 1 29
2 24096 1 29
2 24097 1 29
2 24098 1 29
2 24099 1 29
2 24100 1 29
2 24101 1 29
2 24102 1 29
2 24103 1 29
2 24104 1 29
2 24105 1 29
2 24106 1 29
2 24107 1 29
2 24108 1 29
2 24109 1 29
2 24110 1 29
2 24111 1 29
2 24112 1 29
2 24113 1 29
2 24114 1 29
2 24115 1 29
2 24116 1 29
2 24117 1 29
2 24118 1 29
2 24119 1 29
2 24120 1 29
2 24121 1 29
2 24122 1 29
2 24123 1 29
2 24124 1 29
2 24125 1 29
2 24126 1 29
2 24127 1 29
2 24128 1 29
2 24129 1 29
2 24130 1 29
2 24131 1 29
2 24132 1 29
2 24133 1 29
2 24134 1 29
2 24135 1 30
2 24136 1 30
2 24137 1 30
2 24138 1 30
2 24139 1 30
2 24140 1 30
2 24141 1 30
2 24142 1 30
2 24143 1 30
2 24144 1 30
2 24145 1 30
2 24146 1 30
2 24147 1 30
2 24148 1 30
2 24149 1 30
2 24150 1 30
2 24151 1 30
2 24152 1 30
2 24153 1 30
2 24154 1 30
2 24155 1 30
2 24156 1 30
2 24157 1 30
2 24158 1 30
2 24159 1 30
2 24160 1 30
2 24161 1 30
2 24162 1 30
2 24163 1 30
2 24164 1 30
2 24165 1 30
2 24166 1 30
2 24167 1 30
2 24168 1 30
2 24169 1 30
2 24170 1 30
2 24171 1 30
2 24172 1 30
2 24173 1 30
2 24174 1 30
2 24175 1 30
2 24176 1 30
2 24177 1 30
2 24178 1 30
2 24179 1 30
2 24180 1 30
2 24181 1 31
2 24182 1 31
2 24183 1 31
2 24184 1 31
2 24185 1 31
2 24186 1 31
2 24187 1 31
2 24188 1 31
2 24189 1 31
2 24190 1 31
2 24191 1 31
2 24192 1 31
2 24193 1 31
2 24194 1 31
2 24195 1 31
2 24196 1 31
2 24197 1 31
2 24198 1 31
2 24199 1 31
2 24200 1 31
2 24201 1 31
2 24202 1 31
2 24203 1 31
2 24204 1 31
2 24205 1 31
2 24206 1 31
2 24207 1 31
2 24208 1 31
2 24209 1 31
2 24210 1 31
2 24211 1 31
2 24212 1 31
2 24213 1 31
2 24214 1 31
2 24215 1 31
2 24216 1 31
2 24217 1 31
2 24218 1 31
2 24219 1 31
2 24220 1 31
2 24221 1 31
2 24222 1 31
2 24223 1 31
2 24224 1 31
2 24225 1 31
2 24226 1 31
2 24227 1 31
2 24228 1 31
2 24229 1 31
2 24230 1 31
2 24231 1 31
2 24232 1 31
2 24233 1 31
2 24234 1 31
2 24235 1 31
2 24236 1 31
2 24237 1 31
2 24238 1 31
2 24239 1 31
2 24240 1 31
2 24241 1 31
2 24242 1 31
2 24243 1 31
2 24244 1 31
2 24245 1 31
2 24246 1 31
2 24247 1 31
2 24248 1 31
2 24249 1 31
2 24250 1 31
2 24251 1 31
2 24252 1 31
2 24253 1 31
2 24254 1 31
2 24255 1 32
2 24256 1 32
2 24257 1 32
2 24258 1 32
2 24259 1 32
2 24260 1 32
2 24261 1 32
2 24262 1 32
2 24263 1 32
2 24264 1 32
2 24265 1 32
2 24266 1 32
2 24267 1 32
2 24268 1 32
2 24269 1 32
2 24270 1 32
2 24271 1 32
2 24272 1 32
2 24273 1 32
2 24274 1 32
2 24275 1 32
2 24276 1 32
2 24277 1 32
2 24278 1 32
2 24279 1 32
2 24280 1 32
2 24281 1 32
2 24282 1 32
2 24283 1 32
2 24284 1 32
2 24285 1 32
2 24286 1 32
2 24287 1 32
2 24288 1 32
2 24289 1 32
2 24290 1 32
2 24291 1 32
2 24292 1 32
2 24293 1 32
2 24294 1 32
2 24295 1 32
2 24296 1 32
2 24297 1 32
2 24298 1 32
2 24299 1 32
2 24300 1 33
2 24301 1 33
2 24302 1 33
2 24303 1 33
2 24304 1 33
2 24305 1 33
2 24306 1 33
2 24307 1 33
2 24308 1 33
2 24309 1 33
2 24310 1 33
2 24311 1 33
2 24312 1 33
2 24313 1 33
2 24314 1 33
2 24315 1 33
2 24316 1 33
2 24317 1 33
2 24318 1 33
2 24319 1 33
2 24320 1 33
2 24321 1 33
2 24322 1 33
2 24323 1 33
2 24324 1 33
2 24325 1 33
2 24326 1 33
2 24327 1 33
2 24328 1 33
2 24329 1 33
2 24330 1 33
2 24331 1 33
2 24332 1 33
2 24333 1 33
2 24334 1 33
2 24335 1 33
2 24336 1 33
2 24337 1 33
2 24338 1 33
2 24339 1 33
2 24340 1 33
2 24341 1 33
2 24342 1 33
2 24343 1 33
2 24344 1 33
2 24345 1 33
2 24346 1 33
2 24347 1 33
2 24348 1 33
2 24349 1 33
2 24350 1 33
2 24351 1 33
2 24352 1 33
2 24353 1 33
2 24354 1 33
2 24355 1 33
2 24356 1 34
2 24357 1 34
2 24358 1 34
2 24359 1 34
2 24360 1 34
2 24361 1 34
2 24362 1 34
2 24363 1 34
2 24364 1 34
2 24365 1 34
2 24366 1 34
2 24367 1 34
2 24368 1 34
2 24369 1 34
2 24370 1 34
2 24371 1 34
2 24372 1 34
2 24373 1 34
2 24374 1 34
2 24375 1 34
2 24376 1 34
2 24377 1 34
2 24378 1 34
2 24379 1 34
2 24380 1 34
2 24381 1 34
2 24382 1 34
2 24383 1 34
2 24384 1 34
2 24385 1 34
2 24386 1 34
2 24387 1 34
2 24388 1 34
2 24389 1 34
2 24390 1 34
2 24391 1 34
2 24392 1 34
2 24393 1 34
2 24394 1 34
2 24395 1 34
2 24396 1 34
2 24397 1 34
2 24398 1 34
2 24399 1 34
2 24400 1 34
2 24401 1 34
2 24402 1 34
2 24403 1 34
2 24404 1 34
2 24405 1 34
2 24406 1 34
2 24407 1 34
2 24408 1 34
2 24409 1 34
2 24410 1 34
2 24411 1 34
2 24412 1 34
2 24413 1 34
2 24414 1 34
2 24415 1 34
2 24416 1 34
2 24417 1 34
2 24418 1 34
2 24419 1 34
2 24420 1 34
2 24421 1 34
2 24422 1 34
2 24423 1 34
2 24424 1 34
2 24425 1 34
2 24426 1 34
2 24427 1 35
2 24428 1 35
2 24429 1 35
2 24430 1 35
2 24431 1 35
2 24432 1 35
2 24433 1 35
2 24434 1 35
2 24435 1 35
2 24436 1 35
2 24437 1 35
2 24438 1 35
2 24439 1 35
2 24440 1 35
2 24441 1 35
2 24442 1 35
2 24443 1 35
2 24444 1 35
2 24445 1 35
2 24446 1 35
2 24447 1 35
2 24448 1 35
2 24449 1 35
2 24450 1 35
2 24451 1 35
2 24452 1 35
2 24453 1 35
2 24454 1 35
2 24455 1 35
2 24456 1 35
2 24457 1 35
2 24458 1 35
2 24459 1 35
2 24460 1 35
2 24461 1 35
2 24462 1 35
2 24463 1 35
2 24464 1 35
2 24465 1 35
2 24466 1 35
2 24467 1 35
2 24468 1 35
2 24469 1 35
2 24470 1 35
2 24471 1 35
2 24472 1 35
2 24473 1 35
2 24474 1 35
2 24475 1 35
2 24476 1 35
2 24477 1 35
2 24478 1 35
2 24479 1 35
2 24480 1 35
2 24481 1 35
2 24482 1 35
2 24483 1 35
2 24484 1 35
2 24485 1 35
2 24486 1 35
2 24487 1 35
2 24488 1 35
2 24489 1 36
2 24490 1 36
2 24491 1 36
2 24492 1 36
2 24493 1 36
2 24494 1 36
2 24495 1 36
2 24496 1 36
2 24497 1 36
2 24498 1 36
2 24499 1 36
2 24500 1 36
2 24501 1 36
2 24502 1 36
2 24503 1 36
2 24504 1 36
2 24505 1 36
2 24506 1 36
2 24507 1 36
2 24508 1 36
2 24509 1 36
2 24510 1 36
2 24511 1 36
2 24512 1 36
2 24513 1 36
2 24514 1 36
2 24515 1 36
2 24516 1 36
2 24517 1 36
2 24518 1 36
2 24519 1 36
2 24520 1 36
2 24521 1 36
2 24522 1 36
2 24523 1 36
2 24524 1 36
2 24525 1 36
2 24526 1 36
2 24527 1 36
2 24528 1 36
2 24529 1 36
2 24530 1 36
2 24531 1 36
2 24532 1 36
2 24533 1 36
2 24534 1 36
2 24535 1 36
2 24536 1 36
2 24537 1 36
2 24538 1 36
2 24539 1 36
2 24540 1 36
2 24541 1 36
2 24542 1 36
2 24543 1 36
2 24544 1 36
2 24545 1 36
2 24546 1 36
2 24547 1 36
2 24548 1 36
2 24549 1 37
2 24550 1 37
2 24551 1 37
2 24552 1 37
2 24553 1 37
2 24554 1 37
2 24555 1 37
2 24556 1 37
2 24557 1 37
2 24558 1 37
2 24559 1 37
2 24560 1 37
2 24561 1 37
2 24562 1 37
2 24563 1 37
2 24564 1 37
2 24565 1 37
2 24566 1 37
2 24567 1 37
2 24568 1 37
2 24569 1 37
2 24570 1 37
2 24571 1 37
2 24572 1 37
2 24573 1 37
2 24574 1 37
2 24575 1 37
2 24576 1 37
2 24577 1 37
2 24578 1 37
2 24579 1 37
2 24580 1 37
2 24581 1 37
2 24582 1 37
2 24583 1 37
2 24584 1 37
2 24585 1 37
2 24586 1 37
2 24587 1 37
2 24588 1 37
2 24589 1 37
2 24590 1 37
2 24591 1 37
2 24592 1 37
2 24593 1 37
2 24594 1 37
2 24595 1 37
2 24596 1 37
2 24597 1 37
2 24598 1 37
2 24599 1 37
2 24600 1 37
2 24601 1 37
2 24602 1 37
2 24603 1 37
2 24604 1 37
2 24605 1 37
2 24606 1 37
2 24607 1 37
2 24608 1 37
2 24609 1 37
2 24610 1 37
2 24611 1 37
2 24612 1 37
2 24613 1 37
2 24614 1 37
2 24615 1 37
2 24616 1 37
2 24617 1 37
2 24618 1 37
2 24619 1 37
2 24620 1 37
2 24621 1 37
2 24622 1 37
2 24623 1 37
2 24624 1 37
2 24625 1 37
2 24626 1 37
2 24627 1 37
2 24628 1 37
2 24629 1 37
2 24630 1 37
2 24631 1 37
2 24632 1 37
2 24633 1 37
2 24634 1 37
2 24635 1 38
2 24636 1 38
2 24637 1 38
2 24638 1 38
2 24639 1 38
2 24640 1 38
2 24641 1 38
2 24642 1 38
2 24643 1 38
2 24644 1 38
2 24645 1 38
2 24646 1 38
2 24647 1 38
2 24648 1 38
2 24649 1 38
2 24650 1 38
2 24651 1 38
2 24652 1 38
2 24653 1 38
2 24654 1 38
2 24655 1 38
2 24656 1 38
2 24657 1 38
2 24658 1 38
2 24659 1 38
2 24660 1 38
2 24661 1 38
2 24662 1 38
2 24663 1 38
2 24664 1 38
2 24665 1 39
2 24666 1 39
2 24667 1 39
2 24668 1 39
2 24669 1 39
2 24670 1 39
2 24671 1 39
2 24672 1 39
2 24673 1 39
2 24674 1 39
2 24675 1 39
2 24676 1 39
2 24677 1 39
2 24678 1 39
2 24679 1 39
2 24680 1 39
2 24681 1 39
2 24682 1 39
2 24683 1 39
2 24684 1 39
2 24685 1 39
2 24686 1 39
2 24687 1 39
2 24688 1 39
2 24689 1 39
2 24690 1 39
2 24691 1 39
2 24692 1 39
2 24693 1 39
2 24694 1 39
2 24695 1 39
2 24696 1 39
2 24697 1 39
2 24698 1 39
2 24699 1 39
2 24700 1 39
2 24701 1 39
2 24702 1 39
2 24703 1 39
2 24704 1 39
2 24705 1 39
2 24706 1 39
2 24707 1 39
2 24708 1 39
2 24709 1 39
2 24710 1 39
2 24711 1 39
2 24712 1 39
2 24713 1 39
2 24714 1 39
2 24715 1 39
2 24716 1 39
2 24717 1 39
2 24718 1 39
2 24719 1 39
2 24720 1 39
2 24721 1 39
2 24722 1 39
2 24723 1 39
2 24724 1 39
2 24725 1 39
2 24726 1 39
2 24727 1 39
2 24728 1 39
2 24729 1 39
2 24730 1 40
2 24731 1 40
2 24732 1 40
2 24733 1 40
2 24734 1 40
2 24735 1 40
2 24736 1 40
2 24737 1 40
2 24738 1 40
2 24739 1 40
2 24740 1 40
2 24741 1 40
2 24742 1 40
2 24743 1 40
2 24744 1 40
2 24745 1 40
2 24746 1 40
2 24747 1 40
2 24748 1 40
2 24749 1 40
2 24750 1 40
2 24751 1 40
2 24752 1 40
2 24753 1 40
2 24754 1 40
2 24755 1 40
2 24756 1 40
2 24757 1 40
2 24758 1 40
2 24759 1 40
2 24760 1 40
2 24761 1 40
2 24762 1 40
2 24763 1 40
2 24764 1 40
2 24765 1 40
2 24766 1 40
2 24767 1 40
2 24768 1 40
2 24769 1 41
2 24770 1 41
2 24771 1 41
2 24772 1 41
2 24773 1 41
2 24774 1 41
2 24775 1 41
2 24776 1 41
2 24777 1 41
2 24778 1 41
2 24779 1 41
2 24780 1 41
2 24781 1 41
2 24782 1 41
2 24783 1 41
2 24784 1 41
2 24785 1 41
2 24786 1 41
2 24787 1 41
2 24788 1 41
2 24789 1 41
2 24790 1 41
2 24791 1 41
2 24792 1 41
2 24793 1 41
2 24794 1 41
2 24795 1 41
2 24796 1 41
2 24797 1 41
2 24798 1 41
2 24799 1 41
2 24800 1 41
2 24801 1 41
2 24802 1 41
2 24803 1 41
2 24804 1 41
2 24805 1 41
2 24806 1 41
2 24807 1 41
2 24808 1 41
2 24809 1 41
2 24810 1 41
2 24811 1 41
2 24812 1 41
2 24813 1 41
2 24814 1 41
2 24815 1 41
2 24816 1 41
2 24817 1 41
2 24818 1 41
2 24819 1 41
2 24820 1 41
2 24821 1 41
2 24822 1 41
2 24823 1 41
2 24824 1 41
2 24825 1 41
2 24826 1 41
2 24827 1 42
2 24828 1 42
2 24829 1 42
2 24830 1 42
2 24831 1 42
2 24832 1 42
2 24833 1 42
2 24834 1 42
2 24835 1 42
2 24836 1 42
2 24837 1 42
2 24838 1 42
2 24839 1 42
2 24840 1 42
2 24841 1 42
2 24842 1 42
2 24843 1 42
2 24844 1 42
2 24845 1 42
2 24846 1 42
2 24847 1 42
2 24848 1 42
2 24849 1 42
2 24850 1 42
2 24851 1 42
2 24852 1 42
2 24853 1 42
2 24854 1 42
2 24855 1 42
2 24856 1 42
2 24857 1 42
2 24858 1 42
2 24859 1 42
2 24860 1 42
2 24861 1 42
2 24862 1 42
2 24863 1 42
2 24864 1 42
2 24865 1 42
2 24866 1 42
2 24867 1 42
2 24868 1 42
2 24869 1 42
2 24870 1 42
2 24871 1 42
2 24872 1 42
2 24873 1 42
2 24874 1 42
2 24875 1 42
2 24876 1 42
2 24877 1 42
2 24878 1 42
2 24879 1 42
2 24880 1 42
2 24881 1 42
2 24882 1 42
2 24883 1 42
2 24884 1 42
2 24885 1 42
2 24886 1 42
2 24887 1 42
2 24888 1 43
2 24889 1 43
2 24890 1 43
2 24891 1 43
2 24892 1 43
2 24893 1 43
2 24894 1 43
2 24895 1 43
2 24896 1 43
2 24897 1 43
2 24898 1 43
2 24899 1 43
2 24900 1 43
2 24901 1 43
2 24902 1 43
2 24903 1 43
2 24904 1 43
2 24905 1 43
2 24906 1 43
2 24907 1 43
2 24908 1 43
2 24909 1 43
2 24910 1 43
2 24911 1 43
2 24912 1 43
2 24913 1 43
2 24914 1 43
2 24915 1 43
2 24916 1 43
2 24917 1 43
2 24918 1 43
2 24919 1 43
2 24920 1 43
2 24921 1 43
2 24922 1 43
2 24923 1 43
2 24924 1 43
2 24925 1 43
2 24926 1 43
2 24927 1 43
2 24928 1 43
2 24929 1 43
2 24930 1 43
2 24931 1 43
2 24932 1 43
2 24933 1 43
2 24934 1 43
2 24935 1 43
2 24936 1 43
2 24937 1 43
2 24938 1 43
2 24939 1 43
2 24940 1 43
2 24941 1 43
2 24942 1 43
2 24943 1 43
2 24944 1 43
2 24945 1 43
2 24946 1 43
2 24947 1 43
2 24948 1 43
2 24949 1 43
2 24950 1 43
2 24951 1 43
2 24952 1 43
2 24953 1 43
2 24954 1 43
2 24955 1 43
2 24956 1 43
2 24957 1 43
2 24958 1 43
2 24959 1 43
2 24960 1 43
2 24961 1 43
2 24962 1 43
2 24963 1 43
2 24964 1 43
2 24965 1 43
2 24966 1 43
2 24967 1 43
2 24968 1 43
2 24969 1 43
2 24970 1 43
2 24971 1 43
2 24972 1 43
2 24973 1 43
2 24974 1 43
2 24975 1 43
2 24976 1 43
2 24977 1 43
2 24978 1 43
2 24979 1 43
2 24980 1 43
2 24981 1 43
2 24982 1 43
2 24983 1 43
2 24984 1 43
2 24985 1 43
2 24986 1 43
2 24987 1 43
2 24988 1 43
2 24989 1 43
2 24990 1 43
2 24991 1 43
2 24992 1 43
2 24993 1 43
2 24994 1 43
2 24995 1 43
2 24996 1 44
2 24997 1 44
2 24998 1 44
2 24999 1 44
2 25000 1 44
2 25001 1 44
2 25002 1 44
2 25003 1 44
2 25004 1 44
2 25005 1 44
2 25006 1 44
2 25007 1 44
2 25008 1 44
2 25009 1 44
2 25010 1 44
2 25011 1 44
2 25012 1 44
2 25013 1 44
2 25014 1 44
2 25015 1 44
2 25016 1 44
2 25017 1 44
2 25018 1 44
2 25019 1 44
2 25020 1 44
2 25021 1 44
2 25022 1 44
2 25023 1 44
2 25024 1 44
2 25025 1 44
2 25026 1 44
2 25027 1 44
2 25028 1 44
2 25029 1 44
2 25030 1 44
2 25031 1 44
2 25032 1 44
2 25033 1 44
2 25034 1 44
2 25035 1 44
2 25036 1 44
2 25037 1 44
2 25038 1 44
2 25039 1 44
2 25040 1 44
2 25041 1 44
2 25042 1 44
2 25043 1 44
2 25044 1 44
2 25045 1 44
2 25046 1 44
2 25047 1 44
2 25048 1 44
2 25049 1 44
2 25050 1 44
2 25051 1 44
2 25052 1 44
2 25053 1 44
2 25054 1 44
2 25055 1 44
2 25056 1 44
2 25057 1 44
2 25058 1 44
2 25059 1 44
2 25060 1 44
2 25061 1 44
2 25062 1 44
2 25063 1 44
2 25064 1 44
2 25065 1 44
2 25066 1 44
2 25067 1 44
2 25068 1 44
2 25069 1 44
2 25070 1 44
2 25071 1 44
2 25072 1 44
2 25073 1 44
2 25074 1 44
2 25075 1 44
2 25076 1 44
2 25077 1 44
2 25078 1 44
2 25079 1 44
2 25080 1 44
2 25081 1 44
2 25082 1 44
2 25083 1 44
2 25084 1 44
2 25085 1 44
2 25086 1 44
2 25087 1 44
2 25088 1 44
2 25089 1 44
2 25090 1 44
2 25091 1 44
2 25092 1 44
2 25093 1 44
2 25094 1 44
2 25095 1 44
2 25096 1 44
2 25097 1 44
2 25098 1 44
2 25099 1 44
2 25100 1 44
2 25101 1 44
2 25102 1 44
2 25103 1 44
2 25104 1 44
2 25105 1 44
2 25106 1 44
2 25107 1 44
2 25108 1 44
2 25109 1 44
2 25110 1 44
2 25111 1 44
2 25112 1 44
2 25113 1 44
2 25114 1 44
2 25115 1 44
2 25116 1 45
2 25117 1 45
2 25118 1 45
2 25119 1 45
2 25120 1 45
2 25121 1 45
2 25122 1 45
2 25123 1 45
2 25124 1 45
2 25125 1 45
2 25126 1 45
2 25127 1 45
2 25128 1 45
2 25129 1 45
2 25130 1 45
2 25131 1 45
2 25132 1 45
2 25133 1 45
2 25134 1 45
2 25135 1 45
2 25136 1 45
2 25137 1 45
2 25138 1 45
2 25139 1 45
2 25140 1 45
2 25141 1 45
2 25142 1 45
2 25143 1 45
2 25144 1 45
2 25145 1 45
2 25146 1 45
2 25147 1 45
2 25148 1 45
2 25149 1 45
2 25150 1 45
2 25151 1 45
2 25152 1 45
2 25153 1 45
2 25154 1 45
2 25155 1 45
2 25156 1 45
2 25157 1 45
2 25158 1 45
2 25159 1 45
2 25160 1 45
2 25161 1 45
2 25162 1 45
2 25163 1 45
2 25164 1 45
2 25165 1 45
2 25166 1 45
2 25167 1 45
2 25168 1 45
2 25169 1 45
2 25170 1 45
2 25171 1 45
2 25172 1 45
2 25173 1 45
2 25174 1 45
2 25175 1 45
2 25176 1 45
2 25177 1 45
2 25178 1 45
2 25179 1 45
2 25180 1 45
2 25181 1 45
2 25182 1 45
2 25183 1 45
2 25184 1 45
2 25185 1 45
2 25186 1 45
2 25187 1 45
2 25188 1 45
2 25189 1 45
2 25190 1 45
2 25191 1 45
2 25192 1 45
2 25193 1 45
2 25194 1 45
2 25195 1 45
2 25196 1 45
2 25197 1 46
2 25198 1 46
2 25199 1 46
2 25200 1 46
2 25201 1 46
2 25202 1 46
2 25203 1 46
2 25204 1 46
2 25205 1 46
2 25206 1 46
2 25207 1 46
2 25208 1 46
2 25209 1 46
2 25210 1 46
2 25211 1 46
2 25212 1 46
2 25213 1 46
2 25214 1 46
2 25215 1 46
2 25216 1 46
2 25217 1 46
2 25218 1 46
2 25219 1 46
2 25220 1 46
2 25221 1 46
2 25222 1 46
2 25223 1 46
2 25224 1 46
2 25225 1 46
2 25226 1 46
2 25227 1 46
2 25228 1 46
2 25229 1 46
2 25230 1 46
2 25231 1 46
2 25232 1 46
2 25233 1 46
2 25234 1 46
2 25235 1 46
2 25236 1 46
2 25237 1 46
2 25238 1 46
2 25239 1 46
2 25240 1 46
2 25241 1 46
2 25242 1 46
2 25243 1 46
2 25244 1 46
2 25245 1 46
2 25246 1 46
2 25247 1 46
2 25248 1 46
2 25249 1 46
2 25250 1 46
2 25251 1 46
2 25252 1 46
2 25253 1 46
2 25254 1 46
2 25255 1 46
2 25256 1 46
2 25257 1 46
2 25258 1 46
2 25259 1 46
2 25260 1 46
2 25261 1 46
2 25262 1 46
2 25263 1 46
2 25264 1 46
2 25265 1 46
2 25266 1 46
2 25267 1 46
2 25268 1 46
2 25269 1 46
2 25270 1 46
2 25271 1 46
2 25272 1 46
2 25273 1 46
2 25274 1 46
2 25275 1 46
2 25276 1 46
2 25277 1 46
2 25278 1 46
2 25279 1 46
2 25280 1 46
2 25281 1 46
2 25282 1 46
2 25283 1 46
2 25284 1 46
2 25285 1 46
2 25286 1 46
2 25287 1 46
2 25288 1 46
2 25289 1 46
2 25290 1 46
2 25291 1 46
2 25292 1 47
2 25293 1 47
2 25294 1 47
2 25295 1 47
2 25296 1 47
2 25297 1 47
2 25298 1 47
2 25299 1 47
2 25300 1 47
2 25301 1 47
2 25302 1 47
2 25303 1 47
2 25304 1 47
2 25305 1 47
2 25306 1 47
2 25307 1 47
2 25308 1 47
2 25309 1 47
2 25310 1 47
2 25311 1 47
2 25312 1 47
2 25313 1 47
2 25314 1 47
2 25315 1 47
2 25316 1 47
2 25317 1 47
2 25318 1 47
2 25319 1 47
2 25320 1 47
2 25321 1 47
2 25322 1 47
2 25323 1 47
2 25324 1 47
2 25325 1 47
2 25326 1 47
2 25327 1 47
2 25328 1 47
2 25329 1 47
2 25330 1 47
2 25331 1 47
2 25332 1 47
2 25333 1 47
2 25334 1 47
2 25335 1 47
2 25336 1 47
2 25337 1 47
2 25338 1 47
2 25339 1 47
2 25340 1 47
2 25341 1 47
2 25342 1 47
2 25343 1 47
2 25344 1 47
2 25345 1 47
2 25346 1 47
2 25347 1 47
2 25348 1 47
2 25349 1 47
2 25350 1 47
2 25351 1 47
2 25352 1 47
2 25353 1 47
2 25354 1 47
2 25355 1 47
2 25356 1 47
2 25357 1 47
2 25358 1 47
2 25359 1 47
2 25360 1 47
2 25361 1 47
2 25362 1 48
2 25363 1 48
2 25364 1 48
2 25365 1 48
2 25366 1 48
2 25367 1 48
2 25368 1 48
2 25369 1 48
2 25370 1 48
2 25371 1 48
2 25372 1 48
2 25373 1 48
2 25374 1 48
2 25375 1 48
2 25376 1 48
2 25377 1 48
2 25378 1 48
2 25379 1 48
2 25380 1 48
2 25381 1 48
2 25382 1 48
2 25383 1 48
2 25384 1 48
2 25385 1 48
2 25386 1 48
2 25387 1 48
2 25388 1 48
2 25389 1 48
2 25390 1 48
2 25391 1 48
2 25392 1 48
2 25393 1 48
2 25394 1 48
2 25395 1 48
2 25396 1 48
2 25397 1 48
2 25398 1 48
2 25399 1 48
2 25400 1 48
2 25401 1 48
2 25402 1 48
2 25403 1 48
2 25404 1 48
2 25405 1 48
2 25406 1 48
2 25407 1 48
2 25408 1 48
2 25409 1 48
2 25410 1 48
2 25411 1 48
2 25412 1 48
2 25413 1 48
2 25414 1 48
2 25415 1 48
2 25416 1 48
2 25417 1 48
2 25418 1 48
2 25419 1 48
2 25420 1 48
2 25421 1 48
2 25422 1 48
2 25423 1 48
2 25424 1 48
2 25425 1 48
2 25426 1 48
2 25427 1 48
2 25428 1 48
2 25429 1 48
2 25430 1 48
2 25431 1 48
2 25432 1 49
2 25433 1 49
2 25434 1 49
2 25435 1 49
2 25436 1 49
2 25437 1 49
2 25438 1 49
2 25439 1 49
2 25440 1 49
2 25441 1 49
2 25442 1 49
2 25443 1 49
2 25444 1 49
2 25445 1 49
2 25446 1 49
2 25447 1 49
2 25448 1 49
2 25449 1 49
2 25450 1 49
2 25451 1 49
2 25452 1 49
2 25453 1 49
2 25454 1 49
2 25455 1 49
2 25456 1 49
2 25457 1 49
2 25458 1 49
2 25459 1 49
2 25460 1 49
2 25461 1 49
2 25462 1 49
2 25463 1 49
2 25464 1 49
2 25465 1 49
2 25466 1 49
2 25467 1 49
2 25468 1 49
2 25469 1 49
2 25470 1 49
2 25471 1 49
2 25472 1 49
2 25473 1 49
2 25474 1 49
2 25475 1 49
2 25476 1 49
2 25477 1 49
2 25478 1 49
2 25479 1 49
2 25480 1 49
2 25481 1 49
2 25482 1 49
2 25483 1 49
2 25484 1 49
2 25485 1 49
2 25486 1 49
2 25487 1 49
2 25488 1 49
2 25489 1 49
2 25490 1 49
2 25491 1 49
2 25492 1 49
2 25493 1 49
2 25494 1 49
2 25495 1 49
2 25496 1 49
2 25497 1 49
2 25498 1 49
2 25499 1 49
2 25500 1 49
2 25501 1 49
2 25502 1 49
2 25503 1 49
2 25504 1 49
2 25505 1 49
2 25506 1 49
2 25507 1 49
2 25508 1 49
2 25509 1 49
2 25510 1 49
2 25511 1 49
2 25512 1 49
2 25513 1 49
2 25514 1 49
2 25515 1 49
2 25516 1 49
2 25517 1 49
2 25518 1 49
2 25519 1 49
2 25520 1 49
2 25521 1 49
2 25522 1 49
2 25523 1 49
2 25524 1 49
2 25525 1 49
2 25526 1 49
2 25527 1 49
2 25528 1 49
2 25529 1 49
2 25530 1 49
2 25531 1 49
2 25532 1 49
2 25533 1 49
2 25534 1 49
2 25535 1 49
2 25536 1 49
2 25537 1 49
2 25538 1 50
2 25539 1 50
2 25540 1 50
2 25541 1 50
2 25542 1 50
2 25543 1 50
2 25544 1 50
2 25545 1 50
2 25546 1 50
2 25547 1 50
2 25548 1 50
2 25549 1 50
2 25550 1 50
2 25551 1 50
2 25552 1 50
2 25553 1 50
2 25554 1 50
2 25555 1 50
2 25556 1 50
2 25557 1 50
2 25558 1 50
2 25559 1 50
2 25560 1 50
2 25561 1 50
2 25562 1 50
2 25563 1 50
2 25564 1 50
2 25565 1 50
2 25566 1 50
2 25567 1 50
2 25568 1 50
2 25569 1 50
2 25570 1 50
2 25571 1 50
2 25572 1 50
2 25573 1 50
2 25574 1 50
2 25575 1 50
2 25576 1 50
2 25577 1 50
2 25578 1 50
2 25579 1 50
2 25580 1 50
2 25581 1 50
2 25582 1 50
2 25583 1 50
2 25584 1 50
2 25585 1 50
2 25586 1 50
2 25587 1 50
2 25588 1 50
2 25589 1 50
2 25590 1 50
2 25591 1 50
2 25592 1 50
2 25593 1 50
2 25594 1 50
2 25595 1 50
2 25596 1 50
2 25597 1 50
2 25598 1 50
2 25599 1 50
2 25600 1 50
2 25601 1 50
2 25602 1 50
2 25603 1 50
2 25604 1 50
2 25605 1 50
2 25606 1 50
2 25607 1 50
2 25608 1 50
2 25609 1 50
2 25610 1 50
2 25611 1 50
2 25612 1 50
2 25613 1 50
2 25614 1 50
2 25615 1 50
2 25616 1 50
2 25617 1 50
2 25618 1 50
2 25619 1 50
2 25620 1 50
2 25621 1 50
2 25622 1 50
2 25623 1 50
2 25624 1 50
2 25625 1 50
2 25626 1 50
2 25627 1 50
2 25628 1 50
2 25629 1 50
2 25630 1 50
2 25631 1 50
2 25632 1 50
2 25633 1 50
2 25634 1 50
2 25635 1 50
2 25636 1 50
2 25637 1 50
2 25638 1 51
2 25639 1 51
2 25640 1 51
2 25641 1 51
2 25642 1 51
2 25643 1 51
2 25644 1 51
2 25645 1 51
2 25646 1 51
2 25647 1 51
2 25648 1 51
2 25649 1 51
2 25650 1 51
2 25651 1 51
2 25652 1 51
2 25653 1 51
2 25654 1 51
2 25655 1 51
2 25656 1 51
2 25657 1 51
2 25658 1 51
2 25659 1 51
2 25660 1 51
2 25661 1 51
2 25662 1 51
2 25663 1 51
2 25664 1 51
2 25665 1 51
2 25666 1 51
2 25667 1 51
2 25668 1 51
2 25669 1 51
2 25670 1 51
2 25671 1 51
2 25672 1 51
2 25673 1 51
2 25674 1 51
2 25675 1 51
2 25676 1 51
2 25677 1 51
2 25678 1 51
2 25679 1 51
2 25680 1 51
2 25681 1 51
2 25682 1 51
2 25683 1 51
2 25684 1 51
2 25685 1 51
2 25686 1 51
2 25687 1 51
2 25688 1 52
2 25689 1 52
2 25690 1 54
2 25691 1 54
2 25692 1 54
2 25693 1 54
2 25694 1 54
2 25695 1 56
2 25696 1 56
2 25697 1 57
2 25698 1 57
2 25699 1 57
2 25700 1 57
2 25701 1 57
2 25702 1 57
2 25703 1 57
2 25704 1 57
2 25705 1 57
2 25706 1 57
2 25707 1 57
2 25708 1 57
2 25709 1 57
2 25710 1 57
2 25711 1 57
2 25712 1 57
2 25713 1 57
2 25714 1 57
2 25715 1 57
2 25716 1 57
2 25717 1 57
2 25718 1 57
2 25719 1 57
2 25720 1 57
2 25721 1 57
2 25722 1 57
2 25723 1 57
2 25724 1 57
2 25725 1 57
2 25726 1 57
2 25727 1 57
2 25728 1 57
2 25729 1 57
2 25730 1 57
2 25731 1 57
2 25732 1 57
2 25733 1 57
2 25734 1 57
2 25735 1 57
2 25736 1 57
2 25737 1 57
2 25738 1 58
2 25739 1 58
2 25740 1 58
2 25741 1 58
2 25742 1 58
2 25743 1 58
2 25744 1 58
2 25745 1 58
2 25746 1 58
2 25747 1 58
2 25748 1 58
2 25749 1 58
2 25750 1 58
2 25751 1 58
2 25752 1 58
2 25753 1 58
2 25754 1 58
2 25755 1 58
2 25756 1 58
2 25757 1 58
2 25758 1 58
2 25759 1 58
2 25760 1 58
2 25761 1 58
2 25762 1 58
2 25763 1 58
2 25764 1 58
2 25765 1 58
2 25766 1 58
2 25767 1 60
2 25768 1 60
2 25769 1 60
2 25770 1 60
2 25771 1 60
2 25772 1 60
2 25773 1 60
2 25774 1 60
2 25775 1 61
2 25776 1 61
2 25777 1 61
2 25778 1 61
2 25779 1 61
2 25780 1 61
2 25781 1 62
2 25782 1 62
2 25783 1 62
2 25784 1 62
2 25785 1 62
2 25786 1 62
2 25787 1 62
2 25788 1 62
2 25789 1 62
2 25790 1 63
2 25791 1 63
2 25792 1 64
2 25793 1 64
2 25794 1 65
2 25795 1 65
2 25796 1 65
2 25797 1 65
2 25798 1 65
2 25799 1 65
2 25800 1 65
2 25801 1 65
2 25802 1 65
2 25803 1 65
2 25804 1 65
2 25805 1 65
2 25806 1 65
2 25807 1 65
2 25808 1 65
2 25809 1 65
2 25810 1 66
2 25811 1 66
2 25812 1 66
2 25813 1 66
2 25814 1 66
2 25815 1 66
2 25816 1 66
2 25817 1 66
2 25818 1 66
2 25819 1 66
2 25820 1 67
2 25821 1 67
2 25822 1 68
2 25823 1 68
2 25824 1 68
2 25825 1 68
2 25826 1 68
2 25827 1 71
2 25828 1 71
2 25829 1 71
2 25830 1 71
2 25831 1 71
2 25832 1 71
2 25833 1 71
2 25834 1 71
2 25835 1 71
2 25836 1 71
2 25837 1 71
2 25838 1 71
2 25839 1 71
2 25840 1 71
2 25841 1 71
2 25842 1 71
2 25843 1 71
2 25844 1 71
2 25845 1 71
2 25846 1 71
2 25847 1 71
2 25848 1 71
2 25849 1 71
2 25850 1 71
2 25851 1 71
2 25852 1 71
2 25853 1 71
2 25854 1 71
2 25855 1 71
2 25856 1 71
2 25857 1 71
2 25858 1 71
2 25859 1 71
2 25860 1 71
2 25861 1 71
2 25862 1 71
2 25863 1 71
2 25864 1 71
2 25865 1 71
2 25866 1 71
2 25867 1 71
2 25868 1 71
2 25869 1 71
2 25870 1 71
2 25871 1 72
2 25872 1 72
2 25873 1 72
2 25874 1 73
2 25875 1 73
2 25876 1 73
2 25877 1 73
2 25878 1 73
2 25879 1 75
2 25880 1 75
2 25881 1 75
2 25882 1 75
2 25883 1 75
2 25884 1 75
2 25885 1 75
2 25886 1 75
2 25887 1 75
2 25888 1 75
2 25889 1 75
2 25890 1 77
2 25891 1 77
2 25892 1 77
2 25893 1 77
2 25894 1 78
2 25895 1 78
2 25896 1 78
2 25897 1 78
2 25898 1 78
2 25899 1 78
2 25900 1 78
2 25901 1 78
2 25902 1 78
2 25903 1 78
2 25904 1 78
2 25905 1 78
2 25906 1 78
2 25907 1 78
2 25908 1 78
2 25909 1 78
2 25910 1 78
2 25911 1 78
2 25912 1 78
2 25913 1 78
2 25914 1 78
2 25915 1 78
2 25916 1 78
2 25917 1 78
2 25918 1 78
2 25919 1 78
2 25920 1 78
2 25921 1 78
2 25922 1 78
2 25923 1 78
2 25924 1 78
2 25925 1 78
2 25926 1 78
2 25927 1 78
2 25928 1 78
2 25929 1 78
2 25930 1 78
2 25931 1 78
2 25932 1 78
2 25933 1 78
2 25934 1 78
2 25935 1 78
2 25936 1 78
2 25937 1 78
2 25938 1 78
2 25939 1 78
2 25940 1 78
2 25941 1 78
2 25942 1 78
2 25943 1 78
2 25944 1 78
2 25945 1 78
2 25946 1 78
2 25947 1 78
2 25948 1 78
2 25949 1 78
2 25950 1 78
2 25951 1 78
2 25952 1 78
2 25953 1 78
2 25954 1 78
2 25955 1 78
2 25956 1 78
2 25957 1 78
2 25958 1 78
2 25959 1 78
2 25960 1 78
2 25961 1 78
2 25962 1 78
2 25963 1 78
2 25964 1 79
2 25965 1 79
2 25966 1 81
2 25967 1 81
2 25968 1 82
2 25969 1 82
2 25970 1 83
2 25971 1 83
2 25972 1 83
2 25973 1 83
2 25974 1 83
2 25975 1 83
2 25976 1 83
2 25977 1 83
2 25978 1 83
2 25979 1 86
2 25980 1 86
2 25981 1 86
2 25982 1 86
2 25983 1 86
2 25984 1 86
2 25985 1 86
2 25986 1 86
2 25987 1 86
2 25988 1 86
2 25989 1 86
2 25990 1 86
2 25991 1 86
2 25992 1 86
2 25993 1 86
2 25994 1 86
2 25995 1 86
2 25996 1 87
2 25997 1 87
2 25998 1 87
2 25999 1 87
2 26000 1 87
2 26001 1 87
2 26002 1 87
2 26003 1 87
2 26004 1 87
2 26005 1 87
2 26006 1 89
2 26007 1 89
2 26008 1 89
2 26009 1 89
2 26010 1 89
2 26011 1 89
2 26012 1 89
2 26013 1 89
2 26014 1 89
2 26015 1 89
2 26016 1 89
2 26017 1 89
2 26018 1 89
2 26019 1 89
2 26020 1 89
2 26021 1 89
2 26022 1 89
2 26023 1 89
2 26024 1 89
2 26025 1 89
2 26026 1 90
2 26027 1 90
2 26028 1 90
2 26029 1 90
2 26030 1 91
2 26031 1 91
2 26032 1 91
2 26033 1 98
2 26034 1 98
2 26035 1 98
2 26036 1 98
2 26037 1 98
2 26038 1 98
2 26039 1 98
2 26040 1 98
2 26041 1 98
2 26042 1 100
2 26043 1 100
2 26044 1 101
2 26045 1 101
2 26046 1 101
2 26047 1 101
2 26048 1 101
2 26049 1 101
2 26050 1 101
2 26051 1 101
2 26052 1 101
2 26053 1 101
2 26054 1 101
2 26055 1 101
2 26056 1 101
2 26057 1 101
2 26058 1 101
2 26059 1 101
2 26060 1 101
2 26061 1 101
2 26062 1 101
2 26063 1 101
2 26064 1 101
2 26065 1 101
2 26066 1 101
2 26067 1 101
2 26068 1 101
2 26069 1 101
2 26070 1 101
2 26071 1 101
2 26072 1 101
2 26073 1 101
2 26074 1 101
2 26075 1 101
2 26076 1 101
2 26077 1 101
2 26078 1 101
2 26079 1 101
2 26080 1 101
2 26081 1 101
2 26082 1 101
2 26083 1 101
2 26084 1 101
2 26085 1 101
2 26086 1 101
2 26087 1 101
2 26088 1 101
2 26089 1 101
2 26090 1 101
2 26091 1 101
2 26092 1 101
2 26093 1 101
2 26094 1 101
2 26095 1 101
2 26096 1 101
2 26097 1 101
2 26098 1 101
2 26099 1 102
2 26100 1 102
2 26101 1 103
2 26102 1 103
2 26103 1 103
2 26104 1 103
2 26105 1 103
2 26106 1 103
2 26107 1 103
2 26108 1 103
2 26109 1 103
2 26110 1 103
2 26111 1 103
2 26112 1 103
2 26113 1 103
2 26114 1 103
2 26115 1 103
2 26116 1 103
2 26117 1 103
2 26118 1 103
2 26119 1 103
2 26120 1 103
2 26121 1 103
2 26122 1 103
2 26123 1 103
2 26124 1 103
2 26125 1 103
2 26126 1 103
2 26127 1 103
2 26128 1 103
2 26129 1 104
2 26130 1 104
2 26131 1 104
2 26132 1 104
2 26133 1 104
2 26134 1 104
2 26135 1 104
2 26136 1 104
2 26137 1 104
2 26138 1 104
2 26139 1 105
2 26140 1 105
2 26141 1 105
2 26142 1 113
2 26143 1 113
2 26144 1 113
2 26145 1 113
2 26146 1 113
2 26147 1 113
2 26148 1 113
2 26149 1 113
2 26150 1 113
2 26151 1 113
2 26152 1 113
2 26153 1 113
2 26154 1 113
2 26155 1 113
2 26156 1 113
2 26157 1 113
2 26158 1 113
2 26159 1 113
2 26160 1 113
2 26161 1 113
2 26162 1 114
2 26163 1 114
2 26164 1 114
2 26165 1 114
2 26166 1 114
2 26167 1 114
2 26168 1 114
2 26169 1 114
2 26170 1 114
2 26171 1 114
2 26172 1 114
2 26173 1 114
2 26174 1 114
2 26175 1 114
2 26176 1 114
2 26177 1 114
2 26178 1 114
2 26179 1 114
2 26180 1 114
2 26181 1 114
2 26182 1 114
2 26183 1 114
2 26184 1 115
2 26185 1 115
2 26186 1 115
2 26187 1 115
2 26188 1 115
2 26189 1 124
2 26190 1 124
2 26191 1 124
2 26192 1 124
2 26193 1 124
2 26194 1 124
2 26195 1 124
2 26196 1 124
2 26197 1 124
2 26198 1 124
2 26199 1 124
2 26200 1 124
2 26201 1 124
2 26202 1 124
2 26203 1 124
2 26204 1 124
2 26205 1 124
2 26206 1 124
2 26207 1 124
2 26208 1 124
2 26209 1 124
2 26210 1 124
2 26211 1 124
2 26212 1 124
2 26213 1 124
2 26214 1 124
2 26215 1 124
2 26216 1 124
2 26217 1 124
2 26218 1 125
2 26219 1 125
2 26220 1 125
2 26221 1 125
2 26222 1 125
2 26223 1 125
2 26224 1 125
2 26225 1 125
2 26226 1 125
2 26227 1 125
2 26228 1 125
2 26229 1 125
2 26230 1 125
2 26231 1 125
2 26232 1 125
2 26233 1 126
2 26234 1 126
2 26235 1 126
2 26236 1 126
2 26237 1 126
2 26238 1 126
2 26239 1 126
2 26240 1 128
2 26241 1 128
2 26242 1 128
2 26243 1 128
2 26244 1 128
2 26245 1 130
2 26246 1 130
2 26247 1 132
2 26248 1 132
2 26249 1 132
2 26250 1 132
2 26251 1 132
2 26252 1 132
2 26253 1 132
2 26254 1 132
2 26255 1 132
2 26256 1 132
2 26257 1 132
2 26258 1 132
2 26259 1 132
2 26260 1 132
2 26261 1 132
2 26262 1 132
2 26263 1 132
2 26264 1 132
2 26265 1 132
2 26266 1 132
2 26267 1 132
2 26268 1 132
2 26269 1 132
2 26270 1 132
2 26271 1 132
2 26272 1 133
2 26273 1 133
2 26274 1 133
2 26275 1 134
2 26276 1 134
2 26277 1 134
2 26278 1 134
2 26279 1 135
2 26280 1 135
2 26281 1 137
2 26282 1 137
2 26283 1 137
2 26284 1 137
2 26285 1 137
2 26286 1 137
2 26287 1 137
2 26288 1 137
2 26289 1 145
2 26290 1 145
2 26291 1 146
2 26292 1 146
2 26293 1 148
2 26294 1 148
2 26295 1 149
2 26296 1 149
2 26297 1 149
2 26298 1 149
2 26299 1 149
2 26300 1 149
2 26301 1 149
2 26302 1 149
2 26303 1 149
2 26304 1 149
2 26305 1 149
2 26306 1 149
2 26307 1 149
2 26308 1 149
2 26309 1 149
2 26310 1 149
2 26311 1 149
2 26312 1 149
2 26313 1 150
2 26314 1 150
2 26315 1 151
2 26316 1 151
2 26317 1 151
2 26318 1 151
2 26319 1 152
2 26320 1 152
2 26321 1 152
2 26322 1 154
2 26323 1 154
2 26324 1 154
2 26325 1 154
2 26326 1 155
2 26327 1 155
2 26328 1 160
2 26329 1 160
2 26330 1 161
2 26331 1 161
2 26332 1 161
2 26333 1 162
2 26334 1 162
2 26335 1 162
2 26336 1 162
2 26337 1 162
2 26338 1 162
2 26339 1 162
2 26340 1 162
2 26341 1 162
2 26342 1 162
2 26343 1 162
2 26344 1 164
2 26345 1 164
2 26346 1 164
2 26347 1 164
2 26348 1 164
2 26349 1 164
2 26350 1 164
2 26351 1 164
2 26352 1 164
2 26353 1 164
2 26354 1 165
2 26355 1 165
2 26356 1 173
2 26357 1 173
2 26358 1 173
2 26359 1 173
2 26360 1 173
2 26361 1 173
2 26362 1 176
2 26363 1 176
2 26364 1 176
2 26365 1 177
2 26366 1 177
2 26367 1 177
2 26368 1 177
2 26369 1 177
2 26370 1 177
2 26371 1 181
2 26372 1 181
2 26373 1 184
2 26374 1 184
2 26375 1 184
2 26376 1 184
2 26377 1 184
2 26378 1 184
2 26379 1 184
2 26380 1 184
2 26381 1 184
2 26382 1 184
2 26383 1 184
2 26384 1 184
2 26385 1 184
2 26386 1 184
2 26387 1 185
2 26388 1 185
2 26389 1 185
2 26390 1 186
2 26391 1 186
2 26392 1 186
2 26393 1 187
2 26394 1 187
2 26395 1 187
2 26396 1 187
2 26397 1 188
2 26398 1 188
2 26399 1 188
2 26400 1 188
2 26401 1 188
2 26402 1 188
2 26403 1 188
2 26404 1 188
2 26405 1 188
2 26406 1 188
2 26407 1 188
2 26408 1 188
2 26409 1 188
2 26410 1 188
2 26411 1 188
2 26412 1 188
2 26413 1 188
2 26414 1 188
2 26415 1 188
2 26416 1 188
2 26417 1 188
2 26418 1 189
2 26419 1 189
2 26420 1 189
2 26421 1 190
2 26422 1 190
2 26423 1 190
2 26424 1 190
2 26425 1 190
2 26426 1 190
2 26427 1 190
2 26428 1 190
2 26429 1 190
2 26430 1 191
2 26431 1 191
2 26432 1 191
2 26433 1 204
2 26434 1 204
2 26435 1 204
2 26436 1 204
2 26437 1 204
2 26438 1 204
2 26439 1 204
2 26440 1 205
2 26441 1 205
2 26442 1 206
2 26443 1 206
2 26444 1 206
2 26445 1 206
2 26446 1 212
2 26447 1 212
2 26448 1 212
2 26449 1 212
2 26450 1 212
2 26451 1 212
2 26452 1 212
2 26453 1 212
2 26454 1 212
2 26455 1 213
2 26456 1 213
2 26457 1 213
2 26458 1 221
2 26459 1 221
2 26460 1 221
2 26461 1 221
2 26462 1 221
2 26463 1 223
2 26464 1 223
2 26465 1 223
2 26466 1 225
2 26467 1 225
2 26468 1 225
2 26469 1 225
2 26470 1 225
2 26471 1 228
2 26472 1 228
2 26473 1 228
2 26474 1 228
2 26475 1 228
2 26476 1 228
2 26477 1 228
2 26478 1 228
2 26479 1 228
2 26480 1 228
2 26481 1 229
2 26482 1 229
2 26483 1 231
2 26484 1 231
2 26485 1 234
2 26486 1 234
2 26487 1 234
2 26488 1 234
2 26489 1 234
2 26490 1 234
2 26491 1 234
2 26492 1 234
2 26493 1 234
2 26494 1 234
2 26495 1 241
2 26496 1 241
2 26497 1 241
2 26498 1 241
2 26499 1 241
2 26500 1 241
2 26501 1 241
2 26502 1 241
2 26503 1 242
2 26504 1 242
2 26505 1 242
2 26506 1 242
2 26507 1 242
2 26508 1 242
2 26509 1 249
2 26510 1 249
2 26511 1 250
2 26512 1 250
2 26513 1 250
2 26514 1 250
2 26515 1 250
2 26516 1 250
2 26517 1 251
2 26518 1 251
2 26519 1 251
2 26520 1 251
2 26521 1 251
2 26522 1 251
2 26523 1 251
2 26524 1 251
2 26525 1 251
2 26526 1 251
2 26527 1 251
2 26528 1 251
2 26529 1 251
2 26530 1 251
2 26531 1 251
2 26532 1 251
2 26533 1 251
2 26534 1 251
2 26535 1 251
2 26536 1 251
2 26537 1 251
2 26538 1 251
2 26539 1 251
2 26540 1 251
2 26541 1 251
2 26542 1 251
2 26543 1 251
2 26544 1 251
2 26545 1 251
2 26546 1 251
2 26547 1 251
2 26548 1 251
2 26549 1 251
2 26550 1 251
2 26551 1 251
2 26552 1 251
2 26553 1 251
2 26554 1 251
2 26555 1 251
2 26556 1 251
2 26557 1 251
2 26558 1 251
2 26559 1 251
2 26560 1 251
2 26561 1 251
2 26562 1 251
2 26563 1 251
2 26564 1 251
2 26565 1 253
2 26566 1 253
2 26567 1 253
2 26568 1 253
2 26569 1 253
2 26570 1 253
2 26571 1 253
2 26572 1 253
2 26573 1 253
2 26574 1 253
2 26575 1 253
2 26576 1 253
2 26577 1 253
2 26578 1 253
2 26579 1 253
2 26580 1 253
2 26581 1 253
2 26582 1 253
2 26583 1 253
2 26584 1 254
2 26585 1 254
2 26586 1 254
2 26587 1 256
2 26588 1 256
2 26589 1 263
2 26590 1 263
2 26591 1 263
2 26592 1 263
2 26593 1 263
2 26594 1 264
2 26595 1 264
2 26596 1 265
2 26597 1 265
2 26598 1 265
2 26599 1 265
2 26600 1 265
2 26601 1 265
2 26602 1 267
2 26603 1 267
2 26604 1 275
2 26605 1 275
2 26606 1 278
2 26607 1 278
2 26608 1 278
2 26609 1 278
2 26610 1 279
2 26611 1 279
2 26612 1 279
2 26613 1 279
2 26614 1 279
2 26615 1 279
2 26616 1 279
2 26617 1 279
2 26618 1 279
2 26619 1 288
2 26620 1 288
2 26621 1 288
2 26622 1 288
2 26623 1 288
2 26624 1 290
2 26625 1 290
2 26626 1 290
2 26627 1 290
2 26628 1 290
2 26629 1 290
2 26630 1 290
2 26631 1 290
2 26632 1 290
2 26633 1 290
2 26634 1 290
2 26635 1 290
2 26636 1 290
2 26637 1 290
2 26638 1 290
2 26639 1 290
2 26640 1 290
2 26641 1 290
2 26642 1 290
2 26643 1 290
2 26644 1 291
2 26645 1 291
2 26646 1 297
2 26647 1 297
2 26648 1 297
2 26649 1 297
2 26650 1 297
2 26651 1 297
2 26652 1 297
2 26653 1 297
2 26654 1 297
2 26655 1 297
2 26656 1 297
2 26657 1 297
2 26658 1 297
2 26659 1 297
2 26660 1 297
2 26661 1 297
2 26662 1 297
2 26663 1 297
2 26664 1 297
2 26665 1 297
2 26666 1 297
2 26667 1 297
2 26668 1 297
2 26669 1 297
2 26670 1 297
2 26671 1 297
2 26672 1 297
2 26673 1 297
2 26674 1 297
2 26675 1 297
2 26676 1 297
2 26677 1 297
2 26678 1 297
2 26679 1 297
2 26680 1 298
2 26681 1 298
2 26682 1 298
2 26683 1 306
2 26684 1 306
2 26685 1 306
2 26686 1 306
2 26687 1 306
2 26688 1 306
2 26689 1 306
2 26690 1 306
2 26691 1 306
2 26692 1 306
2 26693 1 306
2 26694 1 306
2 26695 1 306
2 26696 1 306
2 26697 1 306
2 26698 1 306
2 26699 1 306
2 26700 1 306
2 26701 1 306
2 26702 1 306
2 26703 1 306
2 26704 1 306
2 26705 1 308
2 26706 1 308
2 26707 1 309
2 26708 1 309
2 26709 1 309
2 26710 1 309
2 26711 1 309
2 26712 1 309
2 26713 1 323
2 26714 1 323
2 26715 1 323
2 26716 1 323
2 26717 1 323
2 26718 1 323
2 26719 1 323
2 26720 1 325
2 26721 1 325
2 26722 1 325
2 26723 1 325
2 26724 1 325
2 26725 1 325
2 26726 1 325
2 26727 1 325
2 26728 1 325
2 26729 1 325
2 26730 1 325
2 26731 1 325
2 26732 1 325
2 26733 1 325
2 26734 1 325
2 26735 1 325
2 26736 1 325
2 26737 1 325
2 26738 1 325
2 26739 1 325
2 26740 1 325
2 26741 1 325
2 26742 1 325
2 26743 1 327
2 26744 1 327
2 26745 1 327
2 26746 1 330
2 26747 1 330
2 26748 1 330
2 26749 1 330
2 26750 1 330
2 26751 1 331
2 26752 1 331
2 26753 1 342
2 26754 1 342
2 26755 1 342
2 26756 1 342
2 26757 1 342
2 26758 1 342
2 26759 1 342
2 26760 1 342
2 26761 1 342
2 26762 1 342
2 26763 1 342
2 26764 1 342
2 26765 1 342
2 26766 1 342
2 26767 1 342
2 26768 1 342
2 26769 1 342
2 26770 1 342
2 26771 1 342
2 26772 1 342
2 26773 1 342
2 26774 1 342
2 26775 1 342
2 26776 1 342
2 26777 1 342
2 26778 1 342
2 26779 1 342
2 26780 1 343
2 26781 1 343
2 26782 1 343
2 26783 1 343
2 26784 1 343
2 26785 1 343
2 26786 1 343
2 26787 1 343
2 26788 1 343
2 26789 1 343
2 26790 1 343
2 26791 1 343
2 26792 1 343
2 26793 1 343
2 26794 1 343
2 26795 1 343
2 26796 1 343
2 26797 1 343
2 26798 1 343
2 26799 1 343
2 26800 1 343
2 26801 1 343
2 26802 1 343
2 26803 1 343
2 26804 1 343
2 26805 1 343
2 26806 1 343
2 26807 1 343
2 26808 1 343
2 26809 1 343
2 26810 1 343
2 26811 1 344
2 26812 1 344
2 26813 1 344
2 26814 1 344
2 26815 1 344
2 26816 1 344
2 26817 1 344
2 26818 1 344
2 26819 1 344
2 26820 1 344
2 26821 1 344
2 26822 1 344
2 26823 1 344
2 26824 1 345
2 26825 1 345
2 26826 1 346
2 26827 1 346
2 26828 1 353
2 26829 1 353
2 26830 1 353
2 26831 1 353
2 26832 1 354
2 26833 1 354
2 26834 1 354
2 26835 1 354
2 26836 1 354
2 26837 1 354
2 26838 1 355
2 26839 1 355
2 26840 1 355
2 26841 1 359
2 26842 1 359
2 26843 1 359
2 26844 1 360
2 26845 1 360
2 26846 1 360
2 26847 1 366
2 26848 1 366
2 26849 1 366
2 26850 1 366
2 26851 1 368
2 26852 1 368
2 26853 1 368
2 26854 1 369
2 26855 1 369
2 26856 1 369
2 26857 1 369
2 26858 1 369
2 26859 1 369
2 26860 1 369
2 26861 1 369
2 26862 1 369
2 26863 1 369
2 26864 1 369
2 26865 1 369
2 26866 1 370
2 26867 1 370
2 26868 1 373
2 26869 1 373
2 26870 1 373
2 26871 1 373
2 26872 1 373
2 26873 1 373
2 26874 1 374
2 26875 1 374
2 26876 1 374
2 26877 1 374
2 26878 1 375
2 26879 1 375
2 26880 1 375
2 26881 1 375
2 26882 1 375
2 26883 1 383
2 26884 1 383
2 26885 1 383
2 26886 1 383
2 26887 1 383
2 26888 1 383
2 26889 1 384
2 26890 1 384
2 26891 1 384
2 26892 1 384
2 26893 1 384
2 26894 1 385
2 26895 1 385
2 26896 1 385
2 26897 1 385
2 26898 1 385
2 26899 1 385
2 26900 1 389
2 26901 1 389
2 26902 1 389
2 26903 1 390
2 26904 1 390
2 26905 1 390
2 26906 1 390
2 26907 1 390
2 26908 1 390
2 26909 1 390
2 26910 1 390
2 26911 1 390
2 26912 1 390
2 26913 1 390
2 26914 1 390
2 26915 1 390
2 26916 1 390
2 26917 1 390
2 26918 1 390
2 26919 1 390
2 26920 1 391
2 26921 1 391
2 26922 1 391
2 26923 1 391
2 26924 1 391
2 26925 1 391
2 26926 1 391
2 26927 1 391
2 26928 1 391
2 26929 1 391
2 26930 1 391
2 26931 1 392
2 26932 1 392
2 26933 1 392
2 26934 1 392
2 26935 1 402
2 26936 1 402
2 26937 1 402
2 26938 1 403
2 26939 1 403
2 26940 1 403
2 26941 1 403
2 26942 1 403
2 26943 1 403
2 26944 1 403
2 26945 1 403
2 26946 1 403
2 26947 1 404
2 26948 1 404
2 26949 1 404
2 26950 1 404
2 26951 1 404
2 26952 1 405
2 26953 1 405
2 26954 1 413
2 26955 1 413
2 26956 1 413
2 26957 1 413
2 26958 1 413
2 26959 1 413
2 26960 1 413
2 26961 1 413
2 26962 1 413
2 26963 1 413
2 26964 1 413
2 26965 1 413
2 26966 1 413
2 26967 1 413
2 26968 1 413
2 26969 1 413
2 26970 1 413
2 26971 1 413
2 26972 1 413
2 26973 1 413
2 26974 1 414
2 26975 1 414
2 26976 1 414
2 26977 1 415
2 26978 1 415
2 26979 1 415
2 26980 1 415
2 26981 1 415
2 26982 1 415
2 26983 1 416
2 26984 1 416
2 26985 1 416
2 26986 1 417
2 26987 1 417
2 26988 1 417
2 26989 1 417
2 26990 1 418
2 26991 1 418
2 26992 1 427
2 26993 1 427
2 26994 1 430
2 26995 1 430
2 26996 1 430
2 26997 1 432
2 26998 1 432
2 26999 1 432
2 27000 1 432
2 27001 1 433
2 27002 1 433
2 27003 1 434
2 27004 1 434
2 27005 1 434
2 27006 1 437
2 27007 1 437
2 27008 1 437
2 27009 1 437
2 27010 1 444
2 27011 1 444
2 27012 1 444
2 27013 1 444
2 27014 1 444
2 27015 1 444
2 27016 1 444
2 27017 1 444
2 27018 1 444
2 27019 1 444
2 27020 1 444
2 27021 1 444
2 27022 1 444
2 27023 1 444
2 27024 1 444
2 27025 1 461
2 27026 1 461
2 27027 1 461
2 27028 1 461
2 27029 1 461
2 27030 1 461
2 27031 1 461
2 27032 1 461
2 27033 1 461
2 27034 1 461
2 27035 1 461
2 27036 1 461
2 27037 1 461
2 27038 1 463
2 27039 1 463
2 27040 1 463
2 27041 1 463
2 27042 1 463
2 27043 1 463
2 27044 1 463
2 27045 1 464
2 27046 1 464
2 27047 1 464
2 27048 1 465
2 27049 1 465
2 27050 1 465
2 27051 1 465
2 27052 1 468
2 27053 1 468
2 27054 1 468
2 27055 1 470
2 27056 1 470
2 27057 1 470
2 27058 1 470
2 27059 1 470
2 27060 1 470
2 27061 1 470
2 27062 1 470
2 27063 1 473
2 27064 1 473
2 27065 1 473
2 27066 1 473
2 27067 1 473
2 27068 1 473
2 27069 1 473
2 27070 1 473
2 27071 1 474
2 27072 1 474
2 27073 1 474
2 27074 1 475
2 27075 1 475
2 27076 1 485
2 27077 1 485
2 27078 1 486
2 27079 1 486
2 27080 1 486
2 27081 1 486
2 27082 1 487
2 27083 1 487
2 27084 1 487
2 27085 1 487
2 27086 1 489
2 27087 1 489
2 27088 1 489
2 27089 1 489
2 27090 1 489
2 27091 1 489
2 27092 1 490
2 27093 1 490
2 27094 1 490
2 27095 1 490
2 27096 1 490
2 27097 1 490
2 27098 1 491
2 27099 1 491
2 27100 1 493
2 27101 1 493
2 27102 1 493
2 27103 1 493
2 27104 1 493
2 27105 1 493
2 27106 1 493
2 27107 1 493
2 27108 1 493
2 27109 1 493
2 27110 1 493
2 27111 1 493
2 27112 1 493
2 27113 1 493
2 27114 1 496
2 27115 1 496
2 27116 1 496
2 27117 1 496
2 27118 1 496
2 27119 1 496
2 27120 1 496
2 27121 1 496
2 27122 1 496
2 27123 1 496
2 27124 1 496
2 27125 1 496
2 27126 1 496
2 27127 1 496
2 27128 1 496
2 27129 1 496
2 27130 1 496
2 27131 1 496
2 27132 1 496
2 27133 1 496
2 27134 1 496
2 27135 1 496
2 27136 1 496
2 27137 1 496
2 27138 1 496
2 27139 1 496
2 27140 1 496
2 27141 1 496
2 27142 1 496
2 27143 1 496
2 27144 1 496
2 27145 1 496
2 27146 1 496
2 27147 1 496
2 27148 1 496
2 27149 1 496
2 27150 1 496
2 27151 1 496
2 27152 1 496
2 27153 1 496
2 27154 1 496
2 27155 1 496
2 27156 1 496
2 27157 1 496
2 27158 1 497
2 27159 1 497
2 27160 1 497
2 27161 1 497
2 27162 1 497
2 27163 1 497
2 27164 1 497
2 27165 1 497
2 27166 1 497
2 27167 1 497
2 27168 1 497
2 27169 1 497
2 27170 1 497
2 27171 1 497
2 27172 1 497
2 27173 1 497
2 27174 1 497
2 27175 1 497
2 27176 1 497
2 27177 1 497
2 27178 1 497
2 27179 1 497
2 27180 1 497
2 27181 1 497
2 27182 1 497
2 27183 1 497
2 27184 1 497
2 27185 1 497
2 27186 1 497
2 27187 1 497
2 27188 1 497
2 27189 1 497
2 27190 1 497
2 27191 1 497
2 27192 1 497
2 27193 1 497
2 27194 1 497
2 27195 1 497
2 27196 1 497
2 27197 1 497
2 27198 1 497
2 27199 1 497
2 27200 1 497
2 27201 1 497
2 27202 1 497
2 27203 1 498
2 27204 1 498
2 27205 1 498
2 27206 1 498
2 27207 1 498
2 27208 1 498
2 27209 1 498
2 27210 1 498
2 27211 1 498
2 27212 1 498
2 27213 1 498
2 27214 1 498
2 27215 1 499
2 27216 1 499
2 27217 1 499
2 27218 1 499
2 27219 1 499
2 27220 1 499
2 27221 1 499
2 27222 1 499
2 27223 1 520
2 27224 1 520
2 27225 1 526
2 27226 1 526
2 27227 1 529
2 27228 1 529
2 27229 1 537
2 27230 1 537
2 27231 1 537
2 27232 1 537
2 27233 1 537
2 27234 1 537
2 27235 1 537
2 27236 1 537
2 27237 1 537
2 27238 1 537
2 27239 1 537
2 27240 1 539
2 27241 1 539
2 27242 1 539
2 27243 1 540
2 27244 1 540
2 27245 1 540
2 27246 1 540
2 27247 1 540
2 27248 1 540
2 27249 1 540
2 27250 1 540
2 27251 1 541
2 27252 1 541
2 27253 1 542
2 27254 1 542
2 27255 1 547
2 27256 1 547
2 27257 1 548
2 27258 1 548
2 27259 1 548
2 27260 1 548
2 27261 1 548
2 27262 1 548
2 27263 1 548
2 27264 1 548
2 27265 1 548
2 27266 1 548
2 27267 1 548
2 27268 1 548
2 27269 1 548
2 27270 1 548
2 27271 1 550
2 27272 1 550
2 27273 1 550
2 27274 1 552
2 27275 1 552
2 27276 1 552
2 27277 1 552
2 27278 1 552
2 27279 1 552
2 27280 1 552
2 27281 1 552
2 27282 1 552
2 27283 1 552
2 27284 1 552
2 27285 1 552
2 27286 1 552
2 27287 1 552
2 27288 1 552
2 27289 1 552
2 27290 1 552
2 27291 1 552
2 27292 1 553
2 27293 1 553
2 27294 1 553
2 27295 1 553
2 27296 1 553
2 27297 1 553
2 27298 1 553
2 27299 1 553
2 27300 1 553
2 27301 1 553
2 27302 1 553
2 27303 1 553
2 27304 1 553
2 27305 1 553
2 27306 1 553
2 27307 1 553
2 27308 1 553
2 27309 1 553
2 27310 1 553
2 27311 1 553
2 27312 1 553
2 27313 1 553
2 27314 1 553
2 27315 1 553
2 27316 1 553
2 27317 1 553
2 27318 1 553
2 27319 1 553
2 27320 1 562
2 27321 1 562
2 27322 1 562
2 27323 1 562
2 27324 1 565
2 27325 1 565
2 27326 1 565
2 27327 1 565
2 27328 1 565
2 27329 1 565
2 27330 1 565
2 27331 1 566
2 27332 1 566
2 27333 1 566
2 27334 1 567
2 27335 1 567
2 27336 1 567
2 27337 1 568
2 27338 1 568
2 27339 1 568
2 27340 1 569
2 27341 1 569
2 27342 1 569
2 27343 1 569
2 27344 1 570
2 27345 1 570
2 27346 1 570
2 27347 1 570
2 27348 1 570
2 27349 1 570
2 27350 1 570
2 27351 1 570
2 27352 1 570
2 27353 1 570
2 27354 1 570
2 27355 1 570
2 27356 1 570
2 27357 1 570
2 27358 1 571
2 27359 1 571
2 27360 1 571
2 27361 1 571
2 27362 1 571
2 27363 1 572
2 27364 1 572
2 27365 1 572
2 27366 1 580
2 27367 1 580
2 27368 1 580
2 27369 1 581
2 27370 1 581
2 27371 1 581
2 27372 1 581
2 27373 1 581
2 27374 1 581
2 27375 1 581
2 27376 1 581
2 27377 1 581
2 27378 1 581
2 27379 1 581
2 27380 1 581
2 27381 1 581
2 27382 1 581
2 27383 1 581
2 27384 1 581
2 27385 1 581
2 27386 1 581
2 27387 1 582
2 27388 1 582
2 27389 1 582
2 27390 1 583
2 27391 1 583
2 27392 1 583
2 27393 1 583
2 27394 1 583
2 27395 1 583
2 27396 1 583
2 27397 1 583
2 27398 1 583
2 27399 1 583
2 27400 1 583
2 27401 1 583
2 27402 1 583
2 27403 1 583
2 27404 1 583
2 27405 1 583
2 27406 1 583
2 27407 1 583
2 27408 1 583
2 27409 1 583
2 27410 1 583
2 27411 1 583
2 27412 1 583
2 27413 1 583
2 27414 1 591
2 27415 1 591
2 27416 1 591
2 27417 1 591
2 27418 1 591
2 27419 1 591
2 27420 1 591
2 27421 1 591
2 27422 1 591
2 27423 1 591
2 27424 1 591
2 27425 1 591
2 27426 1 591
2 27427 1 591
2 27428 1 591
2 27429 1 591
2 27430 1 591
2 27431 1 591
2 27432 1 591
2 27433 1 591
2 27434 1 591
2 27435 1 591
2 27436 1 591
2 27437 1 591
2 27438 1 591
2 27439 1 591
2 27440 1 591
2 27441 1 591
2 27442 1 591
2 27443 1 591
2 27444 1 591
2 27445 1 591
2 27446 1 591
2 27447 1 591
2 27448 1 591
2 27449 1 591
2 27450 1 591
2 27451 1 591
2 27452 1 591
2 27453 1 591
2 27454 1 591
2 27455 1 591
2 27456 1 591
2 27457 1 591
2 27458 1 591
2 27459 1 591
2 27460 1 591
2 27461 1 591
2 27462 1 591
2 27463 1 591
2 27464 1 591
2 27465 1 591
2 27466 1 591
2 27467 1 591
2 27468 1 591
2 27469 1 591
2 27470 1 591
2 27471 1 591
2 27472 1 591
2 27473 1 591
2 27474 1 592
2 27475 1 592
2 27476 1 592
2 27477 1 592
2 27478 1 592
2 27479 1 592
2 27480 1 592
2 27481 1 592
2 27482 1 592
2 27483 1 592
2 27484 1 592
2 27485 1 592
2 27486 1 592
2 27487 1 592
2 27488 1 592
2 27489 1 592
2 27490 1 592
2 27491 1 592
2 27492 1 592
2 27493 1 592
2 27494 1 592
2 27495 1 592
2 27496 1 592
2 27497 1 592
2 27498 1 592
2 27499 1 592
2 27500 1 592
2 27501 1 592
2 27502 1 592
2 27503 1 592
2 27504 1 592
2 27505 1 592
2 27506 1 592
2 27507 1 592
2 27508 1 592
2 27509 1 592
2 27510 1 592
2 27511 1 592
2 27512 1 592
2 27513 1 592
2 27514 1 592
2 27515 1 592
2 27516 1 592
2 27517 1 592
2 27518 1 592
2 27519 1 592
2 27520 1 592
2 27521 1 592
2 27522 1 592
2 27523 1 592
2 27524 1 592
2 27525 1 592
2 27526 1 592
2 27527 1 592
2 27528 1 592
2 27529 1 592
2 27530 1 592
2 27531 1 592
2 27532 1 592
2 27533 1 592
2 27534 1 592
2 27535 1 592
2 27536 1 592
2 27537 1 592
2 27538 1 592
2 27539 1 593
2 27540 1 593
2 27541 1 593
2 27542 1 593
2 27543 1 593
2 27544 1 594
2 27545 1 594
2 27546 1 594
2 27547 1 594
2 27548 1 594
2 27549 1 594
2 27550 1 595
2 27551 1 595
2 27552 1 595
2 27553 1 598
2 27554 1 598
2 27555 1 598
2 27556 1 598
2 27557 1 598
2 27558 1 598
2 27559 1 598
2 27560 1 598
2 27561 1 598
2 27562 1 598
2 27563 1 598
2 27564 1 598
2 27565 1 598
2 27566 1 598
2 27567 1 605
2 27568 1 605
2 27569 1 605
2 27570 1 605
2 27571 1 606
2 27572 1 606
2 27573 1 606
2 27574 1 606
2 27575 1 606
2 27576 1 607
2 27577 1 607
2 27578 1 607
2 27579 1 607
2 27580 1 608
2 27581 1 608
2 27582 1 624
2 27583 1 624
2 27584 1 624
2 27585 1 624
2 27586 1 624
2 27587 1 624
2 27588 1 624
2 27589 1 624
2 27590 1 624
2 27591 1 624
2 27592 1 624
2 27593 1 624
2 27594 1 624
2 27595 1 624
2 27596 1 624
2 27597 1 624
2 27598 1 624
2 27599 1 624
2 27600 1 625
2 27601 1 625
2 27602 1 625
2 27603 1 625
2 27604 1 625
2 27605 1 625
2 27606 1 625
2 27607 1 625
2 27608 1 625
2 27609 1 625
2 27610 1 625
2 27611 1 625
2 27612 1 625
2 27613 1 625
2 27614 1 625
2 27615 1 628
2 27616 1 628
2 27617 1 628
2 27618 1 628
2 27619 1 628
2 27620 1 628
2 27621 1 628
2 27622 1 628
2 27623 1 628
2 27624 1 628
2 27625 1 628
2 27626 1 628
2 27627 1 628
2 27628 1 629
2 27629 1 629
2 27630 1 629
2 27631 1 629
2 27632 1 631
2 27633 1 631
2 27634 1 632
2 27635 1 632
2 27636 1 632
2 27637 1 633
2 27638 1 633
2 27639 1 633
2 27640 1 634
2 27641 1 634
2 27642 1 638
2 27643 1 638
2 27644 1 640
2 27645 1 640
2 27646 1 641
2 27647 1 641
2 27648 1 641
2 27649 1 641
2 27650 1 641
2 27651 1 642
2 27652 1 642
2 27653 1 643
2 27654 1 643
2 27655 1 643
2 27656 1 643
2 27657 1 644
2 27658 1 644
2 27659 1 644
2 27660 1 644
2 27661 1 644
2 27662 1 644
2 27663 1 644
2 27664 1 645
2 27665 1 645
2 27666 1 645
2 27667 1 645
2 27668 1 645
2 27669 1 647
2 27670 1 647
2 27671 1 648
2 27672 1 648
2 27673 1 648
2 27674 1 648
2 27675 1 648
2 27676 1 648
2 27677 1 649
2 27678 1 649
2 27679 1 649
2 27680 1 649
2 27681 1 649
2 27682 1 649
2 27683 1 649
2 27684 1 649
2 27685 1 650
2 27686 1 650
2 27687 1 650
2 27688 1 650
2 27689 1 650
2 27690 1 650
2 27691 1 650
2 27692 1 650
2 27693 1 650
2 27694 1 650
2 27695 1 650
2 27696 1 650
2 27697 1 650
2 27698 1 652
2 27699 1 652
2 27700 1 652
2 27701 1 652
2 27702 1 654
2 27703 1 654
2 27704 1 659
2 27705 1 659
2 27706 1 660
2 27707 1 660
2 27708 1 660
2 27709 1 660
2 27710 1 660
2 27711 1 660
2 27712 1 660
2 27713 1 660
2 27714 1 660
2 27715 1 660
2 27716 1 660
2 27717 1 660
2 27718 1 660
2 27719 1 660
2 27720 1 660
2 27721 1 661
2 27722 1 661
2 27723 1 661
2 27724 1 661
2 27725 1 662
2 27726 1 662
2 27727 1 662
2 27728 1 662
2 27729 1 662
2 27730 1 662
2 27731 1 662
2 27732 1 662
2 27733 1 662
2 27734 1 662
2 27735 1 662
2 27736 1 662
2 27737 1 662
2 27738 1 662
2 27739 1 662
2 27740 1 662
2 27741 1 662
2 27742 1 662
2 27743 1 662
2 27744 1 663
2 27745 1 663
2 27746 1 665
2 27747 1 665
2 27748 1 665
2 27749 1 665
2 27750 1 665
2 27751 1 665
2 27752 1 665
2 27753 1 665
2 27754 1 665
2 27755 1 665
2 27756 1 665
2 27757 1 665
2 27758 1 665
2 27759 1 665
2 27760 1 665
2 27761 1 665
2 27762 1 665
2 27763 1 665
2 27764 1 665
2 27765 1 665
2 27766 1 665
2 27767 1 665
2 27768 1 665
2 27769 1 665
2 27770 1 665
2 27771 1 665
2 27772 1 665
2 27773 1 665
2 27774 1 665
2 27775 1 665
2 27776 1 665
2 27777 1 665
2 27778 1 665
2 27779 1 665
2 27780 1 665
2 27781 1 665
2 27782 1 665
2 27783 1 665
2 27784 1 665
2 27785 1 665
2 27786 1 665
2 27787 1 665
2 27788 1 665
2 27789 1 665
2 27790 1 665
2 27791 1 665
2 27792 1 666
2 27793 1 666
2 27794 1 666
2 27795 1 668
2 27796 1 668
2 27797 1 676
2 27798 1 676
2 27799 1 683
2 27800 1 683
2 27801 1 683
2 27802 1 691
2 27803 1 691
2 27804 1 693
2 27805 1 693
2 27806 1 693
2 27807 1 694
2 27808 1 694
2 27809 1 694
2 27810 1 700
2 27811 1 700
2 27812 1 702
2 27813 1 702
2 27814 1 703
2 27815 1 703
2 27816 1 703
2 27817 1 703
2 27818 1 703
2 27819 1 703
2 27820 1 703
2 27821 1 703
2 27822 1 703
2 27823 1 703
2 27824 1 703
2 27825 1 703
2 27826 1 703
2 27827 1 704
2 27828 1 704
2 27829 1 704
2 27830 1 704
2 27831 1 704
2 27832 1 704
2 27833 1 704
2 27834 1 704
2 27835 1 704
2 27836 1 704
2 27837 1 704
2 27838 1 704
2 27839 1 704
2 27840 1 704
2 27841 1 704
2 27842 1 704
2 27843 1 704
2 27844 1 704
2 27845 1 704
2 27846 1 704
2 27847 1 704
2 27848 1 705
2 27849 1 705
2 27850 1 705
2 27851 1 710
2 27852 1 710
2 27853 1 710
2 27854 1 711
2 27855 1 711
2 27856 1 711
2 27857 1 711
2 27858 1 711
2 27859 1 711
2 27860 1 711
2 27861 1 712
2 27862 1 712
2 27863 1 712
2 27864 1 712
2 27865 1 729
2 27866 1 729
2 27867 1 729
2 27868 1 729
2 27869 1 729
2 27870 1 729
2 27871 1 729
2 27872 1 729
2 27873 1 729
2 27874 1 729
2 27875 1 729
2 27876 1 730
2 27877 1 730
2 27878 1 730
2 27879 1 730
2 27880 1 730
2 27881 1 730
2 27882 1 730
2 27883 1 730
2 27884 1 730
2 27885 1 730
2 27886 1 730
2 27887 1 731
2 27888 1 731
2 27889 1 731
2 27890 1 731
2 27891 1 731
2 27892 1 731
2 27893 1 732
2 27894 1 732
2 27895 1 732
2 27896 1 732
2 27897 1 732
2 27898 1 732
2 27899 1 732
2 27900 1 732
2 27901 1 732
2 27902 1 732
2 27903 1 732
2 27904 1 732
2 27905 1 732
2 27906 1 732
2 27907 1 732
2 27908 1 732
2 27909 1 732
2 27910 1 732
2 27911 1 732
2 27912 1 732
2 27913 1 732
2 27914 1 741
2 27915 1 741
2 27916 1 744
2 27917 1 744
2 27918 1 744
2 27919 1 745
2 27920 1 745
2 27921 1 746
2 27922 1 746
2 27923 1 748
2 27924 1 748
2 27925 1 754
2 27926 1 754
2 27927 1 754
2 27928 1 754
2 27929 1 754
2 27930 1 754
2 27931 1 754
2 27932 1 754
2 27933 1 755
2 27934 1 755
2 27935 1 755
2 27936 1 755
2 27937 1 755
2 27938 1 757
2 27939 1 757
2 27940 1 757
2 27941 1 757
2 27942 1 758
2 27943 1 758
2 27944 1 758
2 27945 1 758
2 27946 1 758
2 27947 1 758
2 27948 1 758
2 27949 1 760
2 27950 1 760
2 27951 1 760
2 27952 1 760
2 27953 1 760
2 27954 1 769
2 27955 1 769
2 27956 1 769
2 27957 1 769
2 27958 1 769
2 27959 1 769
2 27960 1 769
2 27961 1 769
2 27962 1 769
2 27963 1 769
2 27964 1 769
2 27965 1 769
2 27966 1 769
2 27967 1 769
2 27968 1 769
2 27969 1 770
2 27970 1 770
2 27971 1 770
2 27972 1 770
2 27973 1 770
2 27974 1 770
2 27975 1 772
2 27976 1 772
2 27977 1 772
2 27978 1 772
2 27979 1 772
2 27980 1 782
2 27981 1 782
2 27982 1 782
2 27983 1 782
2 27984 1 783
2 27985 1 783
2 27986 1 783
2 27987 1 784
2 27988 1 784
2 27989 1 791
2 27990 1 791
2 27991 1 791
2 27992 1 792
2 27993 1 792
2 27994 1 792
2 27995 1 792
2 27996 1 792
2 27997 1 792
2 27998 1 793
2 27999 1 793
2 28000 1 797
2 28001 1 797
2 28002 1 797
2 28003 1 798
2 28004 1 798
2 28005 1 799
2 28006 1 799
2 28007 1 806
2 28008 1 806
2 28009 1 806
2 28010 1 807
2 28011 1 807
2 28012 1 807
2 28013 1 807
2 28014 1 807
2 28015 1 807
2 28016 1 808
2 28017 1 808
2 28018 1 809
2 28019 1 809
2 28020 1 809
2 28021 1 809
2 28022 1 809
2 28023 1 809
2 28024 1 809
2 28025 1 823
2 28026 1 823
2 28027 1 823
2 28028 1 824
2 28029 1 824
2 28030 1 824
2 28031 1 826
2 28032 1 826
2 28033 1 827
2 28034 1 827
2 28035 1 827
2 28036 1 827
2 28037 1 827
2 28038 1 828
2 28039 1 828
2 28040 1 828
2 28041 1 828
2 28042 1 829
2 28043 1 829
2 28044 1 829
2 28045 1 829
2 28046 1 829
2 28047 1 829
2 28048 1 829
2 28049 1 839
2 28050 1 839
2 28051 1 840
2 28052 1 840
2 28053 1 840
2 28054 1 840
2 28055 1 840
2 28056 1 840
2 28057 1 840
2 28058 1 849
2 28059 1 849
2 28060 1 849
2 28061 1 849
2 28062 1 849
2 28063 1 863
2 28064 1 863
2 28065 1 864
2 28066 1 864
2 28067 1 864
2 28068 1 864
2 28069 1 864
2 28070 1 864
2 28071 1 865
2 28072 1 865
2 28073 1 865
2 28074 1 865
2 28075 1 873
2 28076 1 873
2 28077 1 873
2 28078 1 874
2 28079 1 874
2 28080 1 874
2 28081 1 874
2 28082 1 874
2 28083 1 882
2 28084 1 882
2 28085 1 882
2 28086 1 883
2 28087 1 883
2 28088 1 883
2 28089 1 883
2 28090 1 883
2 28091 1 884
2 28092 1 884
2 28093 1 899
2 28094 1 899
2 28095 1 899
2 28096 1 902
2 28097 1 902
2 28098 1 911
2 28099 1 911
2 28100 1 912
2 28101 1 912
2 28102 1 917
2 28103 1 917
2 28104 1 930
2 28105 1 930
2 28106 1 930
2 28107 1 930
2 28108 1 930
2 28109 1 930
2 28110 1 930
2 28111 1 930
2 28112 1 931
2 28113 1 931
2 28114 1 932
2 28115 1 932
2 28116 1 932
2 28117 1 932
2 28118 1 932
2 28119 1 932
2 28120 1 932
2 28121 1 932
2 28122 1 932
2 28123 1 932
2 28124 1 932
2 28125 1 932
2 28126 1 932
2 28127 1 932
2 28128 1 932
2 28129 1 932
2 28130 1 932
2 28131 1 932
2 28132 1 936
2 28133 1 936
2 28134 1 951
2 28135 1 951
2 28136 1 951
2 28137 1 951
2 28138 1 951
2 28139 1 951
2 28140 1 951
2 28141 1 951
2 28142 1 951
2 28143 1 951
2 28144 1 951
2 28145 1 951
2 28146 1 952
2 28147 1 952
2 28148 1 952
2 28149 1 959
2 28150 1 959
2 28151 1 959
2 28152 1 960
2 28153 1 960
2 28154 1 966
2 28155 1 966
2 28156 1 967
2 28157 1 967
2 28158 1 968
2 28159 1 968
2 28160 1 968
2 28161 1 968
2 28162 1 968
2 28163 1 970
2 28164 1 970
2 28165 1 970
2 28166 1 971
2 28167 1 971
2 28168 1 971
2 28169 1 972
2 28170 1 972
2 28171 1 973
2 28172 1 973
2 28173 1 973
2 28174 1 973
2 28175 1 973
2 28176 1 973
2 28177 1 973
2 28178 1 973
2 28179 1 973
2 28180 1 973
2 28181 1 973
2 28182 1 973
2 28183 1 973
2 28184 1 975
2 28185 1 975
2 28186 1 975
2 28187 1 975
2 28188 1 975
2 28189 1 975
2 28190 1 980
2 28191 1 980
2 28192 1 1003
2 28193 1 1003
2 28194 1 1004
2 28195 1 1004
2 28196 1 1004
2 28197 1 1004
2 28198 1 1004
2 28199 1 1004
2 28200 1 1004
2 28201 1 1004
2 28202 1 1005
2 28203 1 1005
2 28204 1 1006
2 28205 1 1006
2 28206 1 1007
2 28207 1 1007
2 28208 1 1008
2 28209 1 1008
2 28210 1 1009
2 28211 1 1009
2 28212 1 1009
2 28213 1 1009
2 28214 1 1009
2 28215 1 1009
2 28216 1 1009
2 28217 1 1009
2 28218 1 1009
2 28219 1 1009
2 28220 1 1009
2 28221 1 1009
2 28222 1 1009
2 28223 1 1009
2 28224 1 1009
2 28225 1 1009
2 28226 1 1009
2 28227 1 1009
2 28228 1 1010
2 28229 1 1010
2 28230 1 1010
2 28231 1 1011
2 28232 1 1011
2 28233 1 1011
2 28234 1 1012
2 28235 1 1012
2 28236 1 1014
2 28237 1 1014
2 28238 1 1014
2 28239 1 1014
2 28240 1 1014
2 28241 1 1014
2 28242 1 1026
2 28243 1 1026
2 28244 1 1026
2 28245 1 1026
2 28246 1 1027
2 28247 1 1027
2 28248 1 1027
2 28249 1 1028
2 28250 1 1028
2 28251 1 1028
2 28252 1 1029
2 28253 1 1029
2 28254 1 1029
2 28255 1 1029
2 28256 1 1029
2 28257 1 1029
2 28258 1 1029
2 28259 1 1029
2 28260 1 1029
2 28261 1 1029
2 28262 1 1029
2 28263 1 1029
2 28264 1 1038
2 28265 1 1038
2 28266 1 1038
2 28267 1 1038
2 28268 1 1038
2 28269 1 1038
2 28270 1 1039
2 28271 1 1039
2 28272 1 1039
2 28273 1 1039
2 28274 1 1039
2 28275 1 1039
2 28276 1 1040
2 28277 1 1040
2 28278 1 1040
2 28279 1 1040
2 28280 1 1040
2 28281 1 1041
2 28282 1 1041
2 28283 1 1041
2 28284 1 1041
2 28285 1 1041
2 28286 1 1041
2 28287 1 1041
2 28288 1 1041
2 28289 1 1041
2 28290 1 1041
2 28291 1 1041
2 28292 1 1041
2 28293 1 1041
2 28294 1 1041
2 28295 1 1041
2 28296 1 1041
2 28297 1 1041
2 28298 1 1041
2 28299 1 1041
2 28300 1 1041
2 28301 1 1041
2 28302 1 1041
2 28303 1 1041
2 28304 1 1041
2 28305 1 1041
2 28306 1 1041
2 28307 1 1041
2 28308 1 1043
2 28309 1 1043
2 28310 1 1043
2 28311 1 1043
2 28312 1 1043
2 28313 1 1043
2 28314 1 1044
2 28315 1 1044
2 28316 1 1045
2 28317 1 1045
2 28318 1 1047
2 28319 1 1047
2 28320 1 1047
2 28321 1 1047
2 28322 1 1047
2 28323 1 1047
2 28324 1 1047
2 28325 1 1047
2 28326 1 1050
2 28327 1 1050
2 28328 1 1050
2 28329 1 1050
2 28330 1 1056
2 28331 1 1056
2 28332 1 1059
2 28333 1 1059
2 28334 1 1064
2 28335 1 1064
2 28336 1 1072
2 28337 1 1072
2 28338 1 1072
2 28339 1 1072
2 28340 1 1072
2 28341 1 1073
2 28342 1 1073
2 28343 1 1073
2 28344 1 1077
2 28345 1 1077
2 28346 1 1077
2 28347 1 1077
2 28348 1 1077
2 28349 1 1077
2 28350 1 1077
2 28351 1 1077
2 28352 1 1077
2 28353 1 1085
2 28354 1 1085
2 28355 1 1085
2 28356 1 1085
2 28357 1 1085
2 28358 1 1086
2 28359 1 1086
2 28360 1 1086
2 28361 1 1086
2 28362 1 1086
2 28363 1 1086
2 28364 1 1086
2 28365 1 1086
2 28366 1 1088
2 28367 1 1088
2 28368 1 1106
2 28369 1 1106
2 28370 1 1106
2 28371 1 1108
2 28372 1 1108
2 28373 1 1108
2 28374 1 1108
2 28375 1 1109
2 28376 1 1109
2 28377 1 1109
2 28378 1 1109
2 28379 1 1109
2 28380 1 1110
2 28381 1 1110
2 28382 1 1111
2 28383 1 1111
2 28384 1 1114
2 28385 1 1114
2 28386 1 1114
2 28387 1 1118
2 28388 1 1118
2 28389 1 1118
2 28390 1 1118
2 28391 1 1118
2 28392 1 1118
2 28393 1 1118
2 28394 1 1118
2 28395 1 1119
2 28396 1 1119
2 28397 1 1127
2 28398 1 1127
2 28399 1 1127
2 28400 1 1128
2 28401 1 1128
2 28402 1 1128
2 28403 1 1129
2 28404 1 1129
2 28405 1 1130
2 28406 1 1130
2 28407 1 1130
2 28408 1 1133
2 28409 1 1133
2 28410 1 1133
2 28411 1 1133
2 28412 1 1133
2 28413 1 1133
2 28414 1 1133
2 28415 1 1133
2 28416 1 1134
2 28417 1 1134
2 28418 1 1134
2 28419 1 1135
2 28420 1 1135
2 28421 1 1135
2 28422 1 1135
2 28423 1 1135
2 28424 1 1135
2 28425 1 1135
2 28426 1 1135
2 28427 1 1136
2 28428 1 1136
2 28429 1 1136
2 28430 1 1136
2 28431 1 1136
2 28432 1 1136
2 28433 1 1137
2 28434 1 1137
2 28435 1 1148
2 28436 1 1148
2 28437 1 1148
2 28438 1 1148
2 28439 1 1148
2 28440 1 1148
2 28441 1 1151
2 28442 1 1151
2 28443 1 1151
2 28444 1 1151
2 28445 1 1151
2 28446 1 1151
2 28447 1 1151
2 28448 1 1151
2 28449 1 1151
2 28450 1 1151
2 28451 1 1151
2 28452 1 1151
2 28453 1 1151
2 28454 1 1151
2 28455 1 1151
2 28456 1 1152
2 28457 1 1152
2 28458 1 1152
2 28459 1 1152
2 28460 1 1152
2 28461 1 1152
2 28462 1 1153
2 28463 1 1153
2 28464 1 1153
2 28465 1 1154
2 28466 1 1154
2 28467 1 1154
2 28468 1 1154
2 28469 1 1154
2 28470 1 1163
2 28471 1 1163
2 28472 1 1164
2 28473 1 1164
2 28474 1 1164
2 28475 1 1169
2 28476 1 1169
2 28477 1 1178
2 28478 1 1178
2 28479 1 1178
2 28480 1 1178
2 28481 1 1178
2 28482 1 1178
2 28483 1 1178
2 28484 1 1178
2 28485 1 1178
2 28486 1 1178
2 28487 1 1179
2 28488 1 1179
2 28489 1 1179
2 28490 1 1179
2 28491 1 1180
2 28492 1 1180
2 28493 1 1188
2 28494 1 1188
2 28495 1 1188
2 28496 1 1195
2 28497 1 1195
2 28498 1 1205
2 28499 1 1205
2 28500 1 1205
2 28501 1 1206
2 28502 1 1206
2 28503 1 1206
2 28504 1 1206
2 28505 1 1209
2 28506 1 1209
2 28507 1 1209
2 28508 1 1209
2 28509 1 1209
2 28510 1 1223
2 28511 1 1223
2 28512 1 1223
2 28513 1 1223
2 28514 1 1223
2 28515 1 1223
2 28516 1 1225
2 28517 1 1225
2 28518 1 1225
2 28519 1 1225
2 28520 1 1225
2 28521 1 1225
2 28522 1 1225
2 28523 1 1227
2 28524 1 1227
2 28525 1 1228
2 28526 1 1228
2 28527 1 1228
2 28528 1 1228
2 28529 1 1228
2 28530 1 1228
2 28531 1 1228
2 28532 1 1228
2 28533 1 1228
2 28534 1 1228
2 28535 1 1228
2 28536 1 1228
2 28537 1 1228
2 28538 1 1228
2 28539 1 1228
2 28540 1 1228
2 28541 1 1228
2 28542 1 1228
2 28543 1 1228
2 28544 1 1228
2 28545 1 1228
2 28546 1 1228
2 28547 1 1228
2 28548 1 1229
2 28549 1 1229
2 28550 1 1229
2 28551 1 1230
2 28552 1 1230
2 28553 1 1231
2 28554 1 1231
2 28555 1 1232
2 28556 1 1232
2 28557 1 1232
2 28558 1 1232
2 28559 1 1233
2 28560 1 1233
2 28561 1 1233
2 28562 1 1233
2 28563 1 1234
2 28564 1 1234
2 28565 1 1235
2 28566 1 1235
2 28567 1 1238
2 28568 1 1238
2 28569 1 1238
2 28570 1 1238
2 28571 1 1238
2 28572 1 1238
2 28573 1 1238
2 28574 1 1238
2 28575 1 1238
2 28576 1 1238
2 28577 1 1238
2 28578 1 1238
2 28579 1 1238
2 28580 1 1238
2 28581 1 1238
2 28582 1 1238
2 28583 1 1238
2 28584 1 1238
2 28585 1 1238
2 28586 1 1238
2 28587 1 1238
2 28588 1 1238
2 28589 1 1238
2 28590 1 1238
2 28591 1 1238
2 28592 1 1240
2 28593 1 1240
2 28594 1 1248
2 28595 1 1248
2 28596 1 1248
2 28597 1 1248
2 28598 1 1248
2 28599 1 1248
2 28600 1 1255
2 28601 1 1255
2 28602 1 1255
2 28603 1 1256
2 28604 1 1256
2 28605 1 1257
2 28606 1 1257
2 28607 1 1257
2 28608 1 1259
2 28609 1 1259
2 28610 1 1259
2 28611 1 1259
2 28612 1 1260
2 28613 1 1260
2 28614 1 1272
2 28615 1 1272
2 28616 1 1272
2 28617 1 1272
2 28618 1 1272
2 28619 1 1272
2 28620 1 1272
2 28621 1 1272
2 28622 1 1281
2 28623 1 1281
2 28624 1 1281
2 28625 1 1281
2 28626 1 1281
2 28627 1 1281
2 28628 1 1281
2 28629 1 1281
2 28630 1 1282
2 28631 1 1282
2 28632 1 1290
2 28633 1 1290
2 28634 1 1290
2 28635 1 1290
2 28636 1 1290
2 28637 1 1290
2 28638 1 1290
2 28639 1 1290
2 28640 1 1290
2 28641 1 1290
2 28642 1 1290
2 28643 1 1290
2 28644 1 1290
2 28645 1 1290
2 28646 1 1290
2 28647 1 1290
2 28648 1 1290
2 28649 1 1290
2 28650 1 1290
2 28651 1 1290
2 28652 1 1290
2 28653 1 1292
2 28654 1 1292
2 28655 1 1292
2 28656 1 1292
2 28657 1 1292
2 28658 1 1292
2 28659 1 1292
2 28660 1 1300
2 28661 1 1300
2 28662 1 1300
2 28663 1 1300
2 28664 1 1300
2 28665 1 1300
2 28666 1 1300
2 28667 1 1300
2 28668 1 1300
2 28669 1 1300
2 28670 1 1300
2 28671 1 1300
2 28672 1 1300
2 28673 1 1300
2 28674 1 1300
2 28675 1 1300
2 28676 1 1300
2 28677 1 1300
2 28678 1 1300
2 28679 1 1300
2 28680 1 1300
2 28681 1 1300
2 28682 1 1300
2 28683 1 1301
2 28684 1 1301
2 28685 1 1303
2 28686 1 1303
2 28687 1 1303
2 28688 1 1303
2 28689 1 1304
2 28690 1 1304
2 28691 1 1306
2 28692 1 1306
2 28693 1 1306
2 28694 1 1306
2 28695 1 1306
2 28696 1 1306
2 28697 1 1306
2 28698 1 1308
2 28699 1 1308
2 28700 1 1308
2 28701 1 1309
2 28702 1 1309
2 28703 1 1309
2 28704 1 1309
2 28705 1 1309
2 28706 1 1309
2 28707 1 1309
2 28708 1 1309
2 28709 1 1309
2 28710 1 1309
2 28711 1 1309
2 28712 1 1309
2 28713 1 1309
2 28714 1 1314
2 28715 1 1314
2 28716 1 1314
2 28717 1 1314
2 28718 1 1314
2 28719 1 1314
2 28720 1 1314
2 28721 1 1314
2 28722 1 1314
2 28723 1 1314
2 28724 1 1314
2 28725 1 1314
2 28726 1 1315
2 28727 1 1315
2 28728 1 1315
2 28729 1 1315
2 28730 1 1316
2 28731 1 1316
2 28732 1 1316
2 28733 1 1316
2 28734 1 1316
2 28735 1 1317
2 28736 1 1317
2 28737 1 1317
2 28738 1 1318
2 28739 1 1318
2 28740 1 1328
2 28741 1 1328
2 28742 1 1328
2 28743 1 1328
2 28744 1 1328
2 28745 1 1328
2 28746 1 1329
2 28747 1 1329
2 28748 1 1329
2 28749 1 1330
2 28750 1 1330
2 28751 1 1330
2 28752 1 1333
2 28753 1 1333
2 28754 1 1333
2 28755 1 1333
2 28756 1 1333
2 28757 1 1333
2 28758 1 1333
2 28759 1 1333
2 28760 1 1334
2 28761 1 1334
2 28762 1 1335
2 28763 1 1335
2 28764 1 1335
2 28765 1 1335
2 28766 1 1335
2 28767 1 1342
2 28768 1 1342
2 28769 1 1342
2 28770 1 1342
2 28771 1 1343
2 28772 1 1343
2 28773 1 1350
2 28774 1 1350
2 28775 1 1350
2 28776 1 1350
2 28777 1 1351
2 28778 1 1351
2 28779 1 1351
2 28780 1 1351
2 28781 1 1351
2 28782 1 1351
2 28783 1 1351
2 28784 1 1351
2 28785 1 1351
2 28786 1 1351
2 28787 1 1351
2 28788 1 1351
2 28789 1 1351
2 28790 1 1351
2 28791 1 1351
2 28792 1 1351
2 28793 1 1351
2 28794 1 1351
2 28795 1 1351
2 28796 1 1351
2 28797 1 1351
2 28798 1 1351
2 28799 1 1351
2 28800 1 1351
2 28801 1 1351
2 28802 1 1351
2 28803 1 1351
2 28804 1 1351
2 28805 1 1351
2 28806 1 1351
2 28807 1 1351
2 28808 1 1351
2 28809 1 1351
2 28810 1 1351
2 28811 1 1351
2 28812 1 1351
2 28813 1 1351
2 28814 1 1351
2 28815 1 1351
2 28816 1 1351
2 28817 1 1351
2 28818 1 1351
2 28819 1 1351
2 28820 1 1351
2 28821 1 1351
2 28822 1 1351
2 28823 1 1351
2 28824 1 1351
2 28825 1 1351
2 28826 1 1351
2 28827 1 1351
2 28828 1 1351
2 28829 1 1351
2 28830 1 1351
2 28831 1 1351
2 28832 1 1351
2 28833 1 1351
2 28834 1 1351
2 28835 1 1351
2 28836 1 1351
2 28837 1 1351
2 28838 1 1351
2 28839 1 1351
2 28840 1 1351
2 28841 1 1351
2 28842 1 1351
2 28843 1 1351
2 28844 1 1351
2 28845 1 1351
2 28846 1 1351
2 28847 1 1351
2 28848 1 1351
2 28849 1 1351
2 28850 1 1351
2 28851 1 1351
2 28852 1 1351
2 28853 1 1351
2 28854 1 1351
2 28855 1 1351
2 28856 1 1351
2 28857 1 1351
2 28858 1 1351
2 28859 1 1351
2 28860 1 1351
2 28861 1 1351
2 28862 1 1351
2 28863 1 1351
2 28864 1 1351
2 28865 1 1351
2 28866 1 1352
2 28867 1 1352
2 28868 1 1352
2 28869 1 1352
2 28870 1 1353
2 28871 1 1353
2 28872 1 1353
2 28873 1 1353
2 28874 1 1355
2 28875 1 1355
2 28876 1 1355
2 28877 1 1355
2 28878 1 1355
2 28879 1 1356
2 28880 1 1356
2 28881 1 1356
2 28882 1 1367
2 28883 1 1367
2 28884 1 1367
2 28885 1 1367
2 28886 1 1367
2 28887 1 1368
2 28888 1 1368
2 28889 1 1368
2 28890 1 1368
2 28891 1 1368
2 28892 1 1369
2 28893 1 1369
2 28894 1 1376
2 28895 1 1376
2 28896 1 1376
2 28897 1 1376
2 28898 1 1376
2 28899 1 1377
2 28900 1 1377
2 28901 1 1377
2 28902 1 1377
2 28903 1 1387
2 28904 1 1387
2 28905 1 1387
2 28906 1 1396
2 28907 1 1396
2 28908 1 1396
2 28909 1 1396
2 28910 1 1396
2 28911 1 1396
2 28912 1 1396
2 28913 1 1396
2 28914 1 1396
2 28915 1 1396
2 28916 1 1396
2 28917 1 1396
2 28918 1 1396
2 28919 1 1396
2 28920 1 1396
2 28921 1 1397
2 28922 1 1397
2 28923 1 1397
2 28924 1 1400
2 28925 1 1400
2 28926 1 1400
2 28927 1 1400
2 28928 1 1400
2 28929 1 1400
2 28930 1 1400
2 28931 1 1400
2 28932 1 1400
2 28933 1 1400
2 28934 1 1400
2 28935 1 1400
2 28936 1 1401
2 28937 1 1401
2 28938 1 1401
2 28939 1 1402
2 28940 1 1402
2 28941 1 1406
2 28942 1 1406
2 28943 1 1406
2 28944 1 1409
2 28945 1 1409
2 28946 1 1414
2 28947 1 1414
2 28948 1 1423
2 28949 1 1423
2 28950 1 1423
2 28951 1 1424
2 28952 1 1424
2 28953 1 1424
2 28954 1 1424
2 28955 1 1425
2 28956 1 1425
2 28957 1 1426
2 28958 1 1426
2 28959 1 1426
2 28960 1 1426
2 28961 1 1426
2 28962 1 1427
2 28963 1 1427
2 28964 1 1436
2 28965 1 1436
2 28966 1 1436
2 28967 1 1446
2 28968 1 1446
2 28969 1 1446
2 28970 1 1446
2 28971 1 1446
2 28972 1 1446
2 28973 1 1446
2 28974 1 1446
2 28975 1 1446
2 28976 1 1446
2 28977 1 1446
2 28978 1 1446
2 28979 1 1446
2 28980 1 1446
2 28981 1 1446
2 28982 1 1446
2 28983 1 1446
2 28984 1 1446
2 28985 1 1446
2 28986 1 1446
2 28987 1 1446
2 28988 1 1446
2 28989 1 1446
2 28990 1 1446
2 28991 1 1446
2 28992 1 1446
2 28993 1 1446
2 28994 1 1446
2 28995 1 1446
2 28996 1 1446
2 28997 1 1446
2 28998 1 1447
2 28999 1 1447
2 29000 1 1447
2 29001 1 1447
2 29002 1 1447
2 29003 1 1447
2 29004 1 1447
2 29005 1 1447
2 29006 1 1447
2 29007 1 1447
2 29008 1 1447
2 29009 1 1447
2 29010 1 1447
2 29011 1 1447
2 29012 1 1447
2 29013 1 1449
2 29014 1 1449
2 29015 1 1449
2 29016 1 1449
2 29017 1 1449
2 29018 1 1453
2 29019 1 1453
2 29020 1 1454
2 29021 1 1454
2 29022 1 1456
2 29023 1 1456
2 29024 1 1456
2 29025 1 1460
2 29026 1 1460
2 29027 1 1466
2 29028 1 1466
2 29029 1 1481
2 29030 1 1481
2 29031 1 1481
2 29032 1 1481
2 29033 1 1481
2 29034 1 1481
2 29035 1 1481
2 29036 1 1482
2 29037 1 1482
2 29038 1 1482
2 29039 1 1483
2 29040 1 1483
2 29041 1 1485
2 29042 1 1485
2 29043 1 1486
2 29044 1 1486
2 29045 1 1489
2 29046 1 1489
2 29047 1 1489
2 29048 1 1489
2 29049 1 1489
2 29050 1 1489
2 29051 1 1489
2 29052 1 1489
2 29053 1 1489
2 29054 1 1489
2 29055 1 1489
2 29056 1 1489
2 29057 1 1489
2 29058 1 1489
2 29059 1 1489
2 29060 1 1489
2 29061 1 1489
2 29062 1 1489
2 29063 1 1489
2 29064 1 1489
2 29065 1 1490
2 29066 1 1490
2 29067 1 1491
2 29068 1 1491
2 29069 1 1491
2 29070 1 1492
2 29071 1 1492
2 29072 1 1501
2 29073 1 1501
2 29074 1 1501
2 29075 1 1501
2 29076 1 1501
2 29077 1 1501
2 29078 1 1501
2 29079 1 1501
2 29080 1 1501
2 29081 1 1501
2 29082 1 1501
2 29083 1 1501
2 29084 1 1501
2 29085 1 1501
2 29086 1 1501
2 29087 1 1501
2 29088 1 1501
2 29089 1 1501
2 29090 1 1501
2 29091 1 1501
2 29092 1 1501
2 29093 1 1501
2 29094 1 1501
2 29095 1 1501
2 29096 1 1501
2 29097 1 1501
2 29098 1 1501
2 29099 1 1501
2 29100 1 1501
2 29101 1 1501
2 29102 1 1501
2 29103 1 1502
2 29104 1 1502
2 29105 1 1502
2 29106 1 1502
2 29107 1 1502
2 29108 1 1502
2 29109 1 1502
2 29110 1 1502
2 29111 1 1502
2 29112 1 1502
2 29113 1 1502
2 29114 1 1502
2 29115 1 1502
2 29116 1 1502
2 29117 1 1502
2 29118 1 1502
2 29119 1 1502
2 29120 1 1502
2 29121 1 1503
2 29122 1 1503
2 29123 1 1503
2 29124 1 1503
2 29125 1 1503
2 29126 1 1504
2 29127 1 1504
2 29128 1 1504
2 29129 1 1504
2 29130 1 1504
2 29131 1 1505
2 29132 1 1505
2 29133 1 1506
2 29134 1 1506
2 29135 1 1506
2 29136 1 1506
2 29137 1 1507
2 29138 1 1507
2 29139 1 1507
2 29140 1 1507
2 29141 1 1509
2 29142 1 1509
2 29143 1 1509
2 29144 1 1509
2 29145 1 1509
2 29146 1 1510
2 29147 1 1510
2 29148 1 1510
2 29149 1 1520
2 29150 1 1520
2 29151 1 1523
2 29152 1 1523
2 29153 1 1524
2 29154 1 1524
2 29155 1 1524
2 29156 1 1524
2 29157 1 1524
2 29158 1 1524
2 29159 1 1525
2 29160 1 1525
2 29161 1 1532
2 29162 1 1532
2 29163 1 1532
2 29164 1 1532
2 29165 1 1532
2 29166 1 1532
2 29167 1 1532
2 29168 1 1532
2 29169 1 1540
2 29170 1 1540
2 29171 1 1542
2 29172 1 1542
2 29173 1 1542
2 29174 1 1543
2 29175 1 1543
2 29176 1 1543
2 29177 1 1550
2 29178 1 1550
2 29179 1 1550
2 29180 1 1550
2 29181 1 1551
2 29182 1 1551
2 29183 1 1551
2 29184 1 1552
2 29185 1 1552
2 29186 1 1553
2 29187 1 1553
2 29188 1 1568
2 29189 1 1568
2 29190 1 1574
2 29191 1 1574
2 29192 1 1577
2 29193 1 1577
2 29194 1 1577
2 29195 1 1577
2 29196 1 1580
2 29197 1 1580
2 29198 1 1580
2 29199 1 1580
2 29200 1 1580
2 29201 1 1581
2 29202 1 1581
2 29203 1 1604
2 29204 1 1604
2 29205 1 1604
2 29206 1 1604
2 29207 1 1604
2 29208 1 1604
2 29209 1 1604
2 29210 1 1604
2 29211 1 1604
2 29212 1 1604
2 29213 1 1604
2 29214 1 1604
2 29215 1 1604
2 29216 1 1604
2 29217 1 1604
2 29218 1 1604
2 29219 1 1604
2 29220 1 1604
2 29221 1 1604
2 29222 1 1604
2 29223 1 1604
2 29224 1 1604
2 29225 1 1605
2 29226 1 1605
2 29227 1 1605
2 29228 1 1605
2 29229 1 1605
2 29230 1 1605
2 29231 1 1605
2 29232 1 1606
2 29233 1 1606
2 29234 1 1606
2 29235 1 1607
2 29236 1 1607
2 29237 1 1612
2 29238 1 1612
2 29239 1 1612
2 29240 1 1612
2 29241 1 1612
2 29242 1 1613
2 29243 1 1613
2 29244 1 1613
2 29245 1 1624
2 29246 1 1624
2 29247 1 1624
2 29248 1 1624
2 29249 1 1625
2 29250 1 1625
2 29251 1 1625
2 29252 1 1625
2 29253 1 1625
2 29254 1 1625
2 29255 1 1625
2 29256 1 1625
2 29257 1 1625
2 29258 1 1625
2 29259 1 1626
2 29260 1 1626
2 29261 1 1626
2 29262 1 1633
2 29263 1 1633
2 29264 1 1633
2 29265 1 1634
2 29266 1 1634
2 29267 1 1634
2 29268 1 1643
2 29269 1 1643
2 29270 1 1643
2 29271 1 1643
2 29272 1 1651
2 29273 1 1651
2 29274 1 1654
2 29275 1 1654
2 29276 1 1654
2 29277 1 1654
2 29278 1 1655
2 29279 1 1655
2 29280 1 1656
2 29281 1 1656
2 29282 1 1657
2 29283 1 1657
2 29284 1 1657
2 29285 1 1657
2 29286 1 1657
2 29287 1 1657
2 29288 1 1657
2 29289 1 1657
2 29290 1 1657
2 29291 1 1657
2 29292 1 1657
2 29293 1 1657
2 29294 1 1657
2 29295 1 1657
2 29296 1 1658
2 29297 1 1658
2 29298 1 1659
2 29299 1 1659
2 29300 1 1659
2 29301 1 1659
2 29302 1 1659
2 29303 1 1659
2 29304 1 1659
2 29305 1 1659
2 29306 1 1659
2 29307 1 1660
2 29308 1 1660
2 29309 1 1660
2 29310 1 1660
2 29311 1 1669
2 29312 1 1669
2 29313 1 1669
2 29314 1 1670
2 29315 1 1670
2 29316 1 1670
2 29317 1 1670
2 29318 1 1670
2 29319 1 1671
2 29320 1 1671
2 29321 1 1671
2 29322 1 1671
2 29323 1 1685
2 29324 1 1685
2 29325 1 1685
2 29326 1 1685
2 29327 1 1687
2 29328 1 1687
2 29329 1 1688
2 29330 1 1688
2 29331 1 1688
2 29332 1 1698
2 29333 1 1698
2 29334 1 1698
2 29335 1 1698
2 29336 1 1699
2 29337 1 1699
2 29338 1 1700
2 29339 1 1700
2 29340 1 1700
2 29341 1 1701
2 29342 1 1701
2 29343 1 1701
2 29344 1 1701
2 29345 1 1701
2 29346 1 1701
2 29347 1 1702
2 29348 1 1702
2 29349 1 1702
2 29350 1 1702
2 29351 1 1702
2 29352 1 1702
2 29353 1 1702
2 29354 1 1702
2 29355 1 1702
2 29356 1 1702
2 29357 1 1702
2 29358 1 1702
2 29359 1 1702
2 29360 1 1716
2 29361 1 1716
2 29362 1 1716
2 29363 1 1717
2 29364 1 1717
2 29365 1 1717
2 29366 1 1717
2 29367 1 1718
2 29368 1 1718
2 29369 1 1719
2 29370 1 1719
2 29371 1 1719
2 29372 1 1719
2 29373 1 1719
2 29374 1 1719
2 29375 1 1721
2 29376 1 1721
2 29377 1 1722
2 29378 1 1722
2 29379 1 1722
2 29380 1 1722
2 29381 1 1732
2 29382 1 1732
2 29383 1 1747
2 29384 1 1747
2 29385 1 1747
2 29386 1 1747
2 29387 1 1747
2 29388 1 1747
2 29389 1 1747
2 29390 1 1747
2 29391 1 1747
2 29392 1 1747
2 29393 1 1747
2 29394 1 1747
2 29395 1 1748
2 29396 1 1748
2 29397 1 1749
2 29398 1 1749
2 29399 1 1749
2 29400 1 1749
2 29401 1 1754
2 29402 1 1754
2 29403 1 1754
2 29404 1 1755
2 29405 1 1755
2 29406 1 1755
2 29407 1 1755
2 29408 1 1769
2 29409 1 1769
2 29410 1 1769
2 29411 1 1769
2 29412 1 1769
2 29413 1 1769
2 29414 1 1769
2 29415 1 1769
2 29416 1 1770
2 29417 1 1770
2 29418 1 1770
2 29419 1 1772
2 29420 1 1772
2 29421 1 1772
2 29422 1 1772
2 29423 1 1772
2 29424 1 1772
2 29425 1 1772
2 29426 1 1772
2 29427 1 1772
2 29428 1 1772
2 29429 1 1772
2 29430 1 1772
2 29431 1 1772
2 29432 1 1774
2 29433 1 1774
2 29434 1 1774
2 29435 1 1774
2 29436 1 1775
2 29437 1 1775
2 29438 1 1775
2 29439 1 1775
2 29440 1 1775
2 29441 1 1778
2 29442 1 1778
2 29443 1 1778
2 29444 1 1778
2 29445 1 1778
2 29446 1 1778
2 29447 1 1778
2 29448 1 1778
2 29449 1 1778
2 29450 1 1778
2 29451 1 1778
2 29452 1 1778
2 29453 1 1778
2 29454 1 1778
2 29455 1 1778
2 29456 1 1778
2 29457 1 1778
2 29458 1 1778
2 29459 1 1778
2 29460 1 1778
2 29461 1 1778
2 29462 1 1778
2 29463 1 1778
2 29464 1 1778
2 29465 1 1778
2 29466 1 1778
2 29467 1 1778
2 29468 1 1778
2 29469 1 1779
2 29470 1 1779
2 29471 1 1779
2 29472 1 1779
2 29473 1 1779
2 29474 1 1779
2 29475 1 1779
2 29476 1 1779
2 29477 1 1779
2 29478 1 1779
2 29479 1 1779
2 29480 1 1779
2 29481 1 1779
2 29482 1 1779
2 29483 1 1779
2 29484 1 1779
2 29485 1 1779
2 29486 1 1779
2 29487 1 1779
2 29488 1 1779
2 29489 1 1779
2 29490 1 1779
2 29491 1 1779
2 29492 1 1779
2 29493 1 1779
2 29494 1 1779
2 29495 1 1779
2 29496 1 1779
2 29497 1 1779
2 29498 1 1779
2 29499 1 1779
2 29500 1 1779
2 29501 1 1779
2 29502 1 1779
2 29503 1 1779
2 29504 1 1779
2 29505 1 1779
2 29506 1 1779
2 29507 1 1779
2 29508 1 1779
2 29509 1 1779
2 29510 1 1779
2 29511 1 1779
2 29512 1 1779
2 29513 1 1779
2 29514 1 1779
2 29515 1 1779
2 29516 1 1779
2 29517 1 1779
2 29518 1 1779
2 29519 1 1779
2 29520 1 1779
2 29521 1 1779
2 29522 1 1779
2 29523 1 1779
2 29524 1 1779
2 29525 1 1779
2 29526 1 1780
2 29527 1 1780
2 29528 1 1780
2 29529 1 1781
2 29530 1 1781
2 29531 1 1781
2 29532 1 1781
2 29533 1 1783
2 29534 1 1783
2 29535 1 1784
2 29536 1 1784
2 29537 1 1784
2 29538 1 1784
2 29539 1 1784
2 29540 1 1784
2 29541 1 1785
2 29542 1 1785
2 29543 1 1785
2 29544 1 1785
2 29545 1 1786
2 29546 1 1786
2 29547 1 1792
2 29548 1 1792
2 29549 1 1792
2 29550 1 1792
2 29551 1 1792
2 29552 1 1792
2 29553 1 1792
2 29554 1 1792
2 29555 1 1792
2 29556 1 1792
2 29557 1 1792
2 29558 1 1792
2 29559 1 1792
2 29560 1 1792
2 29561 1 1792
2 29562 1 1792
2 29563 1 1792
2 29564 1 1792
2 29565 1 1792
2 29566 1 1792
2 29567 1 1792
2 29568 1 1792
2 29569 1 1792
2 29570 1 1792
2 29571 1 1792
2 29572 1 1792
2 29573 1 1792
2 29574 1 1792
2 29575 1 1792
2 29576 1 1792
2 29577 1 1792
2 29578 1 1792
2 29579 1 1792
2 29580 1 1792
2 29581 1 1793
2 29582 1 1793
2 29583 1 1793
2 29584 1 1793
2 29585 1 1793
2 29586 1 1793
2 29587 1 1793
2 29588 1 1793
2 29589 1 1793
2 29590 1 1793
2 29591 1 1793
2 29592 1 1793
2 29593 1 1793
2 29594 1 1793
2 29595 1 1793
2 29596 1 1793
2 29597 1 1793
2 29598 1 1793
2 29599 1 1793
2 29600 1 1793
2 29601 1 1793
2 29602 1 1793
2 29603 1 1793
2 29604 1 1793
2 29605 1 1793
2 29606 1 1793
2 29607 1 1793
2 29608 1 1793
2 29609 1 1793
2 29610 1 1793
2 29611 1 1794
2 29612 1 1794
2 29613 1 1795
2 29614 1 1795
2 29615 1 1795
2 29616 1 1795
2 29617 1 1795
2 29618 1 1795
2 29619 1 1796
2 29620 1 1796
2 29621 1 1796
2 29622 1 1796
2 29623 1 1796
2 29624 1 1796
2 29625 1 1796
2 29626 1 1796
2 29627 1 1796
2 29628 1 1796
2 29629 1 1796
2 29630 1 1796
2 29631 1 1796
2 29632 1 1797
2 29633 1 1797
2 29634 1 1797
2 29635 1 1797
2 29636 1 1797
2 29637 1 1800
2 29638 1 1800
2 29639 1 1800
2 29640 1 1800
2 29641 1 1800
2 29642 1 1800
2 29643 1 1800
2 29644 1 1802
2 29645 1 1802
2 29646 1 1802
2 29647 1 1802
2 29648 1 1802
2 29649 1 1802
2 29650 1 1802
2 29651 1 1802
2 29652 1 1802
2 29653 1 1802
2 29654 1 1802
2 29655 1 1803
2 29656 1 1803
2 29657 1 1803
2 29658 1 1804
2 29659 1 1804
2 29660 1 1815
2 29661 1 1815
2 29662 1 1815
2 29663 1 1815
2 29664 1 1815
2 29665 1 1816
2 29666 1 1816
2 29667 1 1817
2 29668 1 1817
2 29669 1 1817
2 29670 1 1817
2 29671 1 1818
2 29672 1 1818
2 29673 1 1818
2 29674 1 1818
2 29675 1 1818
2 29676 1 1818
2 29677 1 1818
2 29678 1 1818
2 29679 1 1818
2 29680 1 1818
2 29681 1 1818
2 29682 1 1819
2 29683 1 1819
2 29684 1 1819
2 29685 1 1821
2 29686 1 1821
2 29687 1 1821
2 29688 1 1821
2 29689 1 1822
2 29690 1 1822
2 29691 1 1835
2 29692 1 1835
2 29693 1 1835
2 29694 1 1835
2 29695 1 1835
2 29696 1 1835
2 29697 1 1835
2 29698 1 1835
2 29699 1 1835
2 29700 1 1835
2 29701 1 1835
2 29702 1 1836
2 29703 1 1836
2 29704 1 1836
2 29705 1 1837
2 29706 1 1837
2 29707 1 1837
2 29708 1 1842
2 29709 1 1842
2 29710 1 1842
2 29711 1 1842
2 29712 1 1842
2 29713 1 1842
2 29714 1 1856
2 29715 1 1856
2 29716 1 1856
2 29717 1 1863
2 29718 1 1863
2 29719 1 1863
2 29720 1 1863
2 29721 1 1863
2 29722 1 1863
2 29723 1 1864
2 29724 1 1864
2 29725 1 1864
2 29726 1 1864
2 29727 1 1864
2 29728 1 1864
2 29729 1 1864
2 29730 1 1865
2 29731 1 1865
2 29732 1 1865
2 29733 1 1865
2 29734 1 1879
2 29735 1 1879
2 29736 1 1879
2 29737 1 1879
2 29738 1 1879
2 29739 1 1879
2 29740 1 1879
2 29741 1 1879
2 29742 1 1879
2 29743 1 1879
2 29744 1 1879
2 29745 1 1879
2 29746 1 1880
2 29747 1 1880
2 29748 1 1880
2 29749 1 1880
2 29750 1 1880
2 29751 1 1880
2 29752 1 1880
2 29753 1 1880
2 29754 1 1880
2 29755 1 1880
2 29756 1 1880
2 29757 1 1880
2 29758 1 1880
2 29759 1 1882
2 29760 1 1882
2 29761 1 1882
2 29762 1 1890
2 29763 1 1890
2 29764 1 1890
2 29765 1 1891
2 29766 1 1891
2 29767 1 1891
2 29768 1 1892
2 29769 1 1892
2 29770 1 1892
2 29771 1 1892
2 29772 1 1893
2 29773 1 1893
2 29774 1 1893
2 29775 1 1898
2 29776 1 1898
2 29777 1 1898
2 29778 1 1898
2 29779 1 1898
2 29780 1 1898
2 29781 1 1898
2 29782 1 1898
2 29783 1 1898
2 29784 1 1898
2 29785 1 1898
2 29786 1 1899
2 29787 1 1899
2 29788 1 1899
2 29789 1 1899
2 29790 1 1899
2 29791 1 1899
2 29792 1 1899
2 29793 1 1899
2 29794 1 1899
2 29795 1 1899
2 29796 1 1899
2 29797 1 1899
2 29798 1 1899
2 29799 1 1899
2 29800 1 1899
2 29801 1 1899
2 29802 1 1899
2 29803 1 1900
2 29804 1 1900
2 29805 1 1900
2 29806 1 1900
2 29807 1 1900
2 29808 1 1900
2 29809 1 1901
2 29810 1 1901
2 29811 1 1901
2 29812 1 1902
2 29813 1 1902
2 29814 1 1902
2 29815 1 1902
2 29816 1 1905
2 29817 1 1905
2 29818 1 1906
2 29819 1 1906
2 29820 1 1906
2 29821 1 1907
2 29822 1 1907
2 29823 1 1907
2 29824 1 1907
2 29825 1 1913
2 29826 1 1913
2 29827 1 1913
2 29828 1 1913
2 29829 1 1914
2 29830 1 1914
2 29831 1 1914
2 29832 1 1914
2 29833 1 1921
2 29834 1 1921
2 29835 1 1921
2 29836 1 1921
2 29837 1 1921
2 29838 1 1921
2 29839 1 1921
2 29840 1 1922
2 29841 1 1922
2 29842 1 1922
2 29843 1 1922
2 29844 1 1923
2 29845 1 1923
2 29846 1 1923
2 29847 1 1925
2 29848 1 1925
2 29849 1 1929
2 29850 1 1929
2 29851 1 1929
2 29852 1 1933
2 29853 1 1933
2 29854 1 1933
2 29855 1 1933
2 29856 1 1933
2 29857 1 1933
2 29858 1 1933
2 29859 1 1935
2 29860 1 1935
2 29861 1 1935
2 29862 1 1937
2 29863 1 1937
2 29864 1 1938
2 29865 1 1938
2 29866 1 1938
2 29867 1 1947
2 29868 1 1947
2 29869 1 1947
2 29870 1 1947
2 29871 1 1947
2 29872 1 1947
2 29873 1 1947
2 29874 1 1947
2 29875 1 1947
2 29876 1 1947
2 29877 1 1947
2 29878 1 1949
2 29879 1 1949
2 29880 1 1949
2 29881 1 1957
2 29882 1 1957
2 29883 1 1957
2 29884 1 1957
2 29885 1 1957
2 29886 1 1957
2 29887 1 1958
2 29888 1 1958
2 29889 1 1958
2 29890 1 1958
2 29891 1 1958
2 29892 1 1958
2 29893 1 1958
2 29894 1 1958
2 29895 1 1958
2 29896 1 1958
2 29897 1 1958
2 29898 1 1958
2 29899 1 1958
2 29900 1 1958
2 29901 1 1958
2 29902 1 1958
2 29903 1 1959
2 29904 1 1959
2 29905 1 1959
2 29906 1 1959
2 29907 1 1959
2 29908 1 1959
2 29909 1 1961
2 29910 1 1961
2 29911 1 1961
2 29912 1 1972
2 29913 1 1972
2 29914 1 1972
2 29915 1 1972
2 29916 1 1972
2 29917 1 1972
2 29918 1 1972
2 29919 1 1972
2 29920 1 1972
2 29921 1 1972
2 29922 1 1972
2 29923 1 1972
2 29924 1 1972
2 29925 1 1972
2 29926 1 1972
2 29927 1 1972
2 29928 1 1972
2 29929 1 1972
2 29930 1 1972
2 29931 1 1972
2 29932 1 1973
2 29933 1 1973
2 29934 1 1973
2 29935 1 1974
2 29936 1 1974
2 29937 1 1974
2 29938 1 1974
2 29939 1 1974
2 29940 1 1975
2 29941 1 1975
2 29942 1 1975
2 29943 1 1975
2 29944 1 1976
2 29945 1 1976
2 29946 1 1981
2 29947 1 1981
2 29948 1 1981
2 29949 1 1981
2 29950 1 1981
2 29951 1 1982
2 29952 1 1982
2 29953 1 1986
2 29954 1 1986
2 29955 1 1987
2 29956 1 1987
2 29957 1 1987
2 29958 1 1987
2 29959 1 1987
2 29960 1 1987
2 29961 1 1987
2 29962 1 1987
2 29963 1 1987
2 29964 1 1988
2 29965 1 1988
2 29966 1 1988
2 29967 1 1988
2 29968 1 1989
2 29969 1 1989
2 29970 1 1989
2 29971 1 1992
2 29972 1 1992
2 29973 1 2001
2 29974 1 2001
2 29975 1 2002
2 29976 1 2002
2 29977 1 2002
2 29978 1 2002
2 29979 1 2003
2 29980 1 2003
2 29981 1 2003
2 29982 1 2004
2 29983 1 2004
2 29984 1 2004
2 29985 1 2004
2 29986 1 2004
2 29987 1 2004
2 29988 1 2004
2 29989 1 2004
2 29990 1 2013
2 29991 1 2013
2 29992 1 2013
2 29993 1 2022
2 29994 1 2022
2 29995 1 2022
2 29996 1 2024
2 29997 1 2024
2 29998 1 2026
2 29999 1 2026
2 30000 1 2026
2 30001 1 2026
2 30002 1 2026
2 30003 1 2026
2 30004 1 2026
2 30005 1 2028
2 30006 1 2028
2 30007 1 2028
2 30008 1 2029
2 30009 1 2029
2 30010 1 2034
2 30011 1 2034
2 30012 1 2034
2 30013 1 2034
2 30014 1 2034
2 30015 1 2035
2 30016 1 2035
2 30017 1 2047
2 30018 1 2047
2 30019 1 2047
2 30020 1 2048
2 30021 1 2048
2 30022 1 2056
2 30023 1 2056
2 30024 1 2056
2 30025 1 2056
2 30026 1 2056
2 30027 1 2056
2 30028 1 2056
2 30029 1 2061
2 30030 1 2061
2 30031 1 2061
2 30032 1 2066
2 30033 1 2066
2 30034 1 2068
2 30035 1 2068
2 30036 1 2068
2 30037 1 2069
2 30038 1 2069
2 30039 1 2069
2 30040 1 2069
2 30041 1 2070
2 30042 1 2070
2 30043 1 2070
2 30044 1 2070
2 30045 1 2070
2 30046 1 2070
2 30047 1 2070
2 30048 1 2071
2 30049 1 2071
2 30050 1 2071
2 30051 1 2073
2 30052 1 2073
2 30053 1 2073
2 30054 1 2073
2 30055 1 2077
2 30056 1 2077
2 30057 1 2077
2 30058 1 2077
2 30059 1 2077
2 30060 1 2080
2 30061 1 2080
2 30062 1 2083
2 30063 1 2083
2 30064 1 2083
2 30065 1 2083
2 30066 1 2083
2 30067 1 2083
2 30068 1 2083
2 30069 1 2084
2 30070 1 2084
2 30071 1 2084
2 30072 1 2085
2 30073 1 2085
2 30074 1 2085
2 30075 1 2093
2 30076 1 2093
2 30077 1 2093
2 30078 1 2093
2 30079 1 2093
2 30080 1 2093
2 30081 1 2093
2 30082 1 2093
2 30083 1 2094
2 30084 1 2094
2 30085 1 2094
2 30086 1 2097
2 30087 1 2097
2 30088 1 2097
2 30089 1 2097
2 30090 1 2097
2 30091 1 2097
2 30092 1 2098
2 30093 1 2098
2 30094 1 2121
2 30095 1 2121
2 30096 1 2121
2 30097 1 2121
2 30098 1 2121
2 30099 1 2121
2 30100 1 2122
2 30101 1 2122
2 30102 1 2122
2 30103 1 2123
2 30104 1 2123
2 30105 1 2123
2 30106 1 2123
2 30107 1 2123
2 30108 1 2123
2 30109 1 2123
2 30110 1 2123
2 30111 1 2123
2 30112 1 2124
2 30113 1 2124
2 30114 1 2124
2 30115 1 2124
2 30116 1 2124
2 30117 1 2124
2 30118 1 2124
2 30119 1 2125
2 30120 1 2125
2 30121 1 2125
2 30122 1 2125
2 30123 1 2125
2 30124 1 2125
2 30125 1 2125
2 30126 1 2126
2 30127 1 2126
2 30128 1 2126
2 30129 1 2126
2 30130 1 2128
2 30131 1 2128
2 30132 1 2129
2 30133 1 2129
2 30134 1 2129
2 30135 1 2129
2 30136 1 2129
2 30137 1 2130
2 30138 1 2130
2 30139 1 2132
2 30140 1 2132
2 30141 1 2132
2 30142 1 2139
2 30143 1 2139
2 30144 1 2139
2 30145 1 2139
2 30146 1 2139
2 30147 1 2139
2 30148 1 2140
2 30149 1 2140
2 30150 1 2149
2 30151 1 2149
2 30152 1 2152
2 30153 1 2152
2 30154 1 2152
2 30155 1 2152
2 30156 1 2152
2 30157 1 2155
2 30158 1 2155
2 30159 1 2155
2 30160 1 2169
2 30161 1 2169
2 30162 1 2169
2 30163 1 2169
2 30164 1 2169
2 30165 1 2169
2 30166 1 2169
2 30167 1 2169
2 30168 1 2169
2 30169 1 2169
2 30170 1 2169
2 30171 1 2169
2 30172 1 2169
2 30173 1 2169
2 30174 1 2169
2 30175 1 2169
2 30176 1 2169
2 30177 1 2169
2 30178 1 2169
2 30179 1 2171
2 30180 1 2171
2 30181 1 2171
2 30182 1 2171
2 30183 1 2172
2 30184 1 2172
2 30185 1 2172
2 30186 1 2173
2 30187 1 2173
2 30188 1 2176
2 30189 1 2176
2 30190 1 2176
2 30191 1 2176
2 30192 1 2179
2 30193 1 2179
2 30194 1 2179
2 30195 1 2182
2 30196 1 2182
2 30197 1 2183
2 30198 1 2183
2 30199 1 2183
2 30200 1 2183
2 30201 1 2186
2 30202 1 2186
2 30203 1 2186
2 30204 1 2190
2 30205 1 2190
2 30206 1 2190
2 30207 1 2190
2 30208 1 2190
2 30209 1 2190
2 30210 1 2190
2 30211 1 2190
2 30212 1 2191
2 30213 1 2191
2 30214 1 2191
2 30215 1 2198
2 30216 1 2198
2 30217 1 2200
2 30218 1 2200
2 30219 1 2200
2 30220 1 2200
2 30221 1 2200
2 30222 1 2200
2 30223 1 2200
2 30224 1 2200
2 30225 1 2200
2 30226 1 2200
2 30227 1 2202
2 30228 1 2202
2 30229 1 2202
2 30230 1 2202
2 30231 1 2203
2 30232 1 2203
2 30233 1 2203
2 30234 1 2217
2 30235 1 2217
2 30236 1 2217
2 30237 1 2217
2 30238 1 2218
2 30239 1 2218
2 30240 1 2218
2 30241 1 2218
2 30242 1 2218
2 30243 1 2218
2 30244 1 2218
2 30245 1 2218
2 30246 1 2218
2 30247 1 2218
2 30248 1 2218
2 30249 1 2218
2 30250 1 2218
2 30251 1 2218
2 30252 1 2218
2 30253 1 2218
2 30254 1 2218
2 30255 1 2219
2 30256 1 2219
2 30257 1 2219
2 30258 1 2219
2 30259 1 2219
2 30260 1 2220
2 30261 1 2220
2 30262 1 2220
2 30263 1 2222
2 30264 1 2222
2 30265 1 2224
2 30266 1 2224
2 30267 1 2224
2 30268 1 2224
2 30269 1 2224
2 30270 1 2224
2 30271 1 2224
2 30272 1 2225
2 30273 1 2225
2 30274 1 2225
2 30275 1 2225
2 30276 1 2225
2 30277 1 2226
2 30278 1 2226
2 30279 1 2229
2 30280 1 2229
2 30281 1 2229
2 30282 1 2229
2 30283 1 2229
2 30284 1 2230
2 30285 1 2230
2 30286 1 2230
2 30287 1 2230
2 30288 1 2230
2 30289 1 2231
2 30290 1 2231
2 30291 1 2231
2 30292 1 2231
2 30293 1 2231
2 30294 1 2232
2 30295 1 2232
2 30296 1 2232
2 30297 1 2240
2 30298 1 2240
2 30299 1 2240
2 30300 1 2240
2 30301 1 2240
2 30302 1 2240
2 30303 1 2240
2 30304 1 2240
2 30305 1 2240
2 30306 1 2240
2 30307 1 2240
2 30308 1 2240
2 30309 1 2240
2 30310 1 2240
2 30311 1 2241
2 30312 1 2241
2 30313 1 2241
2 30314 1 2241
2 30315 1 2241
2 30316 1 2241
2 30317 1 2243
2 30318 1 2243
2 30319 1 2243
2 30320 1 2243
2 30321 1 2243
2 30322 1 2243
2 30323 1 2243
2 30324 1 2244
2 30325 1 2244
2 30326 1 2258
2 30327 1 2258
2 30328 1 2260
2 30329 1 2260
2 30330 1 2260
2 30331 1 2261
2 30332 1 2261
2 30333 1 2261
2 30334 1 2261
2 30335 1 2261
2 30336 1 2261
2 30337 1 2261
2 30338 1 2261
2 30339 1 2261
2 30340 1 2264
2 30341 1 2264
2 30342 1 2264
2 30343 1 2265
2 30344 1 2265
2 30345 1 2267
2 30346 1 2267
2 30347 1 2267
2 30348 1 2267
2 30349 1 2267
2 30350 1 2267
2 30351 1 2274
2 30352 1 2274
2 30353 1 2274
2 30354 1 2277
2 30355 1 2277
2 30356 1 2277
2 30357 1 2277
2 30358 1 2277
2 30359 1 2278
2 30360 1 2278
2 30361 1 2278
2 30362 1 2293
2 30363 1 2293
2 30364 1 2293
2 30365 1 2294
2 30366 1 2294
2 30367 1 2297
2 30368 1 2297
2 30369 1 2301
2 30370 1 2301
2 30371 1 2304
2 30372 1 2304
2 30373 1 2304
2 30374 1 2304
2 30375 1 2312
2 30376 1 2312
2 30377 1 2312
2 30378 1 2312
2 30379 1 2312
2 30380 1 2312
2 30381 1 2321
2 30382 1 2321
2 30383 1 2321
2 30384 1 2322
2 30385 1 2322
2 30386 1 2322
2 30387 1 2323
2 30388 1 2323
2 30389 1 2323
2 30390 1 2323
2 30391 1 2323
2 30392 1 2324
2 30393 1 2324
2 30394 1 2324
2 30395 1 2325
2 30396 1 2325
2 30397 1 2338
2 30398 1 2338
2 30399 1 2338
2 30400 1 2339
2 30401 1 2339
2 30402 1 2339
2 30403 1 2340
2 30404 1 2340
2 30405 1 2340
2 30406 1 2340
2 30407 1 2341
2 30408 1 2341
2 30409 1 2360
2 30410 1 2360
2 30411 1 2361
2 30412 1 2361
2 30413 1 2363
2 30414 1 2363
2 30415 1 2367
2 30416 1 2367
2 30417 1 2367
2 30418 1 2367
2 30419 1 2371
2 30420 1 2371
2 30421 1 2371
2 30422 1 2374
2 30423 1 2374
2 30424 1 2380
2 30425 1 2380
2 30426 1 2387
2 30427 1 2387
2 30428 1 2387
2 30429 1 2388
2 30430 1 2388
2 30431 1 2396
2 30432 1 2396
2 30433 1 2402
2 30434 1 2402
2 30435 1 2402
2 30436 1 2402
2 30437 1 2402
2 30438 1 2402
2 30439 1 2402
2 30440 1 2403
2 30441 1 2403
2 30442 1 2403
2 30443 1 2403
2 30444 1 2403
2 30445 1 2403
2 30446 1 2403
2 30447 1 2407
2 30448 1 2407
2 30449 1 2407
2 30450 1 2407
2 30451 1 2409
2 30452 1 2409
2 30453 1 2410
2 30454 1 2410
2 30455 1 2419
2 30456 1 2419
2 30457 1 2420
2 30458 1 2420
2 30459 1 2421
2 30460 1 2421
2 30461 1 2421
2 30462 1 2421
2 30463 1 2421
2 30464 1 2422
2 30465 1 2422
2 30466 1 2423
2 30467 1 2423
2 30468 1 2423
2 30469 1 2423
2 30470 1 2423
2 30471 1 2423
2 30472 1 2434
2 30473 1 2434
2 30474 1 2435
2 30475 1 2435
2 30476 1 2443
2 30477 1 2443
2 30478 1 2444
2 30479 1 2444
2 30480 1 2444
2 30481 1 2444
2 30482 1 2444
2 30483 1 2445
2 30484 1 2445
2 30485 1 2456
2 30486 1 2456
2 30487 1 2456
2 30488 1 2465
2 30489 1 2465
2 30490 1 2465
2 30491 1 2466
2 30492 1 2466
2 30493 1 2471
2 30494 1 2471
2 30495 1 2471
2 30496 1 2471
2 30497 1 2471
2 30498 1 2471
2 30499 1 2471
2 30500 1 2471
2 30501 1 2488
2 30502 1 2488
2 30503 1 2488
2 30504 1 2507
2 30505 1 2507
2 30506 1 2507
2 30507 1 2507
2 30508 1 2508
2 30509 1 2508
2 30510 1 2509
2 30511 1 2509
2 30512 1 2511
2 30513 1 2511
2 30514 1 2515
2 30515 1 2515
2 30516 1 2515
2 30517 1 2515
2 30518 1 2515
2 30519 1 2515
2 30520 1 2515
2 30521 1 2515
2 30522 1 2515
2 30523 1 2515
2 30524 1 2515
2 30525 1 2515
2 30526 1 2515
2 30527 1 2515
2 30528 1 2515
2 30529 1 2515
2 30530 1 2518
2 30531 1 2518
2 30532 1 2518
2 30533 1 2518
2 30534 1 2530
2 30535 1 2530
2 30536 1 2530
2 30537 1 2530
2 30538 1 2530
2 30539 1 2530
2 30540 1 2530
2 30541 1 2531
2 30542 1 2531
2 30543 1 2531
2 30544 1 2531
2 30545 1 2532
2 30546 1 2532
2 30547 1 2532
2 30548 1 2532
2 30549 1 2532
2 30550 1 2541
2 30551 1 2541
2 30552 1 2541
2 30553 1 2541
2 30554 1 2542
2 30555 1 2542
2 30556 1 2544
2 30557 1 2544
2 30558 1 2545
2 30559 1 2545
2 30560 1 2545
2 30561 1 2549
2 30562 1 2549
2 30563 1 2549
2 30564 1 2549
2 30565 1 2549
2 30566 1 2549
2 30567 1 2549
2 30568 1 2549
2 30569 1 2549
2 30570 1 2549
2 30571 1 2550
2 30572 1 2550
2 30573 1 2550
2 30574 1 2550
2 30575 1 2550
2 30576 1 2550
2 30577 1 2550
2 30578 1 2550
2 30579 1 2550
2 30580 1 2551
2 30581 1 2551
2 30582 1 2551
2 30583 1 2551
2 30584 1 2551
2 30585 1 2563
2 30586 1 2563
2 30587 1 2563
2 30588 1 2564
2 30589 1 2564
2 30590 1 2566
2 30591 1 2566
2 30592 1 2566
2 30593 1 2566
2 30594 1 2579
2 30595 1 2579
2 30596 1 2579
2 30597 1 2579
2 30598 1 2579
2 30599 1 2579
2 30600 1 2580
2 30601 1 2580
2 30602 1 2580
2 30603 1 2580
2 30604 1 2580
2 30605 1 2580
2 30606 1 2580
2 30607 1 2580
2 30608 1 2580
2 30609 1 2580
2 30610 1 2580
2 30611 1 2580
2 30612 1 2580
2 30613 1 2580
2 30614 1 2580
2 30615 1 2580
2 30616 1 2580
2 30617 1 2580
2 30618 1 2580
2 30619 1 2580
2 30620 1 2580
2 30621 1 2581
2 30622 1 2581
2 30623 1 2581
2 30624 1 2581
2 30625 1 2585
2 30626 1 2585
2 30627 1 2585
2 30628 1 2585
2 30629 1 2585
2 30630 1 2585
2 30631 1 2585
2 30632 1 2585
2 30633 1 2585
2 30634 1 2585
2 30635 1 2585
2 30636 1 2585
2 30637 1 2585
2 30638 1 2586
2 30639 1 2586
2 30640 1 2591
2 30641 1 2591
2 30642 1 2594
2 30643 1 2594
2 30644 1 2595
2 30645 1 2595
2 30646 1 2603
2 30647 1 2603
2 30648 1 2603
2 30649 1 2603
2 30650 1 2603
2 30651 1 2604
2 30652 1 2604
2 30653 1 2604
2 30654 1 2605
2 30655 1 2605
2 30656 1 2605
2 30657 1 2605
2 30658 1 2606
2 30659 1 2606
2 30660 1 2609
2 30661 1 2609
2 30662 1 2609
2 30663 1 2609
2 30664 1 2609
2 30665 1 2609
2 30666 1 2609
2 30667 1 2609
2 30668 1 2618
2 30669 1 2618
2 30670 1 2623
2 30671 1 2623
2 30672 1 2623
2 30673 1 2625
2 30674 1 2625
2 30675 1 2626
2 30676 1 2626
2 30677 1 2626
2 30678 1 2638
2 30679 1 2638
2 30680 1 2638
2 30681 1 2638
2 30682 1 2638
2 30683 1 2640
2 30684 1 2640
2 30685 1 2641
2 30686 1 2641
2 30687 1 2642
2 30688 1 2642
2 30689 1 2652
2 30690 1 2652
2 30691 1 2652
2 30692 1 2654
2 30693 1 2654
2 30694 1 2655
2 30695 1 2655
2 30696 1 2655
2 30697 1 2655
2 30698 1 2656
2 30699 1 2656
2 30700 1 2659
2 30701 1 2659
2 30702 1 2668
2 30703 1 2668
2 30704 1 2668
2 30705 1 2668
2 30706 1 2669
2 30707 1 2669
2 30708 1 2669
2 30709 1 2669
2 30710 1 2670
2 30711 1 2670
2 30712 1 2683
2 30713 1 2683
2 30714 1 2683
2 30715 1 2691
2 30716 1 2691
2 30717 1 2691
2 30718 1 2691
2 30719 1 2691
2 30720 1 2691
2 30721 1 2699
2 30722 1 2699
2 30723 1 2699
2 30724 1 2699
2 30725 1 2700
2 30726 1 2700
2 30727 1 2716
2 30728 1 2716
2 30729 1 2716
2 30730 1 2716
2 30731 1 2717
2 30732 1 2717
2 30733 1 2717
2 30734 1 2717
2 30735 1 2720
2 30736 1 2720
2 30737 1 2720
2 30738 1 2720
2 30739 1 2720
2 30740 1 2721
2 30741 1 2721
2 30742 1 2730
2 30743 1 2730
2 30744 1 2730
2 30745 1 2730
2 30746 1 2730
2 30747 1 2730
2 30748 1 2731
2 30749 1 2731
2 30750 1 2743
2 30751 1 2743
2 30752 1 2744
2 30753 1 2744
2 30754 1 2747
2 30755 1 2747
2 30756 1 2747
2 30757 1 2747
2 30758 1 2747
2 30759 1 2748
2 30760 1 2748
2 30761 1 2759
2 30762 1 2759
2 30763 1 2759
2 30764 1 2759
2 30765 1 2759
2 30766 1 2759
2 30767 1 2759
2 30768 1 2769
2 30769 1 2769
2 30770 1 2770
2 30771 1 2770
2 30772 1 2770
2 30773 1 2770
2 30774 1 2770
2 30775 1 2771
2 30776 1 2771
2 30777 1 2772
2 30778 1 2772
2 30779 1 2772
2 30780 1 2772
2 30781 1 2772
2 30782 1 2772
2 30783 1 2772
2 30784 1 2772
2 30785 1 2772
2 30786 1 2773
2 30787 1 2773
2 30788 1 2773
2 30789 1 2786
2 30790 1 2786
2 30791 1 2786
2 30792 1 2787
2 30793 1 2787
2 30794 1 2788
2 30795 1 2788
2 30796 1 2790
2 30797 1 2790
2 30798 1 2799
2 30799 1 2799
2 30800 1 2806
2 30801 1 2806
2 30802 1 2806
2 30803 1 2815
2 30804 1 2815
2 30805 1 2823
2 30806 1 2823
2 30807 1 2823
2 30808 1 2831
2 30809 1 2831
2 30810 1 2831
2 30811 1 2831
2 30812 1 2831
2 30813 1 2851
2 30814 1 2851
2 30815 1 2852
2 30816 1 2852
2 30817 1 2854
2 30818 1 2854
2 30819 1 2856
2 30820 1 2856
2 30821 1 2856
2 30822 1 2856
2 30823 1 2859
2 30824 1 2859
2 30825 1 2859
2 30826 1 2859
2 30827 1 2870
2 30828 1 2870
2 30829 1 2871
2 30830 1 2871
2 30831 1 2871
2 30832 1 2872
2 30833 1 2872
2 30834 1 2872
2 30835 1 2880
2 30836 1 2880
2 30837 1 2881
2 30838 1 2881
2 30839 1 2882
2 30840 1 2882
2 30841 1 2882
2 30842 1 2883
2 30843 1 2883
2 30844 1 2883
2 30845 1 2883
2 30846 1 2886
2 30847 1 2886
2 30848 1 2886
2 30849 1 2887
2 30850 1 2887
2 30851 1 2889
2 30852 1 2889
2 30853 1 2889
2 30854 1 2889
2 30855 1 2889
2 30856 1 2889
2 30857 1 2891
2 30858 1 2891
2 30859 1 2894
2 30860 1 2894
2 30861 1 2895
2 30862 1 2895
2 30863 1 2895
2 30864 1 2895
2 30865 1 2895
2 30866 1 2895
2 30867 1 2895
2 30868 1 2903
2 30869 1 2903
2 30870 1 2903
2 30871 1 2904
2 30872 1 2904
2 30873 1 2905
2 30874 1 2905
2 30875 1 2906
2 30876 1 2906
2 30877 1 2906
2 30878 1 2906
2 30879 1 2917
2 30880 1 2917
2 30881 1 2917
2 30882 1 2925
2 30883 1 2925
2 30884 1 2925
2 30885 1 2933
2 30886 1 2933
2 30887 1 2933
2 30888 1 2933
2 30889 1 2933
2 30890 1 2933
2 30891 1 2933
2 30892 1 2933
2 30893 1 2933
2 30894 1 2934
2 30895 1 2934
2 30896 1 2934
2 30897 1 2934
2 30898 1 2934
2 30899 1 2934
2 30900 1 2934
2 30901 1 2934
2 30902 1 2935
2 30903 1 2935
2 30904 1 2935
2 30905 1 2936
2 30906 1 2936
2 30907 1 2945
2 30908 1 2945
2 30909 1 2945
2 30910 1 2945
2 30911 1 2945
2 30912 1 2945
2 30913 1 2945
2 30914 1 2946
2 30915 1 2946
2 30916 1 2948
2 30917 1 2948
2 30918 1 2948
2 30919 1 2948
2 30920 1 2948
2 30921 1 2948
2 30922 1 2948
2 30923 1 2948
2 30924 1 2948
2 30925 1 2948
2 30926 1 2948
2 30927 1 2948
2 30928 1 2948
2 30929 1 2948
2 30930 1 2948
2 30931 1 2948
2 30932 1 2948
2 30933 1 2948
2 30934 1 2950
2 30935 1 2950
2 30936 1 2951
2 30937 1 2951
2 30938 1 2951
2 30939 1 2951
2 30940 1 2951
2 30941 1 2952
2 30942 1 2952
2 30943 1 2953
2 30944 1 2953
2 30945 1 2956
2 30946 1 2956
2 30947 1 2956
2 30948 1 2965
2 30949 1 2965
2 30950 1 2965
2 30951 1 2965
2 30952 1 2966
2 30953 1 2966
2 30954 1 2966
2 30955 1 2966
2 30956 1 2966
2 30957 1 2969
2 30958 1 2969
2 30959 1 2969
2 30960 1 2969
2 30961 1 2969
2 30962 1 2969
2 30963 1 2969
2 30964 1 2969
2 30965 1 2969
2 30966 1 2970
2 30967 1 2970
2 30968 1 2971
2 30969 1 2971
2 30970 1 2988
2 30971 1 2988
2 30972 1 2988
2 30973 1 2988
2 30974 1 2988
2 30975 1 2988
2 30976 1 2988
2 30977 1 2988
2 30978 1 2990
2 30979 1 2990
2 30980 1 2990
2 30981 1 2992
2 30982 1 2992
2 30983 1 2995
2 30984 1 2995
2 30985 1 2995
2 30986 1 2996
2 30987 1 2996
2 30988 1 2997
2 30989 1 2997
2 30990 1 2998
2 30991 1 2998
2 30992 1 2999
2 30993 1 2999
2 30994 1 3006
2 30995 1 3006
2 30996 1 3007
2 30997 1 3007
2 30998 1 3007
2 30999 1 3007
2 31000 1 3010
2 31001 1 3010
2 31002 1 3014
2 31003 1 3014
2 31004 1 3019
2 31005 1 3019
2 31006 1 3022
2 31007 1 3022
2 31008 1 3038
2 31009 1 3038
2 31010 1 3038
2 31011 1 3040
2 31012 1 3040
2 31013 1 3040
2 31014 1 3040
2 31015 1 3040
2 31016 1 3042
2 31017 1 3042
2 31018 1 3043
2 31019 1 3043
2 31020 1 3043
2 31021 1 3044
2 31022 1 3044
2 31023 1 3052
2 31024 1 3052
2 31025 1 3052
2 31026 1 3052
2 31027 1 3052
2 31028 1 3052
2 31029 1 3053
2 31030 1 3053
2 31031 1 3053
2 31032 1 3053
2 31033 1 3057
2 31034 1 3057
2 31035 1 3058
2 31036 1 3058
2 31037 1 3059
2 31038 1 3059
2 31039 1 3059
2 31040 1 3059
2 31041 1 3060
2 31042 1 3060
2 31043 1 3060
2 31044 1 3060
2 31045 1 3060
2 31046 1 3060
2 31047 1 3060
2 31048 1 3072
2 31049 1 3072
2 31050 1 3075
2 31051 1 3075
2 31052 1 3078
2 31053 1 3078
2 31054 1 3078
2 31055 1 3078
2 31056 1 3079
2 31057 1 3079
2 31058 1 3079
2 31059 1 3079
2 31060 1 3080
2 31061 1 3080
2 31062 1 3080
2 31063 1 3080
2 31064 1 3083
2 31065 1 3083
2 31066 1 3083
2 31067 1 3083
2 31068 1 3083
2 31069 1 3092
2 31070 1 3092
2 31071 1 3092
2 31072 1 3092
2 31073 1 3094
2 31074 1 3094
2 31075 1 3097
2 31076 1 3097
2 31077 1 3100
2 31078 1 3100
2 31079 1 3100
2 31080 1 3100
2 31081 1 3100
2 31082 1 3100
2 31083 1 3102
2 31084 1 3102
2 31085 1 3102
2 31086 1 3104
2 31087 1 3104
2 31088 1 3105
2 31089 1 3105
2 31090 1 3111
2 31091 1 3111
2 31092 1 3111
2 31093 1 3128
2 31094 1 3128
2 31095 1 3156
2 31096 1 3156
2 31097 1 3158
2 31098 1 3158
2 31099 1 3163
2 31100 1 3163
2 31101 1 3163
2 31102 1 3163
2 31103 1 3181
2 31104 1 3181
2 31105 1 3182
2 31106 1 3182
2 31107 1 3201
2 31108 1 3201
2 31109 1 3206
2 31110 1 3206
2 31111 1 3207
2 31112 1 3207
2 31113 1 3207
2 31114 1 3225
2 31115 1 3225
2 31116 1 3234
2 31117 1 3234
2 31118 1 3243
2 31119 1 3243
2 31120 1 3243
2 31121 1 3243
2 31122 1 3258
2 31123 1 3258
2 31124 1 3263
2 31125 1 3263
2 31126 1 3265
2 31127 1 3265
2 31128 1 3271
2 31129 1 3271
2 31130 1 3271
2 31131 1 3271
2 31132 1 3271
2 31133 1 3271
2 31134 1 3272
2 31135 1 3272
2 31136 1 3274
2 31137 1 3274
2 31138 1 3292
2 31139 1 3292
2 31140 1 3292
2 31141 1 3292
2 31142 1 3292
2 31143 1 3292
2 31144 1 3293
2 31145 1 3293
2 31146 1 3294
2 31147 1 3294
2 31148 1 3294
2 31149 1 3295
2 31150 1 3295
2 31151 1 3295
2 31152 1 3296
2 31153 1 3296
2 31154 1 3296
2 31155 1 3299
2 31156 1 3299
2 31157 1 3299
2 31158 1 3299
2 31159 1 3300
2 31160 1 3300
2 31161 1 3300
2 31162 1 3300
2 31163 1 3308
2 31164 1 3308
2 31165 1 3308
2 31166 1 3308
2 31167 1 3308
2 31168 1 3308
2 31169 1 3308
2 31170 1 3308
2 31171 1 3308
2 31172 1 3308
2 31173 1 3308
2 31174 1 3308
2 31175 1 3308
2 31176 1 3308
2 31177 1 3309
2 31178 1 3309
2 31179 1 3319
2 31180 1 3319
2 31181 1 3319
2 31182 1 3319
2 31183 1 3319
2 31184 1 3319
2 31185 1 3319
2 31186 1 3319
2 31187 1 3320
2 31188 1 3320
2 31189 1 3320
2 31190 1 3320
2 31191 1 3320
2 31192 1 3320
2 31193 1 3320
2 31194 1 3320
2 31195 1 3320
2 31196 1 3320
2 31197 1 3320
2 31198 1 3320
2 31199 1 3320
2 31200 1 3320
2 31201 1 3320
2 31202 1 3322
2 31203 1 3322
2 31204 1 3325
2 31205 1 3325
2 31206 1 3328
2 31207 1 3328
2 31208 1 3328
2 31209 1 3329
2 31210 1 3329
2 31211 1 3329
2 31212 1 3329
2 31213 1 3330
2 31214 1 3330
2 31215 1 3330
2 31216 1 3339
2 31217 1 3339
2 31218 1 3339
2 31219 1 3340
2 31220 1 3340
2 31221 1 3341
2 31222 1 3341
2 31223 1 3341
2 31224 1 3341
2 31225 1 3342
2 31226 1 3342
2 31227 1 3348
2 31228 1 3348
2 31229 1 3348
2 31230 1 3348
2 31231 1 3348
2 31232 1 3348
2 31233 1 3349
2 31234 1 3349
2 31235 1 3349
2 31236 1 3349
2 31237 1 3349
2 31238 1 3350
2 31239 1 3350
2 31240 1 3351
2 31241 1 3351
2 31242 1 3351
2 31243 1 3351
2 31244 1 3351
2 31245 1 3351
2 31246 1 3351
2 31247 1 3351
2 31248 1 3351
2 31249 1 3351
2 31250 1 3351
2 31251 1 3351
2 31252 1 3351
2 31253 1 3351
2 31254 1 3351
2 31255 1 3352
2 31256 1 3352
2 31257 1 3352
2 31258 1 3352
2 31259 1 3352
2 31260 1 3353
2 31261 1 3353
2 31262 1 3353
2 31263 1 3353
2 31264 1 3361
2 31265 1 3361
2 31266 1 3361
2 31267 1 3389
2 31268 1 3389
2 31269 1 3389
2 31270 1 3389
2 31271 1 3389
2 31272 1 3389
2 31273 1 3389
2 31274 1 3390
2 31275 1 3390
2 31276 1 3391
2 31277 1 3391
2 31278 1 3391
2 31279 1 3400
2 31280 1 3400
2 31281 1 3400
2 31282 1 3403
2 31283 1 3403
2 31284 1 3403
2 31285 1 3403
2 31286 1 3403
2 31287 1 3404
2 31288 1 3404
2 31289 1 3404
2 31290 1 3404
2 31291 1 3404
2 31292 1 3404
2 31293 1 3404
2 31294 1 3404
2 31295 1 3404
2 31296 1 3404
2 31297 1 3404
2 31298 1 3404
2 31299 1 3404
2 31300 1 3405
2 31301 1 3405
2 31302 1 3405
2 31303 1 3428
2 31304 1 3428
2 31305 1 3428
2 31306 1 3436
2 31307 1 3436
2 31308 1 3436
2 31309 1 3437
2 31310 1 3437
2 31311 1 3437
2 31312 1 3437
2 31313 1 3437
2 31314 1 3437
2 31315 1 3437
2 31316 1 3437
2 31317 1 3440
2 31318 1 3440
2 31319 1 3440
2 31320 1 3440
2 31321 1 3440
2 31322 1 3440
2 31323 1 3440
2 31324 1 3440
2 31325 1 3447
2 31326 1 3447
2 31327 1 3447
2 31328 1 3447
2 31329 1 3447
2 31330 1 3449
2 31331 1 3449
2 31332 1 3449
2 31333 1 3458
2 31334 1 3458
2 31335 1 3460
2 31336 1 3460
2 31337 1 3461
2 31338 1 3461
2 31339 1 3474
2 31340 1 3474
2 31341 1 3474
2 31342 1 3474
2 31343 1 3474
2 31344 1 3474
2 31345 1 3474
2 31346 1 3474
2 31347 1 3474
2 31348 1 3474
2 31349 1 3474
2 31350 1 3474
2 31351 1 3474
2 31352 1 3474
2 31353 1 3476
2 31354 1 3476
2 31355 1 3476
2 31356 1 3476
2 31357 1 3476
2 31358 1 3476
2 31359 1 3476
2 31360 1 3477
2 31361 1 3477
2 31362 1 3477
2 31363 1 3485
2 31364 1 3485
2 31365 1 3486
2 31366 1 3486
2 31367 1 3486
2 31368 1 3487
2 31369 1 3487
2 31370 1 3487
2 31371 1 3487
2 31372 1 3487
2 31373 1 3487
2 31374 1 3487
2 31375 1 3487
2 31376 1 3487
2 31377 1 3497
2 31378 1 3497
2 31379 1 3497
2 31380 1 3497
2 31381 1 3498
2 31382 1 3498
2 31383 1 3498
2 31384 1 3498
2 31385 1 3499
2 31386 1 3499
2 31387 1 3501
2 31388 1 3501
2 31389 1 3501
2 31390 1 3515
2 31391 1 3515
2 31392 1 3529
2 31393 1 3529
2 31394 1 3550
2 31395 1 3550
2 31396 1 3552
2 31397 1 3552
2 31398 1 3559
2 31399 1 3559
2 31400 1 3559
2 31401 1 3560
2 31402 1 3560
2 31403 1 3560
2 31404 1 3564
2 31405 1 3564
2 31406 1 3564
2 31407 1 3565
2 31408 1 3565
2 31409 1 3566
2 31410 1 3566
2 31411 1 3566
2 31412 1 3566
2 31413 1 3566
2 31414 1 3566
2 31415 1 3566
2 31416 1 3566
2 31417 1 3566
2 31418 1 3566
2 31419 1 3566
2 31420 1 3593
2 31421 1 3593
2 31422 1 3612
2 31423 1 3612
2 31424 1 3616
2 31425 1 3616
2 31426 1 3636
2 31427 1 3636
2 31428 1 3636
2 31429 1 3636
2 31430 1 3645
2 31431 1 3645
2 31432 1 3646
2 31433 1 3646
2 31434 1 3646
2 31435 1 3648
2 31436 1 3648
2 31437 1 3649
2 31438 1 3649
2 31439 1 3649
2 31440 1 3649
2 31441 1 3649
2 31442 1 3649
2 31443 1 3649
2 31444 1 3649
2 31445 1 3650
2 31446 1 3650
2 31447 1 3650
2 31448 1 3650
2 31449 1 3650
2 31450 1 3652
2 31451 1 3652
2 31452 1 3669
2 31453 1 3669
2 31454 1 3669
2 31455 1 3670
2 31456 1 3670
2 31457 1 3670
2 31458 1 3670
2 31459 1 3670
2 31460 1 3670
2 31461 1 3670
2 31462 1 3670
2 31463 1 3670
2 31464 1 3670
2 31465 1 3670
2 31466 1 3670
2 31467 1 3670
2 31468 1 3670
2 31469 1 3670
2 31470 1 3670
2 31471 1 3670
2 31472 1 3670
2 31473 1 3670
2 31474 1 3670
2 31475 1 3670
2 31476 1 3671
2 31477 1 3671
2 31478 1 3671
2 31479 1 3672
2 31480 1 3672
2 31481 1 3672
2 31482 1 3672
2 31483 1 3673
2 31484 1 3673
2 31485 1 3685
2 31486 1 3685
2 31487 1 3685
2 31488 1 3692
2 31489 1 3692
2 31490 1 3692
2 31491 1 3692
2 31492 1 3693
2 31493 1 3693
2 31494 1 3693
2 31495 1 3693
2 31496 1 3693
2 31497 1 3693
2 31498 1 3693
2 31499 1 3693
2 31500 1 3693
2 31501 1 3693
2 31502 1 3693
2 31503 1 3694
2 31504 1 3694
2 31505 1 3694
2 31506 1 3708
2 31507 1 3708
2 31508 1 3708
2 31509 1 3730
2 31510 1 3730
2 31511 1 3730
2 31512 1 3730
2 31513 1 3731
2 31514 1 3731
2 31515 1 3731
2 31516 1 3731
2 31517 1 3731
2 31518 1 3731
2 31519 1 3735
2 31520 1 3735
2 31521 1 3743
2 31522 1 3743
2 31523 1 3744
2 31524 1 3744
2 31525 1 3746
2 31526 1 3746
2 31527 1 3746
2 31528 1 3746
2 31529 1 3746
2 31530 1 3746
2 31531 1 3747
2 31532 1 3747
2 31533 1 3747
2 31534 1 3747
2 31535 1 3747
2 31536 1 3747
2 31537 1 3748
2 31538 1 3748
2 31539 1 3748
2 31540 1 3748
2 31541 1 3748
2 31542 1 3757
2 31543 1 3757
2 31544 1 3757
2 31545 1 3760
2 31546 1 3760
2 31547 1 3760
2 31548 1 3760
2 31549 1 3772
2 31550 1 3772
2 31551 1 3785
2 31552 1 3785
2 31553 1 3785
2 31554 1 3785
2 31555 1 3786
2 31556 1 3786
2 31557 1 3800
2 31558 1 3800
2 31559 1 3805
2 31560 1 3805
2 31561 1 3807
2 31562 1 3807
2 31563 1 3816
2 31564 1 3816
2 31565 1 3816
2 31566 1 3830
2 31567 1 3830
2 31568 1 3830
2 31569 1 3830
2 31570 1 3830
2 31571 1 3830
2 31572 1 3838
2 31573 1 3838
2 31574 1 3839
2 31575 1 3839
2 31576 1 3842
2 31577 1 3842
2 31578 1 3843
2 31579 1 3843
2 31580 1 3843
2 31581 1 3845
2 31582 1 3845
2 31583 1 3845
2 31584 1 3845
2 31585 1 3845
2 31586 1 3846
2 31587 1 3846
2 31588 1 3847
2 31589 1 3847
2 31590 1 3847
2 31591 1 3848
2 31592 1 3848
2 31593 1 3849
2 31594 1 3849
2 31595 1 3861
2 31596 1 3861
2 31597 1 3866
2 31598 1 3866
2 31599 1 3873
2 31600 1 3873
2 31601 1 3873
2 31602 1 3873
2 31603 1 3873
2 31604 1 3873
2 31605 1 3873
2 31606 1 3874
2 31607 1 3874
2 31608 1 3874
2 31609 1 3874
2 31610 1 3874
2 31611 1 3874
2 31612 1 3874
2 31613 1 3874
2 31614 1 3875
2 31615 1 3875
2 31616 1 3881
2 31617 1 3881
2 31618 1 3881
2 31619 1 3881
2 31620 1 3881
2 31621 1 3885
2 31622 1 3885
2 31623 1 3886
2 31624 1 3886
2 31625 1 3892
2 31626 1 3892
2 31627 1 3892
2 31628 1 3892
2 31629 1 3892
2 31630 1 3892
2 31631 1 3892
2 31632 1 3892
2 31633 1 3892
2 31634 1 3892
2 31635 1 3892
2 31636 1 3893
2 31637 1 3893
2 31638 1 3893
2 31639 1 3893
2 31640 1 3894
2 31641 1 3894
2 31642 1 3894
2 31643 1 3894
2 31644 1 3894
2 31645 1 3894
2 31646 1 3895
2 31647 1 3895
2 31648 1 3895
2 31649 1 3895
2 31650 1 3915
2 31651 1 3915
2 31652 1 3915
2 31653 1 3915
2 31654 1 3915
2 31655 1 3915
2 31656 1 3915
2 31657 1 3916
2 31658 1 3916
2 31659 1 3917
2 31660 1 3917
2 31661 1 3923
2 31662 1 3923
2 31663 1 3941
2 31664 1 3941
2 31665 1 3941
2 31666 1 3942
2 31667 1 3942
2 31668 1 3961
2 31669 1 3961
2 31670 1 3964
2 31671 1 3964
2 31672 1 3964
2 31673 1 3965
2 31674 1 3965
2 31675 1 3966
2 31676 1 3966
2 31677 1 3966
2 31678 1 3966
2 31679 1 3966
2 31680 1 3973
2 31681 1 3973
2 31682 1 3974
2 31683 1 3974
2 31684 1 3974
2 31685 1 3974
2 31686 1 3975
2 31687 1 3975
2 31688 1 3975
2 31689 1 3975
2 31690 1 3976
2 31691 1 3976
2 31692 1 3977
2 31693 1 3977
2 31694 1 3977
2 31695 1 3986
2 31696 1 3986
2 31697 1 3987
2 31698 1 3987
2 31699 1 3988
2 31700 1 3988
2 31701 1 3988
2 31702 1 3990
2 31703 1 3990
2 31704 1 3990
2 31705 1 3990
2 31706 1 3990
2 31707 1 3991
2 31708 1 3991
2 31709 1 3992
2 31710 1 3992
2 31711 1 3992
2 31712 1 3993
2 31713 1 3993
2 31714 1 3993
2 31715 1 3993
2 31716 1 3993
2 31717 1 4012
2 31718 1 4012
2 31719 1 4013
2 31720 1 4013
2 31721 1 4015
2 31722 1 4015
2 31723 1 4035
2 31724 1 4035
2 31725 1 4036
2 31726 1 4036
2 31727 1 4036
2 31728 1 4036
2 31729 1 4036
2 31730 1 4036
2 31731 1 4037
2 31732 1 4037
2 31733 1 4037
2 31734 1 4041
2 31735 1 4041
2 31736 1 4052
2 31737 1 4052
2 31738 1 4077
2 31739 1 4077
2 31740 1 4077
2 31741 1 4077
2 31742 1 4077
2 31743 1 4077
2 31744 1 4077
2 31745 1 4078
2 31746 1 4078
2 31747 1 4099
2 31748 1 4099
2 31749 1 4099
2 31750 1 4099
2 31751 1 4100
2 31752 1 4100
2 31753 1 4100
2 31754 1 4100
2 31755 1 4112
2 31756 1 4112
2 31757 1 4113
2 31758 1 4113
2 31759 1 4114
2 31760 1 4114
2 31761 1 4114
2 31762 1 4116
2 31763 1 4116
2 31764 1 4137
2 31765 1 4137
2 31766 1 4139
2 31767 1 4139
2 31768 1 4141
2 31769 1 4141
2 31770 1 4151
2 31771 1 4151
2 31772 1 4151
2 31773 1 4160
2 31774 1 4160
2 31775 1 4160
2 31776 1 4160
2 31777 1 4161
2 31778 1 4161
2 31779 1 4172
2 31780 1 4172
2 31781 1 4172
2 31782 1 4172
2 31783 1 4172
2 31784 1 4174
2 31785 1 4174
2 31786 1 4176
2 31787 1 4176
2 31788 1 4177
2 31789 1 4177
2 31790 1 4177
2 31791 1 4177
2 31792 1 4177
2 31793 1 4183
2 31794 1 4183
2 31795 1 4189
2 31796 1 4189
2 31797 1 4193
2 31798 1 4193
2 31799 1 4193
2 31800 1 4203
2 31801 1 4203
2 31802 1 4203
2 31803 1 4204
2 31804 1 4204
2 31805 1 4205
2 31806 1 4205
2 31807 1 4214
2 31808 1 4214
2 31809 1 4214
2 31810 1 4222
2 31811 1 4222
2 31812 1 4222
2 31813 1 4222
2 31814 1 4222
2 31815 1 4230
2 31816 1 4230
2 31817 1 4233
2 31818 1 4233
2 31819 1 4233
2 31820 1 4233
2 31821 1 4233
2 31822 1 4233
2 31823 1 4233
2 31824 1 4233
2 31825 1 4233
2 31826 1 4233
2 31827 1 4233
2 31828 1 4233
2 31829 1 4233
2 31830 1 4233
2 31831 1 4233
2 31832 1 4233
2 31833 1 4233
2 31834 1 4233
2 31835 1 4234
2 31836 1 4234
2 31837 1 4235
2 31838 1 4235
2 31839 1 4235
2 31840 1 4235
2 31841 1 4235
2 31842 1 4236
2 31843 1 4236
2 31844 1 4236
2 31845 1 4237
2 31846 1 4237
2 31847 1 4243
2 31848 1 4243
2 31849 1 4243
2 31850 1 4243
2 31851 1 4244
2 31852 1 4244
2 31853 1 4246
2 31854 1 4246
2 31855 1 4246
2 31856 1 4246
2 31857 1 4246
2 31858 1 4247
2 31859 1 4247
2 31860 1 4264
2 31861 1 4264
2 31862 1 4264
2 31863 1 4264
2 31864 1 4265
2 31865 1 4265
2 31866 1 4266
2 31867 1 4266
2 31868 1 4269
2 31869 1 4269
2 31870 1 4269
2 31871 1 4269
2 31872 1 4269
2 31873 1 4276
2 31874 1 4276
2 31875 1 4277
2 31876 1 4277
2 31877 1 4277
2 31878 1 4277
2 31879 1 4286
2 31880 1 4286
2 31881 1 4286
2 31882 1 4286
2 31883 1 4286
2 31884 1 4287
2 31885 1 4287
2 31886 1 4288
2 31887 1 4288
2 31888 1 4296
2 31889 1 4296
2 31890 1 4296
2 31891 1 4296
2 31892 1 4297
2 31893 1 4297
2 31894 1 4297
2 31895 1 4299
2 31896 1 4299
2 31897 1 4299
2 31898 1 4300
2 31899 1 4300
2 31900 1 4300
2 31901 1 4300
2 31902 1 4300
2 31903 1 4300
2 31904 1 4301
2 31905 1 4301
2 31906 1 4301
2 31907 1 4305
2 31908 1 4305
2 31909 1 4316
2 31910 1 4316
2 31911 1 4316
2 31912 1 4316
2 31913 1 4316
2 31914 1 4316
2 31915 1 4316
2 31916 1 4316
2 31917 1 4316
2 31918 1 4316
2 31919 1 4316
2 31920 1 4316
2 31921 1 4329
2 31922 1 4329
2 31923 1 4329
2 31924 1 4334
2 31925 1 4334
2 31926 1 4334
2 31927 1 4334
2 31928 1 4334
2 31929 1 4343
2 31930 1 4343
2 31931 1 4343
2 31932 1 4343
2 31933 1 4376
2 31934 1 4376
2 31935 1 4376
2 31936 1 4376
2 31937 1 4378
2 31938 1 4378
2 31939 1 4378
2 31940 1 4378
2 31941 1 4378
2 31942 1 4378
2 31943 1 4379
2 31944 1 4379
2 31945 1 4382
2 31946 1 4382
2 31947 1 4382
2 31948 1 4382
2 31949 1 4384
2 31950 1 4384
2 31951 1 4384
2 31952 1 4399
2 31953 1 4399
2 31954 1 4400
2 31955 1 4400
2 31956 1 4400
2 31957 1 4401
2 31958 1 4401
2 31959 1 4401
2 31960 1 4401
2 31961 1 4401
2 31962 1 4402
2 31963 1 4402
2 31964 1 4402
2 31965 1 4410
2 31966 1 4410
2 31967 1 4410
2 31968 1 4410
2 31969 1 4418
2 31970 1 4418
2 31971 1 4418
2 31972 1 4418
2 31973 1 4418
2 31974 1 4418
2 31975 1 4419
2 31976 1 4419
2 31977 1 4419
2 31978 1 4439
2 31979 1 4439
2 31980 1 4441
2 31981 1 4441
2 31982 1 4446
2 31983 1 4446
2 31984 1 4448
2 31985 1 4448
2 31986 1 4448
2 31987 1 4448
2 31988 1 4462
2 31989 1 4462
2 31990 1 4477
2 31991 1 4477
2 31992 1 4484
2 31993 1 4484
2 31994 1 4492
2 31995 1 4492
2 31996 1 4492
2 31997 1 4492
2 31998 1 4492
2 31999 1 4497
2 32000 1 4497
2 32001 1 4523
2 32002 1 4523
2 32003 1 4523
2 32004 1 4532
2 32005 1 4532
2 32006 1 4539
2 32007 1 4539
2 32008 1 4540
2 32009 1 4540
2 32010 1 4542
2 32011 1 4542
2 32012 1 4556
2 32013 1 4556
2 32014 1 4563
2 32015 1 4563
2 32016 1 4563
2 32017 1 4563
2 32018 1 4564
2 32019 1 4564
2 32020 1 4571
2 32021 1 4571
2 32022 1 4571
2 32023 1 4571
2 32024 1 4579
2 32025 1 4579
2 32026 1 4580
2 32027 1 4580
2 32028 1 4580
2 32029 1 4580
2 32030 1 4589
2 32031 1 4589
2 32032 1 4605
2 32033 1 4605
2 32034 1 4633
2 32035 1 4633
2 32036 1 4633
2 32037 1 4633
2 32038 1 4642
2 32039 1 4642
2 32040 1 4642
2 32041 1 4644
2 32042 1 4644
2 32043 1 4644
2 32044 1 4644
2 32045 1 4644
2 32046 1 4644
2 32047 1 4644
2 32048 1 4644
2 32049 1 4644
2 32050 1 4649
2 32051 1 4649
2 32052 1 4649
2 32053 1 4649
2 32054 1 4649
2 32055 1 4649
2 32056 1 4649
2 32057 1 4649
2 32058 1 4650
2 32059 1 4650
2 32060 1 4650
2 32061 1 4651
2 32062 1 4651
2 32063 1 4651
2 32064 1 4659
2 32065 1 4659
2 32066 1 4659
2 32067 1 4663
2 32068 1 4663
2 32069 1 4666
2 32070 1 4666
2 32071 1 4667
2 32072 1 4667
2 32073 1 4668
2 32074 1 4668
2 32075 1 4668
2 32076 1 4669
2 32077 1 4669
2 32078 1 4689
2 32079 1 4689
2 32080 1 4690
2 32081 1 4690
2 32082 1 4690
2 32083 1 4693
2 32084 1 4693
2 32085 1 4693
2 32086 1 4693
2 32087 1 4693
2 32088 1 4693
2 32089 1 4693
2 32090 1 4693
2 32091 1 4693
2 32092 1 4693
2 32093 1 4693
2 32094 1 4693
2 32095 1 4693
2 32096 1 4693
2 32097 1 4694
2 32098 1 4694
2 32099 1 4694
2 32100 1 4694
2 32101 1 4703
2 32102 1 4703
2 32103 1 4732
2 32104 1 4732
2 32105 1 4743
2 32106 1 4743
2 32107 1 4751
2 32108 1 4751
2 32109 1 4752
2 32110 1 4752
2 32111 1 4752
2 32112 1 4753
2 32113 1 4753
2 32114 1 4753
2 32115 1 4764
2 32116 1 4764
2 32117 1 4765
2 32118 1 4765
2 32119 1 4773
2 32120 1 4773
2 32121 1 4774
2 32122 1 4774
2 32123 1 4774
2 32124 1 4782
2 32125 1 4782
2 32126 1 4782
2 32127 1 4782
2 32128 1 4782
2 32129 1 4782
2 32130 1 4795
2 32131 1 4795
2 32132 1 4798
2 32133 1 4798
2 32134 1 4798
2 32135 1 4798
2 32136 1 4798
2 32137 1 4806
2 32138 1 4806
2 32139 1 4811
2 32140 1 4811
2 32141 1 4811
2 32142 1 4812
2 32143 1 4812
2 32144 1 4813
2 32145 1 4813
2 32146 1 4821
2 32147 1 4821
2 32148 1 4822
2 32149 1 4822
2 32150 1 4823
2 32151 1 4823
2 32152 1 4823
2 32153 1 4834
2 32154 1 4834
2 32155 1 4834
2 32156 1 4834
2 32157 1 4834
2 32158 1 4834
2 32159 1 4834
2 32160 1 4835
2 32161 1 4835
2 32162 1 4846
2 32163 1 4846
2 32164 1 4846
2 32165 1 4846
2 32166 1 4847
2 32167 1 4847
2 32168 1 4847
2 32169 1 4848
2 32170 1 4848
2 32171 1 4865
2 32172 1 4865
2 32173 1 4865
2 32174 1 4865
2 32175 1 4865
2 32176 1 4865
2 32177 1 4866
2 32178 1 4866
2 32179 1 4866
2 32180 1 4866
2 32181 1 4869
2 32182 1 4869
2 32183 1 4869
2 32184 1 4879
2 32185 1 4879
2 32186 1 4880
2 32187 1 4880
2 32188 1 4880
2 32189 1 4880
2 32190 1 4880
2 32191 1 4880
2 32192 1 4881
2 32193 1 4881
2 32194 1 4881
2 32195 1 4881
2 32196 1 4882
2 32197 1 4882
2 32198 1 4882
2 32199 1 4906
2 32200 1 4906
2 32201 1 4906
2 32202 1 4918
2 32203 1 4918
2 32204 1 4919
2 32205 1 4919
2 32206 1 4919
2 32207 1 4932
2 32208 1 4932
2 32209 1 4932
2 32210 1 4932
2 32211 1 4932
2 32212 1 4932
2 32213 1 4932
2 32214 1 4932
2 32215 1 4932
2 32216 1 4932
2 32217 1 4932
2 32218 1 4932
2 32219 1 4933
2 32220 1 4933
2 32221 1 4933
2 32222 1 4936
2 32223 1 4936
2 32224 1 4940
2 32225 1 4940
2 32226 1 4941
2 32227 1 4941
2 32228 1 4941
2 32229 1 4951
2 32230 1 4951
2 32231 1 4963
2 32232 1 4963
2 32233 1 4966
2 32234 1 4966
2 32235 1 4966
2 32236 1 4969
2 32237 1 4969
2 32238 1 4980
2 32239 1 4980
2 32240 1 4980
2 32241 1 4981
2 32242 1 4981
2 32243 1 4981
2 32244 1 4981
2 32245 1 4981
2 32246 1 4981
2 32247 1 4981
2 32248 1 4985
2 32249 1 4985
2 32250 1 4986
2 32251 1 4986
2 32252 1 5008
2 32253 1 5008
2 32254 1 5008
2 32255 1 5009
2 32256 1 5009
2 32257 1 5020
2 32258 1 5020
2 32259 1 5020
2 32260 1 5020
2 32261 1 5031
2 32262 1 5031
2 32263 1 5050
2 32264 1 5050
2 32265 1 5050
2 32266 1 5050
2 32267 1 5050
2 32268 1 5050
2 32269 1 5051
2 32270 1 5051
2 32271 1 5052
2 32272 1 5052
2 32273 1 5052
2 32274 1 5052
2 32275 1 5052
2 32276 1 5053
2 32277 1 5053
2 32278 1 5060
2 32279 1 5060
2 32280 1 5060
2 32281 1 5076
2 32282 1 5076
2 32283 1 5077
2 32284 1 5077
2 32285 1 5077
2 32286 1 5078
2 32287 1 5078
2 32288 1 5078
2 32289 1 5078
2 32290 1 5084
2 32291 1 5084
2 32292 1 5084
2 32293 1 5084
2 32294 1 5084
2 32295 1 5084
2 32296 1 5092
2 32297 1 5092
2 32298 1 5094
2 32299 1 5094
2 32300 1 5108
2 32301 1 5108
2 32302 1 5139
2 32303 1 5139
2 32304 1 5141
2 32305 1 5141
2 32306 1 5141
2 32307 1 5141
2 32308 1 5141
2 32309 1 5141
2 32310 1 5141
2 32311 1 5141
2 32312 1 5141
2 32313 1 5141
2 32314 1 5141
2 32315 1 5141
2 32316 1 5142
2 32317 1 5142
2 32318 1 5142
2 32319 1 5164
2 32320 1 5164
2 32321 1 5164
2 32322 1 5164
2 32323 1 5164
2 32324 1 5164
2 32325 1 5164
2 32326 1 5164
2 32327 1 5164
2 32328 1 5164
2 32329 1 5164
2 32330 1 5164
2 32331 1 5164
2 32332 1 5164
2 32333 1 5164
2 32334 1 5164
2 32335 1 5165
2 32336 1 5165
2 32337 1 5168
2 32338 1 5168
2 32339 1 5168
2 32340 1 5168
2 32341 1 5168
2 32342 1 5168
2 32343 1 5168
2 32344 1 5168
2 32345 1 5168
2 32346 1 5168
2 32347 1 5169
2 32348 1 5169
2 32349 1 5169
2 32350 1 5178
2 32351 1 5178
2 32352 1 5178
2 32353 1 5179
2 32354 1 5179
2 32355 1 5179
2 32356 1 5179
2 32357 1 5180
2 32358 1 5180
2 32359 1 5180
2 32360 1 5188
2 32361 1 5188
2 32362 1 5188
2 32363 1 5188
2 32364 1 5188
2 32365 1 5188
2 32366 1 5205
2 32367 1 5205
2 32368 1 5205
2 32369 1 5205
2 32370 1 5205
2 32371 1 5205
2 32372 1 5206
2 32373 1 5206
2 32374 1 5209
2 32375 1 5209
2 32376 1 5210
2 32377 1 5210
2 32378 1 5225
2 32379 1 5225
2 32380 1 5227
2 32381 1 5227
2 32382 1 5227
2 32383 1 5227
2 32384 1 5231
2 32385 1 5231
2 32386 1 5237
2 32387 1 5237
2 32388 1 5237
2 32389 1 5238
2 32390 1 5238
2 32391 1 5238
2 32392 1 5238
2 32393 1 5239
2 32394 1 5239
2 32395 1 5240
2 32396 1 5240
2 32397 1 5240
2 32398 1 5240
2 32399 1 5240
2 32400 1 5249
2 32401 1 5249
2 32402 1 5249
2 32403 1 5252
2 32404 1 5252
2 32405 1 5252
2 32406 1 5256
2 32407 1 5256
2 32408 1 5259
2 32409 1 5259
2 32410 1 5259
2 32411 1 5294
2 32412 1 5294
2 32413 1 5295
2 32414 1 5295
2 32415 1 5298
2 32416 1 5298
2 32417 1 5306
2 32418 1 5306
2 32419 1 5306
2 32420 1 5310
2 32421 1 5310
2 32422 1 5322
2 32423 1 5322
2 32424 1 5337
2 32425 1 5337
2 32426 1 5349
2 32427 1 5349
2 32428 1 5349
2 32429 1 5349
2 32430 1 5364
2 32431 1 5364
2 32432 1 5364
2 32433 1 5364
2 32434 1 5365
2 32435 1 5365
2 32436 1 5367
2 32437 1 5367
2 32438 1 5367
2 32439 1 5367
2 32440 1 5370
2 32441 1 5370
2 32442 1 5370
2 32443 1 5370
2 32444 1 5372
2 32445 1 5372
2 32446 1 5375
2 32447 1 5375
2 32448 1 5375
2 32449 1 5375
2 32450 1 5375
2 32451 1 5375
2 32452 1 5381
2 32453 1 5381
2 32454 1 5409
2 32455 1 5409
2 32456 1 5409
2 32457 1 5409
2 32458 1 5409
2 32459 1 5409
2 32460 1 5410
2 32461 1 5410
2 32462 1 5445
2 32463 1 5445
2 32464 1 5495
2 32465 1 5495
2 32466 1 5495
2 32467 1 5526
2 32468 1 5526
2 32469 1 5526
2 32470 1 5526
2 32471 1 5537
2 32472 1 5537
2 32473 1 5537
2 32474 1 5538
2 32475 1 5538
2 32476 1 5538
2 32477 1 5538
2 32478 1 5538
2 32479 1 5538
2 32480 1 5538
2 32481 1 5538
2 32482 1 5538
2 32483 1 5538
2 32484 1 5538
2 32485 1 5538
2 32486 1 5538
2 32487 1 5538
2 32488 1 5538
2 32489 1 5538
2 32490 1 5538
2 32491 1 5538
2 32492 1 5538
2 32493 1 5538
2 32494 1 5538
2 32495 1 5539
2 32496 1 5539
2 32497 1 5546
2 32498 1 5546
2 32499 1 5546
2 32500 1 5546
2 32501 1 5546
2 32502 1 5546
2 32503 1 5546
2 32504 1 5546
2 32505 1 5546
2 32506 1 5546
2 32507 1 5546
2 32508 1 5546
2 32509 1 5546
2 32510 1 5546
2 32511 1 5546
2 32512 1 5546
2 32513 1 5547
2 32514 1 5547
2 32515 1 5547
2 32516 1 5550
2 32517 1 5550
2 32518 1 5551
2 32519 1 5551
2 32520 1 5551
2 32521 1 5554
2 32522 1 5554
2 32523 1 5554
2 32524 1 5554
2 32525 1 5554
2 32526 1 5554
2 32527 1 5554
2 32528 1 5554
2 32529 1 5554
2 32530 1 5554
2 32531 1 5559
2 32532 1 5559
2 32533 1 5566
2 32534 1 5566
2 32535 1 5566
2 32536 1 5566
2 32537 1 5566
2 32538 1 5567
2 32539 1 5567
2 32540 1 5568
2 32541 1 5568
2 32542 1 5571
2 32543 1 5571
2 32544 1 5571
2 32545 1 5573
2 32546 1 5573
2 32547 1 5574
2 32548 1 5574
2 32549 1 5574
2 32550 1 5575
2 32551 1 5575
2 32552 1 5575
2 32553 1 5578
2 32554 1 5578
2 32555 1 5578
2 32556 1 5583
2 32557 1 5583
2 32558 1 5583
2 32559 1 5584
2 32560 1 5584
2 32561 1 5585
2 32562 1 5585
2 32563 1 5587
2 32564 1 5587
2 32565 1 5593
2 32566 1 5593
2 32567 1 5594
2 32568 1 5594
2 32569 1 5606
2 32570 1 5606
2 32571 1 5607
2 32572 1 5607
2 32573 1 5609
2 32574 1 5609
2 32575 1 5609
2 32576 1 5609
2 32577 1 5609
2 32578 1 5609
2 32579 1 5609
2 32580 1 5609
2 32581 1 5609
2 32582 1 5609
2 32583 1 5609
2 32584 1 5609
2 32585 1 5609
2 32586 1 5609
2 32587 1 5609
2 32588 1 5609
2 32589 1 5609
2 32590 1 5609
2 32591 1 5610
2 32592 1 5610
2 32593 1 5611
2 32594 1 5611
2 32595 1 5618
2 32596 1 5618
2 32597 1 5618
2 32598 1 5618
2 32599 1 5618
2 32600 1 5618
2 32601 1 5619
2 32602 1 5619
2 32603 1 5619
2 32604 1 5642
2 32605 1 5642
2 32606 1 5642
2 32607 1 5642
2 32608 1 5642
2 32609 1 5642
2 32610 1 5642
2 32611 1 5642
2 32612 1 5642
2 32613 1 5644
2 32614 1 5644
2 32615 1 5645
2 32616 1 5645
2 32617 1 5645
2 32618 1 5645
2 32619 1 5645
2 32620 1 5645
2 32621 1 5645
2 32622 1 5645
2 32623 1 5645
2 32624 1 5646
2 32625 1 5646
2 32626 1 5646
2 32627 1 5647
2 32628 1 5647
2 32629 1 5647
2 32630 1 5647
2 32631 1 5647
2 32632 1 5647
2 32633 1 5647
2 32634 1 5647
2 32635 1 5647
2 32636 1 5647
2 32637 1 5647
2 32638 1 5648
2 32639 1 5648
2 32640 1 5654
2 32641 1 5654
2 32642 1 5654
2 32643 1 5654
2 32644 1 5654
2 32645 1 5654
2 32646 1 5654
2 32647 1 5661
2 32648 1 5661
2 32649 1 5664
2 32650 1 5664
2 32651 1 5673
2 32652 1 5673
2 32653 1 5673
2 32654 1 5682
2 32655 1 5682
2 32656 1 5692
2 32657 1 5692
2 32658 1 5741
2 32659 1 5741
2 32660 1 5741
2 32661 1 5741
2 32662 1 5752
2 32663 1 5752
2 32664 1 5760
2 32665 1 5760
2 32666 1 5763
2 32667 1 5763
2 32668 1 5763
2 32669 1 5767
2 32670 1 5767
2 32671 1 5767
2 32672 1 5767
2 32673 1 5767
2 32674 1 5767
2 32675 1 5767
2 32676 1 5767
2 32677 1 5767
2 32678 1 5772
2 32679 1 5772
2 32680 1 5775
2 32681 1 5775
2 32682 1 5775
2 32683 1 5776
2 32684 1 5776
2 32685 1 5779
2 32686 1 5779
2 32687 1 5782
2 32688 1 5782
2 32689 1 5782
2 32690 1 5783
2 32691 1 5783
2 32692 1 5787
2 32693 1 5787
2 32694 1 5787
2 32695 1 5787
2 32696 1 5791
2 32697 1 5791
2 32698 1 5791
2 32699 1 5791
2 32700 1 5792
2 32701 1 5792
2 32702 1 5792
2 32703 1 5792
2 32704 1 5793
2 32705 1 5793
2 32706 1 5794
2 32707 1 5794
2 32708 1 5797
2 32709 1 5797
2 32710 1 5797
2 32711 1 5813
2 32712 1 5813
2 32713 1 5813
2 32714 1 5813
2 32715 1 5815
2 32716 1 5815
2 32717 1 5816
2 32718 1 5816
2 32719 1 5817
2 32720 1 5817
2 32721 1 5818
2 32722 1 5818
2 32723 1 5818
2 32724 1 5818
2 32725 1 5818
2 32726 1 5818
2 32727 1 5818
2 32728 1 5818
2 32729 1 5818
2 32730 1 5818
2 32731 1 5818
2 32732 1 5818
2 32733 1 5818
2 32734 1 5818
2 32735 1 5818
2 32736 1 5818
2 32737 1 5818
2 32738 1 5818
2 32739 1 5818
2 32740 1 5826
2 32741 1 5826
2 32742 1 5837
2 32743 1 5837
2 32744 1 5837
2 32745 1 5846
2 32746 1 5846
2 32747 1 5849
2 32748 1 5849
2 32749 1 5851
2 32750 1 5851
2 32751 1 5852
2 32752 1 5852
2 32753 1 5852
2 32754 1 5852
2 32755 1 5852
2 32756 1 5854
2 32757 1 5854
2 32758 1 5855
2 32759 1 5855
2 32760 1 5857
2 32761 1 5857
2 32762 1 5858
2 32763 1 5858
2 32764 1 5858
2 32765 1 5860
2 32766 1 5860
2 32767 1 5860
2 32768 1 5863
2 32769 1 5863
2 32770 1 5863
2 32771 1 5863
2 32772 1 5878
2 32773 1 5878
2 32774 1 5893
2 32775 1 5893
2 32776 1 5893
2 32777 1 5893
2 32778 1 5893
2 32779 1 5893
2 32780 1 5893
2 32781 1 5893
2 32782 1 5893
2 32783 1 5893
2 32784 1 5893
2 32785 1 5897
2 32786 1 5897
2 32787 1 5897
2 32788 1 5897
2 32789 1 5898
2 32790 1 5898
2 32791 1 5914
2 32792 1 5914
2 32793 1 5914
2 32794 1 5931
2 32795 1 5931
2 32796 1 5932
2 32797 1 5932
2 32798 1 5939
2 32799 1 5939
2 32800 1 5960
2 32801 1 5960
2 32802 1 5963
2 32803 1 5963
2 32804 1 5963
2 32805 1 5963
2 32806 1 5977
2 32807 1 5977
2 32808 1 5978
2 32809 1 5978
2 32810 1 5978
2 32811 1 5978
2 32812 1 5986
2 32813 1 5986
2 32814 1 6000
2 32815 1 6000
2 32816 1 6013
2 32817 1 6013
2 32818 1 6022
2 32819 1 6022
2 32820 1 6025
2 32821 1 6025
2 32822 1 6026
2 32823 1 6026
2 32824 1 6026
2 32825 1 6027
2 32826 1 6027
2 32827 1 6035
2 32828 1 6035
2 32829 1 6035
2 32830 1 6035
2 32831 1 6035
2 32832 1 6035
2 32833 1 6035
2 32834 1 6036
2 32835 1 6036
2 32836 1 6036
2 32837 1 6037
2 32838 1 6037
2 32839 1 6044
2 32840 1 6044
2 32841 1 6045
2 32842 1 6045
2 32843 1 6046
2 32844 1 6046
2 32845 1 6046
2 32846 1 6046
2 32847 1 6046
2 32848 1 6046
2 32849 1 6046
2 32850 1 6047
2 32851 1 6047
2 32852 1 6051
2 32853 1 6051
2 32854 1 6057
2 32855 1 6057
2 32856 1 6057
2 32857 1 6074
2 32858 1 6074
2 32859 1 6082
2 32860 1 6082
2 32861 1 6117
2 32862 1 6117
2 32863 1 6134
2 32864 1 6134
2 32865 1 6134
2 32866 1 6135
2 32867 1 6135
2 32868 1 6147
2 32869 1 6147
2 32870 1 6147
2 32871 1 6147
2 32872 1 6147
2 32873 1 6148
2 32874 1 6148
2 32875 1 6158
2 32876 1 6158
2 32877 1 6159
2 32878 1 6159
2 32879 1 6162
2 32880 1 6162
2 32881 1 6166
2 32882 1 6166
2 32883 1 6167
2 32884 1 6167
2 32885 1 6176
2 32886 1 6176
2 32887 1 6176
2 32888 1 6185
2 32889 1 6185
2 32890 1 6203
2 32891 1 6203
2 32892 1 6232
2 32893 1 6232
2 32894 1 6234
2 32895 1 6234
2 32896 1 6234
2 32897 1 6236
2 32898 1 6236
2 32899 1 6245
2 32900 1 6245
2 32901 1 6245
2 32902 1 6245
2 32903 1 6254
2 32904 1 6254
2 32905 1 6254
2 32906 1 6262
2 32907 1 6262
2 32908 1 6262
2 32909 1 6262
2 32910 1 6262
2 32911 1 6262
2 32912 1 6262
2 32913 1 6262
2 32914 1 6262
2 32915 1 6262
2 32916 1 6262
2 32917 1 6262
2 32918 1 6264
2 32919 1 6264
2 32920 1 6269
2 32921 1 6269
2 32922 1 6269
2 32923 1 6269
2 32924 1 6269
2 32925 1 6269
2 32926 1 6269
2 32927 1 6269
2 32928 1 6269
2 32929 1 6269
2 32930 1 6270
2 32931 1 6270
2 32932 1 6270
2 32933 1 6270
2 32934 1 6270
2 32935 1 6270
2 32936 1 6271
2 32937 1 6271
2 32938 1 6279
2 32939 1 6279
2 32940 1 6280
2 32941 1 6280
2 32942 1 6280
2 32943 1 6281
2 32944 1 6281
2 32945 1 6281
2 32946 1 6288
2 32947 1 6288
2 32948 1 6295
2 32949 1 6295
2 32950 1 6295
2 32951 1 6295
2 32952 1 6295
2 32953 1 6295
2 32954 1 6295
2 32955 1 6295
2 32956 1 6295
2 32957 1 6295
2 32958 1 6295
2 32959 1 6295
2 32960 1 6298
2 32961 1 6298
2 32962 1 6298
2 32963 1 6298
2 32964 1 6298
2 32965 1 6298
2 32966 1 6298
2 32967 1 6298
2 32968 1 6298
2 32969 1 6298
2 32970 1 6298
2 32971 1 6298
2 32972 1 6298
2 32973 1 6298
2 32974 1 6298
2 32975 1 6298
2 32976 1 6298
2 32977 1 6298
2 32978 1 6298
2 32979 1 6298
2 32980 1 6298
2 32981 1 6298
2 32982 1 6298
2 32983 1 6298
2 32984 1 6298
2 32985 1 6298
2 32986 1 6298
2 32987 1 6298
2 32988 1 6298
2 32989 1 6298
2 32990 1 6298
2 32991 1 6298
2 32992 1 6298
2 32993 1 6298
2 32994 1 6298
2 32995 1 6298
2 32996 1 6298
2 32997 1 6299
2 32998 1 6299
2 32999 1 6299
2 33000 1 6300
2 33001 1 6300
2 33002 1 6301
2 33003 1 6301
2 33004 1 6305
2 33005 1 6305
2 33006 1 6305
2 33007 1 6305
2 33008 1 6305
2 33009 1 6305
2 33010 1 6305
2 33011 1 6305
2 33012 1 6305
2 33013 1 6306
2 33014 1 6306
2 33015 1 6315
2 33016 1 6315
2 33017 1 6316
2 33018 1 6316
2 33019 1 6316
2 33020 1 6316
2 33021 1 6317
2 33022 1 6317
2 33023 1 6333
2 33024 1 6333
2 33025 1 6333
2 33026 1 6333
2 33027 1 6333
2 33028 1 6333
2 33029 1 6333
2 33030 1 6333
2 33031 1 6333
2 33032 1 6333
2 33033 1 6333
2 33034 1 6334
2 33035 1 6334
2 33036 1 6334
2 33037 1 6334
2 33038 1 6334
2 33039 1 6334
2 33040 1 6334
2 33041 1 6334
2 33042 1 6334
2 33043 1 6336
2 33044 1 6336
2 33045 1 6336
2 33046 1 6340
2 33047 1 6340
2 33048 1 6340
2 33049 1 6342
2 33050 1 6342
2 33051 1 6345
2 33052 1 6345
2 33053 1 6345
2 33054 1 6345
2 33055 1 6345
2 33056 1 6347
2 33057 1 6347
2 33058 1 6351
2 33059 1 6351
2 33060 1 6368
2 33061 1 6368
2 33062 1 6373
2 33063 1 6373
2 33064 1 6375
2 33065 1 6375
2 33066 1 6375
2 33067 1 6375
2 33068 1 6375
2 33069 1 6386
2 33070 1 6386
2 33071 1 6387
2 33072 1 6387
2 33073 1 6387
2 33074 1 6392
2 33075 1 6392
2 33076 1 6394
2 33077 1 6394
2 33078 1 6394
2 33079 1 6399
2 33080 1 6399
2 33081 1 6415
2 33082 1 6415
2 33083 1 6416
2 33084 1 6416
2 33085 1 6433
2 33086 1 6433
2 33087 1 6435
2 33088 1 6435
2 33089 1 6435
2 33090 1 6437
2 33091 1 6437
2 33092 1 6437
2 33093 1 6437
2 33094 1 6454
2 33095 1 6454
2 33096 1 6455
2 33097 1 6455
2 33098 1 6459
2 33099 1 6459
2 33100 1 6462
2 33101 1 6462
2 33102 1 6468
2 33103 1 6468
2 33104 1 6473
2 33105 1 6473
2 33106 1 6473
2 33107 1 6473
2 33108 1 6473
2 33109 1 6474
2 33110 1 6474
2 33111 1 6484
2 33112 1 6484
2 33113 1 6535
2 33114 1 6535
2 33115 1 6545
2 33116 1 6545
2 33117 1 6546
2 33118 1 6546
2 33119 1 6561
2 33120 1 6561
2 33121 1 6570
2 33122 1 6570
2 33123 1 6570
2 33124 1 6570
2 33125 1 6570
2 33126 1 6572
2 33127 1 6572
2 33128 1 6584
2 33129 1 6584
2 33130 1 6584
2 33131 1 6599
2 33132 1 6599
2 33133 1 6600
2 33134 1 6600
2 33135 1 6600
2 33136 1 6608
2 33137 1 6608
2 33138 1 6629
2 33139 1 6629
2 33140 1 6630
2 33141 1 6630
2 33142 1 6630
2 33143 1 6630
2 33144 1 6642
2 33145 1 6642
2 33146 1 6642
2 33147 1 6655
2 33148 1 6655
2 33149 1 6655
2 33150 1 6655
2 33151 1 6655
2 33152 1 6656
2 33153 1 6656
2 33154 1 6656
2 33155 1 6656
2 33156 1 6656
2 33157 1 6656
2 33158 1 6659
2 33159 1 6659
2 33160 1 6671
2 33161 1 6671
2 33162 1 6671
2 33163 1 6671
2 33164 1 6671
2 33165 1 6675
2 33166 1 6675
2 33167 1 6675
2 33168 1 6675
2 33169 1 6675
2 33170 1 6676
2 33171 1 6676
2 33172 1 6676
2 33173 1 6676
2 33174 1 6676
2 33175 1 6676
2 33176 1 6676
2 33177 1 6676
2 33178 1 6676
2 33179 1 6690
2 33180 1 6690
2 33181 1 6690
2 33182 1 6691
2 33183 1 6691
2 33184 1 6691
2 33185 1 6692
2 33186 1 6692
2 33187 1 6698
2 33188 1 6698
2 33189 1 6706
2 33190 1 6706
2 33191 1 6709
2 33192 1 6709
2 33193 1 6712
2 33194 1 6712
2 33195 1 6745
2 33196 1 6745
2 33197 1 6748
2 33198 1 6748
2 33199 1 6748
2 33200 1 6752
2 33201 1 6752
2 33202 1 6752
2 33203 1 6752
2 33204 1 6752
2 33205 1 6752
2 33206 1 6752
2 33207 1 6756
2 33208 1 6756
2 33209 1 6775
2 33210 1 6775
2 33211 1 6775
2 33212 1 6776
2 33213 1 6776
2 33214 1 6778
2 33215 1 6778
2 33216 1 6778
2 33217 1 6778
2 33218 1 6778
2 33219 1 6780
2 33220 1 6780
2 33221 1 6783
2 33222 1 6783
2 33223 1 6783
2 33224 1 6785
2 33225 1 6785
2 33226 1 6788
2 33227 1 6788
2 33228 1 6788
2 33229 1 6788
2 33230 1 6788
2 33231 1 6788
2 33232 1 6788
2 33233 1 6788
2 33234 1 6790
2 33235 1 6790
2 33236 1 6792
2 33237 1 6792
2 33238 1 6792
2 33239 1 6792
2 33240 1 6806
2 33241 1 6806
2 33242 1 6809
2 33243 1 6809
2 33244 1 6809
2 33245 1 6809
2 33246 1 6809
2 33247 1 6809
2 33248 1 6809
2 33249 1 6809
2 33250 1 6814
2 33251 1 6814
2 33252 1 6814
2 33253 1 6814
2 33254 1 6814
2 33255 1 6814
2 33256 1 6814
2 33257 1 6815
2 33258 1 6815
2 33259 1 6836
2 33260 1 6836
2 33261 1 6836
2 33262 1 6836
2 33263 1 6836
2 33264 1 6837
2 33265 1 6837
2 33266 1 6837
2 33267 1 6848
2 33268 1 6848
2 33269 1 6848
2 33270 1 6851
2 33271 1 6851
2 33272 1 6859
2 33273 1 6859
2 33274 1 6859
2 33275 1 6859
2 33276 1 6861
2 33277 1 6861
2 33278 1 6867
2 33279 1 6867
2 33280 1 6867
2 33281 1 6867
2 33282 1 6867
2 33283 1 6894
2 33284 1 6894
2 33285 1 6894
2 33286 1 6894
2 33287 1 6894
2 33288 1 6894
2 33289 1 6894
2 33290 1 6894
2 33291 1 6894
2 33292 1 6894
2 33293 1 6894
2 33294 1 6894
2 33295 1 6894
2 33296 1 6894
2 33297 1 6894
2 33298 1 6894
2 33299 1 6894
2 33300 1 6894
2 33301 1 6894
2 33302 1 6894
2 33303 1 6894
2 33304 1 6894
2 33305 1 6894
2 33306 1 6894
2 33307 1 6894
2 33308 1 6894
2 33309 1 6894
2 33310 1 6894
2 33311 1 6894
2 33312 1 6894
2 33313 1 6894
2 33314 1 6894
2 33315 1 6894
2 33316 1 6894
2 33317 1 6894
2 33318 1 6894
2 33319 1 6894
2 33320 1 6894
2 33321 1 6894
2 33322 1 6894
2 33323 1 6894
2 33324 1 6894
2 33325 1 6894
2 33326 1 6894
2 33327 1 6894
2 33328 1 6894
2 33329 1 6894
2 33330 1 6894
2 33331 1 6894
2 33332 1 6894
2 33333 1 6894
2 33334 1 6894
2 33335 1 6894
2 33336 1 6898
2 33337 1 6898
2 33338 1 6898
2 33339 1 6898
2 33340 1 6898
2 33341 1 6898
2 33342 1 6898
2 33343 1 6898
2 33344 1 6898
2 33345 1 6898
2 33346 1 6898
2 33347 1 6898
2 33348 1 6898
2 33349 1 6898
2 33350 1 6898
2 33351 1 6898
2 33352 1 6898
2 33353 1 6898
2 33354 1 6898
2 33355 1 6898
2 33356 1 6898
2 33357 1 6898
2 33358 1 6898
2 33359 1 6898
2 33360 1 6898
2 33361 1 6898
2 33362 1 6898
2 33363 1 6898
2 33364 1 6898
2 33365 1 6898
2 33366 1 6898
2 33367 1 6898
2 33368 1 6898
2 33369 1 6898
2 33370 1 6898
2 33371 1 6898
2 33372 1 6898
2 33373 1 6898
2 33374 1 6898
2 33375 1 6898
2 33376 1 6898
2 33377 1 6898
2 33378 1 6898
2 33379 1 6898
2 33380 1 6898
2 33381 1 6898
2 33382 1 6898
2 33383 1 6898
2 33384 1 6898
2 33385 1 6898
2 33386 1 6898
2 33387 1 6898
2 33388 1 6898
2 33389 1 6898
2 33390 1 6898
2 33391 1 6900
2 33392 1 6900
2 33393 1 6900
2 33394 1 6900
2 33395 1 6900
2 33396 1 6901
2 33397 1 6901
2 33398 1 6907
2 33399 1 6907
2 33400 1 6907
2 33401 1 6907
2 33402 1 6907
2 33403 1 6907
2 33404 1 6907
2 33405 1 6907
2 33406 1 6908
2 33407 1 6908
2 33408 1 6908
2 33409 1 6908
2 33410 1 6908
2 33411 1 6908
2 33412 1 6908
2 33413 1 6908
2 33414 1 6908
2 33415 1 6908
2 33416 1 6908
2 33417 1 6908
2 33418 1 6909
2 33419 1 6909
2 33420 1 6910
2 33421 1 6910
2 33422 1 6912
2 33423 1 6912
2 33424 1 6912
2 33425 1 6912
2 33426 1 6912
2 33427 1 6912
2 33428 1 6912
2 33429 1 6913
2 33430 1 6913
2 33431 1 6913
2 33432 1 6913
2 33433 1 6913
2 33434 1 6913
2 33435 1 6914
2 33436 1 6914
2 33437 1 6915
2 33438 1 6915
2 33439 1 6915
2 33440 1 6928
2 33441 1 6928
2 33442 1 6928
2 33443 1 6928
2 33444 1 6928
2 33445 1 6929
2 33446 1 6929
2 33447 1 6929
2 33448 1 6929
2 33449 1 6930
2 33450 1 6930
2 33451 1 6930
2 33452 1 6930
2 33453 1 6930
2 33454 1 6930
2 33455 1 6930
2 33456 1 6930
2 33457 1 6930
2 33458 1 6930
2 33459 1 6930
2 33460 1 6931
2 33461 1 6931
2 33462 1 6939
2 33463 1 6939
2 33464 1 6939
2 33465 1 6939
2 33466 1 6939
2 33467 1 6940
2 33468 1 6940
2 33469 1 6941
2 33470 1 6941
2 33471 1 6941
2 33472 1 6956
2 33473 1 6956
2 33474 1 6956
2 33475 1 6956
2 33476 1 6956
2 33477 1 6956
2 33478 1 6956
2 33479 1 6956
2 33480 1 6957
2 33481 1 6957
2 33482 1 6958
2 33483 1 6958
2 33484 1 6981
2 33485 1 6981
2 33486 1 6981
2 33487 1 6981
2 33488 1 6989
2 33489 1 6989
2 33490 1 6989
2 33491 1 6989
2 33492 1 6990
2 33493 1 6990
2 33494 1 7001
2 33495 1 7001
2 33496 1 7001
2 33497 1 7002
2 33498 1 7002
2 33499 1 7003
2 33500 1 7003
2 33501 1 7003
2 33502 1 7003
2 33503 1 7003
2 33504 1 7003
2 33505 1 7003
2 33506 1 7004
2 33507 1 7004
2 33508 1 7004
2 33509 1 7004
2 33510 1 7004
2 33511 1 7004
2 33512 1 7005
2 33513 1 7005
2 33514 1 7005
2 33515 1 7005
2 33516 1 7005
2 33517 1 7007
2 33518 1 7007
2 33519 1 7007
2 33520 1 7010
2 33521 1 7010
2 33522 1 7010
2 33523 1 7010
2 33524 1 7010
2 33525 1 7010
2 33526 1 7010
2 33527 1 7010
2 33528 1 7010
2 33529 1 7010
2 33530 1 7010
2 33531 1 7010
2 33532 1 7010
2 33533 1 7010
2 33534 1 7010
2 33535 1 7010
2 33536 1 7010
2 33537 1 7011
2 33538 1 7011
2 33539 1 7012
2 33540 1 7012
2 33541 1 7013
2 33542 1 7013
2 33543 1 7014
2 33544 1 7014
2 33545 1 7016
2 33546 1 7016
2 33547 1 7016
2 33548 1 7016
2 33549 1 7060
2 33550 1 7060
2 33551 1 7060
2 33552 1 7067
2 33553 1 7067
2 33554 1 7067
2 33555 1 7068
2 33556 1 7068
2 33557 1 7068
2 33558 1 7069
2 33559 1 7069
2 33560 1 7073
2 33561 1 7073
2 33562 1 7073
2 33563 1 7073
2 33564 1 7073
2 33565 1 7073
2 33566 1 7073
2 33567 1 7073
2 33568 1 7073
2 33569 1 7073
2 33570 1 7073
2 33571 1 7073
2 33572 1 7073
2 33573 1 7073
2 33574 1 7074
2 33575 1 7074
2 33576 1 7076
2 33577 1 7076
2 33578 1 7081
2 33579 1 7081
2 33580 1 7094
2 33581 1 7094
2 33582 1 7094
2 33583 1 7094
2 33584 1 7094
2 33585 1 7095
2 33586 1 7095
2 33587 1 7095
2 33588 1 7096
2 33589 1 7096
2 33590 1 7098
2 33591 1 7098
2 33592 1 7098
2 33593 1 7098
2 33594 1 7098
2 33595 1 7100
2 33596 1 7100
2 33597 1 7100
2 33598 1 7100
2 33599 1 7100
2 33600 1 7100
2 33601 1 7100
2 33602 1 7100
2 33603 1 7100
2 33604 1 7110
2 33605 1 7110
2 33606 1 7110
2 33607 1 7111
2 33608 1 7111
2 33609 1 7113
2 33610 1 7113
2 33611 1 7113
2 33612 1 7114
2 33613 1 7114
2 33614 1 7115
2 33615 1 7115
2 33616 1 7115
2 33617 1 7115
2 33618 1 7115
2 33619 1 7116
2 33620 1 7116
2 33621 1 7116
2 33622 1 7116
2 33623 1 7116
2 33624 1 7116
2 33625 1 7116
2 33626 1 7116
2 33627 1 7116
2 33628 1 7116
2 33629 1 7116
2 33630 1 7116
2 33631 1 7117
2 33632 1 7117
2 33633 1 7117
2 33634 1 7118
2 33635 1 7118
2 33636 1 7121
2 33637 1 7121
2 33638 1 7121
2 33639 1 7121
2 33640 1 7121
2 33641 1 7129
2 33642 1 7129
2 33643 1 7130
2 33644 1 7130
2 33645 1 7130
2 33646 1 7136
2 33647 1 7136
2 33648 1 7147
2 33649 1 7147
2 33650 1 7147
2 33651 1 7147
2 33652 1 7147
2 33653 1 7147
2 33654 1 7148
2 33655 1 7148
2 33656 1 7148
2 33657 1 7148
2 33658 1 7148
2 33659 1 7148
2 33660 1 7148
2 33661 1 7148
2 33662 1 7148
2 33663 1 7148
2 33664 1 7158
2 33665 1 7158
2 33666 1 7158
2 33667 1 7169
2 33668 1 7169
2 33669 1 7169
2 33670 1 7171
2 33671 1 7171
2 33672 1 7171
2 33673 1 7172
2 33674 1 7172
2 33675 1 7174
2 33676 1 7174
2 33677 1 7174
2 33678 1 7174
2 33679 1 7174
2 33680 1 7175
2 33681 1 7175
2 33682 1 7184
2 33683 1 7184
2 33684 1 7184
2 33685 1 7184
2 33686 1 7185
2 33687 1 7185
2 33688 1 7185
2 33689 1 7185
2 33690 1 7188
2 33691 1 7188
2 33692 1 7188
2 33693 1 7188
2 33694 1 7188
2 33695 1 7188
2 33696 1 7189
2 33697 1 7189
2 33698 1 7189
2 33699 1 7189
2 33700 1 7189
2 33701 1 7197
2 33702 1 7197
2 33703 1 7197
2 33704 1 7197
2 33705 1 7207
2 33706 1 7207
2 33707 1 7215
2 33708 1 7215
2 33709 1 7215
2 33710 1 7215
2 33711 1 7215
2 33712 1 7215
2 33713 1 7216
2 33714 1 7216
2 33715 1 7216
2 33716 1 7223
2 33717 1 7223
2 33718 1 7223
2 33719 1 7223
2 33720 1 7223
2 33721 1 7231
2 33722 1 7231
2 33723 1 7233
2 33724 1 7233
2 33725 1 7233
2 33726 1 7233
2 33727 1 7233
2 33728 1 7233
2 33729 1 7233
2 33730 1 7233
2 33731 1 7236
2 33732 1 7236
2 33733 1 7236
2 33734 1 7236
2 33735 1 7236
2 33736 1 7236
2 33737 1 7236
2 33738 1 7236
2 33739 1 7236
2 33740 1 7236
2 33741 1 7236
2 33742 1 7236
2 33743 1 7236
2 33744 1 7237
2 33745 1 7237
2 33746 1 7237
2 33747 1 7237
2 33748 1 7237
2 33749 1 7237
2 33750 1 7237
2 33751 1 7238
2 33752 1 7238
2 33753 1 7251
2 33754 1 7251
2 33755 1 7259
2 33756 1 7259
2 33757 1 7260
2 33758 1 7260
2 33759 1 7261
2 33760 1 7261
2 33761 1 7261
2 33762 1 7261
2 33763 1 7274
2 33764 1 7274
2 33765 1 7283
2 33766 1 7283
2 33767 1 7284
2 33768 1 7284
2 33769 1 7284
2 33770 1 7284
2 33771 1 7285
2 33772 1 7285
2 33773 1 7285
2 33774 1 7297
2 33775 1 7297
2 33776 1 7315
2 33777 1 7315
2 33778 1 7315
2 33779 1 7316
2 33780 1 7316
2 33781 1 7318
2 33782 1 7318
2 33783 1 7323
2 33784 1 7323
2 33785 1 7323
2 33786 1 7324
2 33787 1 7324
2 33788 1 7324
2 33789 1 7324
2 33790 1 7324
2 33791 1 7324
2 33792 1 7324
2 33793 1 7324
2 33794 1 7325
2 33795 1 7325
2 33796 1 7325
2 33797 1 7326
2 33798 1 7326
2 33799 1 7326
2 33800 1 7326
2 33801 1 7326
2 33802 1 7326
2 33803 1 7326
2 33804 1 7326
2 33805 1 7326
2 33806 1 7326
2 33807 1 7326
2 33808 1 7327
2 33809 1 7327
2 33810 1 7330
2 33811 1 7330
2 33812 1 7330
2 33813 1 7330
2 33814 1 7330
2 33815 1 7330
2 33816 1 7333
2 33817 1 7333
2 33818 1 7340
2 33819 1 7340
2 33820 1 7357
2 33821 1 7357
2 33822 1 7357
2 33823 1 7357
2 33824 1 7357
2 33825 1 7357
2 33826 1 7360
2 33827 1 7360
2 33828 1 7360
2 33829 1 7360
2 33830 1 7360
2 33831 1 7360
2 33832 1 7367
2 33833 1 7367
2 33834 1 7367
2 33835 1 7368
2 33836 1 7368
2 33837 1 7376
2 33838 1 7376
2 33839 1 7377
2 33840 1 7377
2 33841 1 7396
2 33842 1 7396
2 33843 1 7405
2 33844 1 7405
2 33845 1 7405
2 33846 1 7406
2 33847 1 7406
2 33848 1 7407
2 33849 1 7407
2 33850 1 7407
2 33851 1 7410
2 33852 1 7410
2 33853 1 7410
2 33854 1 7410
2 33855 1 7410
2 33856 1 7410
2 33857 1 7410
2 33858 1 7410
2 33859 1 7410
2 33860 1 7410
2 33861 1 7410
2 33862 1 7413
2 33863 1 7413
2 33864 1 7416
2 33865 1 7416
2 33866 1 7416
2 33867 1 7416
2 33868 1 7416
2 33869 1 7420
2 33870 1 7420
2 33871 1 7420
2 33872 1 7420
2 33873 1 7420
2 33874 1 7420
2 33875 1 7420
2 33876 1 7420
2 33877 1 7420
2 33878 1 7421
2 33879 1 7421
2 33880 1 7421
2 33881 1 7421
2 33882 1 7421
2 33883 1 7422
2 33884 1 7422
2 33885 1 7422
2 33886 1 7432
2 33887 1 7432
2 33888 1 7433
2 33889 1 7433
2 33890 1 7433
2 33891 1 7438
2 33892 1 7438
2 33893 1 7451
2 33894 1 7451
2 33895 1 7457
2 33896 1 7457
2 33897 1 7457
2 33898 1 7458
2 33899 1 7458
2 33900 1 7458
2 33901 1 7458
2 33902 1 7460
2 33903 1 7460
2 33904 1 7460
2 33905 1 7460
2 33906 1 7464
2 33907 1 7464
2 33908 1 7464
2 33909 1 7464
2 33910 1 7465
2 33911 1 7465
2 33912 1 7465
2 33913 1 7472
2 33914 1 7472
2 33915 1 7472
2 33916 1 7472
2 33917 1 7472
2 33918 1 7472
2 33919 1 7472
2 33920 1 7472
2 33921 1 7472
2 33922 1 7472
2 33923 1 7472
2 33924 1 7472
2 33925 1 7472
2 33926 1 7472
2 33927 1 7472
2 33928 1 7472
2 33929 1 7472
2 33930 1 7472
2 33931 1 7472
2 33932 1 7472
2 33933 1 7472
2 33934 1 7482
2 33935 1 7482
2 33936 1 7494
2 33937 1 7494
2 33938 1 7494
2 33939 1 7494
2 33940 1 7494
2 33941 1 7494
2 33942 1 7494
2 33943 1 7508
2 33944 1 7508
2 33945 1 7508
2 33946 1 7510
2 33947 1 7510
2 33948 1 7510
2 33949 1 7510
2 33950 1 7510
2 33951 1 7510
2 33952 1 7510
2 33953 1 7510
2 33954 1 7510
2 33955 1 7511
2 33956 1 7511
2 33957 1 7514
2 33958 1 7514
2 33959 1 7514
2 33960 1 7515
2 33961 1 7515
2 33962 1 7515
2 33963 1 7517
2 33964 1 7517
2 33965 1 7517
2 33966 1 7517
2 33967 1 7517
2 33968 1 7517
2 33969 1 7517
2 33970 1 7517
2 33971 1 7517
2 33972 1 7517
2 33973 1 7517
2 33974 1 7517
2 33975 1 7517
2 33976 1 7517
2 33977 1 7517
2 33978 1 7517
2 33979 1 7517
2 33980 1 7517
2 33981 1 7517
2 33982 1 7517
2 33983 1 7517
2 33984 1 7517
2 33985 1 7528
2 33986 1 7528
2 33987 1 7528
2 33988 1 7528
2 33989 1 7528
2 33990 1 7529
2 33991 1 7529
2 33992 1 7529
2 33993 1 7530
2 33994 1 7530
2 33995 1 7530
2 33996 1 7531
2 33997 1 7531
2 33998 1 7544
2 33999 1 7544
2 34000 1 7544
2 34001 1 7544
2 34002 1 7545
2 34003 1 7545
2 34004 1 7545
2 34005 1 7545
2 34006 1 7545
2 34007 1 7545
2 34008 1 7545
2 34009 1 7545
2 34010 1 7545
2 34011 1 7546
2 34012 1 7546
2 34013 1 7547
2 34014 1 7547
2 34015 1 7556
2 34016 1 7556
2 34017 1 7556
2 34018 1 7556
2 34019 1 7564
2 34020 1 7564
2 34021 1 7564
2 34022 1 7564
2 34023 1 7564
2 34024 1 7564
2 34025 1 7565
2 34026 1 7565
2 34027 1 7565
2 34028 1 7565
2 34029 1 7566
2 34030 1 7566
2 34031 1 7567
2 34032 1 7567
2 34033 1 7567
2 34034 1 7570
2 34035 1 7570
2 34036 1 7570
2 34037 1 7571
2 34038 1 7571
2 34039 1 7571
2 34040 1 7571
2 34041 1 7571
2 34042 1 7571
2 34043 1 7572
2 34044 1 7572
2 34045 1 7572
2 34046 1 7572
2 34047 1 7572
2 34048 1 7572
2 34049 1 7572
2 34050 1 7572
2 34051 1 7583
2 34052 1 7583
2 34053 1 7583
2 34054 1 7587
2 34055 1 7587
2 34056 1 7587
2 34057 1 7587
2 34058 1 7588
2 34059 1 7588
2 34060 1 7603
2 34061 1 7603
2 34062 1 7603
2 34063 1 7603
2 34064 1 7603
2 34065 1 7603
2 34066 1 7603
2 34067 1 7605
2 34068 1 7605
2 34069 1 7605
2 34070 1 7605
2 34071 1 7605
2 34072 1 7605
2 34073 1 7605
2 34074 1 7605
2 34075 1 7606
2 34076 1 7606
2 34077 1 7606
2 34078 1 7608
2 34079 1 7608
2 34080 1 7608
2 34081 1 7608
2 34082 1 7608
2 34083 1 7608
2 34084 1 7608
2 34085 1 7608
2 34086 1 7610
2 34087 1 7610
2 34088 1 7615
2 34089 1 7615
2 34090 1 7659
2 34091 1 7659
2 34092 1 7659
2 34093 1 7659
2 34094 1 7659
2 34095 1 7660
2 34096 1 7660
2 34097 1 7661
2 34098 1 7661
2 34099 1 7663
2 34100 1 7663
2 34101 1 7663
2 34102 1 7663
2 34103 1 7663
2 34104 1 7663
2 34105 1 7663
2 34106 1 7663
2 34107 1 7663
2 34108 1 7663
2 34109 1 7663
2 34110 1 7663
2 34111 1 7663
2 34112 1 7663
2 34113 1 7663
2 34114 1 7663
2 34115 1 7663
2 34116 1 7663
2 34117 1 7664
2 34118 1 7664
2 34119 1 7664
2 34120 1 7664
2 34121 1 7665
2 34122 1 7665
2 34123 1 7665
2 34124 1 7665
2 34125 1 7665
2 34126 1 7665
2 34127 1 7666
2 34128 1 7666
2 34129 1 7668
2 34130 1 7668
2 34131 1 7669
2 34132 1 7669
2 34133 1 7671
2 34134 1 7671
2 34135 1 7674
2 34136 1 7674
2 34137 1 7674
2 34138 1 7674
2 34139 1 7674
2 34140 1 7674
2 34141 1 7674
2 34142 1 7674
2 34143 1 7674
2 34144 1 7674
2 34145 1 7674
2 34146 1 7674
2 34147 1 7686
2 34148 1 7686
2 34149 1 7689
2 34150 1 7689
2 34151 1 7689
2 34152 1 7694
2 34153 1 7694
2 34154 1 7694
2 34155 1 7694
2 34156 1 7695
2 34157 1 7695
2 34158 1 7708
2 34159 1 7708
2 34160 1 7710
2 34161 1 7710
2 34162 1 7710
2 34163 1 7710
2 34164 1 7723
2 34165 1 7723
2 34166 1 7723
2 34167 1 7731
2 34168 1 7731
2 34169 1 7731
2 34170 1 7731
2 34171 1 7731
2 34172 1 7734
2 34173 1 7734
2 34174 1 7742
2 34175 1 7742
2 34176 1 7742
2 34177 1 7742
2 34178 1 7742
2 34179 1 7742
2 34180 1 7742
2 34181 1 7742
2 34182 1 7742
2 34183 1 7742
2 34184 1 7742
2 34185 1 7743
2 34186 1 7743
2 34187 1 7743
2 34188 1 7743
2 34189 1 7743
2 34190 1 7743
2 34191 1 7743
2 34192 1 7743
2 34193 1 7743
2 34194 1 7744
2 34195 1 7744
2 34196 1 7744
2 34197 1 7744
2 34198 1 7744
2 34199 1 7752
2 34200 1 7752
2 34201 1 7752
2 34202 1 7752
2 34203 1 7753
2 34204 1 7753
2 34205 1 7753
2 34206 1 7753
2 34207 1 7754
2 34208 1 7754
2 34209 1 7754
2 34210 1 7754
2 34211 1 7755
2 34212 1 7755
2 34213 1 7755
2 34214 1 7755
2 34215 1 7755
2 34216 1 7758
2 34217 1 7758
2 34218 1 7758
2 34219 1 7758
2 34220 1 7759
2 34221 1 7759
2 34222 1 7759
2 34223 1 7759
2 34224 1 7760
2 34225 1 7760
2 34226 1 7769
2 34227 1 7769
2 34228 1 7769
2 34229 1 7770
2 34230 1 7770
2 34231 1 7770
2 34232 1 7770
2 34233 1 7779
2 34234 1 7779
2 34235 1 7779
2 34236 1 7779
2 34237 1 7779
2 34238 1 7780
2 34239 1 7780
2 34240 1 7783
2 34241 1 7783
2 34242 1 7783
2 34243 1 7795
2 34244 1 7795
2 34245 1 7795
2 34246 1 7801
2 34247 1 7801
2 34248 1 7828
2 34249 1 7828
2 34250 1 7829
2 34251 1 7829
2 34252 1 7837
2 34253 1 7837
2 34254 1 7837
2 34255 1 7839
2 34256 1 7839
2 34257 1 7839
2 34258 1 7840
2 34259 1 7840
2 34260 1 7843
2 34261 1 7843
2 34262 1 7849
2 34263 1 7849
2 34264 1 7849
2 34265 1 7850
2 34266 1 7850
2 34267 1 7850
2 34268 1 7850
2 34269 1 7850
2 34270 1 7850
2 34271 1 7850
2 34272 1 7850
2 34273 1 7851
2 34274 1 7851
2 34275 1 7866
2 34276 1 7866
2 34277 1 7866
2 34278 1 7866
2 34279 1 7868
2 34280 1 7868
2 34281 1 7868
2 34282 1 7868
2 34283 1 7868
2 34284 1 7868
2 34285 1 7869
2 34286 1 7869
2 34287 1 7869
2 34288 1 7871
2 34289 1 7871
2 34290 1 7871
2 34291 1 7871
2 34292 1 7871
2 34293 1 7871
2 34294 1 7871
2 34295 1 7871
2 34296 1 7871
2 34297 1 7871
2 34298 1 7871
2 34299 1 7871
2 34300 1 7871
2 34301 1 7871
2 34302 1 7871
2 34303 1 7871
2 34304 1 7871
2 34305 1 7871
2 34306 1 7871
2 34307 1 7871
2 34308 1 7871
2 34309 1 7871
2 34310 1 7872
2 34311 1 7872
2 34312 1 7872
2 34313 1 7872
2 34314 1 7872
2 34315 1 7872
2 34316 1 7872
2 34317 1 7872
2 34318 1 7873
2 34319 1 7873
2 34320 1 7873
2 34321 1 7874
2 34322 1 7874
2 34323 1 7877
2 34324 1 7877
2 34325 1 7881
2 34326 1 7881
2 34327 1 7885
2 34328 1 7885
2 34329 1 7885
2 34330 1 7886
2 34331 1 7886
2 34332 1 7887
2 34333 1 7887
2 34334 1 7894
2 34335 1 7894
2 34336 1 7894
2 34337 1 7898
2 34338 1 7898
2 34339 1 7898
2 34340 1 7898
2 34341 1 7898
2 34342 1 7898
2 34343 1 7898
2 34344 1 7904
2 34345 1 7904
2 34346 1 7912
2 34347 1 7912
2 34348 1 7912
2 34349 1 7912
2 34350 1 7912
2 34351 1 7912
2 34352 1 7912
2 34353 1 7912
2 34354 1 7912
2 34355 1 7912
2 34356 1 7912
2 34357 1 7915
2 34358 1 7915
2 34359 1 7915
2 34360 1 7915
2 34361 1 7915
2 34362 1 7915
2 34363 1 7915
2 34364 1 7915
2 34365 1 7915
2 34366 1 7915
2 34367 1 7915
2 34368 1 7915
2 34369 1 7915
2 34370 1 7915
2 34371 1 7915
2 34372 1 7915
2 34373 1 7919
2 34374 1 7919
2 34375 1 7919
2 34376 1 7919
2 34377 1 7919
2 34378 1 7919
2 34379 1 7920
2 34380 1 7920
2 34381 1 7920
2 34382 1 7920
2 34383 1 7920
2 34384 1 7920
2 34385 1 7920
2 34386 1 7920
2 34387 1 7921
2 34388 1 7921
2 34389 1 7921
2 34390 1 7921
2 34391 1 7922
2 34392 1 7922
2 34393 1 7922
2 34394 1 7932
2 34395 1 7932
2 34396 1 7932
2 34397 1 7936
2 34398 1 7936
2 34399 1 7936
2 34400 1 7939
2 34401 1 7939
2 34402 1 7939
2 34403 1 7939
2 34404 1 7939
2 34405 1 7939
2 34406 1 7939
2 34407 1 7939
2 34408 1 7939
2 34409 1 7939
2 34410 1 7939
2 34411 1 7939
2 34412 1 7939
2 34413 1 7939
2 34414 1 7939
2 34415 1 7939
2 34416 1 7939
2 34417 1 7939
2 34418 1 7939
2 34419 1 7939
2 34420 1 7939
2 34421 1 7939
2 34422 1 7939
2 34423 1 7939
2 34424 1 7940
2 34425 1 7940
2 34426 1 7953
2 34427 1 7953
2 34428 1 7953
2 34429 1 7953
2 34430 1 7953
2 34431 1 7953
2 34432 1 7953
2 34433 1 7953
2 34434 1 7954
2 34435 1 7954
2 34436 1 7955
2 34437 1 7955
2 34438 1 7963
2 34439 1 7963
2 34440 1 7963
2 34441 1 7963
2 34442 1 7963
2 34443 1 7963
2 34444 1 7963
2 34445 1 7963
2 34446 1 7972
2 34447 1 7972
2 34448 1 7973
2 34449 1 7973
2 34450 1 7974
2 34451 1 7974
2 34452 1 7974
2 34453 1 7974
2 34454 1 7975
2 34455 1 7975
2 34456 1 7981
2 34457 1 7981
2 34458 1 7997
2 34459 1 7997
2 34460 1 7997
2 34461 1 7997
2 34462 1 7997
2 34463 1 7997
2 34464 1 7997
2 34465 1 8010
2 34466 1 8010
2 34467 1 8011
2 34468 1 8011
2 34469 1 8011
2 34470 1 8015
2 34471 1 8015
2 34472 1 8015
2 34473 1 8015
2 34474 1 8017
2 34475 1 8017
2 34476 1 8036
2 34477 1 8036
2 34478 1 8036
2 34479 1 8036
2 34480 1 8036
2 34481 1 8036
2 34482 1 8037
2 34483 1 8037
2 34484 1 8037
2 34485 1 8037
2 34486 1 8037
2 34487 1 8037
2 34488 1 8037
2 34489 1 8037
2 34490 1 8037
2 34491 1 8038
2 34492 1 8038
2 34493 1 8039
2 34494 1 8039
2 34495 1 8069
2 34496 1 8069
2 34497 1 8070
2 34498 1 8070
2 34499 1 8070
2 34500 1 8070
2 34501 1 8083
2 34502 1 8083
2 34503 1 8093
2 34504 1 8093
2 34505 1 8093
2 34506 1 8093
2 34507 1 8093
2 34508 1 8093
2 34509 1 8093
2 34510 1 8093
2 34511 1 8093
2 34512 1 8094
2 34513 1 8094
2 34514 1 8095
2 34515 1 8095
2 34516 1 8095
2 34517 1 8096
2 34518 1 8096
2 34519 1 8097
2 34520 1 8097
2 34521 1 8104
2 34522 1 8104
2 34523 1 8114
2 34524 1 8114
2 34525 1 8115
2 34526 1 8115
2 34527 1 8116
2 34528 1 8116
2 34529 1 8116
2 34530 1 8141
2 34531 1 8141
2 34532 1 8141
2 34533 1 8148
2 34534 1 8148
2 34535 1 8149
2 34536 1 8149
2 34537 1 8149
2 34538 1 8149
2 34539 1 8149
2 34540 1 8149
2 34541 1 8149
2 34542 1 8150
2 34543 1 8150
2 34544 1 8150
2 34545 1 8165
2 34546 1 8165
2 34547 1 8168
2 34548 1 8168
2 34549 1 8169
2 34550 1 8169
2 34551 1 8176
2 34552 1 8176
2 34553 1 8177
2 34554 1 8177
2 34555 1 8177
2 34556 1 8177
2 34557 1 8181
2 34558 1 8181
2 34559 1 8181
2 34560 1 8181
2 34561 1 8181
2 34562 1 8181
2 34563 1 8181
2 34564 1 8181
2 34565 1 8204
2 34566 1 8204
2 34567 1 8223
2 34568 1 8223
2 34569 1 8223
2 34570 1 8225
2 34571 1 8225
2 34572 1 8228
2 34573 1 8228
2 34574 1 8231
2 34575 1 8231
2 34576 1 8252
2 34577 1 8252
2 34578 1 8253
2 34579 1 8253
2 34580 1 8253
2 34581 1 8253
2 34582 1 8253
2 34583 1 8253
2 34584 1 8253
2 34585 1 8253
2 34586 1 8253
2 34587 1 8253
2 34588 1 8253
2 34589 1 8253
2 34590 1 8253
2 34591 1 8253
2 34592 1 8253
2 34593 1 8253
2 34594 1 8257
2 34595 1 8257
2 34596 1 8257
2 34597 1 8257
2 34598 1 8259
2 34599 1 8259
2 34600 1 8259
2 34601 1 8291
2 34602 1 8291
2 34603 1 8296
2 34604 1 8296
2 34605 1 8296
2 34606 1 8302
2 34607 1 8302
2 34608 1 8314
2 34609 1 8314
2 34610 1 8317
2 34611 1 8317
2 34612 1 8331
2 34613 1 8331
2 34614 1 8340
2 34615 1 8340
2 34616 1 8341
2 34617 1 8341
2 34618 1 8360
2 34619 1 8360
2 34620 1 8376
2 34621 1 8376
2 34622 1 8387
2 34623 1 8387
2 34624 1 8421
2 34625 1 8421
2 34626 1 8434
2 34627 1 8434
2 34628 1 8434
2 34629 1 8439
2 34630 1 8439
2 34631 1 8440
2 34632 1 8440
2 34633 1 8444
2 34634 1 8444
2 34635 1 8444
2 34636 1 8449
2 34637 1 8449
2 34638 1 8449
2 34639 1 8470
2 34640 1 8470
2 34641 1 8470
2 34642 1 8471
2 34643 1 8471
2 34644 1 8494
2 34645 1 8494
2 34646 1 8495
2 34647 1 8495
2 34648 1 8495
2 34649 1 8495
2 34650 1 8505
2 34651 1 8505
2 34652 1 8506
2 34653 1 8506
2 34654 1 8514
2 34655 1 8514
2 34656 1 8529
2 34657 1 8529
2 34658 1 8554
2 34659 1 8554
2 34660 1 8554
2 34661 1 8561
2 34662 1 8561
2 34663 1 8561
2 34664 1 8561
2 34665 1 8561
2 34666 1 8561
2 34667 1 8561
2 34668 1 8572
2 34669 1 8572
2 34670 1 8572
2 34671 1 8575
2 34672 1 8575
2 34673 1 8575
2 34674 1 8579
2 34675 1 8579
2 34676 1 8593
2 34677 1 8593
2 34678 1 8594
2 34679 1 8594
2 34680 1 8596
2 34681 1 8596
2 34682 1 8602
2 34683 1 8602
2 34684 1 8634
2 34685 1 8634
2 34686 1 8634
2 34687 1 8642
2 34688 1 8642
2 34689 1 8648
2 34690 1 8648
2 34691 1 8654
2 34692 1 8654
2 34693 1 8663
2 34694 1 8663
2 34695 1 8673
2 34696 1 8673
2 34697 1 8688
2 34698 1 8688
2 34699 1 8688
2 34700 1 8688
2 34701 1 8691
2 34702 1 8691
2 34703 1 8691
2 34704 1 8701
2 34705 1 8701
2 34706 1 8702
2 34707 1 8702
2 34708 1 8702
2 34709 1 8719
2 34710 1 8719
2 34711 1 8719
2 34712 1 8728
2 34713 1 8728
2 34714 1 8728
2 34715 1 8743
2 34716 1 8743
2 34717 1 8766
2 34718 1 8766
2 34719 1 8822
2 34720 1 8822
2 34721 1 8822
2 34722 1 8822
2 34723 1 8822
2 34724 1 8822
2 34725 1 8822
2 34726 1 8822
2 34727 1 8835
2 34728 1 8835
2 34729 1 8835
2 34730 1 8836
2 34731 1 8836
2 34732 1 8836
2 34733 1 8836
2 34734 1 8836
2 34735 1 8836
2 34736 1 8847
2 34737 1 8847
2 34738 1 8855
2 34739 1 8855
2 34740 1 8857
2 34741 1 8857
2 34742 1 8879
2 34743 1 8879
2 34744 1 8879
2 34745 1 8879
2 34746 1 8888
2 34747 1 8888
2 34748 1 8898
2 34749 1 8898
2 34750 1 8917
2 34751 1 8917
2 34752 1 8917
2 34753 1 8918
2 34754 1 8918
2 34755 1 8928
2 34756 1 8928
2 34757 1 8941
2 34758 1 8941
2 34759 1 8943
2 34760 1 8943
2 34761 1 8943
2 34762 1 8943
2 34763 1 8943
2 34764 1 8943
2 34765 1 8943
2 34766 1 8950
2 34767 1 8950
2 34768 1 8958
2 34769 1 8958
2 34770 1 8958
2 34771 1 8958
2 34772 1 8959
2 34773 1 8959
2 34774 1 8959
2 34775 1 8959
2 34776 1 8972
2 34777 1 8972
2 34778 1 8975
2 34779 1 8975
2 34780 1 8975
2 34781 1 8976
2 34782 1 8976
2 34783 1 8976
2 34784 1 8977
2 34785 1 8977
2 34786 1 8984
2 34787 1 8984
2 34788 1 8984
2 34789 1 8986
2 34790 1 8986
2 34791 1 8993
2 34792 1 8993
2 34793 1 8993
2 34794 1 8993
2 34795 1 8994
2 34796 1 8994
2 34797 1 8994
2 34798 1 8995
2 34799 1 8995
2 34800 1 9012
2 34801 1 9012
2 34802 1 9012
2 34803 1 9035
2 34804 1 9035
2 34805 1 9056
2 34806 1 9056
2 34807 1 9058
2 34808 1 9058
2 34809 1 9061
2 34810 1 9061
2 34811 1 9062
2 34812 1 9062
2 34813 1 9062
2 34814 1 9063
2 34815 1 9063
2 34816 1 9101
2 34817 1 9101
2 34818 1 9101
2 34819 1 9108
2 34820 1 9108
2 34821 1 9108
2 34822 1 9108
2 34823 1 9109
2 34824 1 9109
2 34825 1 9119
2 34826 1 9119
2 34827 1 9119
2 34828 1 9119
2 34829 1 9119
2 34830 1 9119
2 34831 1 9119
2 34832 1 9120
2 34833 1 9120
2 34834 1 9124
2 34835 1 9124
2 34836 1 9132
2 34837 1 9132
2 34838 1 9134
2 34839 1 9134
2 34840 1 9135
2 34841 1 9135
2 34842 1 9139
2 34843 1 9139
2 34844 1 9146
2 34845 1 9146
2 34846 1 9146
2 34847 1 9146
2 34848 1 9146
2 34849 1 9146
2 34850 1 9146
2 34851 1 9146
2 34852 1 9146
2 34853 1 9146
2 34854 1 9146
2 34855 1 9146
2 34856 1 9146
2 34857 1 9146
2 34858 1 9146
2 34859 1 9146
2 34860 1 9146
2 34861 1 9147
2 34862 1 9147
2 34863 1 9151
2 34864 1 9151
2 34865 1 9162
2 34866 1 9162
2 34867 1 9162
2 34868 1 9162
2 34869 1 9162
2 34870 1 9164
2 34871 1 9164
2 34872 1 9168
2 34873 1 9168
2 34874 1 9168
2 34875 1 9168
2 34876 1 9174
2 34877 1 9174
2 34878 1 9191
2 34879 1 9191
2 34880 1 9191
2 34881 1 9191
2 34882 1 9205
2 34883 1 9205
2 34884 1 9221
2 34885 1 9221
2 34886 1 9236
2 34887 1 9236
2 34888 1 9245
2 34889 1 9245
2 34890 1 9256
2 34891 1 9256
2 34892 1 9256
2 34893 1 9269
2 34894 1 9269
2 34895 1 9269
2 34896 1 9269
2 34897 1 9269
2 34898 1 9280
2 34899 1 9280
2 34900 1 9281
2 34901 1 9281
2 34902 1 9281
2 34903 1 9281
2 34904 1 9281
2 34905 1 9281
2 34906 1 9281
2 34907 1 9281
2 34908 1 9281
2 34909 1 9281
2 34910 1 9292
2 34911 1 9292
2 34912 1 9292
2 34913 1 9292
2 34914 1 9315
2 34915 1 9315
2 34916 1 9315
2 34917 1 9315
2 34918 1 9320
2 34919 1 9320
2 34920 1 9329
2 34921 1 9329
2 34922 1 9333
2 34923 1 9333
2 34924 1 9333
2 34925 1 9333
2 34926 1 9333
2 34927 1 9333
2 34928 1 9333
2 34929 1 9333
2 34930 1 9333
2 34931 1 9333
2 34932 1 9333
2 34933 1 9333
2 34934 1 9333
2 34935 1 9333
2 34936 1 9333
2 34937 1 9333
2 34938 1 9333
2 34939 1 9333
2 34940 1 9333
2 34941 1 9333
2 34942 1 9333
2 34943 1 9333
2 34944 1 9333
2 34945 1 9347
2 34946 1 9347
2 34947 1 9347
2 34948 1 9347
2 34949 1 9347
2 34950 1 9347
2 34951 1 9347
2 34952 1 9354
2 34953 1 9354
2 34954 1 9354
2 34955 1 9363
2 34956 1 9363
2 34957 1 9372
2 34958 1 9372
2 34959 1 9438
2 34960 1 9438
2 34961 1 9438
2 34962 1 9438
2 34963 1 9441
2 34964 1 9441
2 34965 1 9474
2 34966 1 9474
2 34967 1 9474
2 34968 1 9478
2 34969 1 9478
2 34970 1 9485
2 34971 1 9485
2 34972 1 9485
2 34973 1 9486
2 34974 1 9486
2 34975 1 9490
2 34976 1 9490
2 34977 1 9490
2 34978 1 9491
2 34979 1 9491
2 34980 1 9518
2 34981 1 9518
2 34982 1 9518
2 34983 1 9527
2 34984 1 9527
2 34985 1 9528
2 34986 1 9528
2 34987 1 9535
2 34988 1 9535
2 34989 1 9544
2 34990 1 9544
2 34991 1 9557
2 34992 1 9557
2 34993 1 9557
2 34994 1 9558
2 34995 1 9558
2 34996 1 9558
2 34997 1 9566
2 34998 1 9566
2 34999 1 9567
2 35000 1 9567
2 35001 1 9579
2 35002 1 9579
2 35003 1 9588
2 35004 1 9588
2 35005 1 9588
2 35006 1 9588
2 35007 1 9588
2 35008 1 9589
2 35009 1 9589
2 35010 1 9589
2 35011 1 9589
2 35012 1 9589
2 35013 1 9590
2 35014 1 9590
2 35015 1 9590
2 35016 1 9591
2 35017 1 9591
2 35018 1 9597
2 35019 1 9597
2 35020 1 9604
2 35021 1 9604
2 35022 1 9607
2 35023 1 9607
2 35024 1 9607
2 35025 1 9607
2 35026 1 9607
2 35027 1 9607
2 35028 1 9628
2 35029 1 9628
2 35030 1 9628
2 35031 1 9631
2 35032 1 9631
2 35033 1 9631
2 35034 1 9631
2 35035 1 9639
2 35036 1 9639
2 35037 1 9642
2 35038 1 9642
2 35039 1 9642
2 35040 1 9642
2 35041 1 9642
2 35042 1 9643
2 35043 1 9643
2 35044 1 9707
2 35045 1 9707
2 35046 1 9710
2 35047 1 9710
2 35048 1 9711
2 35049 1 9711
2 35050 1 9711
2 35051 1 9713
2 35052 1 9713
2 35053 1 9716
2 35054 1 9716
2 35055 1 9737
2 35056 1 9737
2 35057 1 9737
2 35058 1 9746
2 35059 1 9746
2 35060 1 9746
2 35061 1 9757
2 35062 1 9757
2 35063 1 9779
2 35064 1 9779
2 35065 1 9779
2 35066 1 9779
2 35067 1 9794
2 35068 1 9794
2 35069 1 9794
2 35070 1 9794
2 35071 1 9823
2 35072 1 9823
2 35073 1 9825
2 35074 1 9825
2 35075 1 9825
2 35076 1 9825
2 35077 1 9825
2 35078 1 9825
2 35079 1 9825
2 35080 1 9825
2 35081 1 9825
2 35082 1 9825
2 35083 1 9825
2 35084 1 9853
2 35085 1 9853
2 35086 1 9853
2 35087 1 9853
2 35088 1 9853
2 35089 1 9853
2 35090 1 9866
2 35091 1 9866
2 35092 1 9868
2 35093 1 9868
2 35094 1 9868
2 35095 1 9869
2 35096 1 9869
2 35097 1 9876
2 35098 1 9876
2 35099 1 9904
2 35100 1 9904
2 35101 1 9904
2 35102 1 9907
2 35103 1 9907
2 35104 1 9907
2 35105 1 9907
2 35106 1 9907
2 35107 1 9919
2 35108 1 9919
2 35109 1 9919
2 35110 1 9919
2 35111 1 9919
2 35112 1 9919
2 35113 1 9919
2 35114 1 9920
2 35115 1 9920
2 35116 1 9921
2 35117 1 9921
2 35118 1 9930
2 35119 1 9930
2 35120 1 9932
2 35121 1 9932
2 35122 1 9932
2 35123 1 9932
2 35124 1 9933
2 35125 1 9933
2 35126 1 9941
2 35127 1 9941
2 35128 1 9944
2 35129 1 9944
2 35130 1 9944
2 35131 1 9944
2 35132 1 9945
2 35133 1 9945
2 35134 1 9945
2 35135 1 9967
2 35136 1 9967
2 35137 1 9967
2 35138 1 9967
2 35139 1 9967
2 35140 1 9967
2 35141 1 9967
2 35142 1 9968
2 35143 1 9968
2 35144 1 9968
2 35145 1 9969
2 35146 1 9969
2 35147 1 9972
2 35148 1 9972
2 35149 1 9975
2 35150 1 9975
2 35151 1 9998
2 35152 1 9998
2 35153 1 10002
2 35154 1 10002
2 35155 1 10002
2 35156 1 10002
2 35157 1 10002
2 35158 1 10015
2 35159 1 10015
2 35160 1 10020
2 35161 1 10020
2 35162 1 10045
2 35163 1 10045
2 35164 1 10045
2 35165 1 10045
2 35166 1 10047
2 35167 1 10047
2 35168 1 10068
2 35169 1 10068
2 35170 1 10070
2 35171 1 10070
2 35172 1 10103
2 35173 1 10103
2 35174 1 10110
2 35175 1 10110
2 35176 1 10117
2 35177 1 10117
2 35178 1 10118
2 35179 1 10118
2 35180 1 10125
2 35181 1 10125
2 35182 1 10127
2 35183 1 10127
2 35184 1 10141
2 35185 1 10141
2 35186 1 10142
2 35187 1 10142
2 35188 1 10151
2 35189 1 10151
2 35190 1 10152
2 35191 1 10152
2 35192 1 10152
2 35193 1 10155
2 35194 1 10155
2 35195 1 10175
2 35196 1 10175
2 35197 1 10175
2 35198 1 10192
2 35199 1 10192
2 35200 1 10193
2 35201 1 10193
2 35202 1 10197
2 35203 1 10197
2 35204 1 10200
2 35205 1 10200
2 35206 1 10219
2 35207 1 10219
2 35208 1 10239
2 35209 1 10239
2 35210 1 10239
2 35211 1 10239
2 35212 1 10239
2 35213 1 10239
2 35214 1 10240
2 35215 1 10240
2 35216 1 10240
2 35217 1 10247
2 35218 1 10247
2 35219 1 10247
2 35220 1 10247
2 35221 1 10247
2 35222 1 10247
2 35223 1 10247
2 35224 1 10247
2 35225 1 10247
2 35226 1 10249
2 35227 1 10249
2 35228 1 10265
2 35229 1 10265
2 35230 1 10265
2 35231 1 10265
2 35232 1 10265
2 35233 1 10265
2 35234 1 10339
2 35235 1 10339
2 35236 1 10339
2 35237 1 10339
2 35238 1 10364
2 35239 1 10364
2 35240 1 10369
2 35241 1 10369
2 35242 1 10374
2 35243 1 10374
2 35244 1 10374
2 35245 1 10396
2 35246 1 10396
2 35247 1 10442
2 35248 1 10442
2 35249 1 10442
2 35250 1 10444
2 35251 1 10444
2 35252 1 10444
2 35253 1 10463
2 35254 1 10463
2 35255 1 10476
2 35256 1 10476
2 35257 1 10494
2 35258 1 10494
2 35259 1 10495
2 35260 1 10495
2 35261 1 10502
2 35262 1 10502
2 35263 1 10526
2 35264 1 10526
2 35265 1 10535
2 35266 1 10535
2 35267 1 10593
2 35268 1 10593
2 35269 1 10593
2 35270 1 10600
2 35271 1 10600
2 35272 1 10600
2 35273 1 10600
2 35274 1 10626
2 35275 1 10626
2 35276 1 10675
2 35277 1 10675
2 35278 1 10675
2 35279 1 10675
2 35280 1 10710
2 35281 1 10710
2 35282 1 10712
2 35283 1 10712
2 35284 1 10733
2 35285 1 10733
2 35286 1 10743
2 35287 1 10743
2 35288 1 10751
2 35289 1 10751
2 35290 1 10763
2 35291 1 10763
2 35292 1 10763
2 35293 1 10764
2 35294 1 10764
2 35295 1 10764
2 35296 1 10812
2 35297 1 10812
2 35298 1 10820
2 35299 1 10820
2 35300 1 10820
2 35301 1 10829
2 35302 1 10829
2 35303 1 10837
2 35304 1 10837
2 35305 1 10837
2 35306 1 10855
2 35307 1 10855
2 35308 1 10864
2 35309 1 10864
2 35310 1 10887
2 35311 1 10887
2 35312 1 10887
2 35313 1 10915
2 35314 1 10915
2 35315 1 10915
2 35316 1 10916
2 35317 1 10916
2 35318 1 10918
2 35319 1 10918
2 35320 1 10918
2 35321 1 10922
2 35322 1 10922
2 35323 1 10922
2 35324 1 10922
2 35325 1 10927
2 35326 1 10927
2 35327 1 10927
2 35328 1 10927
2 35329 1 10927
2 35330 1 10927
2 35331 1 10927
2 35332 1 10927
2 35333 1 10927
2 35334 1 10928
2 35335 1 10928
2 35336 1 10938
2 35337 1 10938
2 35338 1 10945
2 35339 1 10945
2 35340 1 10945
2 35341 1 10945
2 35342 1 10948
2 35343 1 10948
2 35344 1 10949
2 35345 1 10949
2 35346 1 10960
2 35347 1 10960
2 35348 1 10960
2 35349 1 10978
2 35350 1 10978
2 35351 1 11010
2 35352 1 11010
2 35353 1 11017
2 35354 1 11017
2 35355 1 11023
2 35356 1 11023
2 35357 1 11023
2 35358 1 11030
2 35359 1 11030
2 35360 1 11031
2 35361 1 11031
2 35362 1 11056
2 35363 1 11056
2 35364 1 11056
2 35365 1 11061
2 35366 1 11061
2 35367 1 11074
2 35368 1 11074
2 35369 1 11075
2 35370 1 11075
2 35371 1 11075
2 35372 1 11075
2 35373 1 11076
2 35374 1 11076
2 35375 1 11079
2 35376 1 11079
2 35377 1 11079
2 35378 1 11080
2 35379 1 11080
2 35380 1 11080
2 35381 1 11081
2 35382 1 11081
2 35383 1 11081
2 35384 1 11086
2 35385 1 11086
2 35386 1 11086
2 35387 1 11086
2 35388 1 11089
2 35389 1 11089
2 35390 1 11089
2 35391 1 11089
2 35392 1 11089
2 35393 1 11089
2 35394 1 11089
2 35395 1 11089
2 35396 1 11089
2 35397 1 11090
2 35398 1 11090
2 35399 1 11090
2 35400 1 11090
2 35401 1 11090
2 35402 1 11090
2 35403 1 11102
2 35404 1 11102
2 35405 1 11128
2 35406 1 11128
2 35407 1 11128
2 35408 1 11128
2 35409 1 11128
2 35410 1 11128
2 35411 1 11131
2 35412 1 11131
2 35413 1 11131
2 35414 1 11150
2 35415 1 11150
2 35416 1 11150
2 35417 1 11150
2 35418 1 11150
2 35419 1 11151
2 35420 1 11151
2 35421 1 11152
2 35422 1 11152
2 35423 1 11153
2 35424 1 11153
2 35425 1 11154
2 35426 1 11154
2 35427 1 11156
2 35428 1 11156
2 35429 1 11156
2 35430 1 11157
2 35431 1 11157
2 35432 1 11157
2 35433 1 11157
2 35434 1 11164
2 35435 1 11164
2 35436 1 11165
2 35437 1 11165
2 35438 1 11174
2 35439 1 11174
2 35440 1 11175
2 35441 1 11175
2 35442 1 11175
2 35443 1 11176
2 35444 1 11176
2 35445 1 11184
2 35446 1 11184
2 35447 1 11184
2 35448 1 11184
2 35449 1 11187
2 35450 1 11187
2 35451 1 11190
2 35452 1 11190
2 35453 1 11191
2 35454 1 11191
2 35455 1 11196
2 35456 1 11196
2 35457 1 11214
2 35458 1 11214
2 35459 1 11215
2 35460 1 11215
2 35461 1 11221
2 35462 1 11221
2 35463 1 11232
2 35464 1 11232
2 35465 1 11235
2 35466 1 11235
2 35467 1 11244
2 35468 1 11244
2 35469 1 11251
2 35470 1 11251
2 35471 1 11259
2 35472 1 11259
2 35473 1 11259
2 35474 1 11262
2 35475 1 11262
2 35476 1 11286
2 35477 1 11286
2 35478 1 11286
2 35479 1 11286
2 35480 1 11287
2 35481 1 11287
2 35482 1 11303
2 35483 1 11303
2 35484 1 11303
2 35485 1 11306
2 35486 1 11306
2 35487 1 11313
2 35488 1 11313
2 35489 1 11322
2 35490 1 11322
2 35491 1 11322
2 35492 1 11329
2 35493 1 11329
2 35494 1 11342
2 35495 1 11342
2 35496 1 11361
2 35497 1 11361
2 35498 1 11363
2 35499 1 11363
2 35500 1 11366
2 35501 1 11366
2 35502 1 11366
2 35503 1 11366
2 35504 1 11366
2 35505 1 11366
2 35506 1 11376
2 35507 1 11376
2 35508 1 11379
2 35509 1 11379
2 35510 1 11385
2 35511 1 11385
2 35512 1 11389
2 35513 1 11389
2 35514 1 11389
2 35515 1 11397
2 35516 1 11397
2 35517 1 11409
2 35518 1 11409
2 35519 1 11427
2 35520 1 11427
2 35521 1 11427
2 35522 1 11431
2 35523 1 11431
2 35524 1 11439
2 35525 1 11439
2 35526 1 11439
2 35527 1 11439
2 35528 1 11440
2 35529 1 11440
2 35530 1 11440
2 35531 1 11440
2 35532 1 11452
2 35533 1 11452
2 35534 1 11462
2 35535 1 11462
2 35536 1 11465
2 35537 1 11465
2 35538 1 11476
2 35539 1 11476
2 35540 1 11479
2 35541 1 11479
2 35542 1 11480
2 35543 1 11480
2 35544 1 11480
2 35545 1 11489
2 35546 1 11489
2 35547 1 11496
2 35548 1 11496
2 35549 1 11506
2 35550 1 11506
2 35551 1 11506
2 35552 1 11510
2 35553 1 11510
2 35554 1 11510
2 35555 1 11510
2 35556 1 11525
2 35557 1 11525
2 35558 1 11525
2 35559 1 11525
2 35560 1 11544
2 35561 1 11544
2 35562 1 11610
2 35563 1 11610
2 35564 1 11612
2 35565 1 11612
2 35566 1 11616
2 35567 1 11616
2 35568 1 11619
2 35569 1 11619
2 35570 1 11634
2 35571 1 11634
2 35572 1 11638
2 35573 1 11638
2 35574 1 11642
2 35575 1 11642
2 35576 1 11642
2 35577 1 11650
2 35578 1 11650
2 35579 1 11650
2 35580 1 11653
2 35581 1 11653
2 35582 1 11654
2 35583 1 11654
2 35584 1 11658
2 35585 1 11658
2 35586 1 11658
2 35587 1 11681
2 35588 1 11681
2 35589 1 11681
2 35590 1 11681
2 35591 1 11681
2 35592 1 11684
2 35593 1 11684
2 35594 1 11684
2 35595 1 11684
2 35596 1 11684
2 35597 1 11699
2 35598 1 11699
2 35599 1 11710
2 35600 1 11710
2 35601 1 11711
2 35602 1 11711
2 35603 1 11712
2 35604 1 11712
2 35605 1 11715
2 35606 1 11715
2 35607 1 11726
2 35608 1 11726
2 35609 1 11727
2 35610 1 11727
2 35611 1 11727
2 35612 1 11728
2 35613 1 11728
2 35614 1 11729
2 35615 1 11729
2 35616 1 11737
2 35617 1 11737
2 35618 1 11739
2 35619 1 11739
2 35620 1 11739
2 35621 1 11740
2 35622 1 11740
2 35623 1 11740
2 35624 1 11758
2 35625 1 11758
2 35626 1 11768
2 35627 1 11768
2 35628 1 11768
2 35629 1 11789
2 35630 1 11789
2 35631 1 11798
2 35632 1 11798
2 35633 1 11798
2 35634 1 11798
2 35635 1 11798
2 35636 1 11798
2 35637 1 11799
2 35638 1 11799
2 35639 1 11860
2 35640 1 11860
2 35641 1 11911
2 35642 1 11911
2 35643 1 11914
2 35644 1 11914
2 35645 1 11915
2 35646 1 11915
2 35647 1 11927
2 35648 1 11927
2 35649 1 11964
2 35650 1 11964
2 35651 1 11964
2 35652 1 11964
2 35653 1 11964
2 35654 1 11964
2 35655 1 11975
2 35656 1 11975
2 35657 1 11990
2 35658 1 11990
2 35659 1 12011
2 35660 1 12011
2 35661 1 12011
2 35662 1 12011
2 35663 1 12011
2 35664 1 12025
2 35665 1 12025
2 35666 1 12026
2 35667 1 12026
2 35668 1 12027
2 35669 1 12027
2 35670 1 12027
2 35671 1 12027
2 35672 1 12044
2 35673 1 12044
2 35674 1 12066
2 35675 1 12066
2 35676 1 12069
2 35677 1 12069
2 35678 1 12073
2 35679 1 12073
2 35680 1 12076
2 35681 1 12076
2 35682 1 12076
2 35683 1 12076
2 35684 1 12077
2 35685 1 12077
2 35686 1 12077
2 35687 1 12077
2 35688 1 12078
2 35689 1 12078
2 35690 1 12078
2 35691 1 12094
2 35692 1 12094
2 35693 1 12094
2 35694 1 12094
2 35695 1 12101
2 35696 1 12101
2 35697 1 12101
2 35698 1 12101
2 35699 1 12102
2 35700 1 12102
2 35701 1 12105
2 35702 1 12105
2 35703 1 12105
2 35704 1 12109
2 35705 1 12109
2 35706 1 12109
2 35707 1 12113
2 35708 1 12113
2 35709 1 12118
2 35710 1 12118
2 35711 1 12130
2 35712 1 12130
2 35713 1 12141
2 35714 1 12141
2 35715 1 12142
2 35716 1 12142
2 35717 1 12144
2 35718 1 12144
2 35719 1 12144
2 35720 1 12152
2 35721 1 12152
2 35722 1 12155
2 35723 1 12155
2 35724 1 12178
2 35725 1 12178
2 35726 1 12200
2 35727 1 12200
2 35728 1 12201
2 35729 1 12201
2 35730 1 12204
2 35731 1 12204
2 35732 1 12205
2 35733 1 12205
2 35734 1 12209
2 35735 1 12209
2 35736 1 12229
2 35737 1 12229
2 35738 1 12232
2 35739 1 12232
2 35740 1 12233
2 35741 1 12233
2 35742 1 12282
2 35743 1 12282
2 35744 1 12283
2 35745 1 12283
2 35746 1 12283
2 35747 1 12283
2 35748 1 12283
2 35749 1 12283
2 35750 1 12283
2 35751 1 12296
2 35752 1 12296
2 35753 1 12305
2 35754 1 12305
2 35755 1 12312
2 35756 1 12312
2 35757 1 12313
2 35758 1 12313
2 35759 1 12313
2 35760 1 12313
2 35761 1 12313
2 35762 1 12341
2 35763 1 12341
2 35764 1 12341
2 35765 1 12342
2 35766 1 12342
2 35767 1 12343
2 35768 1 12343
2 35769 1 12344
2 35770 1 12344
2 35771 1 12345
2 35772 1 12345
2 35773 1 12345
2 35774 1 12353
2 35775 1 12353
2 35776 1 12354
2 35777 1 12354
2 35778 1 12354
2 35779 1 12355
2 35780 1 12355
2 35781 1 12360
2 35782 1 12360
2 35783 1 12369
2 35784 1 12369
2 35785 1 12370
2 35786 1 12370
2 35787 1 12370
2 35788 1 12372
2 35789 1 12372
2 35790 1 12373
2 35791 1 12373
2 35792 1 12373
2 35793 1 12373
2 35794 1 12373
2 35795 1 12373
2 35796 1 12373
2 35797 1 12375
2 35798 1 12375
2 35799 1 12380
2 35800 1 12380
2 35801 1 12382
2 35802 1 12382
2 35803 1 12382
2 35804 1 12383
2 35805 1 12383
2 35806 1 12383
2 35807 1 12384
2 35808 1 12384
2 35809 1 12386
2 35810 1 12386
2 35811 1 12386
2 35812 1 12386
2 35813 1 12386
2 35814 1 12387
2 35815 1 12387
2 35816 1 12399
2 35817 1 12399
2 35818 1 12409
2 35819 1 12409
2 35820 1 12412
2 35821 1 12412
2 35822 1 12412
2 35823 1 12428
2 35824 1 12428
2 35825 1 12428
2 35826 1 12428
2 35827 1 12428
2 35828 1 12429
2 35829 1 12429
2 35830 1 12440
2 35831 1 12440
2 35832 1 12440
2 35833 1 12441
2 35834 1 12441
2 35835 1 12456
2 35836 1 12456
2 35837 1 12456
2 35838 1 12459
2 35839 1 12459
2 35840 1 12474
2 35841 1 12474
2 35842 1 12479
2 35843 1 12479
2 35844 1 12501
2 35845 1 12501
2 35846 1 12516
2 35847 1 12516
2 35848 1 12534
2 35849 1 12534
2 35850 1 12534
2 35851 1 12541
2 35852 1 12541
2 35853 1 12541
2 35854 1 12541
2 35855 1 12541
2 35856 1 12541
2 35857 1 12541
2 35858 1 12541
2 35859 1 12541
2 35860 1 12542
2 35861 1 12542
2 35862 1 12549
2 35863 1 12549
2 35864 1 12549
2 35865 1 12549
2 35866 1 12549
2 35867 1 12549
2 35868 1 12549
2 35869 1 12549
2 35870 1 12549
2 35871 1 12549
2 35872 1 12549
2 35873 1 12550
2 35874 1 12550
2 35875 1 12559
2 35876 1 12559
2 35877 1 12560
2 35878 1 12560
2 35879 1 12573
2 35880 1 12573
2 35881 1 12584
2 35882 1 12584
2 35883 1 12612
2 35884 1 12612
2 35885 1 12626
2 35886 1 12626
2 35887 1 12629
2 35888 1 12629
2 35889 1 12629
2 35890 1 12657
2 35891 1 12657
2 35892 1 12666
2 35893 1 12666
2 35894 1 12667
2 35895 1 12667
2 35896 1 12670
2 35897 1 12670
2 35898 1 12677
2 35899 1 12677
2 35900 1 12715
2 35901 1 12715
2 35902 1 12730
2 35903 1 12730
2 35904 1 12730
2 35905 1 12730
2 35906 1 12731
2 35907 1 12731
2 35908 1 12756
2 35909 1 12756
2 35910 1 12756
2 35911 1 12757
2 35912 1 12757
2 35913 1 12766
2 35914 1 12766
2 35915 1 12770
2 35916 1 12770
2 35917 1 12796
2 35918 1 12796
2 35919 1 12796
2 35920 1 12796
2 35921 1 12811
2 35922 1 12811
2 35923 1 12823
2 35924 1 12823
2 35925 1 12826
2 35926 1 12826
2 35927 1 12846
2 35928 1 12846
2 35929 1 12857
2 35930 1 12857
2 35931 1 12857
2 35932 1 12857
2 35933 1 12857
2 35934 1 12866
2 35935 1 12866
2 35936 1 12867
2 35937 1 12867
2 35938 1 12868
2 35939 1 12868
2 35940 1 12887
2 35941 1 12887
2 35942 1 12888
2 35943 1 12888
2 35944 1 12910
2 35945 1 12910
2 35946 1 12910
2 35947 1 12917
2 35948 1 12917
2 35949 1 12924
2 35950 1 12924
2 35951 1 12949
2 35952 1 12949
2 35953 1 12957
2 35954 1 12957
2 35955 1 12968
2 35956 1 12968
2 35957 1 12968
2 35958 1 12977
2 35959 1 12977
2 35960 1 12977
2 35961 1 12977
2 35962 1 12989
2 35963 1 12989
2 35964 1 12990
2 35965 1 12990
2 35966 1 12991
2 35967 1 12991
2 35968 1 13027
2 35969 1 13027
2 35970 1 13028
2 35971 1 13028
2 35972 1 13045
2 35973 1 13045
2 35974 1 13045
2 35975 1 13045
2 35976 1 13047
2 35977 1 13047
2 35978 1 13061
2 35979 1 13061
2 35980 1 13118
2 35981 1 13118
2 35982 1 13151
2 35983 1 13151
2 35984 1 13151
2 35985 1 13152
2 35986 1 13152
2 35987 1 13152
2 35988 1 13154
2 35989 1 13154
2 35990 1 13165
2 35991 1 13165
2 35992 1 13166
2 35993 1 13166
2 35994 1 13168
2 35995 1 13168
2 35996 1 13208
2 35997 1 13208
2 35998 1 13211
2 35999 1 13211
2 36000 1 13219
2 36001 1 13219
2 36002 1 13239
2 36003 1 13239
2 36004 1 13249
2 36005 1 13249
2 36006 1 13284
2 36007 1 13284
2 36008 1 13284
2 36009 1 13284
2 36010 1 13284
2 36011 1 13303
2 36012 1 13303
2 36013 1 13366
2 36014 1 13366
2 36015 1 13367
2 36016 1 13367
2 36017 1 13393
2 36018 1 13393
2 36019 1 13408
2 36020 1 13408
2 36021 1 13409
2 36022 1 13409
2 36023 1 13410
2 36024 1 13410
2 36025 1 13419
2 36026 1 13419
2 36027 1 13419
2 36028 1 13441
2 36029 1 13441
2 36030 1 13445
2 36031 1 13445
2 36032 1 13467
2 36033 1 13467
2 36034 1 13467
2 36035 1 13477
2 36036 1 13477
2 36037 1 13477
2 36038 1 13479
2 36039 1 13479
2 36040 1 13482
2 36041 1 13482
2 36042 1 13486
2 36043 1 13486
2 36044 1 13488
2 36045 1 13488
2 36046 1 13488
2 36047 1 13492
2 36048 1 13492
2 36049 1 13492
2 36050 1 13494
2 36051 1 13494
2 36052 1 13494
2 36053 1 13498
2 36054 1 13498
2 36055 1 13511
2 36056 1 13511
2 36057 1 13512
2 36058 1 13512
2 36059 1 13585
2 36060 1 13585
2 36061 1 13585
2 36062 1 13587
2 36063 1 13587
2 36064 1 13587
2 36065 1 13587
2 36066 1 13587
2 36067 1 13588
2 36068 1 13588
2 36069 1 13592
2 36070 1 13592
2 36071 1 13592
2 36072 1 13609
2 36073 1 13609
2 36074 1 13610
2 36075 1 13610
2 36076 1 13630
2 36077 1 13630
2 36078 1 13651
2 36079 1 13651
2 36080 1 13664
2 36081 1 13664
2 36082 1 13664
2 36083 1 13683
2 36084 1 13683
2 36085 1 13683
2 36086 1 13684
2 36087 1 13684
2 36088 1 13684
2 36089 1 13697
2 36090 1 13697
2 36091 1 13699
2 36092 1 13699
2 36093 1 13699
2 36094 1 13700
2 36095 1 13700
2 36096 1 13701
2 36097 1 13701
2 36098 1 13780
2 36099 1 13780
2 36100 1 13787
2 36101 1 13787
2 36102 1 13788
2 36103 1 13788
2 36104 1 13796
2 36105 1 13796
2 36106 1 13804
2 36107 1 13804
2 36108 1 13866
2 36109 1 13866
2 36110 1 13866
2 36111 1 13883
2 36112 1 13883
2 36113 1 13883
2 36114 1 13892
2 36115 1 13892
2 36116 1 13911
2 36117 1 13911
2 36118 1 13916
2 36119 1 13916
2 36120 1 13916
2 36121 1 13916
2 36122 1 13929
2 36123 1 13929
2 36124 1 13932
2 36125 1 13932
2 36126 1 13932
2 36127 1 13932
2 36128 1 13932
2 36129 1 13932
2 36130 1 13954
2 36131 1 13954
2 36132 1 13954
2 36133 1 13954
2 36134 1 13954
2 36135 1 13954
2 36136 1 13966
2 36137 1 13966
2 36138 1 13967
2 36139 1 13967
2 36140 1 13968
2 36141 1 13968
2 36142 1 13969
2 36143 1 13969
2 36144 1 13970
2 36145 1 13970
2 36146 1 13970
2 36147 1 13980
2 36148 1 13980
2 36149 1 13982
2 36150 1 13982
2 36151 1 13983
2 36152 1 13983
2 36153 1 13984
2 36154 1 13984
2 36155 1 13985
2 36156 1 13985
2 36157 1 13995
2 36158 1 13995
2 36159 1 14017
2 36160 1 14017
2 36161 1 14046
2 36162 1 14046
2 36163 1 14067
2 36164 1 14067
2 36165 1 14076
2 36166 1 14076
2 36167 1 14078
2 36168 1 14078
2 36169 1 14078
2 36170 1 14117
2 36171 1 14117
2 36172 1 14150
2 36173 1 14150
2 36174 1 14162
2 36175 1 14162
2 36176 1 14162
2 36177 1 14164
2 36178 1 14164
2 36179 1 14164
2 36180 1 14173
2 36181 1 14173
2 36182 1 14178
2 36183 1 14178
2 36184 1 14192
2 36185 1 14192
2 36186 1 14193
2 36187 1 14193
2 36188 1 14200
2 36189 1 14200
2 36190 1 14228
2 36191 1 14228
2 36192 1 14271
2 36193 1 14271
2 36194 1 14289
2 36195 1 14289
2 36196 1 14313
2 36197 1 14313
2 36198 1 14313
2 36199 1 14334
2 36200 1 14334
2 36201 1 14352
2 36202 1 14352
2 36203 1 14352
2 36204 1 14356
2 36205 1 14356
2 36206 1 14360
2 36207 1 14360
2 36208 1 14360
2 36209 1 14372
2 36210 1 14372
2 36211 1 14377
2 36212 1 14377
2 36213 1 14381
2 36214 1 14381
2 36215 1 14389
2 36216 1 14389
2 36217 1 14389
2 36218 1 14394
2 36219 1 14394
2 36220 1 14396
2 36221 1 14396
2 36222 1 14415
2 36223 1 14415
2 36224 1 14415
2 36225 1 14417
2 36226 1 14417
2 36227 1 14417
2 36228 1 14424
2 36229 1 14424
2 36230 1 14424
2 36231 1 14424
2 36232 1 14432
2 36233 1 14432
2 36234 1 14435
2 36235 1 14435
2 36236 1 14436
2 36237 1 14436
2 36238 1 14444
2 36239 1 14444
2 36240 1 14445
2 36241 1 14445
2 36242 1 14460
2 36243 1 14460
2 36244 1 14460
2 36245 1 14460
2 36246 1 14460
2 36247 1 14460
2 36248 1 14461
2 36249 1 14461
2 36250 1 14475
2 36251 1 14475
2 36252 1 14476
2 36253 1 14476
2 36254 1 14477
2 36255 1 14477
2 36256 1 14485
2 36257 1 14485
2 36258 1 14505
2 36259 1 14505
2 36260 1 14505
2 36261 1 14506
2 36262 1 14506
2 36263 1 14506
2 36264 1 14511
2 36265 1 14511
2 36266 1 14548
2 36267 1 14548
2 36268 1 14549
2 36269 1 14549
2 36270 1 14565
2 36271 1 14565
2 36272 1 14565
2 36273 1 14571
2 36274 1 14571
2 36275 1 14590
2 36276 1 14590
2 36277 1 14591
2 36278 1 14591
2 36279 1 14593
2 36280 1 14593
2 36281 1 14603
2 36282 1 14603
2 36283 1 14605
2 36284 1 14605
2 36285 1 14636
2 36286 1 14636
2 36287 1 14636
2 36288 1 14636
2 36289 1 14636
2 36290 1 14636
2 36291 1 14636
2 36292 1 14649
2 36293 1 14649
2 36294 1 14669
2 36295 1 14669
2 36296 1 14705
2 36297 1 14705
2 36298 1 14706
2 36299 1 14706
2 36300 1 14706
2 36301 1 14717
2 36302 1 14717
2 36303 1 14728
2 36304 1 14728
2 36305 1 14728
2 36306 1 14728
2 36307 1 14815
2 36308 1 14815
2 36309 1 14820
2 36310 1 14820
2 36311 1 14828
2 36312 1 14828
2 36313 1 14843
2 36314 1 14843
2 36315 1 14843
2 36316 1 14843
2 36317 1 14855
2 36318 1 14855
2 36319 1 14855
2 36320 1 14855
2 36321 1 14855
2 36322 1 14855
2 36323 1 14855
2 36324 1 14855
2 36325 1 14855
2 36326 1 14857
2 36327 1 14857
2 36328 1 14881
2 36329 1 14881
2 36330 1 14881
2 36331 1 14881
2 36332 1 14881
2 36333 1 14881
2 36334 1 14902
2 36335 1 14902
2 36336 1 14932
2 36337 1 14932
2 36338 1 14968
2 36339 1 14968
2 36340 1 15016
2 36341 1 15016
2 36342 1 15037
2 36343 1 15037
2 36344 1 15055
2 36345 1 15055
2 36346 1 15059
2 36347 1 15059
2 36348 1 15092
2 36349 1 15092
2 36350 1 15125
2 36351 1 15125
2 36352 1 15162
2 36353 1 15162
2 36354 1 15165
2 36355 1 15165
2 36356 1 15194
2 36357 1 15194
2 36358 1 15194
2 36359 1 15197
2 36360 1 15197
2 36361 1 15197
2 36362 1 15197
2 36363 1 15205
2 36364 1 15205
2 36365 1 15208
2 36366 1 15208
2 36367 1 15209
2 36368 1 15209
2 36369 1 15221
2 36370 1 15221
2 36371 1 15238
2 36372 1 15238
2 36373 1 15254
2 36374 1 15254
2 36375 1 15254
2 36376 1 15254
2 36377 1 15255
2 36378 1 15255
2 36379 1 15255
2 36380 1 15255
2 36381 1 15255
2 36382 1 15256
2 36383 1 15256
2 36384 1 15264
2 36385 1 15264
2 36386 1 15278
2 36387 1 15278
2 36388 1 15293
2 36389 1 15293
2 36390 1 15293
2 36391 1 15296
2 36392 1 15296
2 36393 1 15296
2 36394 1 15296
2 36395 1 15296
2 36396 1 15296
2 36397 1 15296
2 36398 1 15296
2 36399 1 15296
2 36400 1 15296
2 36401 1 15296
2 36402 1 15296
2 36403 1 15296
2 36404 1 15296
2 36405 1 15296
2 36406 1 15296
2 36407 1 15296
2 36408 1 15296
2 36409 1 15296
2 36410 1 15296
2 36411 1 15296
2 36412 1 15296
2 36413 1 15296
2 36414 1 15296
2 36415 1 15296
2 36416 1 15296
2 36417 1 15296
2 36418 1 15299
2 36419 1 15299
2 36420 1 15299
2 36421 1 15299
2 36422 1 15299
2 36423 1 15299
2 36424 1 15299
2 36425 1 15299
2 36426 1 15299
2 36427 1 15299
2 36428 1 15300
2 36429 1 15300
2 36430 1 15300
2 36431 1 15303
2 36432 1 15303
2 36433 1 15308
2 36434 1 15308
2 36435 1 15311
2 36436 1 15311
2 36437 1 15318
2 36438 1 15318
2 36439 1 15319
2 36440 1 15319
2 36441 1 15319
2 36442 1 15320
2 36443 1 15320
2 36444 1 15328
2 36445 1 15328
2 36446 1 15329
2 36447 1 15329
2 36448 1 15329
2 36449 1 15329
2 36450 1 15329
2 36451 1 15329
2 36452 1 15331
2 36453 1 15331
2 36454 1 15338
2 36455 1 15338
2 36456 1 15354
2 36457 1 15354
2 36458 1 15366
2 36459 1 15366
2 36460 1 15366
2 36461 1 15366
2 36462 1 15379
2 36463 1 15379
2 36464 1 15386
2 36465 1 15386
2 36466 1 15387
2 36467 1 15387
2 36468 1 15387
2 36469 1 15396
2 36470 1 15396
2 36471 1 15398
2 36472 1 15398
2 36473 1 15405
2 36474 1 15405
2 36475 1 15405
2 36476 1 15405
2 36477 1 15405
2 36478 1 15405
2 36479 1 15405
2 36480 1 15409
2 36481 1 15409
2 36482 1 15428
2 36483 1 15428
2 36484 1 15429
2 36485 1 15429
2 36486 1 15442
2 36487 1 15442
2 36488 1 15442
2 36489 1 15442
2 36490 1 15442
2 36491 1 15443
2 36492 1 15443
2 36493 1 15443
2 36494 1 15443
2 36495 1 15445
2 36496 1 15445
2 36497 1 15445
2 36498 1 15445
2 36499 1 15468
2 36500 1 15468
2 36501 1 15469
2 36502 1 15469
2 36503 1 15469
2 36504 1 15471
2 36505 1 15471
2 36506 1 15489
2 36507 1 15489
2 36508 1 15489
2 36509 1 15489
2 36510 1 15489
2 36511 1 15489
2 36512 1 15489
2 36513 1 15489
2 36514 1 15500
2 36515 1 15500
2 36516 1 15500
2 36517 1 15500
2 36518 1 15500
2 36519 1 15502
2 36520 1 15502
2 36521 1 15502
2 36522 1 15502
2 36523 1 15502
2 36524 1 15502
2 36525 1 15502
2 36526 1 15503
2 36527 1 15503
2 36528 1 15531
2 36529 1 15531
2 36530 1 15531
2 36531 1 15547
2 36532 1 15547
2 36533 1 15548
2 36534 1 15548
2 36535 1 15550
2 36536 1 15550
2 36537 1 15550
2 36538 1 15550
2 36539 1 15550
2 36540 1 15564
2 36541 1 15564
2 36542 1 15565
2 36543 1 15565
2 36544 1 15565
2 36545 1 15567
2 36546 1 15567
2 36547 1 15570
2 36548 1 15570
2 36549 1 15570
2 36550 1 15580
2 36551 1 15580
2 36552 1 15595
2 36553 1 15595
2 36554 1 15595
2 36555 1 15595
2 36556 1 15595
2 36557 1 15595
2 36558 1 15595
2 36559 1 15595
2 36560 1 15595
2 36561 1 15595
2 36562 1 15595
2 36563 1 15595
2 36564 1 15595
2 36565 1 15595
2 36566 1 15595
2 36567 1 15595
2 36568 1 15595
2 36569 1 15595
2 36570 1 15595
2 36571 1 15595
2 36572 1 15595
2 36573 1 15595
2 36574 1 15595
2 36575 1 15595
2 36576 1 15595
2 36577 1 15596
2 36578 1 15596
2 36579 1 15600
2 36580 1 15600
2 36581 1 15605
2 36582 1 15605
2 36583 1 15605
2 36584 1 15605
2 36585 1 15605
2 36586 1 15605
2 36587 1 15606
2 36588 1 15606
2 36589 1 15608
2 36590 1 15608
2 36591 1 15612
2 36592 1 15612
2 36593 1 15612
2 36594 1 15613
2 36595 1 15613
2 36596 1 15614
2 36597 1 15614
2 36598 1 15627
2 36599 1 15627
2 36600 1 15629
2 36601 1 15629
2 36602 1 15629
2 36603 1 15630
2 36604 1 15630
2 36605 1 15638
2 36606 1 15638
2 36607 1 15638
2 36608 1 15638
2 36609 1 15638
2 36610 1 15638
2 36611 1 15638
2 36612 1 15638
2 36613 1 15638
2 36614 1 15640
2 36615 1 15640
2 36616 1 15640
2 36617 1 15654
2 36618 1 15654
2 36619 1 15655
2 36620 1 15655
2 36621 1 15658
2 36622 1 15658
2 36623 1 15659
2 36624 1 15659
2 36625 1 15664
2 36626 1 15664
2 36627 1 15667
2 36628 1 15667
2 36629 1 15667
2 36630 1 15675
2 36631 1 15675
2 36632 1 15687
2 36633 1 15687
2 36634 1 15687
2 36635 1 15700
2 36636 1 15700
2 36637 1 15700
2 36638 1 15710
2 36639 1 15710
2 36640 1 15710
2 36641 1 15712
2 36642 1 15712
2 36643 1 15714
2 36644 1 15714
2 36645 1 15725
2 36646 1 15725
2 36647 1 15725
2 36648 1 15725
2 36649 1 15725
2 36650 1 15726
2 36651 1 15726
2 36652 1 15727
2 36653 1 15727
2 36654 1 15728
2 36655 1 15728
2 36656 1 15791
2 36657 1 15791
2 36658 1 15794
2 36659 1 15794
2 36660 1 15808
2 36661 1 15808
2 36662 1 15808
2 36663 1 15808
2 36664 1 15819
2 36665 1 15819
2 36666 1 15819
2 36667 1 15823
2 36668 1 15823
2 36669 1 15823
2 36670 1 15823
2 36671 1 15823
2 36672 1 15823
2 36673 1 15823
2 36674 1 15824
2 36675 1 15824
2 36676 1 15848
2 36677 1 15848
2 36678 1 15868
2 36679 1 15868
2 36680 1 15871
2 36681 1 15871
2 36682 1 15871
2 36683 1 15871
2 36684 1 15871
2 36685 1 15871
2 36686 1 15871
2 36687 1 15872
2 36688 1 15872
2 36689 1 15873
2 36690 1 15873
2 36691 1 15884
2 36692 1 15884
2 36693 1 15887
2 36694 1 15887
2 36695 1 15888
2 36696 1 15888
2 36697 1 15888
2 36698 1 15891
2 36699 1 15891
2 36700 1 15896
2 36701 1 15896
2 36702 1 15915
2 36703 1 15915
2 36704 1 15926
2 36705 1 15926
2 36706 1 15953
2 36707 1 15953
2 36708 1 15954
2 36709 1 15954
2 36710 1 15971
2 36711 1 15971
2 36712 1 16010
2 36713 1 16010
2 36714 1 16010
2 36715 1 16010
2 36716 1 16010
2 36717 1 16011
2 36718 1 16011
2 36719 1 16012
2 36720 1 16012
2 36721 1 16020
2 36722 1 16020
2 36723 1 16022
2 36724 1 16022
2 36725 1 16022
2 36726 1 16022
2 36727 1 16027
2 36728 1 16027
2 36729 1 16028
2 36730 1 16028
2 36731 1 16040
2 36732 1 16040
2 36733 1 16043
2 36734 1 16043
2 36735 1 16044
2 36736 1 16044
2 36737 1 16059
2 36738 1 16059
2 36739 1 16059
2 36740 1 16074
2 36741 1 16074
2 36742 1 16083
2 36743 1 16083
2 36744 1 16113
2 36745 1 16113
2 36746 1 16114
2 36747 1 16114
2 36748 1 16114
2 36749 1 16115
2 36750 1 16115
2 36751 1 16115
2 36752 1 16115
2 36753 1 16115
2 36754 1 16122
2 36755 1 16122
2 36756 1 16123
2 36757 1 16123
2 36758 1 16132
2 36759 1 16132
2 36760 1 16133
2 36761 1 16133
2 36762 1 16134
2 36763 1 16134
2 36764 1 16138
2 36765 1 16138
2 36766 1 16164
2 36767 1 16164
2 36768 1 16164
2 36769 1 16164
2 36770 1 16164
2 36771 1 16167
2 36772 1 16167
2 36773 1 16188
2 36774 1 16188
2 36775 1 16188
2 36776 1 16188
2 36777 1 16219
2 36778 1 16219
2 36779 1 16235
2 36780 1 16235
2 36781 1 16235
2 36782 1 16235
2 36783 1 16235
2 36784 1 16236
2 36785 1 16236
2 36786 1 16236
2 36787 1 16245
2 36788 1 16245
2 36789 1 16259
2 36790 1 16259
2 36791 1 16270
2 36792 1 16270
2 36793 1 16271
2 36794 1 16271
2 36795 1 16271
2 36796 1 16280
2 36797 1 16280
2 36798 1 16286
2 36799 1 16286
2 36800 1 16286
2 36801 1 16289
2 36802 1 16289
2 36803 1 16291
2 36804 1 16291
2 36805 1 16309
2 36806 1 16309
2 36807 1 16336
2 36808 1 16336
2 36809 1 16336
2 36810 1 16336
2 36811 1 16336
2 36812 1 16353
2 36813 1 16353
2 36814 1 16369
2 36815 1 16369
2 36816 1 16450
2 36817 1 16450
2 36818 1 16455
2 36819 1 16455
2 36820 1 16462
2 36821 1 16462
2 36822 1 16462
2 36823 1 16462
2 36824 1 16462
2 36825 1 16471
2 36826 1 16471
2 36827 1 16478
2 36828 1 16478
2 36829 1 16496
2 36830 1 16496
2 36831 1 16496
2 36832 1 16496
2 36833 1 16496
2 36834 1 16501
2 36835 1 16501
2 36836 1 16522
2 36837 1 16522
2 36838 1 16548
2 36839 1 16548
2 36840 1 16566
2 36841 1 16566
2 36842 1 16566
2 36843 1 16574
2 36844 1 16574
2 36845 1 16590
2 36846 1 16590
2 36847 1 16621
2 36848 1 16621
2 36849 1 16702
2 36850 1 16702
2 36851 1 16705
2 36852 1 16705
2 36853 1 16720
2 36854 1 16720
2 36855 1 16721
2 36856 1 16721
2 36857 1 16742
2 36858 1 16742
2 36859 1 16743
2 36860 1 16743
2 36861 1 16750
2 36862 1 16750
2 36863 1 16759
2 36864 1 16759
2 36865 1 16797
2 36866 1 16797
2 36867 1 16818
2 36868 1 16818
2 36869 1 16820
2 36870 1 16820
2 36871 1 16820
2 36872 1 16820
2 36873 1 16820
2 36874 1 16823
2 36875 1 16823
2 36876 1 16830
2 36877 1 16830
2 36878 1 16834
2 36879 1 16834
2 36880 1 16834
2 36881 1 16841
2 36882 1 16841
2 36883 1 16844
2 36884 1 16844
2 36885 1 16845
2 36886 1 16845
2 36887 1 16845
2 36888 1 16852
2 36889 1 16852
2 36890 1 16864
2 36891 1 16864
2 36892 1 16931
2 36893 1 16931
2 36894 1 16931
2 36895 1 16946
2 36896 1 16946
2 36897 1 16946
2 36898 1 16974
2 36899 1 16974
2 36900 1 16992
2 36901 1 16992
2 36902 1 16993
2 36903 1 16993
2 36904 1 17011
2 36905 1 17011
2 36906 1 17066
2 36907 1 17066
2 36908 1 17110
2 36909 1 17110
2 36910 1 17110
2 36911 1 17110
2 36912 1 17121
2 36913 1 17121
2 36914 1 17122
2 36915 1 17122
2 36916 1 17127
2 36917 1 17127
2 36918 1 17130
2 36919 1 17130
2 36920 1 17130
2 36921 1 17130
2 36922 1 17130
2 36923 1 17131
2 36924 1 17131
2 36925 1 17131
2 36926 1 17131
2 36927 1 17132
2 36928 1 17132
2 36929 1 17142
2 36930 1 17142
2 36931 1 17150
2 36932 1 17150
2 36933 1 17173
2 36934 1 17173
2 36935 1 17173
2 36936 1 17175
2 36937 1 17175
2 36938 1 17180
2 36939 1 17180
2 36940 1 17180
2 36941 1 17183
2 36942 1 17183
2 36943 1 17184
2 36944 1 17184
2 36945 1 17199
2 36946 1 17199
2 36947 1 17203
2 36948 1 17203
2 36949 1 17203
2 36950 1 17206
2 36951 1 17206
2 36952 1 17216
2 36953 1 17216
2 36954 1 17260
2 36955 1 17260
2 36956 1 17261
2 36957 1 17261
2 36958 1 17275
2 36959 1 17275
2 36960 1 17275
2 36961 1 17293
2 36962 1 17293
2 36963 1 17293
2 36964 1 17293
2 36965 1 17296
2 36966 1 17296
2 36967 1 17296
2 36968 1 17300
2 36969 1 17300
2 36970 1 17305
2 36971 1 17305
2 36972 1 17305
2 36973 1 17397
2 36974 1 17397
2 36975 1 17414
2 36976 1 17414
2 36977 1 17414
2 36978 1 17476
2 36979 1 17476
2 36980 1 17502
2 36981 1 17502
2 36982 1 17528
2 36983 1 17528
2 36984 1 17569
2 36985 1 17569
2 36986 1 17569
2 36987 1 17577
2 36988 1 17577
2 36989 1 17584
2 36990 1 17584
2 36991 1 17586
2 36992 1 17586
2 36993 1 17588
2 36994 1 17588
2 36995 1 17589
2 36996 1 17589
2 36997 1 17592
2 36998 1 17592
2 36999 1 17592
2 37000 1 17601
2 37001 1 17601
2 37002 1 17604
2 37003 1 17604
2 37004 1 17604
2 37005 1 17660
2 37006 1 17660
2 37007 1 17660
2 37008 1 17665
2 37009 1 17665
2 37010 1 17679
2 37011 1 17679
2 37012 1 17682
2 37013 1 17682
2 37014 1 17682
2 37015 1 17683
2 37016 1 17683
2 37017 1 17711
2 37018 1 17711
2 37019 1 17713
2 37020 1 17713
2 37021 1 17718
2 37022 1 17718
2 37023 1 17766
2 37024 1 17766
2 37025 1 17800
2 37026 1 17800
2 37027 1 17817
2 37028 1 17817
2 37029 1 17824
2 37030 1 17824
2 37031 1 17827
2 37032 1 17827
2 37033 1 17827
2 37034 1 17893
2 37035 1 17893
2 37036 1 17893
2 37037 1 17893
2 37038 1 17899
2 37039 1 17899
2 37040 1 17899
2 37041 1 17900
2 37042 1 17900
2 37043 1 17901
2 37044 1 17901
2 37045 1 17922
2 37046 1 17922
2 37047 1 17931
2 37048 1 17931
2 37049 1 17939
2 37050 1 17939
2 37051 1 18041
2 37052 1 18041
2 37053 1 18061
2 37054 1 18061
2 37055 1 18144
2 37056 1 18144
2 37057 1 18165
2 37058 1 18165
2 37059 1 18186
2 37060 1 18186
2 37061 1 18201
2 37062 1 18201
2 37063 1 18218
2 37064 1 18218
2 37065 1 18226
2 37066 1 18226
2 37067 1 18226
2 37068 1 18226
2 37069 1 18238
2 37070 1 18238
2 37071 1 18238
2 37072 1 18239
2 37073 1 18239
2 37074 1 18239
2 37075 1 18239
2 37076 1 18245
2 37077 1 18245
2 37078 1 18250
2 37079 1 18250
2 37080 1 18253
2 37081 1 18253
2 37082 1 18253
2 37083 1 18262
2 37084 1 18262
2 37085 1 18262
2 37086 1 18263
2 37087 1 18263
2 37088 1 18274
2 37089 1 18274
2 37090 1 18281
2 37091 1 18281
2 37092 1 18293
2 37093 1 18293
2 37094 1 18341
2 37095 1 18341
2 37096 1 18350
2 37097 1 18350
2 37098 1 18361
2 37099 1 18361
2 37100 1 18368
2 37101 1 18368
2 37102 1 18371
2 37103 1 18371
2 37104 1 18376
2 37105 1 18376
2 37106 1 18379
2 37107 1 18379
2 37108 1 18395
2 37109 1 18395
2 37110 1 18395
2 37111 1 18396
2 37112 1 18396
2 37113 1 18436
2 37114 1 18436
2 37115 1 18436
2 37116 1 18437
2 37117 1 18437
2 37118 1 18437
2 37119 1 18437
2 37120 1 18447
2 37121 1 18447
2 37122 1 18453
2 37123 1 18453
2 37124 1 18453
2 37125 1 18453
2 37126 1 18471
2 37127 1 18471
2 37128 1 18478
2 37129 1 18478
2 37130 1 18487
2 37131 1 18487
2 37132 1 18500
2 37133 1 18500
2 37134 1 18546
2 37135 1 18546
2 37136 1 18586
2 37137 1 18586
2 37138 1 18586
2 37139 1 18587
2 37140 1 18587
2 37141 1 18587
2 37142 1 18588
2 37143 1 18588
2 37144 1 18588
2 37145 1 18588
2 37146 1 18591
2 37147 1 18591
2 37148 1 18592
2 37149 1 18592
2 37150 1 18641
2 37151 1 18641
2 37152 1 18645
2 37153 1 18645
2 37154 1 18645
2 37155 1 18648
2 37156 1 18648
2 37157 1 18649
2 37158 1 18649
2 37159 1 18649
2 37160 1 18672
2 37161 1 18672
2 37162 1 18683
2 37163 1 18683
2 37164 1 18684
2 37165 1 18684
2 37166 1 18684
2 37167 1 18684
2 37168 1 18684
2 37169 1 18685
2 37170 1 18685
2 37171 1 18688
2 37172 1 18688
2 37173 1 18709
2 37174 1 18709
2 37175 1 18743
2 37176 1 18743
2 37177 1 18743
2 37178 1 18747
2 37179 1 18747
2 37180 1 18748
2 37181 1 18748
2 37182 1 18749
2 37183 1 18749
2 37184 1 18749
2 37185 1 18766
2 37186 1 18766
2 37187 1 18814
2 37188 1 18814
2 37189 1 18816
2 37190 1 18816
2 37191 1 18842
2 37192 1 18842
2 37193 1 18852
2 37194 1 18852
2 37195 1 18888
2 37196 1 18888
2 37197 1 18897
2 37198 1 18897
2 37199 1 18897
2 37200 1 18898
2 37201 1 18898
2 37202 1 18930
2 37203 1 18930
2 37204 1 18984
2 37205 1 18984
2 37206 1 19001
2 37207 1 19001
2 37208 1 19021
2 37209 1 19021
2 37210 1 19037
2 37211 1 19037
2 37212 1 19054
2 37213 1 19054
2 37214 1 19070
2 37215 1 19070
2 37216 1 19162
2 37217 1 19162
2 37218 1 19163
2 37219 1 19163
2 37220 1 19237
2 37221 1 19237
2 37222 1 19237
2 37223 1 19237
2 37224 1 19280
2 37225 1 19280
2 37226 1 19311
2 37227 1 19311
2 37228 1 19314
2 37229 1 19314
2 37230 1 19381
2 37231 1 19381
2 37232 1 19503
2 37233 1 19503
2 37234 1 19532
2 37235 1 19532
2 37236 1 19566
2 37237 1 19566
2 37238 1 19581
2 37239 1 19581
2 37240 1 19591
2 37241 1 19591
2 37242 1 19600
2 37243 1 19600
2 37244 1 19616
2 37245 1 19616
2 37246 1 19663
2 37247 1 19663
2 37248 1 19669
2 37249 1 19669
2 37250 1 19696
2 37251 1 19696
2 37252 1 19699
2 37253 1 19699
2 37254 1 19702
2 37255 1 19702
2 37256 1 19720
2 37257 1 19720
2 37258 1 19729
2 37259 1 19729
2 37260 1 19738
2 37261 1 19738
2 37262 1 19775
2 37263 1 19775
2 37264 1 19816
2 37265 1 19816
2 37266 1 19824
2 37267 1 19824
2 37268 1 19828
2 37269 1 19828
2 37270 1 19856
2 37271 1 19856
2 37272 1 20036
2 37273 1 20036
2 37274 1 20063
2 37275 1 20063
2 37276 1 20091
2 37277 1 20091
2 37278 1 20120
2 37279 1 20120
2 37280 1 20144
2 37281 1 20144
2 37282 1 20172
2 37283 1 20172
2 37284 1 20178
2 37285 1 20178
2 37286 1 20246
2 37287 1 20246
2 37288 1 20287
2 37289 1 20287
2 37290 1 20287
2 37291 1 20287
2 37292 1 20287
2 37293 1 20287
2 37294 1 20287
2 37295 1 20287
2 37296 1 20287
2 37297 1 20295
2 37298 1 20295
2 37299 1 20295
2 37300 1 20367
2 37301 1 20367
2 37302 1 20372
2 37303 1 20372
2 37304 1 20378
2 37305 1 20378
2 37306 1 20386
2 37307 1 20386
2 37308 1 20386
2 37309 1 20386
2 37310 1 20390
2 37311 1 20390
2 37312 1 20390
2 37313 1 20390
2 37314 1 20430
2 37315 1 20430
2 37316 1 20446
2 37317 1 20446
2 37318 1 20446
2 37319 1 20450
2 37320 1 20450
2 37321 1 20478
2 37322 1 20478
2 37323 1 20481
2 37324 1 20481
2 37325 1 20481
2 37326 1 20481
2 37327 1 20482
2 37328 1 20482
2 37329 1 20520
2 37330 1 20520
2 37331 1 20526
2 37332 1 20526
2 37333 1 20526
2 37334 1 20530
2 37335 1 20530
2 37336 1 20533
2 37337 1 20533
2 37338 1 20552
2 37339 1 20552
2 37340 1 20596
2 37341 1 20596
2 37342 1 20605
2 37343 1 20605
2 37344 1 20605
2 37345 1 20606
2 37346 1 20606
2 37347 1 20606
2 37348 1 20608
2 37349 1 20608
2 37350 1 20608
2 37351 1 20612
2 37352 1 20612
2 37353 1 20614
2 37354 1 20614
2 37355 1 20615
2 37356 1 20615
2 37357 1 20623
2 37358 1 20623
2 37359 1 20626
2 37360 1 20626
2 37361 1 20630
2 37362 1 20630
2 37363 1 20630
2 37364 1 20630
2 37365 1 20630
2 37366 1 20641
2 37367 1 20641
2 37368 1 20650
2 37369 1 20650
2 37370 1 20676
2 37371 1 20676
2 37372 1 20721
2 37373 1 20721
2 37374 1 20721
2 37375 1 20740
2 37376 1 20740
2 37377 1 20758
2 37378 1 20758
2 37379 1 20759
2 37380 1 20759
2 37381 1 20764
2 37382 1 20764
2 37383 1 20779
2 37384 1 20779
2 37385 1 20782
2 37386 1 20782
2 37387 1 20788
2 37388 1 20788
2 37389 1 20790
2 37390 1 20790
2 37391 1 20790
2 37392 1 20814
2 37393 1 20814
2 37394 1 20821
2 37395 1 20821
2 37396 1 20847
2 37397 1 20847
2 37398 1 20880
2 37399 1 20880
2 37400 1 20887
2 37401 1 20887
2 37402 1 20948
2 37403 1 20948
2 37404 1 21097
2 37405 1 21097
2 37406 1 21124
2 37407 1 21124
2 37408 1 21135
2 37409 1 21135
2 37410 1 21174
2 37411 1 21174
2 37412 1 21196
2 37413 1 21196
2 37414 1 21200
2 37415 1 21200
2 37416 1 21212
2 37417 1 21212
2 37418 1 21225
2 37419 1 21225
2 37420 1 21245
2 37421 1 21245
2 37422 1 21261
2 37423 1 21261
2 37424 1 21261
2 37425 1 21262
2 37426 1 21262
2 37427 1 21271
2 37428 1 21271
2 37429 1 21279
2 37430 1 21279
2 37431 1 21280
2 37432 1 21280
2 37433 1 21335
2 37434 1 21335
2 37435 1 21337
2 37436 1 21337
2 37437 1 21453
2 37438 1 21453
2 37439 1 21475
2 37440 1 21475
2 37441 1 21496
2 37442 1 21496
2 37443 1 21511
2 37444 1 21511
2 37445 1 21518
2 37446 1 21518
2 37447 1 21574
2 37448 1 21574
2 37449 1 21603
2 37450 1 21603
2 37451 1 21634
2 37452 1 21634
2 37453 1 21634
2 37454 1 21636
2 37455 1 21636
2 37456 1 21691
2 37457 1 21691
2 37458 1 21693
2 37459 1 21693
0 27 5 120 1 25
0 28 5 115 1 21854
0 29 5 128 1 21972
0 30 5 46 1 22115
0 31 5 74 1 22166
0 32 5 45 1 22241
0 33 5 56 1 22281
0 34 5 71 1 22349
0 35 5 62 1 22428
0 36 5 60 1 22493
0 37 5 86 1 22586
0 38 5 30 1 22687
0 39 5 65 1 22726
0 40 5 39 1 22785
0 41 5 58 1 22822
0 42 5 61 1 22885
0 43 5 108 1 22955
0 44 5 120 1 23033
0 45 5 81 1 23156
0 46 5 95 1 23241
0 47 5 70 1 23331
0 48 5 70 1 23394
0 49 5 106 1 23482
0 50 5 100 1 23591
0 51 5 50 1 23701
0 52 7 2 2 24255 22786
0 53 5 1 1 25688
0 54 7 5 2 22242 24730
0 55 5 1 1 25690
0 56 7 2 2 53 55
0 57 5 41 1 25695
0 58 7 29 2 24181 24665
0 59 5 1 1 25738
0 60 7 8 2 24769 24827
0 61 7 6 2 25638 25767
0 62 7 9 2 24300 24356
0 63 7 2 2 24888 25781
0 64 7 2 2 25775 25790
0 65 7 16 2 25197 23332
0 66 7 10 2 24996 25116
0 67 5 2 1 25810
0 68 7 5 2 25794 25811
0 69 7 1 2 25792 25822
0 70 5 1 1 69
0 71 7 44 2 22282 22823
0 72 5 3 1 25827
0 73 7 5 2 24357 22886
0 74 5 1 1 25874
0 75 7 11 2 22350 24828
0 76 5 1 1 25879
0 77 7 4 2 74 76
0 78 5 70 1 25890
0 79 7 2 2 25828 25894
0 80 5 1 1 25964
0 81 7 2 2 22351 24770
0 82 7 2 2 24301 22887
0 83 7 9 2 25966 25968
0 84 5 1 1 25970
0 85 7 1 2 80 84
0 86 5 17 1 85
0 87 7 10 2 23702 25979
0 88 5 1 1 25996
0 89 7 20 2 23242 25292
0 90 7 4 2 22956 23157
0 91 7 3 2 26006 26026
0 92 7 1 2 25997 26030
0 93 5 1 1 92
0 94 7 1 2 70 93
0 95 5 1 1 94
0 96 7 1 2 24427 95
0 97 5 1 1 96
0 98 7 9 2 22429 22957
0 99 5 1 1 26033
0 100 7 2 2 25639 26034
0 101 7 55 2 24302 24771
0 102 5 2 1 26044
0 103 7 28 2 24358 24829
0 104 5 10 1 26101
0 105 7 3 2 26045 26102
0 106 7 1 2 26139 25823
0 107 7 1 2 26042 106
0 108 5 1 1 107
0 109 7 1 2 97 108
0 110 5 1 1 109
0 111 7 1 2 24549 110
0 112 5 1 1 111
0 113 7 20 2 24428 22958
0 114 5 22 1 26142
0 115 7 5 2 25117 25795
0 116 5 1 1 26184
0 117 7 1 2 26143 26185
0 118 7 1 2 25998 117
0 119 5 1 1 118
0 120 7 1 2 112 119
0 121 5 1 1 120
0 122 7 1 2 25538 121
0 123 5 1 1 122
0 124 7 29 2 22352 22888
0 125 5 15 1 26189
0 126 7 7 2 22959 23592
0 127 5 1 1 26233
0 128 7 5 2 26190 26234
0 129 5 1 1 26240
0 130 7 2 2 25829 26241
0 131 5 1 1 26245
0 132 7 25 2 24550 23158
0 133 5 3 1 26247
0 134 7 4 2 26248 26007
0 135 5 2 1 26275
0 136 7 1 2 116 26279
0 137 5 8 1 136
0 138 7 1 2 23703 26281
0 139 7 1 2 26246 138
0 140 5 1 1 139
0 141 7 1 2 123 140
0 142 5 1 1 141
0 143 7 1 2 22116 142
0 144 5 1 1 143
0 145 7 2 2 24135 25118
0 146 5 2 1 26289
0 147 7 1 2 26008 26290
0 148 5 2 1 147
0 149 7 18 2 22587 25119
0 150 5 2 1 26295
0 151 7 4 2 25796 26296
0 152 5 3 1 26315
0 153 7 1 2 26280 26319
0 154 5 4 1 153
0 155 7 2 2 24997 26322
0 156 5 1 1 26326
0 157 7 1 2 24889 26327
0 158 5 1 1 157
0 159 7 1 2 26293 158
0 160 5 2 1 159
0 161 7 3 2 23704 25830
0 162 7 11 2 23593 26191
0 163 5 1 1 26333
0 164 7 10 2 26330 26334
0 165 5 2 1 26344
0 166 7 1 2 24429 26345
0 167 7 1 2 26328 166
0 168 5 1 1 167
0 169 7 1 2 144 168
0 170 5 1 1 169
0 171 7 1 2 22688 170
0 172 5 1 1 171
0 173 7 6 2 24635 25120
0 174 5 1 1 26356
0 175 7 1 2 25539 25891
0 176 5 3 1 175
0 177 7 6 2 22960 25540
0 178 5 1 1 26365
0 179 7 1 2 26218 178
0 180 5 1 1 179
0 181 7 2 2 26362 180
0 182 7 1 2 26357 26371
0 183 5 1 1 182
0 184 7 14 2 24890 24998
0 185 5 3 1 26373
0 186 7 3 2 26249 26374
0 187 5 4 1 26390
0 188 7 21 2 22889 23594
0 189 5 3 1 26397
0 190 7 9 2 22353 26398
0 191 5 3 1 26421
0 192 7 1 2 26391 26422
0 193 5 1 1 192
0 194 7 1 2 183 193
0 195 5 1 1 194
0 196 7 1 2 24430 195
0 197 5 1 1 196
0 198 7 1 2 26358 26242
0 199 5 1 1 198
0 200 7 1 2 197 199
0 201 5 1 1 200
0 202 7 1 2 25831 201
0 203 5 1 1 202
0 204 7 7 2 22354 24431
0 205 7 2 2 26046 26433
0 206 7 4 2 22890 26366
0 207 7 1 2 26359 26442
0 208 7 1 2 26440 207
0 209 5 1 1 208
0 210 7 1 2 203 209
0 211 5 1 1 210
0 212 7 9 2 25198 25293
0 213 7 3 2 23705 26446
0 214 7 1 2 24136 26455
0 215 7 1 2 211 214
0 216 5 1 1 215
0 217 7 1 2 172 216
0 218 5 1 1 217
0 219 7 1 2 23395 218
0 220 5 1 1 219
0 221 7 5 2 22891 25541
0 222 5 1 1 26458
0 223 7 3 2 24830 23595
0 224 5 1 1 26463
0 225 7 5 2 222 224
0 226 7 1 2 22430 127
0 227 5 1 1 226
0 228 7 10 2 24891 25542
0 229 5 2 1 26471
0 230 7 1 2 227 26481
0 231 7 2 2 26466 230
0 232 7 1 2 22355 26483
0 233 5 1 1 232
0 234 7 10 2 24359 24432
0 235 7 1 2 26485 26443
0 236 5 1 1 235
0 237 7 1 2 233 236
0 238 5 1 1 237
0 239 7 1 2 25832 238
0 240 5 1 1 239
0 241 7 8 2 24772 22892
0 242 7 6 2 24303 26495
0 243 5 1 1 26503
0 244 7 1 2 26367 26434
0 245 7 1 2 26504 244
0 246 5 1 1 245
0 247 7 1 2 240 246
0 248 5 1 1 247
0 249 7 2 2 23706 248
0 250 7 6 2 23243 26250
0 251 7 48 2 24137 24636
0 252 5 1 1 26517
0 253 7 19 2 23333 25362
0 254 7 3 2 26518 26565
0 255 5 1 1 26584
0 256 7 2 2 26511 26585
0 257 7 1 2 26509 26587
0 258 5 1 1 257
0 259 7 1 2 220 258
0 260 5 1 1 259
0 261 7 1 2 25739 260
0 262 5 1 1 261
0 263 7 5 2 22167 23334
0 264 7 2 2 26519 26589
0 265 7 6 2 22727 23396
0 266 7 1 2 26596 26512
0 267 7 2 2 26594 266
0 268 7 1 2 26510 26602
0 269 5 1 1 268
0 270 7 1 2 262 269
0 271 5 1 1 270
0 272 7 1 2 25432 271
0 273 5 1 1 272
0 274 7 1 2 26294 156
0 275 5 2 1 274
0 276 7 1 2 26399 26604
0 277 5 1 1 276
0 278 7 4 2 22117 25543
0 279 7 9 2 24831 22961
0 280 7 1 2 24433 26610
0 281 7 1 2 26606 280
0 282 7 1 2 26282 281
0 283 5 1 1 282
0 284 7 1 2 277 283
0 285 5 1 1 284
0 286 7 1 2 22689 285
0 287 5 1 1 286
0 288 7 5 2 24138 26360
0 289 5 1 1 26619
0 290 7 20 2 24832 25544
0 291 7 2 2 26144 26624
0 292 5 1 1 26644
0 293 7 1 2 26620 26645
0 294 5 1 1 293
0 295 7 1 2 26393 289
0 296 5 1 1 295
0 297 7 34 2 22118 22690
0 298 5 3 1 26646
0 299 7 1 2 26680 26400
0 300 7 1 2 296 299
0 301 5 1 1 300
0 302 7 1 2 294 301
0 303 5 1 1 302
0 304 7 1 2 25199 303
0 305 5 1 1 304
0 306 7 22 2 25121 23244
0 307 5 1 1 26683
0 308 7 2 2 24999 26684
0 309 7 6 2 22588 24637
0 310 7 1 2 26401 26707
0 311 7 1 2 26705 310
0 312 5 1 1 311
0 313 7 1 2 305 312
0 314 5 1 1 313
0 315 7 1 2 25294 314
0 316 5 1 1 315
0 317 7 1 2 287 316
0 318 5 1 1 317
0 319 7 1 2 22356 318
0 320 5 1 1 319
0 321 7 1 2 26647 26283
0 322 5 1 1 321
0 323 7 7 2 25295 26520
0 324 5 1 1 26713
0 325 7 23 2 25122 25200
0 326 5 1 1 26720
0 327 7 3 2 26714 26721
0 328 5 1 1 26743
0 329 7 1 2 322 328
0 330 5 5 1 329
0 331 7 2 2 26746 26444
0 332 7 1 2 26486 26751
0 333 5 1 1 332
0 334 7 1 2 320 333
0 335 5 1 1 334
0 336 7 1 2 25833 335
0 337 5 1 1 336
0 338 7 1 2 26441 26752
0 339 5 1 1 338
0 340 7 1 2 337 339
0 341 5 1 1 340
0 342 7 27 2 22168 22728
0 343 7 31 2 25363 23483
0 344 7 13 2 26753 26780
0 345 5 2 1 26811
0 346 7 2 2 23707 26812
0 347 7 1 2 341 26826
0 348 5 1 1 347
0 349 7 1 2 273 348
0 350 5 1 1 349
0 351 7 1 2 23772 350
0 352 5 1 1 351
0 353 7 4 2 23245 23397
0 354 7 6 2 23335 25433
0 355 7 3 2 26828 26832
0 356 7 1 2 24551 26027
0 357 7 1 2 26838 356
0 358 5 1 1 357
0 359 7 3 2 25296 26781
0 360 7 3 2 26722 26841
0 361 5 1 1 26844
0 362 7 1 2 358 361
0 363 5 1 1 362
0 364 7 1 2 26754 363
0 365 5 1 1 364
0 366 7 4 2 23246 26566
0 367 7 1 2 26251 26847
0 368 5 3 1 367
0 369 7 12 2 25297 23398
0 370 7 2 2 26723 26854
0 371 5 1 1 26866
0 372 7 1 2 26851 371
0 373 5 6 1 372
0 374 7 4 2 24666 25434
0 375 7 5 2 24182 22962
0 376 7 1 2 26874 26878
0 377 7 1 2 26868 376
0 378 5 1 1 377
0 379 7 1 2 365 378
0 380 5 1 1 379
0 381 7 1 2 24139 380
0 382 5 1 1 381
0 383 7 6 2 22589 26685
0 384 5 5 1 26883
0 385 7 6 2 25201 26252
0 386 7 1 2 24892 26894
0 387 5 1 1 386
0 388 7 1 2 26889 387
0 389 5 3 1 388
0 390 7 17 2 25364 26755
0 391 7 11 2 25298 23484
0 392 7 4 2 26903 26920
0 393 7 1 2 25000 26931
0 394 7 1 2 26900 393
0 395 5 1 1 394
0 396 7 1 2 382 395
0 397 5 1 1 396
0 398 7 1 2 24638 397
0 399 5 1 1 398
0 400 7 1 2 26813 26605
0 401 5 1 1 400
0 402 7 3 2 24667 26284
0 403 7 9 2 22963 25435
0 404 7 5 2 22119 24183
0 405 7 2 2 23399 26947
0 406 7 1 2 26938 26952
0 407 7 1 2 26935 406
0 408 5 1 1 407
0 409 7 1 2 401 408
0 410 5 1 1 409
0 411 7 1 2 22691 410
0 412 5 1 1 411
0 413 7 20 2 25001 23159
0 414 5 3 1 26954
0 415 7 6 2 24893 26955
0 416 5 3 1 26977
0 417 7 4 2 24552 25202
0 418 7 2 2 24140 26986
0 419 7 1 2 26978 26990
0 420 7 1 2 26932 419
0 421 5 1 1 420
0 422 7 1 2 412 421
0 423 7 1 2 399 422
0 424 5 1 1 423
0 425 7 1 2 24434 424
0 426 5 1 1 425
0 427 7 2 2 22692 25002
0 428 7 1 2 26276 26992
0 429 5 1 1 428
0 430 7 3 2 24639 23247
0 431 5 1 1 26994
0 432 7 4 2 22693 25203
0 433 5 2 1 26997
0 434 7 3 2 431 27001
0 435 7 1 2 24141 27003
0 436 5 1 1 435
0 437 7 4 2 25003 23248
0 438 7 1 2 26708 27006
0 439 5 1 1 438
0 440 7 1 2 436 439
0 441 5 1 1 440
0 442 7 1 2 25299 441
0 443 5 1 1 442
0 444 7 15 2 22590 25004
0 445 7 1 2 23336 27010
0 446 7 1 2 26998 445
0 447 5 1 1 446
0 448 7 1 2 443 447
0 449 5 1 1 448
0 450 7 1 2 25123 449
0 451 5 1 1 450
0 452 7 1 2 429 451
0 453 5 1 1 452
0 454 7 1 2 22964 26814
0 455 7 1 2 453 454
0 456 5 1 1 455
0 457 7 1 2 426 456
0 458 5 1 1 457
0 459 7 1 2 26346 458
0 460 5 1 1 459
0 461 7 13 2 23400 25545
0 462 5 1 1 27025
0 463 7 7 2 25436 25640
0 464 7 3 2 27026 27038
0 465 7 4 2 23337 27045
0 466 7 1 2 24435 25204
0 467 7 1 2 26648 466
0 468 7 3 2 26 25124
0 469 5 1 1 27052
0 470 7 8 2 24553 25005
0 471 7 1 2 27053 27055
0 472 7 1 2 467 471
0 473 7 8 2 24668 24773
0 474 7 3 2 24184 27063
0 475 7 2 2 26611 25782
0 476 7 1 2 27071 27074
0 477 7 1 2 472 476
0 478 7 1 2 27048 477
0 479 5 1 1 478
0 480 7 1 2 460 479
0 481 7 1 2 352 480
0 482 5 1 1 481
0 483 7 1 2 23892 482
0 484 5 1 1 483
0 485 7 2 2 26347 26815
0 486 7 4 2 24640 25300
0 487 7 4 2 24142 27078
0 488 5 1 1 27082
0 489 7 6 2 22694 23338
0 490 7 6 2 22120 27086
0 491 5 2 1 27092
0 492 7 1 2 488 27098
0 493 5 14 1 492
0 494 7 1 2 24554 27100
0 495 5 1 1 494
0 496 7 44 2 23773 24436
0 497 5 45 1 27114
0 498 7 12 2 22965 27115
0 499 5 8 1 27203
0 500 7 1 2 27087 27011
0 501 5 1 1 500
0 502 7 1 2 324 501
0 503 5 1 1 502
0 504 7 1 2 27204 503
0 505 5 1 1 504
0 506 7 1 2 495 505
0 507 5 1 1 506
0 508 7 1 2 25125 507
0 509 5 1 1 508
0 510 7 1 2 24894 26715
0 511 5 1 1 510
0 512 7 1 2 27099 511
0 513 5 1 1 512
0 514 7 1 2 26956 513
0 515 5 1 1 514
0 516 7 1 2 509 515
0 517 5 1 1 516
0 518 7 1 2 25205 517
0 519 5 1 1 518
0 520 7 2 2 24555 26957
0 521 5 1 1 27223
0 522 7 1 2 26291 521
0 523 5 1 1 522
0 524 7 1 2 22695 523
0 525 5 1 1 524
0 526 7 2 2 26361 27012
0 527 5 1 1 27225
0 528 7 1 2 525 527
0 529 5 2 1 528
0 530 7 1 2 26009 27205
0 531 7 1 2 27227 530
0 532 5 1 1 531
0 533 7 1 2 519 532
0 534 5 1 1 533
0 535 7 1 2 27076 534
0 536 5 1 1 535
0 537 7 11 2 24895 23160
0 538 7 1 2 22591 27229
0 539 5 3 1 538
0 540 7 8 2 24556 25126
0 541 5 2 1 27243
0 542 7 2 2 22431 27244
0 543 5 1 1 27253
0 544 7 1 2 27240 543
0 545 5 1 1 544
0 546 7 1 2 21756 545
0 547 5 2 1 546
0 548 7 14 2 22966 25127
0 549 5 1 1 27257
0 550 7 3 2 27258 27116
0 551 5 1 1 27271
0 552 7 18 2 22432 24896
0 553 5 28 1 27274
0 554 7 1 2 23161 27275
0 555 5 1 1 554
0 556 7 1 2 551 555
0 557 5 1 1 556
0 558 7 1 2 22592 557
0 559 5 1 1 558
0 560 7 1 2 27255 559
0 561 5 1 1 560
0 562 7 4 2 24360 26625
0 563 7 1 2 561 27320
0 564 5 1 1 563
0 565 7 7 2 24557 22967
0 566 5 3 1 27324
0 567 7 3 2 23774 27292
0 568 5 3 1 27334
0 569 7 4 2 26162 27337
0 570 5 14 1 27340
0 571 7 5 2 27331 27344
0 572 7 3 2 25128 23596
0 573 7 1 2 25895 27363
0 574 7 1 2 27358 573
0 575 5 1 1 574
0 576 7 1 2 564 575
0 577 5 1 1 576
0 578 7 1 2 25641 577
0 579 5 1 1 578
0 580 7 3 2 21757 27276
0 581 5 18 1 27366
0 582 7 3 2 25129 26192
0 583 7 24 2 25546 23708
0 584 7 1 2 27387 27390
0 585 7 1 2 27369 584
0 586 5 1 1 585
0 587 7 1 2 579 586
0 588 5 1 1 587
0 589 7 1 2 26047 588
0 590 5 1 1 589
0 591 7 60 2 21758 22433
0 592 5 65 1 27414
0 593 7 5 2 22593 24833
0 594 7 6 2 24361 25642
0 595 7 3 2 27539 27544
0 596 7 1 2 26235 27550
0 597 5 1 1 596
0 598 7 14 2 25547 25896
0 599 7 1 2 23709 27553
0 600 5 1 1 599
0 601 7 1 2 597 600
0 602 5 1 1 601
0 603 7 1 2 27474 602
0 604 5 1 1 603
0 605 7 4 2 23775 26487
0 606 7 5 2 24834 24897
0 607 7 4 2 25643 27571
0 608 7 2 2 27567 27576
0 609 5 1 1 27580
0 610 7 1 2 23597 27581
0 611 5 1 1 610
0 612 7 1 2 23710 26372
0 613 5 1 1 612
0 614 7 1 2 611 613
0 615 7 1 2 604 614
0 616 5 1 1 615
0 617 7 1 2 25130 25834
0 618 7 1 2 616 617
0 619 5 1 1 618
0 620 7 1 2 590 619
0 621 5 1 1 620
0 622 7 1 2 25797 621
0 623 5 1 1 622
0 624 7 18 2 23598 25644
0 625 7 15 2 26048 27582
0 626 7 1 2 27345 27600
0 627 5 1 1 626
0 628 7 13 2 25835 27391
0 629 5 4 1 27615
0 630 7 1 2 27293 27616
0 631 5 2 1 630
0 632 7 3 2 23776 22283
0 633 7 3 2 22824 27634
0 634 7 2 2 27392 27637
0 635 5 1 1 27640
0 636 7 1 2 27632 635
0 637 7 1 2 627 636
0 638 5 2 1 637
0 639 7 1 2 25897 27642
0 640 5 2 1 639
0 641 7 5 2 24304 22357
0 642 7 2 2 24774 27646
0 643 7 4 2 22893 27393
0 644 7 7 2 27651 27653
0 645 5 5 1 27657
0 646 7 1 2 27294 27658
0 647 5 2 1 646
0 648 7 6 2 22284 24362
0 649 7 8 2 22825 24835
0 650 7 13 2 27671 27677
0 651 5 1 1 27685
0 652 7 4 2 23599 27686
0 653 5 1 1 27698
0 654 7 2 2 23777 27699
0 655 5 1 1 27702
0 656 7 1 2 25645 27295
0 657 7 1 2 27703 656
0 658 5 1 1 657
0 659 7 2 2 27669 658
0 660 7 15 2 23600 25836
0 661 5 4 1 27706
0 662 7 19 2 25646 26103
0 663 7 2 2 26145 27725
0 664 5 1 1 27744
0 665 7 46 2 23711 26193
0 666 5 3 1 27746
0 667 7 1 2 664 27792
0 668 5 2 1 667
0 669 7 1 2 27707 27795
0 670 5 1 1 669
0 671 7 1 2 23778 27659
0 672 5 1 1 671
0 673 7 1 2 670 672
0 674 7 1 2 27704 673
0 675 7 1 2 27644 674
0 676 5 2 1 675
0 677 7 1 2 26277 27797
0 678 5 1 1 677
0 679 7 1 2 623 678
0 680 5 1 1 679
0 681 7 1 2 26649 680
0 682 5 1 1 681
0 683 7 3 2 22594 22968
0 684 5 1 1 27799
0 685 7 1 2 27601 27800
0 686 5 1 1 685
0 687 7 1 2 27628 686
0 688 5 1 1 687
0 689 7 1 2 27475 688
0 690 5 1 1 689
0 691 7 2 2 22969 27617
0 692 5 1 1 27802
0 693 7 3 2 24898 27583
0 694 7 3 2 26049 27804
0 695 5 1 1 27807
0 696 7 1 2 27117 27808
0 697 5 1 1 696
0 698 7 1 2 692 697
0 699 7 1 2 690 698
0 700 5 2 1 699
0 701 7 1 2 25898 27810
0 702 5 2 1 701
0 703 7 13 2 22894 23712
0 704 7 21 2 22358 27814
0 705 5 3 1 27827
0 706 7 1 2 609 27848
0 707 5 1 1 706
0 708 7 1 2 27708 707
0 709 5 1 1 708
0 710 7 3 2 27672 27584
0 711 7 7 2 22970 27476
0 712 5 4 1 27854
0 713 7 1 2 22826 27540
0 714 7 1 2 27855 713
0 715 7 1 2 27851 714
0 716 5 1 1 715
0 717 7 1 2 27370 27660
0 718 5 1 1 717
0 719 7 1 2 716 718
0 720 7 1 2 709 719
0 721 7 1 2 27812 720
0 722 5 1 1 721
0 723 7 1 2 26744 722
0 724 5 1 1 723
0 725 7 1 2 682 724
0 726 5 1 1 725
0 727 7 1 2 25740 726
0 728 5 1 1 727
0 729 7 11 2 22827 23601
0 730 7 11 2 22285 27865
0 731 5 6 1 27876
0 732 7 21 2 25548 26050
0 733 7 1 2 23779 27893
0 734 5 1 1 733
0 735 7 1 2 27887 734
0 736 5 1 1 735
0 737 7 1 2 27796 736
0 738 5 1 1 737
0 739 7 1 2 27705 738
0 740 7 1 2 27645 739
0 741 5 2 1 740
0 742 7 1 2 24558 27914
0 743 5 1 1 742
0 744 7 3 2 22286 22895
0 745 7 2 2 27916 27866
0 746 7 2 2 23780 22359
0 747 7 1 2 26146 27921
0 748 7 2 2 27919 747
0 749 5 1 1 27923
0 750 7 1 2 23713 27924
0 751 5 1 1 750
0 752 7 1 2 743 751
0 753 5 1 1 752
0 754 7 8 2 23249 23339
0 755 7 5 2 23162 27925
0 756 5 1 1 27933
0 757 7 4 2 22169 24641
0 758 7 7 2 24143 27938
0 759 5 1 1 27942
0 760 7 5 2 22729 27943
0 761 5 1 1 27949
0 762 7 1 2 27934 27950
0 763 7 1 2 753 762
0 764 5 1 1 763
0 765 7 1 2 728 764
0 766 5 1 1 765
0 767 7 1 2 23401 766
0 768 5 1 1 767
0 769 7 15 2 23163 23250
0 770 7 6 2 26567 27954
0 771 5 1 1 27969
0 772 7 5 2 24185 24559
0 773 7 1 2 24669 26521
0 774 7 1 2 27975 773
0 775 7 1 2 27970 774
0 776 7 1 2 27798 775
0 777 5 1 1 776
0 778 7 1 2 768 777
0 779 5 1 1 778
0 780 7 1 2 25437 779
0 781 5 1 1 780
0 782 7 4 2 22828 27673
0 783 7 3 2 27572 27585
0 784 7 2 2 27980 27984
0 785 7 1 2 24437 27987
0 786 5 1 1 785
0 787 7 1 2 27664 786
0 788 5 1 1 787
0 789 7 1 2 23781 788
0 790 5 1 1 789
0 791 7 3 2 24305 24438
0 792 7 6 2 24775 25549
0 793 7 2 2 27989 27992
0 794 5 1 1 27998
0 795 7 1 2 27888 794
0 796 5 1 1 795
0 797 7 3 2 24363 22595
0 798 7 2 2 23782 28000
0 799 7 2 2 25647 26612
0 800 7 1 2 28003 28005
0 801 5 1 1 800
0 802 7 1 2 27793 801
0 803 5 1 1 802
0 804 7 1 2 796 803
0 805 5 1 1 804
0 806 7 3 2 24439 22596
0 807 7 6 2 22287 23602
0 808 7 2 2 27545 27678
0 809 7 7 2 28010 28016
0 810 5 1 1 28018
0 811 7 1 2 28007 28019
0 812 5 1 1 811
0 813 7 1 2 27665 812
0 814 5 1 1 813
0 815 7 1 2 22971 814
0 816 5 1 1 815
0 817 7 1 2 805 816
0 818 7 1 2 790 817
0 819 7 1 2 27813 818
0 820 5 1 1 819
0 821 7 1 2 27101 820
0 822 5 1 1 821
0 823 7 3 2 22896 22972
0 824 7 3 2 22829 28025
0 825 7 1 2 24144 27635
0 826 7 2 2 28028 825
0 827 7 5 2 23603 23714
0 828 7 4 2 22360 28033
0 829 7 7 2 24440 24560
0 830 5 1 1 28042
0 831 7 1 2 25301 28043
0 832 7 1 2 28038 831
0 833 7 1 2 28031 832
0 834 5 1 1 833
0 835 7 1 2 822 834
0 836 5 1 1 835
0 837 7 1 2 25131 836
0 838 5 1 1 837
0 839 7 2 2 24441 22696
0 840 7 7 2 23164 25302
0 841 7 1 2 28049 28051
0 842 7 1 2 28039 841
0 843 7 1 2 28032 842
0 844 5 1 1 843
0 845 7 1 2 838 844
0 846 5 1 1 845
0 847 7 1 2 25206 846
0 848 5 1 1 847
0 849 7 5 2 25303 26650
0 850 7 1 2 26513 28058
0 851 7 1 2 27915 850
0 852 5 1 1 851
0 853 7 1 2 848 852
0 854 5 1 1 853
0 855 7 1 2 26816 854
0 856 5 1 1 855
0 857 7 1 2 781 856
0 858 5 1 1 857
0 859 7 1 2 23893 858
0 860 5 1 1 859
0 861 7 1 2 27118 25999
0 862 5 1 1 861
0 863 7 2 2 24561 25783
0 864 7 6 2 24836 25648
0 865 7 4 2 21855 24776
0 866 7 1 2 28065 28071
0 867 7 1 2 28063 866
0 868 5 1 1 867
0 869 7 1 2 862 868
0 870 5 1 1 869
0 871 7 1 2 25132 870
0 872 5 1 1 871
0 873 7 3 2 24777 23165
0 874 7 5 2 24306 27415
0 875 7 1 2 28075 28078
0 876 7 1 2 27551 875
0 877 5 1 1 876
0 878 7 1 2 872 877
0 879 5 1 1 878
0 880 7 1 2 25798 879
0 881 5 1 1 880
0 882 7 3 2 25304 27955
0 883 7 5 2 23783 28044
0 884 5 2 1 28086
0 885 7 1 2 28083 28087
0 886 7 1 2 26000 885
0 887 5 1 1 886
0 888 7 1 2 881 887
0 889 5 1 1 888
0 890 7 1 2 25550 889
0 891 5 1 1 890
0 892 7 1 2 26348 27477
0 893 7 1 2 26285 892
0 894 5 1 1 893
0 895 7 1 2 891 894
0 896 5 1 1 895
0 897 7 1 2 26651 896
0 898 5 1 1 897
0 899 7 3 2 25551 27158
0 900 5 1 1 28093
0 901 7 1 2 27478 26467
0 902 7 2 2 900 901
0 903 7 1 2 22361 28096
0 904 5 1 1 903
0 905 7 1 2 26459 27568
0 906 5 1 1 905
0 907 7 1 2 904 906
0 908 5 1 1 907
0 909 7 1 2 25837 908
0 910 5 1 1 909
0 911 7 2 2 23784 26435
0 912 7 2 2 26051 26460
0 913 7 1 2 28098 28100
0 914 5 1 1 913
0 915 7 1 2 910 914
0 916 5 1 1 915
0 917 7 2 2 23715 916
0 918 7 1 2 26745 28102
0 919 5 1 1 918
0 920 7 1 2 898 919
0 921 5 1 1 920
0 922 7 1 2 23402 921
0 923 5 1 1 922
0 924 7 1 2 26588 28103
0 925 5 1 1 924
0 926 7 1 2 923 925
0 927 5 1 1 926
0 928 7 1 2 25741 927
0 929 5 1 1 928
0 930 7 8 2 25838 26335
0 931 5 2 1 28104
0 932 7 18 2 25552 25980
0 933 7 1 2 27119 28114
0 934 5 1 1 933
0 935 7 1 2 28112 934
0 936 5 2 1 935
0 937 7 1 2 23716 26603
0 938 7 1 2 28132 937
0 939 5 1 1 938
0 940 7 1 2 929 939
0 941 5 1 1 940
0 942 7 1 2 25438 941
0 943 5 1 1 942
0 944 7 1 2 26747 26827
0 945 7 1 2 28133 944
0 946 5 1 1 945
0 947 7 1 2 943 946
0 948 5 1 1 947
0 949 7 1 2 22973 948
0 950 5 1 1 949
0 951 7 12 2 23403 25742
0 952 7 3 2 24442 25439
0 953 5 1 1 28146
0 954 7 1 2 28134 28147
0 955 5 1 1 954
0 956 7 1 2 26824 955
0 957 5 1 1 956
0 958 7 1 2 23785 957
0 959 5 3 1 958
0 960 7 2 2 24443 26817
0 961 5 1 1 28152
0 962 7 1 2 28149 961
0 963 5 1 1 962
0 964 7 1 2 26748 963
0 965 5 1 1 964
0 966 7 2 2 24642 23340
0 967 7 2 2 24145 28154
0 968 7 5 2 23251 25440
0 969 7 1 2 26253 28158
0 970 7 3 2 28156 969
0 971 7 3 2 22170 26597
0 972 5 2 1 28166
0 973 7 13 2 24670 25365
0 974 5 1 1 28171
0 975 7 6 2 24186 28172
0 976 5 1 1 28184
0 977 7 1 2 24444 28185
0 978 5 1 1 977
0 979 7 1 2 28169 978
0 980 5 2 1 979
0 981 7 1 2 23786 28190
0 982 5 1 1 981
0 983 7 1 2 24445 28167
0 984 5 1 1 983
0 985 7 1 2 982 984
0 986 5 1 1 985
0 987 7 1 2 28163 986
0 988 5 1 1 987
0 989 7 1 2 965 988
0 990 5 1 1 989
0 991 7 1 2 26349 990
0 992 5 1 1 991
0 993 7 1 2 950 992
0 994 7 1 2 860 993
0 995 5 1 1 994
0 996 7 1 2 23034 995
0 997 5 1 1 996
0 998 7 1 2 536 997
0 999 7 1 2 484 998
0 1000 5 1 1 999
0 1001 7 1 2 24489 1000
0 1002 5 1 1 1001
0 1003 7 2 2 21856 26163
0 1004 5 8 1 28192
0 1005 7 2 2 23894 27296
0 1006 5 2 1 28202
0 1007 7 2 2 21759 28204
0 1008 5 2 1 28206
0 1009 7 18 2 28194 28208
0 1010 5 3 1 28210
0 1011 7 3 2 22697 24671
0 1012 7 2 2 26948 28231
0 1013 5 1 1 28234
0 1014 7 6 2 22494 25133
0 1015 7 1 2 28236 26987
0 1016 7 1 2 26140 1015
0 1017 7 1 2 28235 1016
0 1018 7 1 2 27049 1017
0 1019 5 1 1 1018
0 1020 7 1 2 26782 26749
0 1021 5 1 1 1020
0 1022 7 1 2 23404 28164
0 1023 5 1 1 1022
0 1024 7 1 2 1021 1023
0 1025 5 1 1 1024
0 1026 7 4 2 22288 22730
0 1027 7 3 2 22171 22362
0 1028 7 3 2 28242 28246
0 1029 7 12 2 22830 22897
0 1030 7 1 2 28034 28252
0 1031 7 1 2 28249 1030
0 1032 7 1 2 1025 1031
0 1033 5 1 1 1032
0 1034 7 1 2 1019 1033
0 1035 5 1 1 1034
0 1036 7 1 2 28211 1035
0 1037 5 1 1 1036
0 1038 7 6 2 24187 22289
0 1039 7 6 2 22363 24672
0 1040 7 5 2 28264 28270
0 1041 7 27 2 23405 25441
0 1042 5 1 1 28281
0 1043 7 6 2 23604 28282
0 1044 7 2 2 28253 28308
0 1045 7 2 2 28276 28314
0 1046 5 1 1 28316
0 1047 7 8 2 25442 28135
0 1048 5 1 1 28318
0 1049 7 1 2 26825 1048
0 1050 5 4 1 1049
0 1051 7 1 2 24446 28326
0 1052 7 1 2 28115 1051
0 1053 5 1 1 1052
0 1054 7 1 2 1046 1053
0 1055 5 1 1 1054
0 1056 7 2 2 23787 1055
0 1057 5 1 1 28330
0 1058 7 1 2 24447 28317
0 1059 5 2 1 1058
0 1060 7 1 2 24899 28332
0 1061 5 1 1 1060
0 1062 7 1 2 28331 1061
0 1063 5 1 1 1062
0 1064 7 2 2 28309 28029
0 1065 7 1 2 24448 28277
0 1066 7 1 2 28334 1065
0 1067 5 1 1 1066
0 1068 7 1 2 1063 1067
0 1069 5 1 1 1068
0 1070 7 1 2 26750 1069
0 1071 5 1 1 1070
0 1072 7 5 2 22898 25366
0 1073 7 3 2 27867 28336
0 1074 7 1 2 28278 28341
0 1075 5 1 1 1074
0 1076 7 1 2 28170 976
0 1077 5 9 1 1076
0 1078 7 1 2 26368 28344
0 1079 7 1 2 25981 1078
0 1080 5 1 1 1079
0 1081 7 1 2 1075 1080
0 1082 5 1 1 1081
0 1083 7 1 2 27120 1082
0 1084 5 1 1 1083
0 1085 7 5 2 24673 28265
0 1086 7 8 2 22974 25367
0 1087 5 1 1 28358
0 1088 7 2 2 27868 28359
0 1089 7 1 2 26194 28366
0 1090 7 1 2 28353 1089
0 1091 5 1 1 1090
0 1092 7 1 2 1084 1091
0 1093 5 1 1 1092
0 1094 7 1 2 28165 27479
0 1095 7 1 2 1093 1094
0 1096 5 1 1 1095
0 1097 7 1 2 1071 1096
0 1098 5 1 1 1097
0 1099 7 1 2 23895 23717
0 1100 7 1 2 1098 1099
0 1101 5 1 1 1100
0 1102 7 1 2 1037 1101
0 1103 5 1 1 1102
0 1104 7 1 2 23035 1103
0 1105 5 1 1 1104
0 1106 7 3 2 22121 23166
0 1107 5 1 1 28368
0 1108 7 4 2 28035 26783
0 1109 7 5 2 22364 22831
0 1110 7 2 2 28375 27917
0 1111 7 2 2 28371 28380
0 1112 7 1 2 26756 28382
0 1113 5 1 1 1112
0 1114 7 3 2 22597 24674
0 1115 7 1 2 24778 28384
0 1116 7 1 2 26613 26488
0 1117 7 1 2 1115 1116
0 1118 7 8 2 24188 24307
0 1119 7 2 2 23788 28387
0 1120 7 1 2 28395 27046
0 1121 7 1 2 1117 1120
0 1122 5 1 1 1121
0 1123 7 1 2 1113 1122
0 1124 5 1 1 1123
0 1125 7 1 2 23896 1124
0 1126 5 1 1 1125
0 1127 7 3 2 24900 28283
0 1128 7 3 2 23789 24675
0 1129 7 2 2 24189 24449
0 1130 7 3 2 28400 28403
0 1131 7 1 2 28397 28405
0 1132 5 1 1 1131
0 1133 7 8 2 21760 24901
0 1134 5 3 1 28408
0 1135 7 8 2 22434 28409
0 1136 5 6 1 28419
0 1137 7 2 2 26904 28427
0 1138 7 1 2 23485 28433
0 1139 5 1 1 1138
0 1140 7 1 2 1132 1139
0 1141 5 1 1 1140
0 1142 7 1 2 1141 26350
0 1143 5 1 1 1142
0 1144 7 1 2 1126 1143
0 1145 5 1 1 1144
0 1146 7 1 2 28369 1145
0 1147 5 1 1 1146
0 1148 7 6 2 22365 22598
0 1149 7 1 2 27259 28254
0 1150 7 1 2 28435 1149
0 1151 7 15 2 23790 23897
0 1152 7 6 2 24450 28441
0 1153 5 3 1 28456
0 1154 7 5 2 22172 28243
0 1155 7 1 2 28372 28465
0 1156 7 1 2 28457 1155
0 1157 7 1 2 1150 1156
0 1158 5 1 1 1157
0 1159 7 1 2 1147 1158
0 1160 5 1 1 1159
0 1161 7 1 2 25006 1160
0 1162 5 1 1 1161
0 1163 7 2 2 21857 27277
0 1164 5 3 1 28470
0 1165 7 1 2 26818 28472
0 1166 5 1 1 1165
0 1167 7 1 2 28150 1166
0 1168 5 1 1 1167
0 1169 7 2 2 22122 27245
0 1170 7 1 2 26351 28475
0 1171 7 1 2 1168 1170
0 1172 5 1 1 1171
0 1173 7 1 2 1162 1172
0 1174 5 1 1 1173
0 1175 7 1 2 27088 1174
0 1176 5 1 1 1175
0 1177 7 1 2 27251 26983
0 1178 5 10 1 1177
0 1179 7 4 2 21858 22435
0 1180 5 2 1 28487
0 1181 7 1 2 26819 28491
0 1182 5 1 1 1181
0 1183 7 1 2 28151 1182
0 1184 5 1 1 1183
0 1185 7 1 2 28477 1184
0 1186 5 1 1 1185
0 1187 7 1 2 23898 27272
0 1188 5 3 1 1187
0 1189 7 1 2 26394 28493
0 1190 5 1 1 1189
0 1191 7 1 2 26820 1190
0 1192 5 1 1 1191
0 1193 7 1 2 1186 1192
0 1194 5 1 1 1193
0 1195 7 2 2 22290 23718
0 1196 7 1 2 22832 28496
0 1197 7 1 2 26336 1196
0 1198 7 1 2 26716 1197
0 1199 7 1 2 1194 1198
0 1200 5 1 1 1199
0 1201 7 1 2 1176 1200
0 1202 5 1 1 1201
0 1203 7 1 2 25207 1202
0 1204 5 1 1 1203
0 1205 7 3 2 28442 26147
0 1206 5 4 1 28498
0 1207 7 1 2 27228 28499
0 1208 5 1 1 1207
0 1209 7 5 2 22599 25812
0 1210 7 1 2 26522 28505
0 1211 5 1 1 1210
0 1212 7 1 2 1208 1211
0 1213 5 1 1 1212
0 1214 7 1 2 26010 27077
0 1215 7 1 2 1213 1214
0 1216 5 1 1 1215
0 1217 7 1 2 1204 1216
0 1218 7 1 2 1105 1217
0 1219 7 1 2 1002 1218
0 1220 5 1 1 1219
0 1221 7 1 2 24007 1220
0 1222 5 1 1 1221
0 1223 7 6 2 22173 24676
0 1224 5 1 1 28510
0 1225 7 7 2 24190 22731
0 1226 5 1 1 28516
0 1227 7 2 2 1224 1226
0 1228 5 23 1 28523
0 1229 7 3 2 24146 23406
0 1230 7 2 2 23341 28548
0 1231 7 2 2 25007 27159
0 1232 5 4 1 28553
0 1233 7 4 2 25134 23486
0 1234 7 2 2 27815 28559
0 1235 7 2 2 28555 28563
0 1236 7 1 2 28376 28565
0 1237 5 1 1 1236
0 1238 7 25 2 24779 25443
0 1239 5 1 1 28567
0 1240 7 2 2 22600 27278
0 1241 5 1 1 28592
0 1242 7 1 2 23167 28593
0 1243 5 1 1 1242
0 1244 7 1 2 27256 1243
0 1245 5 1 1 1244
0 1246 7 1 2 27726 1245
0 1247 5 1 1 1246
0 1248 7 6 2 25135 27480
0 1249 7 1 2 27747 28594
0 1250 5 1 1 1249
0 1251 7 1 2 1247 1250
0 1252 5 1 1 1251
0 1253 7 1 2 23036 1252
0 1254 5 1 1 1253
0 1255 7 3 2 24562 25813
0 1256 5 2 1 28600
0 1257 7 3 2 24451 24902
0 1258 5 1 1 28605
0 1259 7 4 2 23791 28606
0 1260 5 2 1 28608
0 1261 7 1 2 27727 28609
0 1262 7 1 2 28601 1261
0 1263 5 1 1 1262
0 1264 7 1 2 1254 1263
0 1265 5 1 1 1264
0 1266 7 1 2 28568 1265
0 1267 5 1 1 1266
0 1268 7 1 2 1237 1267
0 1269 5 1 1 1268
0 1270 7 1 2 24308 1269
0 1271 5 1 1 1270
0 1272 7 8 2 22291 24780
0 1273 5 1 1 28614
0 1274 7 1 2 22366 28615
0 1275 7 1 2 28566 1274
0 1276 5 1 1 1275
0 1277 7 1 2 1271 1276
0 1278 5 1 1 1277
0 1279 7 1 2 25553 1278
0 1280 5 1 1 1279
0 1281 7 8 2 24903 23037
0 1282 7 2 2 27121 28622
0 1283 5 1 1 28630
0 1284 7 1 2 27728 28631
0 1285 5 1 1 1284
0 1286 7 1 2 27828 28556
0 1287 5 1 1 1286
0 1288 7 1 2 1285 1287
0 1289 5 1 1 1288
0 1290 7 21 2 25444 23605
0 1291 5 1 1 28632
0 1292 7 7 2 25839 28633
0 1293 7 1 2 25136 28653
0 1294 7 1 2 1289 1293
0 1295 5 1 1 1294
0 1296 7 1 2 1280 1295
0 1297 5 1 1 1296
0 1298 7 1 2 24643 1297
0 1299 5 1 1 1298
0 1300 7 23 2 23487 25554
0 1301 7 2 2 24781 28660
0 1302 5 1 1 28683
0 1303 7 4 2 22833 28634
0 1304 5 2 1 28685
0 1305 7 1 2 1302 28689
0 1306 5 7 1 1305
0 1307 7 1 2 22292 28691
0 1308 5 3 1 1307
0 1309 7 13 2 24309 22834
0 1310 5 1 1 28701
0 1311 7 1 2 28702 28661
0 1312 5 1 1 1311
0 1313 7 1 2 28698 1312
0 1314 5 12 1 1313
0 1315 7 4 2 22899 24904
0 1316 7 5 2 23719 28726
0 1317 7 3 2 24452 25008
0 1318 7 2 2 23792 28735
0 1319 7 1 2 22367 26254
0 1320 7 1 2 28738 1319
0 1321 7 1 2 28730 1320
0 1322 7 1 2 28714 1321
0 1323 5 1 1 1322
0 1324 7 1 2 1299 1323
0 1325 5 1 1 1324
0 1326 7 1 2 28551 1325
0 1327 5 1 1 1326
0 1328 7 6 2 23038 25555
0 1329 7 3 2 24782 28740
0 1330 7 3 2 22123 24310
0 1331 7 1 2 28746 28749
0 1332 5 1 1 1331
0 1333 7 8 2 25009 23606
0 1334 7 2 2 24905 28752
0 1335 7 5 2 22601 25840
0 1336 7 1 2 28760 28762
0 1337 5 1 1 1336
0 1338 7 1 2 1332 1337
0 1339 5 1 1 1338
0 1340 7 1 2 27481 1339
0 1341 5 1 1 1340
0 1342 7 4 2 22124 23039
0 1343 5 2 1 28767
0 1344 7 1 2 27877 28768
0 1345 5 1 1 1344
0 1346 7 1 2 1341 1345
0 1347 5 1 1 1346
0 1348 7 1 2 23488 1347
0 1349 5 1 1 1348
0 1350 7 4 2 1273 1310
0 1351 5 89 1 28773
0 1352 7 4 2 23607 28777
0 1353 7 4 2 25445 28866
0 1354 5 1 1 28870
0 1355 7 5 2 22602 24906
0 1356 7 3 2 25010 28874
0 1357 7 1 2 27122 28879
0 1358 5 1 1 1357
0 1359 7 1 2 28771 1358
0 1360 5 1 1 1359
0 1361 7 1 2 28871 1360
0 1362 5 1 1 1361
0 1363 7 1 2 1349 1362
0 1364 5 1 1 1363
0 1365 7 1 2 27748 1364
0 1366 5 1 1 1365
0 1367 7 5 2 24453 23040
0 1368 7 5 2 23793 28882
0 1369 5 2 1 28887
0 1370 7 1 2 22125 23489
0 1371 7 1 2 28888 1370
0 1372 7 1 2 27988 1371
0 1373 5 1 1 1372
0 1374 7 1 2 1366 1373
0 1375 5 1 1 1374
0 1376 7 5 2 22698 25368
0 1377 7 4 2 25137 25305
0 1378 7 1 2 28894 28899
0 1379 7 1 2 1375 1378
0 1380 5 1 1 1379
0 1381 7 1 2 1327 1380
0 1382 5 1 1 1381
0 1383 7 1 2 24490 1382
0 1384 5 1 1 1383
0 1385 7 1 2 28383 28059
0 1386 5 1 1 1385
0 1387 7 3 2 22495 25768
0 1388 7 1 2 26523 28064
0 1389 7 1 2 28903 1388
0 1390 7 1 2 27050 1389
0 1391 5 1 1 1390
0 1392 7 1 2 1386 1391
0 1393 5 1 1 1392
0 1394 7 1 2 27482 1393
0 1395 5 1 1 1394
0 1396 7 15 2 23342 23407
0 1397 7 3 2 28906 28662
0 1398 7 1 2 26524 28921
0 1399 5 1 1 1398
0 1400 7 12 2 25369 23608
0 1401 7 3 2 25306 28924
0 1402 7 2 2 26652 28936
0 1403 7 1 2 25446 28939
0 1404 5 1 1 1403
0 1405 7 1 2 1399 1404
0 1406 5 3 1 1405
0 1407 7 1 2 28778 28941
0 1408 5 1 1 1407
0 1409 7 2 2 28284 27709
0 1410 7 1 2 28157 28944
0 1411 5 1 1 1410
0 1412 7 1 2 1408 1411
0 1413 5 1 1 1412
0 1414 7 2 2 24454 1413
0 1415 5 1 1 28946
0 1416 7 1 2 23794 27829
0 1417 7 1 2 28947 1416
0 1418 5 1 1 1417
0 1419 7 1 2 1395 1418
0 1420 5 1 1 1419
0 1421 7 1 2 23041 1420
0 1422 5 1 1 1421
0 1423 7 3 2 22293 22368
0 1424 7 4 2 22126 28948
0 1425 7 2 2 28373 28951
0 1426 7 5 2 22900 25307
0 1427 7 2 2 22699 22835
0 1428 7 1 2 24563 28962
0 1429 7 1 2 28957 1428
0 1430 7 1 2 28955 1429
0 1431 5 1 1 1430
0 1432 7 1 2 1422 1431
0 1433 5 1 1 1432
0 1434 7 1 2 25138 1433
0 1435 5 1 1 1434
0 1436 7 3 2 22700 28255
0 1437 7 1 2 26375 28052
0 1438 7 1 2 28964 1437
0 1439 7 1 2 28956 1438
0 1440 5 1 1 1439
0 1441 7 1 2 1435 1440
0 1442 7 1 2 1384 1441
0 1443 5 1 1 1442
0 1444 7 1 2 23899 1443
0 1445 5 1 1 1444
0 1446 7 31 2 24491 23042
0 1447 5 15 1 28967
0 1448 7 1 2 22603 28998
0 1449 5 5 1 1448
0 1450 7 1 2 25139 29013
0 1451 5 1 1 1450
0 1452 7 1 2 26984 1451
0 1453 5 2 1 1452
0 1454 7 2 2 26784 28060
0 1455 5 1 1 29020
0 1456 7 3 2 27710 29021
0 1457 5 1 1 29022
0 1458 7 1 2 1415 1457
0 1459 5 1 1 1458
0 1460 7 2 2 23795 1459
0 1461 5 1 1 29025
0 1462 7 1 2 29018 29026
0 1463 5 1 1 1462
0 1464 7 1 2 24455 29019
0 1465 5 1 1 1464
0 1466 7 2 2 24492 28478
0 1467 5 1 1 29027
0 1468 7 1 2 26395 1467
0 1469 7 1 2 1465 1468
0 1470 5 1 1 1469
0 1471 7 1 2 29023 1470
0 1472 5 1 1 1471
0 1473 7 1 2 1463 1472
0 1474 5 1 1 1473
0 1475 7 1 2 27749 1474
0 1476 5 1 1 1475
0 1477 7 1 2 1445 1476
0 1478 5 1 1 1477
0 1479 7 1 2 24008 1478
0 1480 5 1 1 1479
0 1481 7 7 2 25447 26052
0 1482 7 3 2 22436 24493
0 1483 7 2 2 23043 29036
0 1484 5 1 1 29039
0 1485 7 2 2 21761 29040
0 1486 5 2 1 29041
0 1487 7 1 2 23168 29042
0 1488 5 1 1 1487
0 1489 7 20 2 23044 25140
0 1490 5 2 1 29045
0 1491 7 3 2 24494 29046
0 1492 5 2 1 29067
0 1493 7 1 2 26974 29070
0 1494 5 1 1 1493
0 1495 7 1 2 28458 1494
0 1496 5 1 1 1495
0 1497 7 1 2 1488 1496
0 1498 5 1 1 1497
0 1499 7 1 2 27552 1498
0 1500 5 1 1 1499
0 1501 7 31 2 22496 25011
0 1502 5 18 1 29072
0 1503 7 5 2 23900 29103
0 1504 5 5 1 29121
0 1505 7 2 2 28999 29126
0 1506 5 4 1 29131
0 1507 7 4 2 25141 29133
0 1508 5 1 1 29137
0 1509 7 5 2 23901 28968
0 1510 5 3 1 29141
0 1511 7 1 2 27160 29146
0 1512 5 1 1 1511
0 1513 7 1 2 27750 1512
0 1514 7 1 2 29138 1513
0 1515 5 1 1 1514
0 1516 7 1 2 1500 1515
0 1517 5 1 1 1516
0 1518 7 1 2 29029 1517
0 1519 5 1 1 1518
0 1520 7 2 2 27483 29134
0 1521 7 1 2 27751 29149
0 1522 5 1 1 1521
0 1523 7 2 2 23902 28066
0 1524 7 6 2 24495 22604
0 1525 7 2 2 23045 29153
0 1526 5 1 1 29159
0 1527 7 1 2 27569 29160
0 1528 7 1 2 29151 1527
0 1529 5 1 1 1528
0 1530 7 1 2 1522 1529
0 1531 5 1 1 1530
0 1532 7 8 2 23490 28779
0 1533 7 1 2 25142 29161
0 1534 7 1 2 1531 1533
0 1535 5 1 1 1534
0 1536 7 1 2 1519 1535
0 1537 5 1 1 1536
0 1538 7 1 2 25556 1537
0 1539 5 1 1 1538
0 1540 7 2 2 27830 29104
0 1541 5 1 1 29169
0 1542 7 3 2 24837 23046
0 1543 7 3 2 27546 29171
0 1544 7 1 2 29154 29174
0 1545 5 1 1 1544
0 1546 7 1 2 1541 1545
0 1547 5 1 1 1546
0 1548 7 1 2 23903 1547
0 1549 5 1 1 1548
0 1550 7 4 2 22901 23047
0 1551 7 3 2 22369 24496
0 1552 7 2 2 29177 29181
0 1553 7 2 2 23720 29184
0 1554 5 1 1 29186
0 1555 7 1 2 1549 1554
0 1556 5 1 1 1555
0 1557 7 1 2 28595 28654
0 1558 7 1 2 1556 1557
0 1559 5 1 1 1558
0 1560 7 1 2 1539 1559
0 1561 5 1 1 1560
0 1562 7 1 2 26525 28907
0 1563 7 1 2 1561 1562
0 1564 5 1 1 1563
0 1565 7 1 2 27123 27894
0 1566 5 1 1 1565
0 1567 7 1 2 27721 1566
0 1568 5 2 1 1567
0 1569 7 1 2 23491 29188
0 1570 5 1 1 1569
0 1571 7 1 2 27484 28872
0 1572 5 1 1 1571
0 1573 7 1 2 1570 1572
0 1574 5 2 1 1573
0 1575 7 1 2 29105 29190
0 1576 5 1 1 1575
0 1577 7 4 2 24311 24497
0 1578 7 1 2 28747 29192
0 1579 5 1 1 1578
0 1580 7 5 2 23609 27124
0 1581 7 2 2 25841 29196
0 1582 5 1 1 29201
0 1583 7 1 2 1579 1582
0 1584 5 1 1 1583
0 1585 7 1 2 23492 1584
0 1586 5 1 1 1585
0 1587 7 1 2 1576 1586
0 1588 5 1 1 1587
0 1589 7 1 2 27752 1588
0 1590 5 1 1 1589
0 1591 7 1 2 25448 28774
0 1592 5 1 1 1591
0 1593 7 1 2 25871 953
0 1594 5 1 1 1593
0 1595 7 1 2 23610 1594
0 1596 7 1 2 1592 1595
0 1597 5 1 1 1596
0 1598 7 1 2 23493 27999
0 1599 5 1 1 1598
0 1600 7 1 2 1597 1599
0 1601 5 1 1 1600
0 1602 7 1 2 23796 1601
0 1603 5 1 1 1602
0 1604 7 22 2 22836 23494
0 1605 5 7 1 29203
0 1606 7 3 2 22294 24456
0 1607 7 2 2 23611 29232
0 1608 7 1 2 29204 29235
0 1609 5 1 1 1608
0 1610 7 1 2 1603 1609
0 1611 5 1 1 1610
0 1612 7 5 2 24498 24838
0 1613 7 3 2 23048 25649
0 1614 7 1 2 28001 29242
0 1615 7 1 2 29237 1614
0 1616 7 1 2 1611 1615
0 1617 5 1 1 1616
0 1618 7 1 2 1590 1617
0 1619 5 1 1 1618
0 1620 7 1 2 23904 1619
0 1621 5 1 1 1620
0 1622 7 1 2 23049 29191
0 1623 5 1 1 1622
0 1624 7 4 2 23797 29233
0 1625 7 10 2 23495 23612
0 1626 7 3 2 22837 29249
0 1627 7 1 2 29245 29259
0 1628 5 1 1 1627
0 1629 7 1 2 1623 1628
0 1630 5 1 1 1629
0 1631 7 1 2 24499 1630
0 1632 5 1 1 1631
0 1633 7 3 2 23050 23613
0 1634 7 3 2 29205 29262
0 1635 7 1 2 29246 29265
0 1636 5 1 1 1635
0 1637 7 1 2 1632 1636
0 1638 5 1 1 1637
0 1639 7 1 2 27753 1638
0 1640 5 1 1 1639
0 1641 7 1 2 1621 1640
0 1642 5 1 1 1641
0 1643 7 4 2 25143 25370
0 1644 7 1 2 28061 29268
0 1645 7 1 2 1642 1644
0 1646 5 1 1 1645
0 1647 7 1 2 1564 1646
0 1648 5 1 1 1647
0 1649 7 1 2 24009 1648
0 1650 5 1 1 1649
0 1651 7 2 2 28952 28965
0 1652 7 1 2 28374 28053
0 1653 7 1 2 29272 1652
0 1654 5 4 1 1653
0 1655 7 2 2 25144 25769
0 1656 7 2 2 27051 29278
0 1657 7 14 2 23905 24010
0 1658 5 2 1 29282
0 1659 7 9 2 24364 24500
0 1660 7 4 2 29283 29298
0 1661 7 1 2 26526 27990
0 1662 7 1 2 29307 1661
0 1663 7 1 2 29280 1662
0 1664 5 1 1 1663
0 1665 7 1 2 29274 1664
0 1666 5 1 1 1665
0 1667 7 1 2 21762 1666
0 1668 5 1 1 1667
0 1669 7 3 2 23906 24147
0 1670 7 5 2 23798 24011
0 1671 7 4 2 29311 29314
0 1672 7 1 2 24312 24644
0 1673 7 1 2 29299 1672
0 1674 7 1 2 29319 1673
0 1675 7 1 2 29281 1674
0 1676 5 1 1 1675
0 1677 7 1 2 29275 1676
0 1678 5 1 1 1677
0 1679 7 1 2 22437 1678
0 1680 5 1 1 1679
0 1681 7 1 2 1668 1680
0 1682 5 1 1 1681
0 1683 7 1 2 25012 1682
0 1684 5 1 1 1683
0 1685 7 4 2 25145 23343
0 1686 7 1 2 29172 29323
0 1687 7 2 2 27047 1686
0 1688 7 3 2 24148 26053
0 1689 7 1 2 24012 24645
0 1690 7 1 2 29300 1689
0 1691 7 1 2 29329 1690
0 1692 7 1 2 29327 1691
0 1693 5 1 1 1692
0 1694 7 1 2 29276 1693
0 1695 5 1 1 1694
0 1696 7 1 2 21859 1695
0 1697 5 1 1 1696
0 1698 7 4 2 24646 24783
0 1699 7 2 2 25784 29332
0 1700 7 3 2 24013 24149
0 1701 7 6 2 21860 27161
0 1702 5 13 1 29341
0 1703 7 1 2 29338 29347
0 1704 7 1 2 29336 1703
0 1705 7 1 2 29328 1704
0 1706 5 1 1 1705
0 1707 7 1 2 29277 1706
0 1708 5 1 1 1707
0 1709 7 1 2 22497 1708
0 1710 5 1 1 1709
0 1711 7 1 2 1697 1710
0 1712 7 1 2 1684 1711
0 1713 5 1 1 1712
0 1714 7 1 2 24564 1713
0 1715 5 1 1 1714
0 1716 7 3 2 22295 23496
0 1717 7 4 2 22127 28895
0 1718 7 2 2 29360 29363
0 1719 7 6 2 25308 23721
0 1720 7 1 2 29068 29369
0 1721 7 2 2 28443 26436
0 1722 7 4 2 23614 28256
0 1723 7 1 2 29375 29377
0 1724 7 1 2 1720 1723
0 1725 7 1 2 29367 1724
0 1726 5 1 1 1725
0 1727 7 1 2 1715 1726
0 1728 7 1 2 1650 1727
0 1729 5 1 1 1728
0 1730 7 1 2 22975 1729
0 1731 5 1 1 1730
0 1732 7 2 2 25309 29250
0 1733 7 1 2 22838 29234
0 1734 7 1 2 29364 1733
0 1735 7 1 2 29381 1734
0 1736 5 1 1 1735
0 1737 7 1 2 1461 1736
0 1738 5 1 1 1737
0 1739 7 1 2 29028 1738
0 1740 5 1 1 1739
0 1741 7 1 2 26392 29024
0 1742 5 1 1 1741
0 1743 7 1 2 1740 1742
0 1744 5 1 1 1743
0 1745 7 1 2 23907 1744
0 1746 5 1 1 1745
0 1747 7 12 2 22976 25013
0 1748 5 2 1 29383
0 1749 7 4 2 22839 25310
0 1750 5 1 1 29397
0 1751 7 1 2 26255 29398
0 1752 7 1 2 29395 1751
0 1753 7 1 2 27416 29073
0 1754 5 3 1 1753
0 1755 7 4 2 23615 29000
0 1756 7 1 2 29401 29404
0 1757 7 1 2 1752 1756
0 1758 7 1 2 29368 1757
0 1759 5 1 1 1758
0 1760 7 1 2 1746 1759
0 1761 5 1 1 1760
0 1762 7 1 2 27754 1761
0 1763 5 1 1 1762
0 1764 7 1 2 1731 1763
0 1765 7 1 2 1480 1764
0 1766 5 1 1 1765
0 1767 7 1 2 25208 1766
0 1768 5 1 1 1767
0 1769 7 8 2 23051 25449
0 1770 7 3 2 24784 29408
0 1771 5 1 1 29416
0 1772 7 13 2 21763 21861
0 1773 5 1 1 29419
0 1774 7 4 2 22498 29420
0 1775 7 5 2 27279 29432
0 1776 7 1 2 29417 29436
0 1777 5 1 1 1776
0 1778 7 28 2 23908 24501
0 1779 5 57 1 29441
0 1780 7 3 2 21764 26035
0 1781 5 4 1 29526
0 1782 7 1 2 29469 29527
0 1783 5 2 1 1782
0 1784 7 6 2 21973 22438
0 1785 7 4 2 29421 29535
0 1786 5 2 1 29541
0 1787 7 1 2 22605 29545
0 1788 5 1 1 1787
0 1789 7 1 2 25014 1788
0 1790 7 1 2 29533 1789
0 1791 5 1 1 1790
0 1792 7 34 2 21862 22499
0 1793 5 30 1 29547
0 1794 7 2 2 24565 29581
0 1795 5 6 1 29611
0 1796 7 13 2 24907 27162
0 1797 5 5 1 29619
0 1798 7 1 2 29613 29620
0 1799 5 1 1 1798
0 1800 7 7 2 22439 22500
0 1801 5 1 1 29637
0 1802 7 11 2 29638 29422
0 1803 5 3 1 29644
0 1804 7 2 2 23052 29655
0 1805 5 1 1 29658
0 1806 7 1 2 1799 29659
0 1807 5 1 1 1806
0 1808 7 1 2 29206 1807
0 1809 7 1 2 1791 1808
0 1810 5 1 1 1809
0 1811 7 1 2 1777 1810
0 1812 5 1 1 1811
0 1813 7 1 2 28940 1812
0 1814 5 1 1 1813
0 1815 7 5 2 23909 24457
0 1816 5 2 1 29660
0 1817 7 4 2 29315 29661
0 1818 7 11 2 24502 29667
0 1819 7 3 2 22701 29671
0 1820 5 1 1 29682
0 1821 7 4 2 24647 27417
0 1822 7 2 2 28623 29548
0 1823 5 1 1 29689
0 1824 7 1 2 29685 29690
0 1825 5 1 1 1824
0 1826 7 1 2 1820 1825
0 1827 5 1 1 1826
0 1828 7 1 2 28552 28692
0 1829 7 1 2 1827 1828
0 1830 5 1 1 1829
0 1831 7 1 2 1814 1830
0 1832 5 1 1 1831
0 1833 7 1 2 22296 1832
0 1834 5 1 1 1833
0 1835 7 11 2 22440 29423
0 1836 5 3 1 29691
0 1837 7 3 2 22501 28624
0 1838 7 1 2 29692 29705
0 1839 7 1 2 28942 1838
0 1840 5 1 1 1839
0 1841 7 1 2 24150 28444
0 1842 7 6 2 24014 24503
0 1843 7 1 2 28050 29708
0 1844 7 1 2 1841 1843
0 1845 7 1 2 28922 1844
0 1846 5 1 1 1845
0 1847 7 1 2 1840 1846
0 1848 5 1 1 1847
0 1849 7 1 2 28703 1848
0 1850 5 1 1 1849
0 1851 7 1 2 1834 1850
0 1852 5 1 1 1851
0 1853 7 1 2 23722 27388
0 1854 7 1 2 1852 1853
0 1855 5 1 1 1854
0 1856 7 3 2 24785 26369
0 1857 7 1 2 23497 29714
0 1858 5 1 1 1857
0 1859 7 1 2 28690 1858
0 1860 5 1 1 1859
0 1861 7 1 2 22297 1860
0 1862 5 1 1 1861
0 1863 7 6 2 24313 25557
0 1864 7 7 2 22977 23498
0 1865 7 4 2 22840 29723
0 1866 5 1 1 29730
0 1867 7 1 2 29717 29731
0 1868 5 1 1 1867
0 1869 7 1 2 1862 1868
0 1870 5 1 1 1869
0 1871 7 1 2 27125 1870
0 1872 5 1 1 1871
0 1873 7 1 2 26939 27711
0 1874 5 1 1 1873
0 1875 7 1 2 1872 1874
0 1876 5 1 1 1875
0 1877 7 1 2 27102 1876
0 1878 5 1 1 1877
0 1879 7 12 2 23799 26148
0 1880 5 13 1 29734
0 1881 7 1 2 22702 28569
0 1882 7 3 2 23344 25558
0 1883 7 1 2 28750 29759
0 1884 7 1 2 1881 1883
0 1885 7 1 2 29735 1884
0 1886 5 1 1 1885
0 1887 7 1 2 1878 1886
0 1888 5 1 1 1887
0 1889 7 1 2 23408 29308
0 1890 7 3 2 23053 27485
0 1891 5 3 1 29762
0 1892 7 4 2 24566 24839
0 1893 7 3 2 25650 29768
0 1894 7 1 2 29763 29772
0 1895 7 1 2 1889 1894
0 1896 7 1 2 1888 1895
0 1897 5 1 1 1896
0 1898 7 11 2 23800 22978
0 1899 5 17 1 29775
0 1900 7 6 2 24458 24504
0 1901 7 3 2 29776 29803
0 1902 5 4 1 29809
0 1903 7 1 2 21974 29812
0 1904 5 1 1 1903
0 1905 7 2 2 28410 29639
0 1906 5 3 1 29816
0 1907 7 4 2 1904 29818
0 1908 5 1 1 29821
0 1909 7 1 2 23910 29822
0 1910 5 1 1 1909
0 1911 7 1 2 22502 29746
0 1912 5 1 1 1911
0 1913 7 4 2 27371 1912
0 1914 5 4 1 29825
0 1915 7 1 2 24015 29826
0 1916 5 1 1 1915
0 1917 7 1 2 1910 1916
0 1918 5 1 1 1917
0 1919 7 1 2 23054 1918
0 1920 5 1 1 1919
0 1921 7 7 2 24505 22979
0 1922 5 4 1 29833
0 1923 7 3 2 29284 29834
0 1924 5 1 1 29844
0 1925 7 2 2 27486 29845
0 1926 5 1 1 29847
0 1927 7 1 2 1920 1926
0 1928 5 1 1 1927
0 1929 7 3 2 24567 23345
0 1930 7 1 2 28285 29849
0 1931 7 1 2 1928 1930
0 1932 5 1 1 1931
0 1933 7 7 2 22441 25015
0 1934 5 1 1 29852
0 1935 7 3 2 21765 29853
0 1936 5 1 1 29859
0 1937 7 2 2 22503 26164
0 1938 5 3 1 29862
0 1939 7 1 2 27338 29863
0 1940 5 1 1 1939
0 1941 7 1 2 1936 1940
0 1942 5 1 1 1941
0 1943 7 1 2 21863 1942
0 1944 5 1 1 1943
0 1945 7 1 2 29402 1944
0 1946 5 1 1 1945
0 1947 7 11 2 25311 25371
0 1948 5 1 1 29867
0 1949 7 3 2 23499 29868
0 1950 7 1 2 22606 29878
0 1951 7 1 2 1946 1950
0 1952 5 1 1 1951
0 1953 7 1 2 1932 1952
0 1954 5 1 1 1953
0 1955 7 1 2 22128 1954
0 1956 5 1 1 1955
0 1957 7 6 2 23346 28286
0 1958 7 16 2 22980 23055
0 1959 5 6 1 29887
0 1960 7 1 2 22607 29903
0 1961 5 3 1 1960
0 1962 7 1 2 24568 26387
0 1963 5 1 1 1962
0 1964 7 1 2 29909 1963
0 1965 7 1 2 29881 1964
0 1966 7 1 2 29672 1965
0 1967 5 1 1 1966
0 1968 7 1 2 1956 1967
0 1969 5 1 1 1968
0 1970 7 1 2 22703 1969
0 1971 5 1 1 1970
0 1972 7 20 2 24016 24569
0 1973 5 3 1 29912
0 1974 7 5 2 25016 29470
0 1975 5 4 1 29935
0 1976 7 2 2 27346 29582
0 1977 5 1 1 29944
0 1978 7 1 2 29940 29945
0 1979 5 1 1 1978
0 1980 7 1 2 29147 1979
0 1981 5 5 1 1980
0 1982 7 2 2 29913 29946
0 1983 5 1 1 29951
0 1984 7 1 2 25312 1983
0 1985 5 1 1 1984
0 1986 7 2 2 28287 26527
0 1987 7 9 2 21864 27418
0 1988 5 4 1 29955
0 1989 7 3 2 22504 28875
0 1990 7 1 2 29956 29968
0 1991 5 1 1 1990
0 1992 7 2 2 23347 1991
0 1993 5 1 1 29971
0 1994 7 1 2 29953 1993
0 1995 7 1 2 1985 1994
0 1996 5 1 1 1995
0 1997 7 1 2 1971 1996
0 1998 5 1 1 1997
0 1999 7 1 2 22841 1998
0 2000 5 1 1 1999
0 2001 7 2 2 28570 29869
0 2002 7 4 2 28411 28488
0 2003 5 3 1 29975
0 2004 7 8 2 22505 22608
0 2005 7 1 2 26653 29982
0 2006 7 1 2 29976 2005
0 2007 7 1 2 29973 2006
0 2008 5 1 1 2007
0 2009 7 1 2 2000 2008
0 2010 5 1 1 2009
0 2011 7 1 2 23616 2010
0 2012 5 1 1 2011
0 2013 7 3 2 24151 26709
0 2014 7 1 2 29645 29990
0 2015 5 1 1 2014
0 2016 7 1 2 27056 29683
0 2017 5 1 1 2016
0 2018 7 1 2 2015 2017
0 2019 5 1 1 2018
0 2020 7 1 2 24908 2019
0 2021 5 1 1 2020
0 2022 7 3 2 22981 29442
0 2023 5 1 1 29993
0 2024 7 2 2 27487 29994
0 2025 5 1 1 29996
0 2026 7 7 2 27163 27861
0 2027 7 1 2 29471 29998
0 2028 5 3 1 2027
0 2029 7 2 2 29583 30005
0 2030 5 1 1 30008
0 2031 7 1 2 23056 30009
0 2032 5 1 1 2031
0 2033 7 1 2 2025 2032
0 2034 5 5 1 2033
0 2035 7 2 2 29914 30010
0 2036 5 1 1 30015
0 2037 7 1 2 26654 30016
0 2038 5 1 1 2037
0 2039 7 1 2 2021 2038
0 2040 5 1 1 2039
0 2041 7 1 2 23348 2040
0 2042 5 1 1 2041
0 2043 7 1 2 27083 29952
0 2044 5 1 1 2043
0 2045 7 1 2 2042 2044
0 2046 5 1 1 2045
0 2047 7 3 2 24786 23409
0 2048 7 2 2 28663 30017
0 2049 7 1 2 2046 30020
0 2050 5 1 1 2049
0 2051 7 1 2 22298 2050
0 2052 7 1 2 2012 2051
0 2053 5 1 1 2052
0 2054 7 1 2 27103 30011
0 2055 5 1 1 2054
0 2056 7 7 2 28445 29804
0 2057 7 1 2 26717 30022
0 2058 5 1 1 2057
0 2059 7 1 2 2055 2058
0 2060 5 1 1 2059
0 2061 7 3 2 23410 28664
0 2062 7 1 2 22842 30029
0 2063 7 1 2 2060 2062
0 2064 5 1 1 2063
0 2065 7 1 2 27297 28969
0 2066 5 2 1 2065
0 2067 7 1 2 21766 30032
0 2068 5 3 1 2067
0 2069 7 4 2 25017 26165
0 2070 5 7 1 30037
0 2071 7 3 2 29864 30041
0 2072 5 1 1 30048
0 2073 7 4 2 29106 30049
0 2074 5 1 1 30051
0 2075 7 1 2 30033 2074
0 2076 5 1 1 2075
0 2077 7 5 2 30034 2076
0 2078 7 1 2 23911 30055
0 2079 5 1 1 2078
0 2080 7 2 2 28970 29736
0 2081 5 1 1 30060
0 2082 7 1 2 2079 2081
0 2083 5 7 1 2082
0 2084 7 3 2 25450 30062
0 2085 7 3 2 25559 30018
0 2086 7 1 2 27104 30072
0 2087 7 1 2 30069 2086
0 2088 5 1 1 2087
0 2089 7 1 2 2064 2088
0 2090 5 1 1 2089
0 2091 7 1 2 29915 2090
0 2092 5 1 1 2091
0 2093 7 8 2 22843 24909
0 2094 7 3 2 29983 29957
0 2095 7 1 2 28943 30083
0 2096 5 1 1 2095
0 2097 7 6 2 24506 24570
0 2098 5 2 1 30086
0 2099 7 1 2 26993 30087
0 2100 7 1 2 28923 2099
0 2101 7 1 2 29668 2100
0 2102 5 1 1 2101
0 2103 7 1 2 2096 2102
0 2104 5 1 1 2103
0 2105 7 1 2 30075 2104
0 2106 5 1 1 2105
0 2107 7 1 2 24314 2106
0 2108 7 1 2 2092 2107
0 2109 5 1 1 2108
0 2110 7 1 2 27755 2109
0 2111 7 1 2 2053 2110
0 2112 5 1 1 2111
0 2113 7 1 2 1897 2112
0 2114 5 1 1 2113
0 2115 7 1 2 23169 2114
0 2116 5 1 1 2115
0 2117 7 1 2 1855 2116
0 2118 5 1 1 2117
0 2119 7 1 2 23252 2118
0 2120 5 1 1 2119
0 2121 7 6 2 23500 27586
0 2122 7 3 2 28908 30094
0 2123 7 9 2 22609 23170
0 2124 5 7 1 30103
0 2125 7 7 2 24910 25146
0 2126 7 4 2 24571 30119
0 2127 5 1 1 30126
0 2128 7 2 2 30112 2127
0 2129 5 5 1 30130
0 2130 7 2 2 22442 30132
0 2131 5 1 1 30137
0 2132 7 3 2 22443 23171
0 2133 7 1 2 29549 30139
0 2134 5 1 1 2133
0 2135 7 1 2 2131 2134
0 2136 5 1 1 2135
0 2137 7 1 2 21767 2136
0 2138 5 1 1 2137
0 2139 7 6 2 26272 26313
0 2140 7 2 2 29472 30142
0 2141 7 1 2 469 29612
0 2142 5 1 1 2141
0 2143 7 1 2 30148 2142
0 2144 5 1 1 2143
0 2145 7 1 2 2138 2144
0 2146 5 1 1 2145
0 2147 7 1 2 25018 2146
0 2148 5 1 1 2147
0 2149 7 2 2 21865 29984
0 2150 7 1 2 23172 30150
0 2151 5 1 1 2150
0 2152 7 5 2 21866 24572
0 2153 7 1 2 28237 30152
0 2154 5 1 1 2153
0 2155 7 3 2 23801 25147
0 2156 5 1 1 30157
0 2157 7 1 2 22444 2156
0 2158 7 1 2 30149 2157
0 2159 5 1 1 2158
0 2160 7 1 2 2154 2159
0 2161 5 1 1 2160
0 2162 7 1 2 24911 2161
0 2163 5 1 1 2162
0 2164 7 1 2 2151 2163
0 2165 7 1 2 2148 2164
0 2166 5 1 1 2165
0 2167 7 1 2 23253 2166
0 2168 5 1 1 2167
0 2169 7 19 2 23173 25209
0 2170 5 1 1 30160
0 2171 7 4 2 24573 30161
0 2172 5 3 1 30179
0 2173 7 2 2 23802 30180
0 2174 5 1 1 30186
0 2175 7 1 2 26890 2174
0 2176 5 4 1 2175
0 2177 7 1 2 22982 30188
0 2178 5 1 1 2177
0 2179 7 3 2 26686 29155
0 2180 5 1 1 30192
0 2181 7 1 2 2178 2180
0 2182 5 2 1 2181
0 2183 7 4 2 23912 25019
0 2184 7 1 2 30195 30197
0 2185 5 1 1 2184
0 2186 7 3 2 22506 29342
0 2187 5 1 1 30201
0 2188 7 1 2 22983 30202
0 2189 5 1 1 2188
0 2190 7 8 2 23913 24912
0 2191 5 3 1 30204
0 2192 7 1 2 22610 30205
0 2193 5 1 1 2192
0 2194 7 1 2 2189 2193
0 2195 5 1 1 2194
0 2196 7 1 2 26687 2195
0 2197 5 1 1 2196
0 2198 7 2 2 30162 30088
0 2199 5 1 1 30215
0 2200 7 10 2 22611 23254
0 2201 5 1 1 30217
0 2202 7 4 2 27260 30218
0 2203 5 3 1 30227
0 2204 7 1 2 2199 30231
0 2205 5 1 1 2204
0 2206 7 1 2 28462 2205
0 2207 5 1 1 2206
0 2208 7 1 2 2197 2207
0 2209 5 1 1 2208
0 2210 7 1 2 23057 2209
0 2211 5 1 1 2210
0 2212 7 1 2 2185 2211
0 2213 7 1 2 2168 2212
0 2214 5 1 1 2213
0 2215 7 1 2 30100 2214
0 2216 5 1 1 2215
0 2217 7 4 2 25148 26447
0 2218 7 17 2 25372 25451
0 2219 7 5 2 27394 30238
0 2220 7 3 2 30234 30255
0 2221 5 1 1 30260
0 2222 7 2 2 27013 30261
0 2223 5 1 1 30263
0 2224 7 7 2 21867 24913
0 2225 5 5 1 30265
0 2226 7 2 2 30266 29640
0 2227 7 1 2 30264 30277
0 2228 5 1 1 2227
0 2229 7 5 2 23411 23617
0 2230 7 5 2 23501 25651
0 2231 7 5 2 30279 30284
0 2232 7 3 2 27926 30289
0 2233 7 1 2 21768 30104
0 2234 5 1 1 2233
0 2235 7 1 2 28603 2234
0 2236 5 1 1 2235
0 2237 7 1 2 29473 2236
0 2238 7 1 2 30294 2237
0 2239 5 1 1 2238
0 2240 7 14 2 25452 25560
0 2241 7 6 2 23723 30297
0 2242 7 1 2 30311 29870
0 2243 7 7 2 25020 25210
0 2244 7 2 2 26297 30317
0 2245 7 1 2 29433 30324
0 2246 7 1 2 2242 2245
0 2247 5 1 1 2246
0 2248 7 1 2 2239 2247
0 2249 5 1 1 2248
0 2250 7 1 2 26166 2249
0 2251 5 1 1 2250
0 2252 7 1 2 2228 2251
0 2253 7 1 2 2216 2252
0 2254 5 1 1 2253
0 2255 7 1 2 26528 2254
0 2256 5 1 1 2255
0 2257 7 1 2 25824 30151
0 2258 5 2 1 2257
0 2259 7 1 2 25149 29904
0 2260 5 3 1 2259
0 2261 7 9 2 26273 30328
0 2262 7 1 2 29474 30331
0 2263 5 1 1 2262
0 2264 7 3 2 26958 29550
0 2265 5 2 1 30340
0 2266 7 1 2 2263 30343
0 2267 5 6 1 2266
0 2268 7 1 2 26011 30345
0 2269 5 1 1 2268
0 2270 7 1 2 30326 2269
0 2271 5 1 1 2270
0 2272 7 1 2 27419 2271
0 2273 5 1 1 2272
0 2274 7 3 2 23174 26012
0 2275 5 1 1 30351
0 2276 7 1 2 26320 2275
0 2277 5 5 1 2276
0 2278 7 3 2 26376 30354
0 2279 7 1 2 30203 30359
0 2280 5 1 1 2279
0 2281 7 1 2 2273 2280
0 2282 5 1 1 2281
0 2283 7 1 2 26655 30256
0 2284 7 1 2 2282 2283
0 2285 5 1 1 2284
0 2286 7 1 2 2256 2285
0 2287 5 1 1 2286
0 2288 7 1 2 28780 2287
0 2289 5 1 1 2288
0 2290 7 1 2 23349 29954
0 2291 5 1 1 2290
0 2292 7 1 2 1455 2291
0 2293 5 3 1 2292
0 2294 7 2 2 23255 30362
0 2295 7 1 2 27280 27602
0 2296 5 1 1 2295
0 2297 7 2 2 26167 27395
0 2298 7 1 2 25842 30367
0 2299 5 1 1 2298
0 2300 7 1 2 2296 2299
0 2301 5 2 1 2300
0 2302 7 1 2 29074 30369
0 2303 5 1 1 2302
0 2304 7 4 2 22445 22612
0 2305 5 1 1 30371
0 2306 7 1 2 27618 30372
0 2307 5 1 1 2306
0 2308 7 1 2 2303 2307
0 2309 5 1 1 2308
0 2310 7 1 2 23175 2309
0 2311 5 1 1 2310
0 2312 7 6 2 25150 29888
0 2313 5 1 1 30375
0 2314 7 1 2 22446 27619
0 2315 7 1 2 30376 2314
0 2316 5 1 1 2315
0 2317 7 1 2 2311 2316
0 2318 5 1 1 2317
0 2319 7 1 2 21769 2318
0 2320 5 1 1 2319
0 2321 7 3 2 22507 25843
0 2322 7 3 2 22447 26377
0 2323 5 5 1 30384
0 2324 7 3 2 23176 23724
0 2325 7 2 2 25561 30392
0 2326 7 1 2 30385 30395
0 2327 7 1 2 30381 2326
0 2328 5 1 1 2327
0 2329 7 1 2 2320 2328
0 2330 5 1 1 2329
0 2331 7 1 2 30365 2330
0 2332 5 1 1 2331
0 2333 7 1 2 21770 30370
0 2334 5 1 1 2333
0 2335 7 1 2 27281 27620
0 2336 5 1 1 2335
0 2337 7 1 2 2334 2336
0 2338 5 3 1 2337
0 2339 7 3 2 25211 25373
0 2340 7 4 2 23502 30400
0 2341 7 2 2 28238 27014
0 2342 7 1 2 30403 30407
0 2343 7 1 2 27105 2342
0 2344 7 1 2 30397 2343
0 2345 5 1 1 2344
0 2346 7 1 2 2332 2345
0 2347 5 1 1 2346
0 2348 7 1 2 21868 2347
0 2349 5 1 1 2348
0 2350 7 1 2 27420 27396
0 2351 7 1 2 30382 2350
0 2352 7 1 2 30332 2351
0 2353 7 1 2 30366 2352
0 2354 5 1 1 2353
0 2355 7 1 2 2349 2354
0 2356 7 1 2 2289 2355
0 2357 5 1 1 2356
0 2358 7 1 2 21975 2357
0 2359 5 1 1 2358
0 2360 7 2 2 25212 27359
0 2361 7 2 2 29709 30409
0 2362 5 1 1 30411
0 2363 7 2 2 29047 30412
0 2364 5 1 1 30413
0 2365 7 1 2 26036 30189
0 2366 5 1 1 2365
0 2367 7 4 2 24914 26688
0 2368 5 1 1 30415
0 2369 7 1 2 28008 30416
0 2370 5 1 1 2369
0 2371 7 3 2 28045 30163
0 2372 5 1 1 30419
0 2373 7 1 2 26891 2372
0 2374 5 2 1 2373
0 2375 7 1 2 28416 29786
0 2376 7 1 2 30422 2375
0 2377 5 1 1 2376
0 2378 7 1 2 2370 2377
0 2379 7 1 2 2366 2378
0 2380 5 2 1 2379
0 2381 7 1 2 29075 30424
0 2382 5 1 1 2381
0 2383 7 1 2 2364 2382
0 2384 5 1 1 2383
0 2385 7 1 2 26529 2384
0 2386 5 1 1 2385
0 2387 7 3 2 24017 23256
0 2388 7 2 2 26256 30426
0 2389 7 1 2 26656 30429
0 2390 7 1 2 30056 2389
0 2391 5 1 1 2390
0 2392 7 1 2 2386 2391
0 2393 5 1 1 2392
0 2394 7 1 2 23914 2393
0 2395 5 1 1 2394
0 2396 7 2 2 26298 27206
0 2397 5 1 1 30431
0 2398 7 1 2 21771 30138
0 2399 5 1 1 2398
0 2400 7 1 2 2397 2399
0 2401 5 1 1 2400
0 2402 7 7 2 21869 29076
0 2403 5 7 1 30433
0 2404 7 1 2 26530 30434
0 2405 7 1 2 2401 2404
0 2406 5 1 1 2405
0 2407 7 4 2 23058 23177
0 2408 5 1 1 30447
0 2409 7 2 2 29737 30448
0 2410 7 2 2 24574 29710
0 2411 5 1 1 30453
0 2412 7 1 2 26657 30454
0 2413 7 1 2 30451 2412
0 2414 5 1 1 2413
0 2415 7 1 2 2406 2414
0 2416 5 1 1 2415
0 2417 7 1 2 23257 2416
0 2418 5 1 1 2417
0 2419 7 2 2 21870 29001
0 2420 5 2 1 30455
0 2421 7 5 2 29107 30457
0 2422 5 2 1 30459
0 2423 7 6 2 30164 29916
0 2424 5 1 1 30466
0 2425 7 1 2 21772 26531
0 2426 7 1 2 30467 2425
0 2427 7 1 2 30464 2426
0 2428 5 1 1 2427
0 2429 7 1 2 2418 2428
0 2430 7 1 2 2395 2429
0 2431 5 1 1 2430
0 2432 7 1 2 23350 2431
0 2433 5 1 1 2432
0 2434 7 2 2 28084 27347
0 2435 7 2 2 26532 29917
0 2436 7 1 2 29142 30474
0 2437 7 1 2 30472 2436
0 2438 5 1 1 2437
0 2439 7 1 2 2433 2438
0 2440 5 1 1 2439
0 2441 7 1 2 30290 2440
0 2442 5 1 1 2441
0 2443 7 2 2 27397 30063
0 2444 7 5 2 24018 22129
0 2445 7 2 2 30239 30478
0 2446 7 1 2 26999 28900
0 2447 7 1 2 30483 2446
0 2448 7 1 2 30476 2447
0 2449 5 1 1 2448
0 2450 7 1 2 2442 2449
0 2451 5 1 1 2450
0 2452 7 1 2 28781 2451
0 2453 5 1 1 2452
0 2454 7 1 2 27643 28971
0 2455 5 1 1 2454
0 2456 7 3 2 22844 22984
0 2457 7 1 2 27398 29108
0 2458 7 1 2 30485 2457
0 2459 7 1 2 29247 2458
0 2460 5 1 1 2459
0 2461 7 1 2 2455 2460
0 2462 5 1 1 2461
0 2463 7 1 2 23915 2462
0 2464 5 1 1 2463
0 2465 7 3 2 26149 27641
0 2466 5 2 1 30488
0 2467 7 1 2 28972 30489
0 2468 5 1 1 2467
0 2469 7 1 2 2464 2468
0 2470 5 1 1 2469
0 2471 7 8 2 24575 27956
0 2472 7 1 2 28288 30493
0 2473 7 1 2 27106 2472
0 2474 7 1 2 2470 2473
0 2475 5 1 1 2474
0 2476 7 1 2 23059 27811
0 2477 5 1 1 2476
0 2478 7 1 2 30491 2477
0 2479 5 1 1 2478
0 2480 7 1 2 24507 2479
0 2481 5 1 1 2480
0 2482 7 1 2 27803 28889
0 2483 5 1 1 2482
0 2484 7 1 2 2481 2483
0 2485 5 1 1 2484
0 2486 7 1 2 23916 2485
0 2487 5 1 1 2486
0 2488 7 3 2 23060 30486
0 2489 7 1 2 27399 27636
0 2490 7 1 2 29805 2489
0 2491 7 1 2 30501 2490
0 2492 5 1 1 2491
0 2493 7 1 2 2487 2492
0 2494 5 1 1 2493
0 2495 7 1 2 26724 30363
0 2496 7 1 2 2494 2495
0 2497 5 1 1 2496
0 2498 7 1 2 2475 2497
0 2499 5 1 1 2498
0 2500 7 1 2 24019 2499
0 2501 5 1 1 2500
0 2502 7 1 2 2453 2501
0 2503 7 1 2 2359 2502
0 2504 5 1 1 2503
0 2505 7 1 2 25899 2504
0 2506 5 1 1 2505
0 2507 7 4 2 22299 24840
0 2508 7 2 2 27547 30504
0 2509 7 2 2 23618 29207
0 2510 7 1 2 30508 30510
0 2511 7 2 2 29437 2510
0 2512 5 1 1 30512
0 2513 7 1 2 25021 30513
0 2514 5 1 1 2513
0 2515 7 16 2 25453 28782
0 2516 7 1 2 28753 30514
0 2517 5 1 1 2516
0 2518 7 4 2 25022 25562
0 2519 7 1 2 26054 30530
0 2520 5 1 1 2519
0 2521 7 1 2 27722 2520
0 2522 5 1 1 2521
0 2523 7 1 2 21773 23503
0 2524 7 1 2 2522 2523
0 2525 5 1 1 2524
0 2526 7 1 2 2517 2525
0 2527 5 1 1 2526
0 2528 7 1 2 29551 2527
0 2529 5 1 1 2528
0 2530 7 7 2 23504 25844
0 2531 5 4 1 30534
0 2532 7 5 2 21774 29475
0 2533 5 1 1 30545
0 2534 7 1 2 28754 30546
0 2535 7 1 2 30535 2534
0 2536 5 1 1 2535
0 2537 7 1 2 2529 2536
0 2538 5 1 1 2537
0 2539 7 1 2 26168 2538
0 2540 5 1 1 2539
0 2541 7 4 2 23061 27298
0 2542 5 2 1 30550
0 2543 7 1 2 24508 27299
0 2544 5 2 1 2543
0 2545 7 3 2 30554 30556
0 2546 5 1 1 30558
0 2547 7 1 2 30456 30559
0 2548 5 1 1 2547
0 2549 7 10 2 22508 24915
0 2550 5 9 1 30561
0 2551 7 5 2 25023 30562
0 2552 7 1 2 22448 30580
0 2553 5 1 1 2552
0 2554 7 1 2 2548 2553
0 2555 5 1 1 2554
0 2556 7 1 2 21775 30515
0 2557 5 1 1 2556
0 2558 7 1 2 30541 2557
0 2559 5 1 1 2558
0 2560 7 1 2 23619 2559
0 2561 7 1 2 2555 2560
0 2562 5 1 1 2561
0 2563 7 3 2 24315 29552
0 2564 7 2 2 24787 27282
0 2565 5 1 1 30588
0 2566 7 4 2 25024 28665
0 2567 7 1 2 30589 30590
0 2568 7 1 2 30585 2567
0 2569 5 1 1 2568
0 2570 7 1 2 2562 2569
0 2571 7 1 2 2540 2570
0 2572 5 1 1 2571
0 2573 7 1 2 27756 2572
0 2574 5 1 1 2573
0 2575 7 1 2 2514 2574
0 2576 5 1 1 2575
0 2577 7 1 2 30355 2576
0 2578 5 1 1 2577
0 2579 7 6 2 29065 30113
0 2580 5 21 1 30594
0 2581 7 4 2 23620 30600
0 2582 7 1 2 24788 29738
0 2583 5 1 1 2582
0 2584 7 1 2 29225 1239
0 2585 5 13 1 2584
0 2586 7 2 2 22300 30625
0 2587 5 1 1 30638
0 2588 7 1 2 29476 30639
0 2589 7 1 2 2583 2588
0 2590 5 1 1 2589
0 2591 7 2 2 27164 30536
0 2592 7 1 2 27862 30640
0 2593 5 1 1 2592
0 2594 7 2 2 27372 29584
0 2595 5 2 1 30642
0 2596 7 1 2 30516 30644
0 2597 5 1 1 2596
0 2598 7 1 2 2593 2597
0 2599 7 1 2 2590 2598
0 2600 5 1 1 2599
0 2601 7 1 2 30621 2600
0 2602 5 1 1 2601
0 2603 7 5 2 22449 24789
0 2604 7 3 2 21776 30646
0 2605 7 4 2 25563 30333
0 2606 7 2 2 23505 30654
0 2607 7 1 2 30651 30658
0 2608 5 1 1 2607
0 2609 7 8 2 22845 25454
0 2610 5 1 1 30660
0 2611 7 1 2 27215 30661
0 2612 7 1 2 30622 2611
0 2613 5 1 1 2612
0 2614 7 1 2 2608 2613
0 2615 5 1 1 2614
0 2616 7 1 2 24316 29477
0 2617 7 1 2 2615 2616
0 2618 5 2 1 2617
0 2619 7 1 2 2602 30668
0 2620 5 1 1 2619
0 2621 7 1 2 23258 2620
0 2622 5 1 1 2621
0 2623 7 3 2 22985 25213
0 2624 5 1 1 30670
0 2625 7 2 2 26257 30671
0 2626 7 3 2 28011 29208
0 2627 7 1 2 30673 30675
0 2628 5 1 1 2627
0 2629 7 1 2 2622 2628
0 2630 5 1 1 2629
0 2631 7 1 2 26195 29370
0 2632 7 1 2 2630 2631
0 2633 5 1 1 2632
0 2634 7 1 2 2578 2633
0 2635 5 1 1 2634
0 2636 7 1 2 22704 2635
0 2637 5 1 1 2636
0 2638 7 5 2 22613 23062
0 2639 7 1 2 30417 30678
0 2640 5 2 1 2639
0 2641 7 2 2 24648 25025
0 2642 7 2 2 25214 30685
0 2643 7 1 2 23178 30687
0 2644 5 1 1 2643
0 2645 7 1 2 30683 2644
0 2646 5 1 1 2645
0 2647 7 1 2 30641 2646
0 2648 5 1 1 2647
0 2649 7 1 2 24916 30517
0 2650 5 1 1 2649
0 2651 7 1 2 30542 2650
0 2652 5 3 1 2651
0 2653 7 1 2 24649 30165
0 2654 5 2 1 2653
0 2655 7 4 2 23063 23259
0 2656 7 2 2 26299 30694
0 2657 5 1 1 30698
0 2658 7 1 2 30692 2657
0 2659 5 2 1 2658
0 2660 7 1 2 27421 30700
0 2661 7 1 2 30689 2660
0 2662 5 1 1 2661
0 2663 7 1 2 2648 2662
0 2664 5 1 1 2663
0 2665 7 1 2 29553 2664
0 2666 5 1 1 2665
0 2667 7 1 2 28763 30547
0 2668 7 4 2 22450 29384
0 2669 7 4 2 23260 23506
0 2670 7 2 2 25151 30706
0 2671 7 1 2 30702 30710
0 2672 7 1 2 2667 2671
0 2673 5 1 1 2672
0 2674 7 1 2 2666 2673
0 2675 5 1 1 2674
0 2676 7 1 2 26337 29371
0 2677 7 1 2 2675 2676
0 2678 5 1 1 2677
0 2679 7 1 2 2637 2678
0 2680 5 1 1 2679
0 2681 7 1 2 22130 2680
0 2682 5 1 1 2681
0 2683 7 3 2 24152 30518
0 2684 5 1 1 30712
0 2685 7 1 2 29361 30487
0 2686 5 1 1 2685
0 2687 7 1 2 2684 2686
0 2688 5 1 1 2687
0 2689 7 1 2 23621 2688
0 2690 5 1 1 2689
0 2691 7 6 2 24917 23507
0 2692 7 1 2 24153 30715
0 2693 7 1 2 27895 2692
0 2694 5 1 1 2693
0 2695 7 1 2 2690 2694
0 2696 5 1 1 2695
0 2697 7 1 2 30688 2696
0 2698 5 1 1 2697
0 2699 7 4 2 24918 23261
0 2700 7 2 2 22705 23064
0 2701 7 1 2 30721 30725
0 2702 7 1 2 30676 2701
0 2703 5 1 1 2702
0 2704 7 1 2 2698 2703
0 2705 5 1 1 2704
0 2706 7 1 2 26300 2705
0 2707 5 1 1 2706
0 2708 7 1 2 27000 28012
0 2709 7 1 2 27224 2708
0 2710 7 1 2 29732 2709
0 2711 5 1 1 2710
0 2712 7 1 2 2707 2711
0 2713 5 1 1 2712
0 2714 7 1 2 27165 2713
0 2715 5 1 1 2714
0 2716 7 4 2 26725 26710
0 2717 7 4 2 24317 30662
0 2718 5 1 1 30731
0 2719 7 1 2 2587 2718
0 2720 5 5 1 2719
0 2721 7 2 2 23622 30735
0 2722 7 1 2 28625 30740
0 2723 5 1 1 2722
0 2724 7 1 2 29330 30591
0 2725 5 1 1 2724
0 2726 7 1 2 2723 2725
0 2727 5 1 1 2726
0 2728 7 1 2 27422 2727
0 2729 5 1 1 2728
0 2730 7 6 2 24154 25026
0 2731 5 2 1 30742
0 2732 7 1 2 24919 30743
0 2733 7 1 2 30741 2732
0 2734 5 1 1 2733
0 2735 7 1 2 2729 2734
0 2736 5 1 1 2735
0 2737 7 1 2 30727 2736
0 2738 5 1 1 2737
0 2739 7 1 2 2715 2738
0 2740 5 1 1 2739
0 2741 7 1 2 29554 2740
0 2742 5 1 1 2741
0 2743 7 2 2 22706 22986
0 2744 7 2 2 23262 29209
0 2745 7 1 2 30750 30752
0 2746 5 1 1 2745
0 2747 7 5 2 24920 25215
0 2748 7 2 2 26533 30754
0 2749 7 1 2 30626 30759
0 2750 5 1 1 2749
0 2751 7 1 2 2746 2750
0 2752 5 1 1 2751
0 2753 7 1 2 22301 2752
0 2754 5 1 1 2753
0 2755 7 1 2 30732 30760
0 2756 5 1 1 2755
0 2757 7 1 2 2754 2756
0 2758 5 1 1 2757
0 2759 7 7 2 22451 30548
0 2760 5 1 1 30761
0 2761 7 1 2 27015 27364
0 2762 7 1 2 30762 2761
0 2763 7 1 2 2758 2762
0 2764 5 1 1 2763
0 2765 7 1 2 2742 2764
0 2766 5 1 1 2765
0 2767 7 1 2 27757 2766
0 2768 5 1 1 2767
0 2769 7 2 2 27852 29646
0 2770 7 5 2 24841 25027
0 2771 7 2 2 30076 30770
0 2772 7 9 2 22614 25216
0 2773 7 3 2 23508 30777
0 2774 7 1 2 26621 30786
0 2775 7 1 2 30775 2774
0 2776 7 1 2 30768 2775
0 2777 5 1 1 2776
0 2778 7 1 2 2768 2777
0 2779 5 1 1 2778
0 2780 7 1 2 25313 2779
0 2781 5 1 1 2780
0 2782 7 1 2 2682 2781
0 2783 5 1 1 2782
0 2784 7 1 2 25374 2783
0 2785 5 1 1 2784
0 2786 7 3 2 28412 29854
0 2787 5 2 1 30789
0 2788 7 2 2 24576 30792
0 2789 5 1 1 30794
0 2790 7 2 2 27216 2789
0 2791 7 1 2 23179 30796
0 2792 5 1 1 2791
0 2793 7 1 2 29048 29747
0 2794 5 1 1 2793
0 2795 7 1 2 2792 2794
0 2796 5 1 1 2795
0 2797 7 1 2 28715 2796
0 2798 5 1 1 2797
0 2799 7 2 2 28079 28571
0 2800 7 1 2 30655 30798
0 2801 5 1 1 2800
0 2802 7 1 2 2798 2801
0 2803 5 1 1 2802
0 2804 7 1 2 29478 2803
0 2805 5 1 1 2804
0 2806 7 3 2 27896 29999
0 2807 7 1 2 25455 30800
0 2808 5 1 1 2807
0 2809 7 1 2 28716 29748
0 2810 5 1 1 2809
0 2811 7 1 2 2808 2810
0 2812 5 1 1 2811
0 2813 7 1 2 30341 2812
0 2814 5 1 1 2813
0 2815 7 2 2 30601 30645
0 2816 7 1 2 28717 30803
0 2817 5 1 1 2816
0 2818 7 1 2 2814 2817
0 2819 7 1 2 2805 2818
0 2820 5 1 1 2819
0 2821 7 1 2 24155 2820
0 2822 5 1 1 2821
0 2823 7 3 2 26258 28626
0 2824 7 1 2 29647 30805
0 2825 7 1 2 28718 2824
0 2826 5 1 1 2825
0 2827 7 1 2 2822 2826
0 2828 5 1 1 2827
0 2829 7 1 2 27758 2828
0 2830 5 1 1 2829
0 2831 7 5 2 23180 25456
0 2832 7 1 2 24156 30808
0 2833 7 1 2 30776 2832
0 2834 7 1 2 30769 2833
0 2835 5 1 1 2834
0 2836 7 1 2 2830 2835
0 2837 5 1 1 2836
0 2838 7 1 2 26995 28909
0 2839 7 1 2 2837 2838
0 2840 5 1 1 2839
0 2841 7 1 2 2785 2840
0 2842 5 1 1 2841
0 2843 7 1 2 21976 2842
0 2844 5 1 1 2843
0 2845 7 1 2 2506 2844
0 2846 7 1 2 2120 2845
0 2847 7 1 2 1768 2846
0 2848 5 1 1 2847
0 2849 7 1 2 28525 2848
0 2850 5 1 1 2849
0 2851 7 2 2 27927 30030
0 2852 7 2 2 26259 30813
0 2853 5 1 1 30815
0 2854 7 2 2 26534 30816
0 2855 5 1 1 30817
0 2856 7 4 2 23623 30240
0 2857 7 1 2 26658 26323
0 2858 5 1 1 2857
0 2859 7 4 2 25314 30778
0 2860 7 1 2 26622 30823
0 2861 5 1 1 2860
0 2862 7 1 2 2858 2861
0 2863 5 1 1 2862
0 2864 7 1 2 30819 2863
0 2865 5 1 1 2864
0 2866 7 1 2 2855 2865
0 2867 5 1 1 2866
0 2868 7 1 2 27207 2867
0 2869 5 1 1 2868
0 2870 7 2 2 26659 28635
0 2871 7 3 2 26568 30827
0 2872 7 3 2 25217 27166
0 2873 7 1 2 30127 30832
0 2874 7 1 2 30829 2873
0 2875 5 1 1 2874
0 2876 7 1 2 2869 2875
0 2877 5 1 1 2876
0 2878 7 1 2 23917 2877
0 2879 5 1 1 2878
0 2880 7 2 2 23918 29632
0 2881 5 2 1 30835
0 2882 7 3 2 27488 30836
0 2883 5 4 1 30839
0 2884 7 1 2 30105 30842
0 2885 5 1 1 2884
0 2886 7 3 2 21871 27489
0 2887 5 2 1 30846
0 2888 7 1 2 29529 30849
0 2889 5 6 1 2888
0 2890 7 1 2 27246 30851
0 2891 5 2 1 2890
0 2892 7 1 2 2885 30857
0 2893 5 1 1 2892
0 2894 7 2 2 25218 27093
0 2895 7 7 2 25375 28636
0 2896 7 1 2 30859 30861
0 2897 7 1 2 2893 2896
0 2898 5 1 1 2897
0 2899 7 1 2 2879 2898
0 2900 5 1 1 2899
0 2901 7 1 2 23065 2900
0 2902 5 1 1 2901
0 2903 7 3 2 23624 27373
0 2904 7 2 2 23919 22131
0 2905 7 2 2 25457 30871
0 2906 7 4 2 25028 25799
0 2907 5 1 1 30875
0 2908 7 1 2 28896 30106
0 2909 7 1 2 30876 2908
0 2910 7 1 2 30873 2909
0 2911 7 1 2 30868 2910
0 2912 5 1 1 2911
0 2913 7 1 2 2902 2912
0 2914 5 1 1 2913
0 2915 7 1 2 24509 2914
0 2916 5 1 1 2915
0 2917 7 3 2 23263 26301
0 2918 5 1 1 30879
0 2919 7 1 2 26037 26895
0 2920 5 1 1 2919
0 2921 7 1 2 2918 2920
0 2922 5 1 1 2921
0 2923 7 1 2 21777 2922
0 2924 5 1 1 2923
0 2925 7 3 2 26689 28876
0 2926 5 1 1 30882
0 2927 7 1 2 2924 2926
0 2928 5 1 1 2927
0 2929 7 1 2 21872 2928
0 2930 5 1 1 2929
0 2931 7 1 2 25152 28091
0 2932 5 1 1 2931
0 2933 7 9 2 23920 22987
0 2934 5 8 1 30885
0 2935 7 3 2 27490 30886
0 2936 5 2 1 30902
0 2937 7 1 2 25219 26274
0 2938 7 1 2 30903 2937
0 2939 7 1 2 2932 2938
0 2940 5 1 1 2939
0 2941 7 1 2 2930 2940
0 2942 5 1 1 2941
0 2943 7 1 2 25029 2942
0 2944 5 1 1 2943
0 2945 7 7 2 30272 30000
0 2946 5 2 1 30907
0 2947 7 1 2 30850 30914
0 2948 5 18 1 2947
0 2949 7 1 2 25030 30916
0 2950 5 2 1 2949
0 2951 7 5 2 22452 23066
0 2952 5 2 1 30936
0 2953 7 2 2 29424 30937
0 2954 5 1 1 30943
0 2955 7 1 2 30934 2954
0 2956 5 3 1 2955
0 2957 7 1 2 24577 30945
0 2958 5 1 1 2957
0 2959 7 1 2 29348 30679
0 2960 5 1 1 2959
0 2961 7 1 2 2958 2960
0 2962 5 1 1 2961
0 2963 7 1 2 30166 2962
0 2964 5 1 1 2963
0 2965 7 4 2 21873 25031
0 2966 5 5 1 30948
0 2967 7 1 2 29777 30952
0 2968 5 1 1 2967
0 2969 7 9 2 23921 23067
0 2970 5 2 1 30957
0 2971 7 2 2 22615 30966
0 2972 5 1 1 30968
0 2973 7 1 2 26690 30969
0 2974 7 1 2 2968 2973
0 2975 5 1 1 2974
0 2976 7 1 2 2964 2975
0 2977 5 1 1 2976
0 2978 7 1 2 22509 2977
0 2979 5 1 1 2978
0 2980 7 1 2 2944 2979
0 2981 5 1 1 2980
0 2982 7 1 2 30830 2981
0 2983 5 1 1 2982
0 2984 7 1 2 2916 2983
0 2985 5 1 1 2984
0 2986 7 1 2 24020 2985
0 2987 5 1 1 2986
0 2988 7 8 2 25220 26855
0 2989 7 1 2 26302 30970
0 2990 5 3 1 2989
0 2991 7 1 2 771 30978
0 2992 5 2 1 2991
0 2993 7 1 2 29438 30981
0 2994 5 1 1 2993
0 2995 7 3 2 23922 24578
0 2996 5 2 1 30983
0 2997 7 2 2 27374 29865
0 2998 7 2 2 30984 30988
0 2999 7 2 2 26569 30167
0 3000 7 1 2 30990 30992
0 3001 5 1 1 3000
0 3002 7 1 2 2994 3001
0 3003 5 1 1 3002
0 3004 7 1 2 25032 3003
0 3005 5 1 1 3004
0 3006 7 2 2 24579 2187
0 3007 7 4 2 27491 29633
0 3008 5 1 1 30996
0 3009 7 1 2 24510 30997
0 3010 5 2 1 3009
0 3011 7 1 2 30994 31000
0 3012 5 1 1 3011
0 3013 7 1 2 29156 30840
0 3014 5 2 1 3013
0 3015 7 1 2 3012 31002
0 3016 5 1 1 3015
0 3017 7 1 2 23181 3016
0 3018 5 1 1 3017
0 3019 7 2 2 24580 27261
0 3020 5 1 1 31004
0 3021 7 1 2 30023 31005
0 3022 5 2 1 3021
0 3023 7 1 2 3018 31006
0 3024 5 1 1 3023
0 3025 7 1 2 25221 3024
0 3026 5 1 1 3025
0 3027 7 1 2 29749 30193
0 3028 5 1 1 3027
0 3029 7 1 2 3026 3028
0 3030 5 1 1 3029
0 3031 7 1 2 23068 26570
0 3032 7 1 2 3030 3031
0 3033 5 1 1 3032
0 3034 7 1 2 3005 3033
0 3035 5 1 1 3034
0 3036 7 1 2 21977 3035
0 3037 5 1 1 3036
0 3038 7 3 2 23923 22510
0 3039 5 1 1 31008
0 3040 7 5 2 25033 31009
0 3041 7 1 2 26150 31011
0 3042 5 2 1 3041
0 3043 7 3 2 21874 28973
0 3044 5 2 1 31018
0 3045 7 1 2 27283 31019
0 3046 5 1 1 3045
0 3047 7 1 2 31016 3046
0 3048 5 1 1 3047
0 3049 7 1 2 21778 3048
0 3050 5 1 1 3049
0 3051 7 1 2 99 1258
0 3052 5 6 1 3051
0 3053 7 4 2 23803 31023
0 3054 5 1 1 31029
0 3055 7 1 2 31012 31030
0 3056 5 1 1 3055
0 3057 7 2 2 3050 3056
0 3058 5 2 1 31033
0 3059 7 4 2 23351 26303
0 3060 7 7 2 23264 25376
0 3061 7 1 2 31037 31041
0 3062 7 1 2 31035 3061
0 3063 5 1 1 3062
0 3064 7 1 2 3037 3063
0 3065 5 1 1 3064
0 3066 7 1 2 30828 3065
0 3067 5 1 1 3066
0 3068 7 1 2 2987 3067
0 3069 5 1 1 3068
0 3070 7 1 2 27729 3069
0 3071 5 1 1 3070
0 3072 7 2 2 23182 30949
0 3073 5 1 1 31048
0 3074 7 1 2 30595 3073
0 3075 5 2 1 3074
0 3076 7 1 2 29829 31050
0 3077 5 1 1 3076
0 3078 7 4 2 24921 27423
0 3079 7 4 2 22511 26959
0 3080 5 4 1 31056
0 3081 7 1 2 31052 31057
0 3082 5 1 1 3081
0 3083 7 5 2 21875 30602
0 3084 5 1 1 31064
0 3085 7 1 2 29813 31065
0 3086 5 1 1 3085
0 3087 7 1 2 3082 3086
0 3088 7 1 2 3077 3087
0 3089 5 1 1 3088
0 3090 7 1 2 21978 3089
0 3091 5 1 1 3090
0 3092 7 4 2 29555 30603
0 3093 5 1 1 31069
0 3094 7 2 2 28420 31070
0 3095 5 1 1 31073
0 3096 7 1 2 3091 3095
0 3097 5 2 1 3096
0 3098 7 1 2 23265 31075
0 3099 5 1 1 3098
0 3100 7 6 2 23804 29806
0 3101 5 1 1 31077
0 3102 7 3 2 25222 31078
0 3103 5 1 1 31083
0 3104 7 2 2 23924 31084
0 3105 7 2 2 28479 31086
0 3106 5 1 1 31088
0 3107 7 1 2 3099 3106
0 3108 5 1 1 3107
0 3109 7 1 2 27107 3108
0 3110 5 1 1 3109
0 3111 7 3 2 24157 25315
0 3112 7 1 2 26979 29443
0 3113 5 1 1 3112
0 3114 7 1 2 174 3113
0 3115 5 1 1 3114
0 3116 7 1 2 24581 3115
0 3117 5 1 1 3116
0 3118 7 1 2 26985 1508
0 3119 5 1 1 3118
0 3120 7 1 2 24650 3119
0 3121 5 1 1 3120
0 3122 7 1 2 3117 3121
0 3123 5 1 1 3122
0 3124 7 1 2 31090 3123
0 3125 5 1 1 3124
0 3126 7 1 2 22132 29014
0 3127 5 1 1 3126
0 3128 7 2 2 24511 24922
0 3129 7 1 2 27016 31093
0 3130 5 1 1 3129
0 3131 7 1 2 28772 3130
0 3132 5 1 1 3131
0 3133 7 1 2 23925 3132
0 3134 5 1 1 3133
0 3135 7 1 2 3127 3134
0 3136 5 1 1 3135
0 3137 7 1 2 25153 3136
0 3138 5 1 1 3137
0 3139 7 1 2 22133 26980
0 3140 5 1 1 3139
0 3141 7 1 2 3138 3140
0 3142 5 1 1 3141
0 3143 7 1 2 27089 3142
0 3144 5 1 1 3143
0 3145 7 1 2 3125 3144
0 3146 5 1 1 3145
0 3147 7 1 2 24459 3146
0 3148 5 1 1 3147
0 3149 7 1 2 22988 27108
0 3150 7 1 2 29139 3149
0 3151 5 1 1 3150
0 3152 7 1 2 3148 3151
0 3153 5 1 1 3152
0 3154 7 1 2 23805 3153
0 3155 5 1 1 3154
0 3156 7 2 2 25154 27109
0 3157 5 1 1 31095
0 3158 7 2 2 26151 28974
0 3159 5 1 1 31097
0 3160 7 1 2 23926 30052
0 3161 5 1 1 3160
0 3162 7 1 2 3159 3161
0 3163 5 4 1 3162
0 3164 7 1 2 31096 31099
0 3165 5 1 1 3164
0 3166 7 1 2 3155 3165
0 3167 5 1 1 3166
0 3168 7 1 2 25223 3167
0 3169 5 1 1 3168
0 3170 7 1 2 22134 30053
0 3171 5 1 1 3170
0 3172 7 1 2 24158 26388
0 3173 5 1 1 3172
0 3174 7 1 2 23806 3173
0 3175 7 1 2 2546 3174
0 3176 5 1 1 3175
0 3177 7 1 2 3171 3176
0 3178 5 1 1 3177
0 3179 7 1 2 23927 3178
0 3180 5 1 1 3179
0 3181 7 2 2 27492 28975
0 3182 7 2 2 29634 31103
0 3183 7 1 2 22135 31105
0 3184 5 1 1 3183
0 3185 7 1 2 3180 3184
0 3186 5 1 1 3185
0 3187 7 1 2 26260 3186
0 3188 5 1 1 3187
0 3189 7 1 2 29312 29807
0 3190 7 1 2 30158 3189
0 3191 5 1 1 3190
0 3192 7 1 2 3188 3191
0 3193 5 1 1 3192
0 3194 7 1 2 22707 26013
0 3195 7 1 2 3193 3194
0 3196 5 1 1 3195
0 3197 7 1 2 24021 3196
0 3198 7 1 2 3169 3197
0 3199 5 1 1 3198
0 3200 7 1 2 30728 30744
0 3201 5 2 1 3200
0 3202 7 1 2 28370 27004
0 3203 5 1 1 3202
0 3204 7 1 2 24159 23266
0 3205 5 1 1 3204
0 3206 7 2 2 27002 3205
0 3207 7 3 2 25155 30680
0 3208 7 1 2 31109 31111
0 3209 5 1 1 3208
0 3210 7 1 2 3203 3209
0 3211 5 1 1 3210
0 3212 7 1 2 27284 3211
0 3213 5 1 1 3212
0 3214 7 1 2 31107 3213
0 3215 5 1 1 3214
0 3216 7 1 2 21779 3215
0 3217 5 1 1 3216
0 3218 7 1 2 26535 26169
0 3219 7 1 2 30325 3218
0 3220 5 1 1 3219
0 3221 7 1 2 3217 3220
0 3222 5 1 1 3221
0 3223 7 1 2 23352 3222
0 3224 5 1 1 3223
0 3225 7 2 2 27079 30494
0 3226 5 1 1 31114
0 3227 7 1 2 23069 28421
0 3228 7 1 2 31115 3227
0 3229 5 1 1 3228
0 3230 7 1 2 3224 3229
0 3231 5 1 1 3230
0 3232 7 1 2 22512 3231
0 3233 5 1 1 3232
0 3234 7 2 2 21780 24160
0 3235 7 1 2 26711 31116
0 3236 7 1 2 26186 3235
0 3237 7 1 2 30386 3236
0 3238 5 1 1 3237
0 3239 7 1 2 3233 3238
0 3240 5 1 1 3239
0 3241 7 1 2 21876 3240
0 3242 5 1 1 3241
0 3243 7 4 2 29077 30373
0 3244 7 1 2 28413 25800
0 3245 7 1 2 26623 3244
0 3246 7 1 2 31118 3245
0 3247 5 1 1 3246
0 3248 7 1 2 21979 3247
0 3249 7 1 2 3242 3248
0 3250 5 1 1 3249
0 3251 7 1 2 3199 3250
0 3252 5 1 1 3251
0 3253 7 1 2 3110 3252
0 3254 5 1 1 3253
0 3255 7 1 2 25377 3254
0 3256 5 1 1 3255
0 3257 7 1 2 28422 29078
0 3258 5 2 1 3257
0 3259 7 1 2 21781 30560
0 3260 5 1 1 3259
0 3261 7 1 2 22513 30038
0 3262 5 1 1 3261
0 3263 7 2 2 3260 3262
0 3264 5 1 1 31124
0 3265 7 2 2 29002 3264
0 3266 5 1 1 31126
0 3267 7 1 2 21877 31127
0 3268 5 1 1 3267
0 3269 7 1 2 31122 3268
0 3270 5 1 1 3269
0 3271 7 6 2 21980 22616
0 3272 5 2 1 31128
0 3273 7 1 2 26660 31129
0 3274 7 2 2 3270 3273
0 3275 7 1 2 26867 31136
0 3276 5 1 1 3275
0 3277 7 1 2 3256 3276
0 3278 5 1 1 3277
0 3279 7 1 2 28637 3278
0 3280 5 1 1 3279
0 3281 7 1 2 24022 30818
0 3282 7 1 2 29947 3281
0 3283 5 1 1 3282
0 3284 7 1 2 3280 3283
0 3285 5 1 1 3284
0 3286 7 1 2 27759 3285
0 3287 5 1 1 3286
0 3288 7 1 2 3071 3287
0 3289 5 1 1 3288
0 3290 7 1 2 26757 3289
0 3291 5 1 1 3290
0 3292 7 6 2 25034 29556
0 3293 5 2 1 31138
0 3294 7 3 2 30356 31139
0 3295 7 3 2 25458 27400
0 3296 7 3 2 30001 31149
0 3297 7 1 2 26905 31152
0 3298 5 1 1 3297
0 3299 7 4 2 22453 24677
0 3300 7 4 2 24191 31155
0 3301 7 1 2 28414 30291
0 3302 7 1 2 31159 3301
0 3303 5 1 1 3302
0 3304 7 1 2 3298 3303
0 3305 5 1 1 3304
0 3306 7 1 2 31146 3305
0 3307 5 1 1 3306
0 3308 7 14 2 22732 25316
0 3309 7 2 2 22174 31163
0 3310 7 1 2 31042 31177
0 3311 7 1 2 30312 3310
0 3312 7 1 2 30334 30763
0 3313 7 1 2 3311 3312
0 3314 5 1 1 3313
0 3315 7 1 2 3307 3314
0 3316 5 1 1 3315
0 3317 7 1 2 21981 3316
0 3318 5 1 1 3317
0 3319 7 8 2 24023 29585
0 3320 5 15 1 31179
0 3321 7 1 2 26261 30295
0 3322 5 2 1 3321
0 3323 7 1 2 2221 31202
0 3324 5 1 1 3323
0 3325 7 2 2 26758 3324
0 3326 5 1 1 31204
0 3327 7 1 2 26852 30979
0 3328 5 3 1 3327
0 3329 7 4 2 24192 25652
0 3330 7 3 2 24678 23509
0 3331 7 1 2 26236 31213
0 3332 7 1 2 31209 3331
0 3333 7 1 2 31206 3332
0 3334 5 1 1 3333
0 3335 7 1 2 3326 3334
0 3336 5 1 1 3335
0 3337 7 1 2 27493 3336
0 3338 5 1 1 3337
0 3339 7 3 2 25653 29251
0 3340 7 2 2 23412 26726
0 3341 7 4 2 24923 25317
0 3342 7 2 2 31219 31221
0 3343 5 1 1 31225
0 3344 7 1 2 26853 3343
0 3345 5 1 1 3344
0 3346 7 1 2 28406 3345
0 3347 5 1 1 3346
0 3348 7 6 2 22175 24582
0 3349 7 5 2 27957 31227
0 3350 5 2 1 31233
0 3351 7 15 2 22733 23353
0 3352 5 5 1 31240
0 3353 7 4 2 22989 23413
0 3354 7 1 2 31241 31260
0 3355 7 1 2 31234 3354
0 3356 5 1 1 3355
0 3357 7 1 2 3347 3356
0 3358 5 1 1 3357
0 3359 7 1 2 31216 3358
0 3360 5 1 1 3359
0 3361 7 3 2 26448 30257
0 3362 7 1 2 26759 27262
0 3363 7 1 2 31264 3362
0 3364 5 1 1 3363
0 3365 7 1 2 3360 3364
0 3366 7 1 2 3338 3365
0 3367 5 1 1 3366
0 3368 7 1 2 29143 3367
0 3369 5 1 1 3368
0 3370 7 1 2 27208 29941
0 3371 7 1 2 31205 3370
0 3372 5 1 1 3371
0 3373 7 1 2 3369 3372
0 3374 5 1 1 3373
0 3375 7 1 2 31180 3374
0 3376 5 1 1 3375
0 3377 7 1 2 3318 3376
0 3378 5 1 1 3377
0 3379 7 1 2 26536 3378
0 3380 5 1 1 3379
0 3381 7 1 2 22514 30425
0 3382 5 1 1 3381
0 3383 7 1 2 21982 30196
0 3384 5 1 1 3383
0 3385 7 1 2 3382 3384
0 3386 5 1 1 3385
0 3387 7 1 2 25035 3386
0 3388 5 1 1 3387
0 3389 7 7 2 21983 24924
0 3390 5 2 1 31267
0 3391 7 3 2 22617 31268
0 3392 7 1 2 23267 31276
0 3393 5 1 1 3392
0 3394 7 1 2 2362 3393
0 3395 5 1 1 3394
0 3396 7 1 2 29049 3395
0 3397 5 1 1 3396
0 3398 7 1 2 3388 3397
0 3399 5 1 1 3398
0 3400 7 3 2 28136 30095
0 3401 7 1 2 3399 31279
0 3402 5 1 1 3401
0 3403 7 5 2 22734 25224
0 3404 7 13 2 24024 22176
0 3405 7 3 2 31282 31287
0 3406 7 1 2 29269 30313
0 3407 7 1 2 31300 3406
0 3408 7 1 2 30057 3407
0 3409 5 1 1 3408
0 3410 7 1 2 3402 3409
0 3411 5 1 1 3410
0 3412 7 1 2 23354 3411
0 3413 5 1 1 3412
0 3414 7 1 2 27348 31280
0 3415 5 1 1 3414
0 3416 7 1 2 28434 31150
0 3417 5 1 1 3416
0 3418 7 1 2 3415 3417
0 3419 5 1 1 3418
0 3420 7 1 2 28976 3419
0 3421 5 1 1 3420
0 3422 7 1 2 26906 29109
0 3423 7 1 2 27209 30314
0 3424 7 1 2 3422 3423
0 3425 5 1 1 3424
0 3426 7 1 2 3421 3425
0 3427 5 1 1 3426
0 3428 7 3 2 24025 25318
0 3429 7 1 2 30495 31303
0 3430 7 1 2 3427 3429
0 3431 5 1 1 3430
0 3432 7 1 2 3413 3431
0 3433 5 1 1 3432
0 3434 7 1 2 23928 3433
0 3435 5 1 1 3434
0 3436 7 3 2 23268 29479
0 3437 7 8 2 21984 27424
0 3438 7 1 2 31306 31309
0 3439 5 1 1 3438
0 3440 7 8 2 24026 25225
0 3441 7 1 2 31079 31317
0 3442 5 1 1 3441
0 3443 7 1 2 3439 3442
0 3444 5 1 1 3443
0 3445 7 1 2 29324 3444
0 3446 5 1 1 3445
0 3447 7 5 2 24027 23183
0 3448 5 1 1 31325
0 3449 7 3 2 24583 31326
0 3450 7 1 2 26014 31080
0 3451 7 1 2 31330 3450
0 3452 5 1 1 3451
0 3453 7 1 2 3446 3452
0 3454 5 1 1 3453
0 3455 7 1 2 29889 3454
0 3456 5 1 1 3455
0 3457 7 1 2 22618 29480
0 3458 5 2 1 3457
0 3459 7 1 2 31333 31144
0 3460 5 2 1 3459
0 3461 7 2 2 27425 31335
0 3462 5 1 1 31337
0 3463 7 1 2 30435 29621
0 3464 5 1 1 3463
0 3465 7 1 2 3462 3464
0 3466 5 1 1 3465
0 3467 7 1 2 21985 27935
0 3468 7 1 2 3466 3467
0 3469 5 1 1 3468
0 3470 7 1 2 3456 3469
0 3471 5 1 1 3470
0 3472 7 1 2 25378 3471
0 3473 5 1 1 3472
0 3474 7 14 2 21878 21986
0 3475 5 1 1 31339
0 3476 7 7 2 22515 31340
0 3477 7 3 2 28506 31353
0 3478 7 1 2 30002 30971
0 3479 7 1 2 31360 3478
0 3480 5 1 1 3479
0 3481 7 1 2 3473 3480
0 3482 5 1 1 3481
0 3483 7 1 2 26760 3482
0 3484 5 1 1 3483
0 3485 7 2 2 25379 26449
0 3486 7 3 2 28385 25814
0 3487 7 9 2 21987 24193
0 3488 7 1 2 29557 31368
0 3489 7 1 2 31365 3488
0 3490 7 1 2 31363 3489
0 3491 7 1 2 30003 3490
0 3492 5 1 1 3491
0 3493 7 1 2 3484 3492
0 3494 5 1 1 3493
0 3495 7 1 2 30315 3494
0 3496 5 1 1 3495
0 3497 7 4 2 23929 27126
0 3498 5 4 1 31377
0 3499 7 2 2 26691 29079
0 3500 5 1 1 31385
0 3501 7 3 2 23070 30168
0 3502 7 1 2 24512 31387
0 3503 5 1 1 3502
0 3504 7 1 2 3500 3503
0 3505 5 1 1 3504
0 3506 7 1 2 24584 3505
0 3507 5 1 1 3506
0 3508 7 1 2 29890 30880
0 3509 5 1 1 3508
0 3510 7 1 2 3507 3509
0 3511 5 1 1 3510
0 3512 7 1 2 31381 3511
0 3513 5 1 1 3512
0 3514 7 1 2 27241 28604
0 3515 5 2 1 3514
0 3516 7 1 2 21879 31390
0 3517 5 1 1 3516
0 3518 7 1 2 21880 30377
0 3519 5 1 1 3518
0 3520 7 1 2 27242 3519
0 3521 5 1 1 3520
0 3522 7 1 2 22516 3521
0 3523 5 1 1 3522
0 3524 7 1 2 3517 3523
0 3525 5 1 1 3524
0 3526 7 1 2 27167 3525
0 3527 5 1 1 3526
0 3528 7 1 2 29080 30133
0 3529 5 2 1 3528
0 3530 7 1 2 30131 31060
0 3531 5 1 1 3530
0 3532 7 1 2 29958 3531
0 3533 5 1 1 3532
0 3534 7 1 2 31392 3533
0 3535 7 1 2 3527 3534
0 3536 5 1 1 3535
0 3537 7 1 2 23269 3536
0 3538 5 1 1 3537
0 3539 7 1 2 3513 3538
0 3540 5 1 1 3539
0 3541 7 1 2 21988 3540
0 3542 5 1 1 3541
0 3543 7 1 2 23270 28489
0 3544 7 1 2 30134 3543
0 3545 5 1 1 3544
0 3546 7 1 2 2424 3545
0 3547 5 1 1 3546
0 3548 7 1 2 21782 3547
0 3549 5 1 1 3548
0 3550 7 2 2 21881 24460
0 3551 5 1 1 31394
0 3552 7 2 2 23807 31395
0 3553 7 1 2 30228 31396
0 3554 5 1 1 3553
0 3555 7 1 2 3549 3554
0 3556 5 1 1 3555
0 3557 7 1 2 29081 3556
0 3558 5 1 1 3557
0 3559 7 3 2 21783 24028
0 3560 7 3 2 21882 31398
0 3561 5 1 1 31401
0 3562 7 1 2 30181 31402
0 3563 5 1 1 3562
0 3564 7 3 2 21989 23271
0 3565 7 2 2 23930 27494
0 3566 5 11 1 31407
0 3567 7 1 2 31404 31409
0 3568 7 1 2 30135 3567
0 3569 5 1 1 3568
0 3570 7 1 2 3563 3569
0 3571 5 1 1 3570
0 3572 7 1 2 29003 3571
0 3573 5 1 1 3572
0 3574 7 1 2 3558 3573
0 3575 7 1 2 3542 3574
0 3576 5 1 1 3575
0 3577 7 1 2 23355 31281
0 3578 7 1 2 3576 3577
0 3579 5 1 1 3578
0 3580 7 1 2 3496 3579
0 3581 7 1 2 3435 3580
0 3582 5 1 1 3581
0 3583 7 1 2 26661 3582
0 3584 5 1 1 3583
0 3585 7 1 2 3380 3584
0 3586 5 1 1 3585
0 3587 7 1 2 25900 3586
0 3588 5 1 1 3587
0 3589 7 1 2 25319 2036
0 3590 5 1 1 3589
0 3591 7 1 2 22619 29814
0 3592 5 1 1 3591
0 3593 7 2 2 29819 3592
0 3594 5 1 1 31420
0 3595 7 1 2 21883 3594
0 3596 5 1 1 3595
0 3597 7 1 2 24585 30953
0 3598 5 1 1 3597
0 3599 7 1 2 29830 3598
0 3600 5 1 1 3599
0 3601 7 1 2 31123 3600
0 3602 7 1 2 3596 3601
0 3603 5 1 1 3602
0 3604 7 1 2 21990 3603
0 3605 5 1 1 3604
0 3606 7 1 2 29972 3605
0 3607 5 1 1 3606
0 3608 7 1 2 23184 3607
0 3609 7 1 2 3590 3608
0 3610 5 1 1 3609
0 3611 7 1 2 21991 29831
0 3612 5 2 1 3611
0 3613 7 1 2 29823 31422
0 3614 5 1 1 3613
0 3615 7 1 2 23931 31423
0 3616 5 2 1 3615
0 3617 7 1 2 23071 29325
0 3618 7 1 2 31424 3617
0 3619 7 1 2 3614 3618
0 3620 5 1 1 3619
0 3621 7 1 2 3610 3620
0 3622 5 1 1 3621
0 3623 7 1 2 22136 3622
0 3624 5 1 1 3623
0 3625 7 1 2 28901 29808
0 3626 7 1 2 29320 3625
0 3627 5 1 1 3626
0 3628 7 1 2 3624 3627
0 3629 5 1 1 3628
0 3630 7 1 2 22708 3629
0 3631 5 1 1 3630
0 3632 7 1 2 26718 31076
0 3633 5 1 1 3632
0 3634 7 1 2 22137 29326
0 3635 7 1 2 30938 3634
0 3636 7 4 2 21784 31341
0 3637 7 1 2 29969 31426
0 3638 7 1 2 3635 3637
0 3639 5 1 1 3638
0 3640 7 1 2 23272 3639
0 3641 7 1 2 3633 3640
0 3642 7 1 2 3631 3641
0 3643 5 1 1 3642
0 3644 7 1 2 24029 31100
0 3645 5 2 1 3644
0 3646 7 3 2 24030 22990
0 3647 7 1 2 29135 31432
0 3648 5 2 1 3647
0 3649 7 8 2 24031 23072
0 3650 5 5 1 31437
0 3651 7 1 2 30092 31445
0 3652 5 2 1 3651
0 3653 7 1 2 23932 31450
0 3654 5 1 1 3653
0 3655 7 1 2 24032 29015
0 3656 5 1 1 3655
0 3657 7 1 2 3654 3656
0 3658 5 1 1 3657
0 3659 7 1 2 24461 3658
0 3660 5 1 1 3659
0 3661 7 1 2 31435 3660
0 3662 5 1 1 3661
0 3663 7 1 2 23808 3662
0 3664 5 1 1 3663
0 3665 7 1 2 31430 3664
0 3666 5 1 1 3665
0 3667 7 1 2 27094 3666
0 3668 5 1 1 3667
0 3669 7 3 2 21992 29481
0 3670 5 21 1 31452
0 3671 7 3 2 24462 31455
0 3672 7 4 2 24033 29110
0 3673 5 2 1 31479
0 3674 7 1 2 30458 31480
0 3675 5 1 1 3674
0 3676 7 1 2 22620 3675
0 3677 5 1 1 3676
0 3678 7 1 2 31476 3677
0 3679 5 1 1 3678
0 3680 7 1 2 31436 3679
0 3681 5 1 1 3680
0 3682 7 1 2 23809 3681
0 3683 5 1 1 3682
0 3684 7 1 2 31431 3683
0 3685 5 3 1 3684
0 3686 7 1 2 25320 31485
0 3687 5 1 1 3686
0 3688 7 1 2 21884 29832
0 3689 5 1 1 3688
0 3690 7 1 2 29820 3689
0 3691 5 1 1 3690
0 3692 7 4 2 22621 23356
0 3693 7 11 2 21993 25036
0 3694 5 3 1 31492
0 3695 7 1 2 31488 31493
0 3696 7 1 2 3691 3695
0 3697 5 1 1 3696
0 3698 7 1 2 3687 3697
0 3699 5 1 1 3698
0 3700 7 1 2 26537 3699
0 3701 5 1 1 3700
0 3702 7 1 2 3668 3701
0 3703 5 1 1 3702
0 3704 7 1 2 25156 3703
0 3705 5 1 1 3704
0 3706 7 1 2 27110 31456
0 3707 5 1 1 3706
0 3708 7 3 2 23933 29339
0 3709 7 1 2 25321 30089
0 3710 7 1 2 31506 3709
0 3711 5 1 1 3710
0 3712 7 1 2 3707 3711
0 3713 5 1 1 3712
0 3714 7 1 2 28739 3713
0 3715 5 1 1 3714
0 3716 7 1 2 21994 22138
0 3717 7 1 2 28155 3716
0 3718 7 1 2 29648 3717
0 3719 5 1 1 3718
0 3720 7 1 2 3715 3719
0 3721 5 1 1 3720
0 3722 7 1 2 27230 3721
0 3723 5 1 1 3722
0 3724 7 1 2 25226 3723
0 3725 7 1 2 3705 3724
0 3726 5 1 1 3725
0 3727 7 1 2 27831 3726
0 3728 7 1 2 3643 3727
0 3729 5 1 1 3728
0 3730 7 4 2 22370 24925
0 3731 7 6 2 27816 31509
0 3732 5 1 1 31513
0 3733 7 1 2 25037 31514
0 3734 5 1 1 3733
0 3735 7 2 2 22991 29243
0 3736 7 1 2 22139 26104
0 3737 7 1 2 31519 3736
0 3738 5 1 1 3737
0 3739 7 1 2 3734 3738
0 3740 5 1 1 3739
0 3741 7 1 2 29684 3740
0 3742 5 1 1 3741
0 3743 7 2 2 21785 30267
0 3744 5 2 1 31521
0 3745 7 1 2 27817 29536
0 3746 7 6 2 22517 23073
0 3747 5 6 1 31525
0 3748 7 5 2 22371 24651
0 3749 7 1 2 31526 31537
0 3750 7 1 2 3745 3749
0 3751 7 1 2 31522 3750
0 3752 5 1 1 3751
0 3753 7 1 2 3742 3752
0 3754 5 1 1 3753
0 3755 7 1 2 26324 3754
0 3756 5 1 1 3755
0 3757 7 3 2 24463 24652
0 3758 7 1 2 25322 29835
0 3759 7 1 2 31542 3758
0 3760 7 4 2 22622 26727
0 3761 7 1 2 29175 29321
0 3762 7 1 2 31545 3761
0 3763 7 1 2 3759 3762
0 3764 5 1 1 3763
0 3765 7 1 2 3756 3764
0 3766 7 1 2 3729 3765
0 3767 5 1 1 3766
0 3768 7 1 2 23414 3767
0 3769 5 1 1 3768
0 3770 7 1 2 27832 29948
0 3771 5 1 1 3770
0 3772 7 2 2 26489 28446
0 3773 7 1 2 29238 31520
0 3774 7 1 2 31549 3773
0 3775 5 1 1 3774
0 3776 7 1 2 3771 3775
0 3777 5 1 1 3776
0 3778 7 1 2 27971 30475
0 3779 7 1 2 3777 3778
0 3780 5 1 1 3779
0 3781 7 1 2 3769 3780
0 3782 5 1 1 3781
0 3783 7 1 2 28666 3782
0 3784 5 1 1 3783
0 3785 7 4 2 28638 29871
0 3786 7 2 2 23725 26728
0 3787 7 1 2 26196 31555
0 3788 7 1 2 31551 3787
0 3789 7 1 2 31137 3788
0 3790 5 1 1 3789
0 3791 7 1 2 3784 3790
0 3792 5 1 1 3791
0 3793 7 1 2 25743 3792
0 3794 5 1 1 3793
0 3795 7 1 2 3588 3794
0 3796 7 1 2 3291 3795
0 3797 5 1 1 3796
0 3798 7 1 2 28783 3797
0 3799 5 1 1 3798
0 3800 7 2 2 22992 29482
0 3801 5 1 1 31557
0 3802 7 1 2 31531 3801
0 3803 5 1 1 3802
0 3804 7 1 2 24586 3803
0 3805 5 2 1 3804
0 3806 7 1 2 27495 31334
0 3807 5 2 1 3806
0 3808 7 1 2 29614 31561
0 3809 5 1 1 3808
0 3810 7 1 2 26378 3809
0 3811 5 1 1 3810
0 3812 7 1 2 31559 3811
0 3813 5 1 1 3812
0 3814 7 1 2 30169 3813
0 3815 5 1 1 3814
0 3816 7 3 2 27017 26692
0 3817 7 1 2 29964 31563
0 3818 5 1 1 3817
0 3819 7 1 2 26896 29385
0 3820 5 1 1 3819
0 3821 7 1 2 30684 3820
0 3822 5 1 1 3821
0 3823 7 1 2 27168 3822
0 3824 5 1 1 3823
0 3825 7 1 2 3818 3824
0 3826 7 1 2 3815 3825
0 3827 5 1 1 3826
0 3828 7 1 2 24653 3827
0 3829 5 1 1 3828
0 3830 7 6 2 24587 23273
0 3831 7 1 2 26960 30751
0 3832 7 1 2 31566 3831
0 3833 5 1 1 3832
0 3834 7 1 2 3829 3833
0 3835 5 1 1 3834
0 3836 7 1 2 31091 3835
0 3837 5 1 1 3836
0 3838 7 2 2 27496 29444
0 3839 5 2 1 31572
0 3840 7 1 2 26961 31573
0 3841 5 1 1 3840
0 3842 7 2 2 27252 26975
0 3843 5 3 1 31576
0 3844 7 1 2 22518 27169
0 3845 5 5 1 3844
0 3846 7 2 2 29349 31581
0 3847 7 3 2 29586 31586
0 3848 7 2 2 22993 31588
0 3849 7 2 2 31578 31591
0 3850 5 1 1 31593
0 3851 7 1 2 3841 3850
0 3852 5 1 1 3851
0 3853 7 1 2 3852 30860
0 3854 5 1 1 3853
0 3855 7 1 2 3837 3854
0 3856 5 1 1 3855
0 3857 7 1 2 26821 3856
0 3858 5 1 1 3857
0 3859 7 1 2 26822 26170
0 3860 5 1 1 3859
0 3861 7 2 2 28398 31160
0 3862 5 1 1 31595
0 3863 7 1 2 3860 3862
0 3864 5 1 1 3863
0 3865 7 1 2 21786 3864
0 3866 5 2 1 3865
0 3867 7 1 2 26823 27285
0 3868 5 1 1 3867
0 3869 7 1 2 31597 3868
0 3870 5 1 1 3869
0 3871 7 1 2 29558 3870
0 3872 5 1 1 3871
0 3873 7 7 2 22735 26785
0 3874 7 8 2 22177 31599
0 3875 5 2 1 31606
0 3876 7 1 2 29855 30549
0 3877 7 1 2 31607 3876
0 3878 5 1 1 3877
0 3879 7 1 2 3872 3878
0 3880 5 1 1 3879
0 3881 7 5 2 23185 23357
0 3882 7 1 2 27005 31616
0 3883 7 1 2 3880 3882
0 3884 5 1 1 3883
0 3885 7 2 2 21885 24194
0 3886 7 2 2 27426 31621
0 3887 7 1 2 28173 30563
0 3888 7 1 2 31623 3887
0 3889 5 1 1 3888
0 3890 7 1 2 30006 31145
0 3891 5 1 1 3890
0 3892 7 11 2 22178 23415
0 3893 7 4 2 22736 31625
0 3894 7 6 2 23074 29587
0 3895 5 4 1 31640
0 3896 7 1 2 31636 31646
0 3897 7 1 2 3891 3896
0 3898 5 1 1 3897
0 3899 7 1 2 3889 3898
0 3900 5 1 1 3899
0 3901 7 1 2 22623 22709
0 3902 7 1 2 26729 3901
0 3903 7 1 2 26921 3902
0 3904 7 1 2 3900 3903
0 3905 5 1 1 3904
0 3906 7 1 2 3884 3905
0 3907 5 1 1 3906
0 3908 7 1 2 22140 3907
0 3909 5 1 1 3908
0 3910 7 1 2 31110 31038
0 3911 5 1 1 3910
0 3912 7 1 2 3911 3226
0 3913 5 1 1 3912
0 3914 7 1 2 29396 31532
0 3915 5 7 1 3914
0 3916 7 2 2 29127 31650
0 3917 7 2 2 22454 31657
0 3918 5 1 1 31659
0 3919 7 1 2 1823 3918
0 3920 5 1 1 3919
0 3921 7 1 2 31608 3920
0 3922 5 1 1 3921
0 3923 7 2 2 21886 31527
0 3924 5 1 1 31661
0 3925 7 1 2 27286 31662
0 3926 7 1 2 28319 3925
0 3927 5 1 1 3926
0 3928 7 1 2 3922 3927
0 3929 5 1 1 3928
0 3930 7 1 2 21787 3929
0 3931 5 1 1 3930
0 3932 7 1 2 23075 30278
0 3933 7 1 2 31609 3932
0 3934 5 1 1 3933
0 3935 7 1 2 3931 3934
0 3936 5 1 1 3935
0 3937 7 1 2 3913 3936
0 3938 5 1 1 3937
0 3939 7 1 2 29588 29635
0 3940 5 1 1 3939
0 3941 7 3 2 29483 3940
0 3942 7 2 2 25815 31489
0 3943 7 1 2 31663 31666
0 3944 5 1 1 3943
0 3945 7 1 2 27325 28054
0 3946 5 1 1 3945
0 3947 7 1 2 3944 3946
0 3948 5 1 1 3947
0 3949 7 1 2 27951 30404
0 3950 7 1 2 3948 3949
0 3951 5 1 1 3950
0 3952 7 1 2 3938 3951
0 3953 7 1 2 3909 3952
0 3954 5 1 1 3953
0 3955 7 1 2 21995 3954
0 3956 5 1 1 3955
0 3957 7 1 2 3858 3956
0 3958 5 1 1 3957
0 3959 7 1 2 26402 3958
0 3960 5 1 1 3959
0 3961 7 2 2 23416 28062
0 3962 5 1 1 31668
0 3963 7 1 2 255 3962
0 3964 5 3 1 3963
0 3965 7 2 2 27339 30039
0 3966 5 5 1 31673
0 3967 7 1 2 31670 31674
0 3968 5 1 1 3967
0 3969 7 1 2 31669 31053
0 3970 5 1 1 3969
0 3971 7 1 2 3968 3970
0 3972 5 1 1 3971
0 3973 7 2 2 26730 3972
0 3974 7 4 2 22179 22624
0 3975 7 4 2 22519 22737
0 3976 7 2 2 31682 31686
0 3977 7 3 2 24842 31342
0 3978 7 1 2 28667 31692
0 3979 7 1 2 31690 3978
0 3980 7 1 2 31680 3979
0 3981 5 1 1 3980
0 3982 7 1 2 3960 3981
0 3983 5 1 1 3982
0 3984 7 1 2 22372 3983
0 3985 5 1 1 3984
0 3986 7 2 2 22902 28668
0 3987 7 2 2 31681 31695
0 3988 7 3 2 21996 22520
0 3989 5 1 1 31699
0 3990 7 5 2 21887 31700
0 3991 5 2 1 31702
0 3992 7 3 2 22625 22738
0 3993 7 5 2 22180 24365
0 3994 7 1 2 31709 31712
0 3995 7 1 2 31703 3994
0 3996 7 1 2 31697 3995
0 3997 5 1 1 3996
0 3998 7 1 2 3985 3997
0 3999 5 1 1 3998
0 4000 7 1 2 25845 3999
0 4001 5 1 1 4000
0 4002 7 1 2 21997 31596
0 4003 5 1 1 4002
0 4004 7 1 2 2305 31274
0 4005 5 1 1 4004
0 4006 7 1 2 31610 4005
0 4007 5 1 1 4006
0 4008 7 1 2 4003 4007
0 4009 5 1 1 4008
0 4010 7 1 2 25038 4009
0 4011 5 1 1 4010
0 4012 7 2 2 25459 28386
0 4013 7 2 2 23417 31717
0 4014 7 1 2 31369 31719
0 4015 5 2 1 4014
0 4016 7 1 2 4011 31721
0 4017 5 1 1 4016
0 4018 7 1 2 21788 4017
0 4019 5 1 1 4018
0 4020 7 1 2 24588 30387
0 4021 5 1 1 4020
0 4022 7 1 2 31611 4021
0 4023 5 1 1 4022
0 4024 7 1 2 24195 26171
0 4025 7 1 2 31720 4024
0 4026 5 1 1 4025
0 4027 7 1 2 4023 4026
0 4028 5 1 1 4027
0 4029 7 1 2 21998 4028
0 4030 5 1 1 4029
0 4031 7 1 2 4019 4030
0 4032 5 1 1 4031
0 4033 7 1 2 29484 4032
0 4034 5 1 1 4033
0 4035 7 2 2 22455 22739
0 4036 7 6 2 22181 31723
0 4037 7 3 2 24926 26786
0 4038 7 1 2 31725 31731
0 4039 5 1 1 4038
0 4040 7 1 2 31598 4039
0 4041 5 2 1 4040
0 4042 7 1 2 31734 31130
0 4043 5 1 1 4042
0 4044 7 1 2 1241 31503
0 4045 5 1 1 4044
0 4046 7 1 2 21789 28320
0 4047 5 1 1 4046
0 4048 7 1 2 31614 4047
0 4049 5 1 1 4048
0 4050 7 1 2 4045 4049
0 4051 5 1 1 4050
0 4052 7 2 2 21790 31683
0 4053 7 1 2 31600 31736
0 4054 5 1 1 4053
0 4055 7 1 2 28321 31494
0 4056 5 1 1 4055
0 4057 7 1 2 4054 4056
0 4058 5 1 1 4057
0 4059 7 1 2 26172 4058
0 4060 5 1 1 4059
0 4061 7 1 2 31722 4060
0 4062 7 1 2 4051 4061
0 4063 5 1 1 4062
0 4064 7 1 2 29559 4063
0 4065 5 1 1 4064
0 4066 7 1 2 4043 4065
0 4067 7 1 2 4034 4066
0 4068 5 1 1 4067
0 4069 7 1 2 23274 4068
0 4070 5 1 1 4069
0 4071 7 1 2 26379 28322
0 4072 7 1 2 31087 4071
0 4073 5 1 1 4072
0 4074 7 1 2 23186 4073
0 4075 7 1 2 4070 4074
0 4076 5 1 1 4075
0 4077 7 7 2 21999 23076
0 4078 5 2 1 31738
0 4079 7 1 2 28323 31739
0 4080 5 1 1 4079
0 4081 7 1 2 30703 31612
0 4082 5 1 1 4081
0 4083 7 1 2 4080 4082
0 4084 5 1 1 4083
0 4085 7 1 2 21791 4084
0 4086 5 1 1 4085
0 4087 7 1 2 26173 28324
0 4088 5 1 1 4087
0 4089 7 1 2 31615 4088
0 4090 5 1 1 4089
0 4091 7 1 2 31740 4090
0 4092 5 1 1 4091
0 4093 7 1 2 4086 4092
0 4094 5 1 1 4093
0 4095 7 1 2 29485 4094
0 4096 5 1 1 4095
0 4097 7 1 2 31735 31187
0 4098 5 1 1 4097
0 4099 7 4 2 21888 31370
0 4100 7 4 2 22521 24679
0 4101 7 1 2 28289 31751
0 4102 7 1 2 31747 4101
0 4103 5 1 1 4102
0 4104 7 1 2 4098 4103
0 4105 5 1 1 4104
0 4106 7 1 2 23077 4105
0 4107 5 1 1 4106
0 4108 7 1 2 4096 4107
0 4109 5 1 1 4108
0 4110 7 1 2 23275 4109
0 4111 5 1 1 4110
0 4112 7 2 2 25227 29445
0 4113 7 2 2 24464 29891
0 4114 5 3 1 31757
0 4115 7 1 2 22626 31759
0 4116 5 2 1 4115
0 4117 7 1 2 31613 31762
0 4118 5 1 1 4117
0 4119 7 1 2 28325 28046
0 4120 5 1 1 4119
0 4121 7 1 2 4118 4120
0 4122 5 1 1 4121
0 4123 7 1 2 23810 4122
0 4124 5 1 1 4123
0 4125 7 1 2 24589 28153
0 4126 5 1 1 4125
0 4127 7 1 2 4124 4126
0 4128 5 1 1 4127
0 4129 7 1 2 31755 4128
0 4130 5 1 1 4129
0 4131 7 1 2 25157 4130
0 4132 7 1 2 4111 4131
0 4133 5 1 1 4132
0 4134 7 1 2 28105 4133
0 4135 7 1 2 4076 4134
0 4136 5 1 1 4135
0 4137 7 2 2 22456 30346
0 4138 5 1 1 31764
0 4139 7 2 2 26962 30564
0 4140 5 1 1 31766
0 4141 7 2 2 21889 31767
0 4142 5 1 1 31768
0 4143 7 1 2 4138 4142
0 4144 5 1 1 4143
0 4145 7 1 2 21792 4144
0 4146 5 1 1 4145
0 4147 7 1 2 27287 30342
0 4148 5 1 1 4147
0 4149 7 1 2 4146 4148
0 4150 5 1 1 4149
0 4151 7 3 2 22000 28116
0 4152 7 1 2 23276 28327
0 4153 7 1 2 31770 4152
0 4154 7 1 2 4150 4153
0 4155 5 1 1 4154
0 4156 7 1 2 4136 4155
0 4157 5 1 1 4156
0 4158 7 1 2 27111 4157
0 4159 5 1 1 4158
0 4160 7 4 2 21890 22373
0 4161 7 2 2 31701 31773
0 4162 7 1 2 22182 26055
0 4163 7 1 2 31710 4162
0 4164 7 1 2 31777 4163
0 4165 7 1 2 31698 4164
0 4166 5 1 1 4165
0 4167 7 1 2 4159 4166
0 4168 7 1 2 4001 4167
0 4169 5 1 1 4168
0 4170 7 1 2 23726 4169
0 4171 5 1 1 4170
0 4172 7 5 2 23934 22183
0 4173 7 1 2 27638 31779
0 4174 7 2 2 24465 30090
0 4175 7 1 2 28040 31784
0 4176 7 2 2 22903 29892
0 4177 7 5 2 22740 27958
0 4178 5 1 1 31788
0 4179 7 1 2 31786 31789
0 4180 7 1 2 4175 4179
0 4181 7 1 2 4173 4180
0 4182 5 1 1 4181
0 4183 7 2 2 21793 27897
0 4184 5 1 1 31793
0 4185 7 1 2 27723 4184
0 4186 5 1 1 4185
0 4187 7 1 2 26174 4186
0 4188 5 1 1 4187
0 4189 7 2 2 26056 26472
0 4190 5 1 1 31795
0 4191 7 1 2 22457 31796
0 4192 5 1 1 4191
0 4193 7 3 2 21794 22302
0 4194 7 1 2 27869 31797
0 4195 5 1 1 4194
0 4196 7 1 2 4192 4195
0 4197 7 1 2 4188 4196
0 4198 5 1 1 4197
0 4199 7 1 2 27760 4198
0 4200 5 1 1 4199
0 4201 7 1 2 25901 30398
0 4202 5 1 1 4201
0 4203 7 3 2 22458 31798
0 4204 7 2 2 24366 22846
0 4205 7 2 2 24843 31803
0 4206 7 1 2 27805 31805
0 4207 7 1 2 31800 4206
0 4208 5 1 1 4207
0 4209 7 1 2 4202 4208
0 4210 7 1 2 4200 4209
0 4211 5 1 1 4210
0 4212 7 1 2 29560 4211
0 4213 5 1 1 4212
0 4214 7 3 2 24927 23727
0 4215 7 1 2 22374 29486
0 4216 7 1 2 31807 4215
0 4217 7 1 2 29378 31801
0 4218 7 1 2 4216 4217
0 4219 5 1 1 4218
0 4220 7 1 2 4213 4219
0 4221 5 1 1 4220
0 4222 7 5 2 25228 31371
0 4223 7 1 2 31810 31366
0 4224 7 1 2 4221 4223
0 4225 5 1 1 4224
0 4226 7 1 2 4182 4225
0 4227 5 1 1 4226
0 4228 7 1 2 30364 4227
0 4229 5 1 1 4228
0 4230 7 2 2 26057 25902
0 4231 5 1 1 31815
0 4232 7 1 2 651 4231
0 4233 5 18 1 4232
0 4234 7 2 2 22459 29985
0 4235 7 5 2 22184 31427
0 4236 7 3 2 31835 31837
0 4237 7 2 2 30120 30318
0 4238 7 1 2 22741 30096
0 4239 7 1 2 31845 4238
0 4240 7 1 2 31671 4239
0 4241 7 1 2 31842 4240
0 4242 5 1 1 4241
0 4243 7 4 2 21795 29537
0 4244 7 2 2 31769 31847
0 4245 5 1 1 31851
0 4246 7 5 2 23277 23625
0 4247 7 2 2 25654 31853
0 4248 7 1 2 27112 31858
0 4249 7 1 2 28328 4248
0 4250 7 1 2 31852 4249
0 4251 5 1 1 4250
0 4252 7 1 2 4242 4251
0 4253 5 1 1 4252
0 4254 7 1 2 31817 4253
0 4255 5 1 1 4254
0 4256 7 1 2 4229 4255
0 4257 7 1 2 4171 4256
0 4258 7 1 2 3799 4257
0 4259 7 1 2 2850 4258
0 4260 7 1 2 1222 4259
0 4261 5 1 1 4260
0 4262 7 1 2 25697 4261
0 4263 5 1 1 4262
0 4264 7 4 2 24928 23418
0 4265 7 2 2 28388 31156
0 4266 7 2 2 31860 31864
0 4267 7 1 2 27587 31866
0 4268 5 1 1 4267
0 4269 7 5 2 22303 26907
0 4270 7 1 2 30368 31868
0 4271 5 1 1 4270
0 4272 7 1 2 4268 4271
0 4273 5 1 1 4272
0 4274 7 1 2 21796 4273
0 4275 5 1 1 4274
0 4276 7 2 2 22460 28466
0 4277 7 4 2 25380 27401
0 4278 7 1 2 24929 31875
0 4279 7 1 2 31873 4278
0 4280 5 1 1 4279
0 4281 7 1 2 4275 4280
0 4282 5 1 1 4281
0 4283 7 1 2 25903 4282
0 4284 5 1 1 4283
0 4285 7 1 2 24844 27853
0 4286 7 5 2 22742 24930
0 4287 7 2 2 22185 31879
0 4288 7 2 2 25381 27427
0 4289 7 1 2 31884 31886
0 4290 7 1 2 4285 4289
0 4291 5 1 1 4290
0 4292 7 1 2 4284 4291
0 4293 5 1 1 4292
0 4294 7 1 2 30627 4293
0 4295 5 1 1 4294
0 4296 7 4 2 24680 23419
0 4297 7 3 2 28266 31888
0 4298 5 1 1 31892
0 4299 7 3 2 22186 24318
0 4300 7 6 2 22743 25382
0 4301 7 3 2 31895 31898
0 4302 5 1 1 31904
0 4303 7 1 2 4298 4302
0 4304 5 1 1 4303
0 4305 7 2 2 24367 27428
0 4306 7 1 2 27577 31907
0 4307 5 1 1 4306
0 4308 7 1 2 27833 29750
0 4309 5 1 1 4308
0 4310 7 1 2 4307 4309
0 4311 5 1 1 4310
0 4312 7 1 2 28686 4311
0 4313 5 1 1 4312
0 4314 7 1 2 22847 31153
0 4315 5 1 1 4314
0 4316 7 12 2 24790 23510
0 4317 5 1 1 31909
0 4318 7 1 2 27588 31910
0 4319 7 1 2 28423 4318
0 4320 5 1 1 4319
0 4321 7 1 2 4315 4320
0 4322 5 1 1 4321
0 4323 7 1 2 25904 4322
0 4324 5 1 1 4323
0 4325 7 1 2 4313 4324
0 4326 5 1 1 4325
0 4327 7 1 2 4304 4326
0 4328 5 1 1 4327
0 4329 7 3 2 28137 28669
0 4330 5 1 1 31921
0 4331 7 1 2 26908 28639
0 4332 5 1 1 4331
0 4333 7 1 2 4330 4332
0 4334 5 5 1 4333
0 4335 7 1 2 28616 31924
0 4336 5 1 1 4335
0 4337 7 1 2 28704 31922
0 4338 5 1 1 4337
0 4339 7 1 2 4336 4338
0 4340 5 1 1 4339
0 4341 7 1 2 29751 4340
0 4342 5 1 1 4341
0 4343 7 4 2 26909 30677
0 4344 5 1 1 31929
0 4345 7 1 2 28329 30801
0 4346 5 1 1 4345
0 4347 7 1 2 4344 4346
0 4348 7 1 2 4342 4347
0 4349 5 1 1 4348
0 4350 7 1 2 27761 4349
0 4351 5 1 1 4350
0 4352 7 1 2 4328 4351
0 4353 7 1 2 4295 4352
0 4354 5 1 1 4353
0 4355 7 1 2 29561 4354
0 4356 5 1 1 4355
0 4357 7 1 2 27170 31930
0 4358 5 1 1 4357
0 4359 7 1 2 28784 31925
0 4360 5 1 1 4359
0 4361 7 1 2 28687 31893
0 4362 5 1 1 4361
0 4363 7 1 2 4360 4362
0 4364 5 1 1 4363
0 4365 7 1 2 27429 4364
0 4366 5 1 1 4365
0 4367 7 1 2 4358 4366
0 4368 5 1 1 4367
0 4369 7 1 2 29487 31515
0 4370 7 1 2 4368 4369
0 4371 5 1 1 4370
0 4372 7 1 2 4356 4371
0 4373 5 1 1 4372
0 4374 7 1 2 31564 4373
0 4375 5 1 1 4374
0 4376 7 4 2 24681 22848
0 4377 5 1 1 31933
0 4378 7 6 2 24196 31934
0 4379 7 2 2 26963 31861
0 4380 7 1 2 31937 31943
0 4381 5 1 1 4380
0 4382 7 4 2 24791 25383
0 4383 5 1 1 31945
0 4384 7 3 2 26761 31946
0 4385 5 1 1 31949
0 4386 7 1 2 30335 31950
0 4387 5 1 1 4386
0 4388 7 1 2 4381 4387
0 4389 5 1 1 4388
0 4390 7 1 2 24319 4389
0 4391 5 1 1 4390
0 4392 7 1 2 24792 28354
0 4393 7 1 2 31944 4392
0 4394 5 1 1 4393
0 4395 7 1 2 4391 4394
0 4396 5 1 1 4395
0 4397 7 1 2 22904 4396
0 4398 5 1 1 4397
0 4399 7 2 2 25384 30336
0 4400 7 3 2 22744 22849
0 4401 7 5 2 22187 22304
0 4402 7 3 2 31954 31957
0 4403 7 1 2 24845 31962
0 4404 7 1 2 31952 4403
0 4405 5 1 1 4404
0 4406 7 1 2 4398 4405
0 4407 5 1 1 4406
0 4408 7 1 2 22375 4407
0 4409 5 1 1 4408
0 4410 7 4 2 24368 28257
0 4411 7 1 2 28467 31965
0 4412 7 1 2 31953 4411
0 4413 5 1 1 4412
0 4414 7 1 2 4409 4413
0 4415 5 1 1 4414
0 4416 7 1 2 27430 4415
0 4417 5 1 1 4416
0 4418 7 6 2 23420 28785
0 4419 7 3 2 26197 25744
0 4420 7 1 2 27217 30604
0 4421 7 1 2 31975 4420
0 4422 7 1 2 31969 4421
0 4423 5 1 1 4422
0 4424 7 1 2 4417 4423
0 4425 5 1 1 4424
0 4426 7 1 2 25564 4425
0 4427 5 1 1 4426
0 4428 7 1 2 26964 29622
0 4429 5 1 1 4428
0 4430 7 1 2 30596 4429
0 4431 5 1 1 4430
0 4432 7 1 2 28250 28342
0 4433 7 1 2 4431 4432
0 4434 5 1 1 4433
0 4435 7 1 2 4427 4434
0 4436 5 1 1 4435
0 4437 7 1 2 21891 4436
0 4438 5 1 1 4437
0 4439 7 2 2 26910 27870
0 4440 5 1 1 31978
0 4441 7 2 2 27027 30647
0 4442 7 1 2 25745 31980
0 4443 5 1 1 4442
0 4444 7 1 2 4440 4443
0 4445 5 1 1 4444
0 4446 7 2 2 24931 4445
0 4447 5 1 1 31982
0 4448 7 4 2 22850 28925
0 4449 7 1 2 31726 31984
0 4450 5 1 1 4449
0 4451 7 1 2 4447 4450
0 4452 5 1 1 4451
0 4453 7 1 2 22305 4452
0 4454 5 1 1 4453
0 4455 7 1 2 27028 30077
0 4456 7 1 2 31865 4455
0 4457 5 1 1 4456
0 4458 7 1 2 4454 4457
0 4459 5 1 1 4458
0 4460 7 1 2 21797 4459
0 4461 5 1 1 4460
0 4462 7 2 2 28926 30078
0 4463 7 1 2 31988 31874
0 4464 5 1 1 4463
0 4465 7 1 2 4461 4464
0 4466 5 1 1 4465
0 4467 7 1 2 26198 30605
0 4468 7 1 2 4466 4467
0 4469 5 1 1 4468
0 4470 7 1 2 4438 4469
0 4471 5 1 1 4470
0 4472 7 1 2 23728 4471
0 4473 5 1 1 4472
0 4474 7 1 2 22461 28020
0 4475 5 1 1 4474
0 4476 7 1 2 27666 4475
0 4477 5 2 1 4476
0 4478 7 1 2 21892 31990
0 4479 5 1 1 4478
0 4480 7 1 2 26354 4479
0 4481 5 1 1 4480
0 4482 7 1 2 26911 4481
0 4483 5 1 1 4482
0 4484 7 2 2 27402 31970
0 4485 7 1 2 22462 31976
0 4486 7 1 2 31992 4485
0 4487 5 1 1 4486
0 4488 7 1 2 4483 4487
0 4489 5 1 1 4488
0 4490 7 1 2 21798 4489
0 4491 5 1 1 4490
0 4492 7 5 2 28138 28786
0 4493 5 1 1 31994
0 4494 7 1 2 21893 25565
0 4495 7 1 2 31995 4494
0 4496 5 1 1 4495
0 4497 7 2 2 28072 29718
0 4498 5 1 1 31999
0 4499 7 1 2 27889 4498
0 4500 5 1 1 4499
0 4501 7 1 2 22188 22463
0 4502 7 1 2 31899 4501
0 4503 7 1 2 4500 4502
0 4504 5 1 1 4503
0 4505 7 1 2 4496 4504
0 4506 5 1 1 4505
0 4507 7 1 2 27762 4506
0 4508 5 1 1 4507
0 4509 7 1 2 4491 4508
0 4510 5 1 1 4509
0 4511 7 1 2 24932 4510
0 4512 5 1 1 4511
0 4513 7 1 2 28080 27993
0 4514 5 1 1 4513
0 4515 7 1 2 27724 4514
0 4516 5 1 1 4515
0 4517 7 1 2 26912 4516
0 4518 5 1 1 4517
0 4519 7 1 2 28094 31996
0 4520 5 1 1 4519
0 4521 7 1 2 4518 4520
0 4522 5 1 1 4521
0 4523 7 3 2 27818 31774
0 4524 5 1 1 32001
0 4525 7 1 2 4522 32002
0 4526 5 1 1 4525
0 4527 7 1 2 4512 4526
0 4528 5 1 1 4527
0 4529 7 1 2 25039 4528
0 4530 5 1 1 4529
0 4531 7 1 2 28501 31997
0 4532 5 2 1 4531
0 4533 7 1 2 30652 31905
0 4534 5 1 1 4533
0 4535 7 1 2 32004 4534
0 4536 5 1 1 4535
0 4537 7 1 2 25566 4536
0 4538 5 1 1 4537
0 4539 7 2 2 26913 27878
0 4540 5 2 1 32006
0 4541 7 1 2 4538 32008
0 4542 5 2 1 4541
0 4543 7 1 2 22627 27763
0 4544 7 1 2 32010 4543
0 4545 5 1 1 4544
0 4546 7 1 2 4530 4545
0 4547 5 1 1 4546
0 4548 7 1 2 23187 4547
0 4549 5 1 1 4548
0 4550 7 1 2 25746 27589
0 4551 7 1 2 31862 4550
0 4552 7 1 2 28787 4551
0 4553 5 1 1 4552
0 4554 7 1 2 27629 695
0 4555 5 1 1 4554
0 4556 7 2 2 25385 4555
0 4557 7 1 2 26762 32012
0 4558 5 1 1 4557
0 4559 7 1 2 4553 4558
0 4560 5 1 1 4559
0 4561 7 1 2 30950 4560
0 4562 5 1 1 4561
0 4563 7 4 2 22851 27403
0 4564 7 2 2 22628 32014
0 4565 7 1 2 32018 31869
0 4566 5 1 1 4565
0 4567 7 1 2 4562 4566
0 4568 5 1 1 4567
0 4569 7 1 2 23188 4568
0 4570 5 1 1 4569
0 4571 7 4 2 22994 29050
0 4572 7 1 2 32020 32015
0 4573 7 1 2 31870 4572
0 4574 5 1 1 4573
0 4575 7 1 2 4570 4574
0 4576 5 1 1 4575
0 4577 7 1 2 27431 4576
0 4578 5 1 1 4577
0 4579 7 2 2 31876 31963
0 4580 7 4 2 24933 29343
0 4581 5 1 1 32026
0 4582 7 1 2 26965 32027
0 4583 7 1 2 32024 4582
0 4584 5 1 1 4583
0 4585 7 1 2 4578 4584
0 4586 5 1 1 4585
0 4587 7 1 2 25905 4586
0 4588 5 1 1 4587
0 4589 7 2 2 27764 29051
0 4590 7 1 2 24934 32009
0 4591 7 1 2 32005 4590
0 4592 5 1 1 4591
0 4593 7 1 2 32030 4592
0 4594 7 1 2 32011 4593
0 4595 5 1 1 4594
0 4596 7 1 2 4588 4595
0 4597 7 1 2 4549 4596
0 4598 5 1 1 4597
0 4599 7 1 2 22522 4598
0 4600 5 1 1 4599
0 4601 7 1 2 23511 4600
0 4602 7 1 2 4473 4601
0 4603 5 1 1 4602
0 4604 7 1 2 24320 29301
0 4605 7 2 2 25776 4604
0 4606 7 1 2 26380 32032
0 4607 5 1 1 4606
0 4608 7 1 2 24793 25040
0 4609 7 1 2 25655 4608
0 4610 7 1 2 27075 4609
0 4611 5 1 1 4610
0 4612 7 1 2 88 4611
0 4613 5 1 1 4612
0 4614 7 1 2 22464 4613
0 4615 5 1 1 4614
0 4616 7 1 2 4607 4615
0 4617 5 1 1 4616
0 4618 7 1 2 21799 4617
0 4619 5 1 1 4618
0 4620 7 1 2 24513 29856
0 4621 7 1 2 25793 4620
0 4622 5 1 1 4621
0 4623 7 1 2 4619 4622
0 4624 5 1 1 4623
0 4625 7 1 2 23189 4624
0 4626 5 1 1 4625
0 4627 7 1 2 30378 32033
0 4628 5 1 1 4627
0 4629 7 1 2 4626 4628
0 4630 5 1 1 4629
0 4631 7 1 2 28139 4630
0 4632 5 1 1 4631
0 4633 7 4 2 25906 28788
0 4634 7 1 2 26763 30393
0 4635 7 1 2 31887 4634
0 4636 7 1 2 32034 4635
0 4637 5 1 1 4636
0 4638 7 1 2 4632 4637
0 4639 5 1 1 4638
0 4640 7 1 2 25567 4639
0 4641 5 1 1 4640
0 4642 7 3 2 26914 28789
0 4643 5 1 1 32038
0 4644 7 9 2 22852 23421
0 4645 5 1 1 32041
0 4646 7 1 2 28355 32042
0 4647 5 1 1 4646
0 4648 7 1 2 4643 4647
0 4649 5 8 1 4648
0 4650 7 3 2 27834 32050
0 4651 7 3 2 23626 27218
0 4652 7 1 2 23190 32061
0 4653 7 1 2 32058 4652
0 4654 5 1 1 4653
0 4655 7 1 2 4641 4654
0 4656 5 1 1 4655
0 4657 7 1 2 21894 4656
0 4658 5 1 1 4657
0 4659 7 3 2 28036 26199
0 4660 7 1 2 27231 32064
0 4661 7 1 2 32051 4660
0 4662 5 1 1 4661
0 4663 7 2 2 25568 28389
0 4664 7 1 2 24682 29446
0 4665 7 1 2 32067 4664
0 4666 7 2 2 24369 24794
0 4667 7 2 2 25656 32069
0 4668 7 3 2 24846 23422
0 4669 7 2 2 29052 32073
0 4670 7 1 2 32071 32076
0 4671 7 1 2 4665 4670
0 4672 5 1 1 4671
0 4673 7 1 2 4662 4672
0 4674 5 1 1 4673
0 4675 7 1 2 27432 4674
0 4676 5 1 1 4675
0 4677 7 1 2 4658 4676
0 4678 5 1 1 4677
0 4679 7 1 2 22629 4678
0 4680 5 1 1 4679
0 4681 7 1 2 27819 32052
0 4682 5 1 1 4681
0 4683 7 1 2 25777 31867
0 4684 5 1 1 4683
0 4685 7 1 2 4682 4684
0 4686 5 1 1 4685
0 4687 7 1 2 22376 4686
0 4688 5 1 1 4687
0 4689 7 2 2 24370 31161
0 4690 7 3 2 22306 27679
0 4691 5 1 1 32080
0 4692 7 1 2 243 4691
0 4693 5 14 1 4692
0 4694 7 4 2 23423 25657
0 4695 7 1 2 24935 32097
0 4696 7 1 2 32083 4695
0 4697 7 1 2 32078 4696
0 4698 5 1 1 4697
0 4699 7 1 2 4688 4698
0 4700 5 1 1 4699
0 4701 7 1 2 21800 4700
0 4702 5 1 1 4701
0 4703 7 2 2 26175 27835
0 4704 7 1 2 32053 32101
0 4705 5 1 1 4704
0 4706 7 1 2 4702 4705
0 4707 5 1 1 4706
0 4708 7 1 2 25041 4707
0 4709 5 1 1 4708
0 4710 7 1 2 22630 32059
0 4711 5 1 1 4710
0 4712 7 1 2 4709 4711
0 4713 5 1 1 4712
0 4714 7 1 2 21895 4713
0 4715 5 1 1 4714
0 4716 7 1 2 30797 32060
0 4717 5 1 1 4716
0 4718 7 1 2 4715 4717
0 4719 5 1 1 4718
0 4720 7 1 2 23191 4719
0 4721 5 1 1 4720
0 4722 7 1 2 28502 32031
0 4723 7 1 2 32054 4722
0 4724 5 1 1 4723
0 4725 7 1 2 23627 4724
0 4726 7 1 2 4721 4725
0 4727 5 1 1 4726
0 4728 7 1 2 26966 30908
0 4729 5 1 1 4728
0 4730 7 1 2 23192 32028
0 4731 5 1 1 4730
0 4732 7 2 2 25158 28195
0 4733 7 1 2 28209 32103
0 4734 5 1 1 4733
0 4735 7 1 2 4731 4734
0 4736 5 1 1 4735
0 4737 7 1 2 23078 4736
0 4738 5 1 1 4737
0 4739 7 1 2 4729 4738
0 4740 5 1 1 4739
0 4741 7 1 2 27730 4740
0 4742 5 1 1 4741
0 4743 7 2 2 21801 30140
0 4744 7 1 2 27836 32105
0 4745 5 1 1 4744
0 4746 7 1 2 4742 4745
0 4747 5 1 1 4746
0 4748 7 1 2 22631 4747
0 4749 5 1 1 4748
0 4750 7 1 2 27433 32021
0 4751 5 2 1 4750
0 4752 7 3 2 21896 27341
0 4753 5 3 1 32109
0 4754 7 1 2 26967 32110
0 4755 5 1 1 4754
0 4756 7 1 2 32107 4755
0 4757 5 1 1 4756
0 4758 7 1 2 27765 4757
0 4759 5 1 1 4758
0 4760 7 1 2 4749 4759
0 4761 5 1 1 4760
0 4762 7 1 2 26058 4761
0 4763 5 1 1 4762
0 4764 7 2 2 22632 27434
0 4765 5 2 1 32115
0 4766 7 1 2 25042 32111
0 4767 5 1 1 4766
0 4768 7 1 2 32117 4767
0 4769 5 1 1 4768
0 4770 7 1 2 23193 4769
0 4771 5 1 1 4770
0 4772 7 1 2 4771 32108
0 4773 5 2 1 4772
0 4774 7 3 2 26331 25907
0 4775 5 1 1 32121
0 4776 7 1 2 32119 32122
0 4777 5 1 1 4776
0 4778 7 1 2 4763 4777
0 4779 5 1 1 4778
0 4780 7 1 2 28140 4779
0 4781 5 1 1 4780
0 4782 7 6 2 23729 25908
0 4783 7 1 2 32039 32124
0 4784 7 1 2 32120 4783
0 4785 5 1 1 4784
0 4786 7 1 2 25569 4785
0 4787 7 1 2 4781 4786
0 4788 5 1 1 4787
0 4789 7 1 2 22523 4788
0 4790 7 1 2 4727 4789
0 4791 5 1 1 4790
0 4792 7 1 2 26038 26626
0 4793 5 1 1 4792
0 4794 7 1 2 26418 4793
0 4795 5 2 1 4794
0 4796 7 1 2 22377 32130
0 4797 5 1 1 4796
0 4798 7 5 2 24371 22465
0 4799 7 1 2 26445 32132
0 4800 5 1 1 4799
0 4801 7 1 2 4797 4800
0 4802 5 1 1 4801
0 4803 7 1 2 21802 4802
0 4804 5 1 1 4803
0 4805 7 1 2 26176 26423
0 4806 5 2 1 4805
0 4807 7 1 2 4804 32137
0 4808 5 1 1 4807
0 4809 7 1 2 29053 4808
0 4810 5 1 1 4809
0 4811 7 3 2 26968 27435
0 4812 5 2 1 32139
0 4813 7 2 2 26403 31510
0 4814 5 1 1 32144
0 4815 7 1 2 32140 32145
0 4816 5 1 1 4815
0 4817 7 1 2 4810 4816
0 4818 5 1 1 4817
0 4819 7 1 2 21897 4818
0 4820 5 1 1 4819
0 4821 7 2 2 22378 22466
0 4822 7 2 2 21803 32146
0 4823 7 3 2 24936 29054
0 4824 5 1 1 32150
0 4825 7 1 2 26404 32151
0 4826 7 1 2 32148 4825
0 4827 5 1 1 4826
0 4828 7 1 2 4820 4827
0 4829 5 1 1 4828
0 4830 7 1 2 32055 4829
0 4831 5 1 1 4830
0 4832 7 1 2 27263 25747
0 4833 7 1 2 28748 4832
0 4834 7 7 2 22905 23424
0 4835 7 2 2 27647 32153
0 4836 7 1 2 29693 32160
0 4837 7 1 2 4833 4836
0 4838 5 1 1 4837
0 4839 7 1 2 4831 4838
0 4840 5 1 1 4839
0 4841 7 1 2 23730 4840
0 4842 5 1 1 4841
0 4843 7 1 2 25770 29302
0 4844 7 1 2 29719 31210
0 4845 7 1 2 4843 4844
0 4846 7 4 2 23425 29425
0 4847 7 3 2 24683 24937
0 4848 7 2 2 25043 32166
0 4849 7 1 2 27254 32169
0 4850 7 1 2 32162 4849
0 4851 7 1 2 4845 4850
0 4852 5 1 1 4851
0 4853 7 1 2 25460 4852
0 4854 7 1 2 4842 4853
0 4855 7 1 2 4791 4854
0 4856 7 1 2 4680 4855
0 4857 5 1 1 4856
0 4858 7 1 2 25229 4857
0 4859 7 1 2 4603 4858
0 4860 5 1 1 4859
0 4861 7 1 2 4375 4860
0 4862 5 1 1 4861
0 4863 7 1 2 22001 4862
0 4864 5 1 1 4863
0 4865 7 6 2 24938 25461
0 4866 7 4 2 24795 32171
0 4867 5 1 1 32177
0 4868 7 1 2 29226 4867
0 4869 5 3 1 4868
0 4870 7 1 2 26915 32181
0 4871 5 1 1 4870
0 4872 7 1 2 28399 31938
0 4873 5 1 1 4872
0 4874 7 1 2 4871 4873
0 4875 5 1 1 4874
0 4876 7 1 2 31071 4875
0 4877 5 1 1 4876
0 4878 7 1 2 549 30114
0 4879 5 2 1 4878
0 4880 7 6 2 22853 25044
0 4881 7 4 2 23512 32186
0 4882 7 3 2 32184 32192
0 4883 7 1 2 26916 29488
0 4884 7 1 2 32196 4883
0 4885 5 1 1 4884
0 4886 7 1 2 4877 4885
0 4887 5 1 1 4886
0 4888 7 1 2 23628 4887
0 4889 5 1 1 4888
0 4890 7 1 2 24796 30565
0 4891 7 1 2 31066 4890
0 4892 7 1 2 31923 4891
0 4893 5 1 1 4892
0 4894 7 1 2 4889 4893
0 4895 5 1 1 4894
0 4896 7 1 2 22307 4895
0 4897 5 1 1 4896
0 4898 7 1 2 30079 30586
0 4899 7 1 2 30606 4898
0 4900 7 1 2 31926 4899
0 4901 5 1 1 4900
0 4902 7 1 2 4897 4901
0 4903 5 1 1 4902
0 4904 7 1 2 27436 4903
0 4905 5 1 1 4904
0 4906 7 3 2 21898 22189
0 4907 7 1 2 30383 32199
0 4908 7 1 2 29623 31601
0 4909 7 1 2 4907 4908
0 4910 7 1 2 30623 4909
0 4911 5 1 1 4910
0 4912 7 1 2 4905 4911
0 4913 5 1 1 4912
0 4914 7 1 2 27766 4913
0 4915 5 1 1 4914
0 4916 7 1 2 29426 31211
0 4917 7 1 2 31836 4916
0 4918 7 2 2 25785 27064
0 4919 7 3 2 24034 30298
0 4920 7 1 2 32202 32204
0 4921 7 1 2 32077 4920
0 4922 7 1 2 4917 4921
0 4923 5 1 1 4922
0 4924 7 1 2 4915 4923
0 4925 5 1 1 4924
0 4926 7 1 2 25230 4925
0 4927 5 1 1 4926
0 4928 7 1 2 4864 4927
0 4929 5 1 1 4928
0 4930 7 1 2 23358 4929
0 4931 5 1 1 4930
0 4932 7 12 2 23935 22002
0 4933 5 3 1 32207
0 4934 7 1 2 30935 32219
0 4935 5 1 1 4934
0 4936 7 2 2 22633 30262
0 4937 5 1 1 32222
0 4938 7 1 2 4935 32223
0 4939 5 1 1 4938
0 4940 7 2 2 22003 27219
0 4941 5 3 1 32224
0 4942 7 1 2 25045 32225
0 4943 5 1 1 4942
0 4944 7 1 2 26177 27375
0 4945 5 1 1 4944
0 4946 7 1 2 23079 4945
0 4947 5 1 1 4946
0 4948 7 1 2 25159 4947
0 4949 7 1 2 4943 4948
0 4950 5 1 1 4949
0 4951 7 2 2 23194 29857
0 4952 5 1 1 32229
0 4953 7 1 2 2313 4952
0 4954 5 1 1 4953
0 4955 7 1 2 21804 4954
0 4956 5 1 1 4955
0 4957 7 1 2 22004 30329
0 4958 5 1 1 4957
0 4959 7 1 2 23936 4958
0 4960 7 1 2 4956 4959
0 4961 7 1 2 4950 4960
0 4962 5 1 1 4961
0 4963 7 2 2 23195 30388
0 4964 5 1 1 32231
0 4965 7 1 2 23080 29636
0 4966 5 3 1 4965
0 4967 7 1 2 32232 32233
0 4968 5 1 1 4967
0 4969 7 2 2 26152 29055
0 4970 5 1 1 32236
0 4971 7 1 2 26976 4970
0 4972 5 1 1 4971
0 4973 7 1 2 23811 4972
0 4974 5 1 1 4973
0 4975 7 1 2 21899 4974
0 4976 7 1 2 4968 4975
0 4977 5 1 1 4976
0 4978 7 1 2 4962 4977
0 4979 5 1 1 4978
0 4980 7 3 2 24035 27376
0 4981 5 7 1 32238
0 4982 7 1 2 25816 32239
0 4983 5 1 1 4982
0 4984 7 1 2 24036 30121
0 4985 5 2 1 4984
0 4986 7 2 2 22005 23196
0 4987 5 1 1 32250
0 4988 7 1 2 32248 4987
0 4989 5 1 1 4988
0 4990 7 1 2 23081 4989
0 4991 5 1 1 4990
0 4992 7 1 2 4983 4991
0 4993 7 1 2 4979 4992
0 4994 5 1 1 4993
0 4995 7 1 2 24590 4994
0 4996 5 1 1 4995
0 4997 7 1 2 3448 30967
0 4998 5 1 1 4997
0 4999 7 1 2 22634 4998
0 5000 5 1 1 4999
0 5001 7 1 2 24591 25820
0 5002 5 1 1 5001
0 5003 7 1 2 27127 30954
0 5004 7 1 2 5002 5003
0 5005 5 1 1 5004
0 5006 7 1 2 5000 5005
0 5007 5 1 1 5006
0 5008 7 3 2 22006 25160
0 5009 5 2 1 32252
0 5010 7 1 2 22995 32255
0 5011 7 1 2 5007 5010
0 5012 5 1 1 5011
0 5013 7 1 2 30115 32249
0 5014 5 1 1 5013
0 5015 7 1 2 27497 30958
0 5016 7 1 2 5014 5015
0 5017 5 1 1 5016
0 5018 7 1 2 25046 29694
0 5019 5 1 1 5018
0 5020 7 4 2 24037 22635
0 5021 5 1 1 32257
0 5022 7 1 2 23197 32258
0 5023 7 1 2 5019 5022
0 5024 5 1 1 5023
0 5025 7 1 2 5017 5024
0 5026 7 1 2 5012 5025
0 5027 7 1 2 4996 5026
0 5028 5 1 1 5027
0 5029 7 1 2 23278 5028
0 5030 5 1 1 5029
0 5031 7 2 2 24592 29285
0 5032 5 1 1 32261
0 5033 7 1 2 31388 32262
0 5034 7 1 2 27349 5033
0 5035 5 1 1 5034
0 5036 7 1 2 5030 5035
0 5037 5 1 1 5036
0 5038 7 1 2 30101 5037
0 5039 5 1 1 5038
0 5040 7 1 2 4939 5039
0 5041 5 1 1 5040
0 5042 7 1 2 24514 5041
0 5043 5 1 1 5042
0 5044 7 1 2 23082 29979
0 5045 5 1 1 5044
0 5046 7 1 2 28228 5045
0 5047 5 1 1 5046
0 5048 7 1 2 23198 5047
0 5049 5 1 1 5048
0 5050 7 6 2 24466 30887
0 5051 5 2 1 32263
0 5052 7 5 2 23812 23083
0 5053 5 2 1 32271
0 5054 7 1 2 32264 32272
0 5055 5 1 1 5054
0 5056 7 1 2 5049 5055
0 5057 5 1 1 5056
0 5058 7 1 2 22636 5057
0 5059 5 1 1 5058
0 5060 7 3 2 23084 29965
0 5061 5 1 1 32278
0 5062 7 1 2 30128 32279
0 5063 5 1 1 5062
0 5064 7 1 2 5059 5063
0 5065 5 1 1 5064
0 5066 7 1 2 24038 5065
0 5067 5 1 1 5066
0 5068 7 1 2 30093 30959
0 5069 7 1 2 29739 5068
0 5070 7 1 2 30143 5069
0 5071 5 1 1 5070
0 5072 7 1 2 5067 5071
0 5073 5 1 1 5072
0 5074 7 1 2 30296 5073
0 5075 5 1 1 5074
0 5076 7 2 2 25658 28212
0 5077 7 3 2 24039 23426
0 5078 7 4 2 23359 23629
0 5079 7 1 2 30707 32286
0 5080 7 1 2 32283 5079
0 5081 7 1 2 32281 5080
0 5082 5 1 1 5081
0 5083 7 1 2 24040 4581
0 5084 5 6 1 5083
0 5085 7 1 2 22524 31265
0 5086 7 1 2 32290 5085
0 5087 5 1 1 5086
0 5088 7 1 2 5082 5087
0 5089 5 1 1 5088
0 5090 7 1 2 24593 5089
0 5091 5 1 1 5090
0 5092 7 2 2 30219 31704
0 5093 5 1 1 32296
0 5094 7 2 2 29872 31154
0 5095 7 1 2 32297 32298
0 5096 5 1 1 5095
0 5097 7 1 2 5091 5096
0 5098 5 1 1 5097
0 5099 7 1 2 25161 5098
0 5100 5 1 1 5099
0 5101 7 1 2 30170 31354
0 5102 7 1 2 32299 5101
0 5103 5 1 1 5102
0 5104 7 1 2 5100 5103
0 5105 5 1 1 5104
0 5106 7 1 2 25047 5105
0 5107 5 1 1 5106
0 5108 7 2 2 22007 30337
0 5109 5 1 1 32300
0 5110 7 1 2 22637 30379
0 5111 5 1 1 5110
0 5112 7 1 2 5109 5111
0 5113 5 1 1 5112
0 5114 7 1 2 31266 5113
0 5115 5 1 1 5114
0 5116 7 1 2 23085 27959
0 5117 7 1 2 27326 28910
0 5118 7 1 2 5116 5117
0 5119 7 1 2 31217 5118
0 5120 5 1 1 5119
0 5121 7 1 2 5115 5120
0 5122 5 1 1 5121
0 5123 7 1 2 27437 5122
0 5124 5 1 1 5123
0 5125 7 1 2 2408 31567
0 5126 7 1 2 30330 5125
0 5127 7 1 2 30102 5126
0 5128 5 1 1 5127
0 5129 7 1 2 2223 5128
0 5130 5 1 1 5129
0 5131 7 1 2 24041 5130
0 5132 5 1 1 5131
0 5133 7 1 2 5124 5132
0 5134 5 1 1 5133
0 5135 7 1 2 29489 5134
0 5136 5 1 1 5135
0 5137 7 1 2 31203 4937
0 5138 5 1 1 5137
0 5139 7 2 2 25048 28213
0 5140 5 1 1 32302
0 5141 7 12 2 21900 24042
0 5142 5 3 1 32304
0 5143 7 1 2 30837 32280
0 5144 5 1 1 5143
0 5145 7 1 2 32316 5144
0 5146 7 1 2 5140 5145
0 5147 5 1 1 5146
0 5148 7 1 2 22525 5147
0 5149 5 1 1 5148
0 5150 7 1 2 22008 30960
0 5151 5 1 1 5150
0 5152 7 1 2 5149 5151
0 5153 5 1 1 5152
0 5154 7 1 2 5138 5153
0 5155 5 1 1 5154
0 5156 7 1 2 5136 5155
0 5157 7 1 2 5107 5156
0 5158 7 1 2 5075 5157
0 5159 7 1 2 5043 5158
0 5160 5 1 1 5159
0 5161 7 1 2 28790 5160
0 5162 5 1 1 5161
0 5163 7 1 2 307 30183
0 5164 5 16 1 5163
0 5165 7 2 2 27621 32319
0 5166 5 1 1 32335
0 5167 7 1 2 26892 30184
0 5168 5 10 1 5167
0 5169 7 3 2 25659 32337
0 5170 7 1 2 26059 26237
0 5171 7 1 2 32347 5170
0 5172 5 1 1 5171
0 5173 7 1 2 5166 5172
0 5174 5 1 1 5173
0 5175 7 1 2 27498 5174
0 5176 5 1 1 5175
0 5177 7 1 2 2368 30185
0 5178 5 3 1 5177
0 5179 7 4 2 25660 32350
0 5180 7 3 2 27128 26060
0 5181 7 1 2 23630 32357
0 5182 7 1 2 32353 5181
0 5183 5 1 1 5182
0 5184 7 1 2 5176 5183
0 5185 5 1 1 5184
0 5186 7 1 2 23086 5185
0 5187 5 1 1 5186
0 5188 7 6 2 22996 28557
0 5189 5 1 1 32360
0 5190 7 1 2 32361 32336
0 5191 5 1 1 5190
0 5192 7 1 2 5187 5191
0 5193 5 1 1 5192
0 5194 7 1 2 29447 5193
0 5195 5 1 1 5194
0 5196 7 1 2 23087 32320
0 5197 7 1 2 30490 5196
0 5198 5 1 1 5197
0 5199 7 1 2 5195 5198
0 5200 5 1 1 5199
0 5201 7 1 2 29882 31181
0 5202 7 1 2 5200 5201
0 5203 5 1 1 5202
0 5204 7 1 2 26893 2170
0 5205 5 6 1 5204
0 5206 7 2 2 31140 32366
0 5207 7 1 2 30399 32372
0 5208 5 1 1 5207
0 5209 7 2 2 22854 29490
0 5210 7 2 2 25231 23731
0 5211 7 1 2 31802 32376
0 5212 7 1 2 32374 5211
0 5213 7 1 2 30656 5212
0 5214 5 1 1 5213
0 5215 7 1 2 5208 5214
0 5216 5 1 1 5215
0 5217 7 1 2 22009 29879
0 5218 7 1 2 5216 5217
0 5219 5 1 1 5218
0 5220 7 1 2 5203 5219
0 5221 7 1 2 5162 5220
0 5222 5 1 1 5221
0 5223 7 1 2 25909 5222
0 5224 5 1 1 5223
0 5225 7 2 2 22997 28719
0 5226 5 1 1 32378
0 5227 7 4 2 24043 32321
0 5228 7 1 2 32379 32380
0 5229 5 1 1 5228
0 5230 7 1 2 27960 28640
0 5231 7 2 2 28764 5230
0 5232 5 1 1 32384
0 5233 7 1 2 5229 5232
0 5234 5 1 1 5233
0 5235 7 1 2 27499 5234
0 5236 5 1 1 5235
0 5237 7 3 2 25462 31854
0 5238 7 4 2 24467 22855
0 5239 5 2 1 32389
0 5240 7 5 2 22308 24594
0 5241 7 1 2 30159 32395
0 5242 7 1 2 32390 5241
0 5243 7 1 2 32386 5242
0 5244 5 1 1 5243
0 5245 7 1 2 5236 5244
0 5246 5 1 1 5245
0 5247 7 1 2 29589 5246
0 5248 5 1 1 5247
0 5249 7 3 2 24797 26940
0 5250 5 1 1 32400
0 5251 7 1 2 29227 5250
0 5252 5 3 1 5251
0 5253 7 1 2 29720 32403
0 5254 5 1 1 5253
0 5255 7 1 2 28699 5254
0 5256 5 2 1 5255
0 5257 7 1 2 27129 32406
0 5258 5 1 1 5257
0 5259 7 3 2 25570 28572
0 5260 7 1 2 29193 32408
0 5261 5 1 1 5260
0 5262 7 1 2 5258 5261
0 5263 5 1 1 5262
0 5264 7 1 2 27500 32381
0 5265 7 1 2 5263 5264
0 5266 5 1 1 5265
0 5267 7 1 2 27327 28596
0 5268 5 1 1 5267
0 5269 7 1 2 23199 29157
0 5270 5 1 1 5269
0 5271 7 1 2 5268 5270
0 5272 5 1 1 5271
0 5273 7 1 2 25846 32387
0 5274 7 1 2 5272 5273
0 5275 5 1 1 5274
0 5276 7 1 2 5266 5275
0 5277 5 1 1 5276
0 5278 7 1 2 23937 5277
0 5279 5 1 1 5278
0 5280 7 1 2 22998 32385
0 5281 5 1 1 5280
0 5282 7 1 2 24515 32382
0 5283 7 1 2 32407 5282
0 5284 5 1 1 5283
0 5285 7 1 2 5281 5284
0 5286 7 1 2 5279 5285
0 5287 5 1 1 5286
0 5288 7 1 2 29350 5287
0 5289 5 1 1 5288
0 5290 7 1 2 5248 5289
0 5291 5 1 1 5290
0 5292 7 1 2 23088 5291
0 5293 5 1 1 5292
0 5294 7 2 2 28480 31457
0 5295 5 2 1 32411
0 5296 7 1 2 24468 32412
0 5297 5 1 1 5296
0 5298 7 2 2 24516 27264
0 5299 5 1 1 32415
0 5300 7 1 2 29286 32416
0 5301 5 1 1 5300
0 5302 7 1 2 5297 5301
0 5303 5 1 1 5302
0 5304 7 1 2 28720 5303
0 5305 5 1 1 5304
0 5306 7 3 2 24595 25847
0 5307 7 1 2 27232 28755
0 5308 7 1 2 32417 5307
0 5309 5 1 1 5308
0 5310 7 2 2 29194 29287
0 5311 7 1 2 27265 27994
0 5312 7 1 2 32420 5311
0 5313 5 1 1 5312
0 5314 7 1 2 5309 5313
0 5315 5 1 1 5314
0 5316 7 1 2 28148 5315
0 5317 5 1 1 5316
0 5318 7 1 2 5305 5317
0 5319 5 1 1 5318
0 5320 7 1 2 23813 5319
0 5321 5 1 1 5320
0 5322 7 2 2 24044 27266
0 5323 7 1 2 29662 32422
0 5324 7 1 2 28721 5323
0 5325 5 1 1 5324
0 5326 7 1 2 25049 31382
0 5327 5 1 1 5326
0 5328 7 1 2 24045 5327
0 5329 5 1 1 5328
0 5330 7 1 2 26262 28655
0 5331 7 1 2 5329 5330
0 5332 5 1 1 5331
0 5333 7 1 2 5325 5332
0 5334 5 1 1 5333
0 5335 7 1 2 24517 5334
0 5336 5 1 1 5335
0 5337 7 2 2 22526 23200
0 5338 7 1 2 24046 27057
0 5339 7 1 2 32424 5338
0 5340 7 1 2 28656 5339
0 5341 5 1 1 5340
0 5342 7 1 2 5336 5341
0 5343 7 1 2 5321 5342
0 5344 5 1 1 5343
0 5345 7 1 2 23279 5344
0 5346 5 1 1 5345
0 5347 7 1 2 27501 28722
0 5348 5 1 1 5347
0 5349 7 4 2 25571 27130
0 5350 7 1 2 29030 32426
0 5351 5 1 1 5350
0 5352 7 1 2 5348 5351
0 5353 5 1 1 5352
0 5354 7 1 2 26897 29846
0 5355 7 1 2 5353 5354
0 5356 5 1 1 5355
0 5357 7 1 2 5346 5356
0 5358 7 1 2 5293 5357
0 5359 5 1 1 5358
0 5360 7 1 2 27767 5359
0 5361 5 1 1 5360
0 5362 7 1 2 27131 32351
0 5363 5 1 1 5362
0 5364 7 4 2 27856 32338
0 5365 5 2 1 32430
0 5366 7 1 2 5363 32434
0 5367 5 4 1 5366
0 5368 7 1 2 28657 32436
0 5369 5 1 1 5368
0 5370 7 4 2 22309 31911
0 5371 5 1 1 32440
0 5372 7 2 2 24321 30628
0 5373 5 1 1 32444
0 5374 7 1 2 5371 5373
0 5375 5 6 1 5374
0 5376 7 1 2 32446 32427
0 5377 7 1 2 32431 5376
0 5378 5 1 1 5377
0 5379 7 1 2 5369 5378
0 5380 5 1 1 5379
0 5381 7 2 2 24847 29244
0 5382 7 1 2 29309 32452
0 5383 7 1 2 5380 5382
0 5384 5 1 1 5383
0 5385 7 1 2 5361 5384
0 5386 5 1 1 5385
0 5387 7 1 2 28911 5386
0 5388 5 1 1 5387
0 5389 7 1 2 27220 28873
0 5390 5 1 1 5389
0 5391 7 1 2 23513 30802
0 5392 5 1 1 5391
0 5393 7 1 2 5390 5392
0 5394 5 1 1 5393
0 5395 7 1 2 29562 5394
0 5396 5 1 1 5395
0 5397 7 1 2 28867 32172
0 5398 7 1 2 30764 5397
0 5399 5 1 1 5398
0 5400 7 1 2 5396 5399
0 5401 5 1 1 5400
0 5402 7 1 2 27768 5401
0 5403 5 1 1 5402
0 5404 7 1 2 2512 5403
0 5405 5 1 1 5404
0 5406 7 1 2 32367 5405
0 5407 5 1 1 5406
0 5408 7 1 2 29590 2760
0 5409 5 6 1 5408
0 5410 7 2 2 24939 32454
0 5411 5 1 1 32460
0 5412 7 1 2 22638 27171
0 5413 5 1 1 5412
0 5414 7 1 2 5411 5413
0 5415 5 1 1 5414
0 5416 7 1 2 30171 5415
0 5417 5 1 1 5416
0 5418 7 1 2 30220 29624
0 5419 5 1 1 5418
0 5420 7 1 2 2624 5419
0 5421 5 1 1 5420
0 5422 7 1 2 29491 5421
0 5423 5 1 1 5422
0 5424 7 1 2 30221 29563
0 5425 5 1 1 5424
0 5426 7 1 2 22999 30833
0 5427 5 1 1 5426
0 5428 7 1 2 5425 5427
0 5429 7 1 2 5423 5428
0 5430 5 1 1 5429
0 5431 7 1 2 25162 5430
0 5432 5 1 1 5431
0 5433 7 1 2 5417 5432
0 5434 5 1 1 5433
0 5435 7 1 2 23514 26352
0 5436 7 1 2 5434 5435
0 5437 5 1 1 5436
0 5438 7 1 2 5407 5437
0 5439 5 1 1 5438
0 5440 7 1 2 25050 5439
0 5441 5 1 1 5440
0 5442 7 1 2 29210 30107
0 5443 5 1 1 5442
0 5444 7 1 2 28573 30607
0 5445 5 2 1 5444
0 5446 7 1 2 29056 29211
0 5447 5 1 1 5446
0 5448 7 1 2 32462 5447
0 5449 5 1 1 5448
0 5450 7 1 2 29752 5449
0 5451 5 1 1 5450
0 5452 7 1 2 5443 5451
0 5453 5 1 1 5452
0 5454 7 1 2 29492 5453
0 5455 5 1 1 5454
0 5456 7 1 2 30116 4824
0 5457 5 1 1 5456
0 5458 7 1 2 27438 5457
0 5459 5 1 1 5458
0 5460 7 1 2 684 3924
0 5461 5 1 1 5460
0 5462 7 1 2 25163 5461
0 5463 5 1 1 5462
0 5464 7 1 2 5459 5463
0 5465 5 1 1 5464
0 5466 7 1 2 29212 5465
0 5467 5 1 1 5466
0 5468 7 1 2 5455 5467
0 5469 5 1 1 5468
0 5470 7 1 2 22310 5469
0 5471 5 1 1 5470
0 5472 7 1 2 30519 30804
0 5473 5 1 1 5472
0 5474 7 1 2 5471 5473
0 5475 5 1 1 5474
0 5476 7 1 2 23631 5475
0 5477 5 1 1 5476
0 5478 7 1 2 30669 5477
0 5479 5 1 1 5478
0 5480 7 1 2 26200 32377
0 5481 7 1 2 5479 5480
0 5482 5 1 1 5481
0 5483 7 1 2 5441 5482
0 5484 5 1 1 5483
0 5485 7 1 2 22010 5484
0 5486 5 1 1 5485
0 5487 7 1 2 30520 30608
0 5488 5 1 1 5487
0 5489 7 1 2 29057 30537
0 5490 5 1 1 5489
0 5491 7 1 2 5488 5490
0 5492 5 1 1 5491
0 5493 7 1 2 24940 5492
0 5494 5 1 1 5493
0 5495 7 3 2 22639 30538
0 5496 5 1 1 32464
0 5497 7 1 2 23201 32465
0 5498 5 1 1 5497
0 5499 7 1 2 5494 5498
0 5500 5 1 1 5499
0 5501 7 1 2 27439 5500
0 5502 5 1 1 5501
0 5503 7 1 2 22311 27172
0 5504 7 1 2 32197 5503
0 5505 5 1 1 5504
0 5506 7 1 2 5502 5505
0 5507 5 1 1 5506
0 5508 7 1 2 22527 5507
0 5509 5 1 1 5508
0 5510 7 1 2 28560 29386
0 5511 7 1 2 28765 5510
0 5512 5 1 1 5511
0 5513 7 1 2 5509 5512
0 5514 5 1 1 5513
0 5515 7 1 2 21901 5514
0 5516 5 1 1 5515
0 5517 7 1 2 28424 31355
0 5518 5 1 1 5517
0 5519 7 1 2 22312 26304
0 5520 7 1 2 29753 5519
0 5521 7 1 2 32193 5520
0 5522 7 1 2 5518 5521
0 5523 5 1 1 5522
0 5524 7 1 2 5516 5523
0 5525 5 1 1 5524
0 5526 7 4 2 25232 23632
0 5527 7 1 2 27769 32467
0 5528 7 1 2 5525 5527
0 5529 5 1 1 5528
0 5530 7 1 2 5486 5529
0 5531 5 1 1 5530
0 5532 7 1 2 29873 5531
0 5533 5 1 1 5532
0 5534 7 1 2 28239 30319
0 5535 7 1 2 31552 5534
0 5536 5 1 1 5535
0 5537 7 3 2 24518 30695
0 5538 7 21 2 23427 23515
0 5539 7 2 2 31617 32474
0 5540 7 1 2 25572 32495
0 5541 7 1 2 32471 5540
0 5542 5 1 1 5541
0 5543 7 1 2 5536 5542
0 5544 5 1 1 5543
0 5545 7 1 2 21902 27863
0 5546 5 16 1 5545
0 5547 7 3 2 22640 32497
0 5548 7 1 2 27770 32513
0 5549 5 1 1 5548
0 5550 7 2 2 25661 30917
0 5551 7 3 2 22011 24596
0 5552 5 1 1 32518
0 5553 7 1 2 5552 5021
0 5554 5 10 1 5553
0 5555 7 1 2 26105 32521
0 5556 7 1 2 32516 5555
0 5557 5 1 1 5556
0 5558 7 1 2 5549 5557
0 5559 5 2 1 5558
0 5560 7 1 2 5544 32531
0 5561 5 1 1 5560
0 5562 7 1 2 31546 31553
0 5563 5 1 1 5562
0 5564 7 1 2 2853 5563
0 5565 5 1 1 5564
0 5566 7 5 2 22012 24519
0 5567 5 2 1 32533
0 5568 7 2 2 24047 30571
0 5569 5 1 1 32540
0 5570 7 1 2 28214 32541
0 5571 5 3 1 5570
0 5572 7 1 2 23089 32542
0 5573 5 2 1 5572
0 5574 7 3 2 32538 32545
0 5575 5 3 1 32547
0 5576 7 1 2 27771 32550
0 5577 5 1 1 5576
0 5578 7 3 2 24048 24372
0 5579 7 1 2 29649 32553
0 5580 7 1 2 32453 5579
0 5581 5 1 1 5580
0 5582 7 1 2 5577 5581
0 5583 7 3 2 23000 25662
0 5584 7 2 2 22013 32556
0 5585 7 2 2 23938 32559
0 5586 7 1 2 26106 32561
0 5587 5 2 1 5586
0 5588 7 1 2 3732 32563
0 5589 5 1 1 5588
0 5590 7 1 2 27132 5589
0 5591 5 1 1 5590
0 5592 7 1 2 22528 27837
0 5593 5 2 1 5592
0 5594 7 2 2 24373 29427
0 5595 7 1 2 24848 26043
0 5596 7 1 2 32567 5595
0 5597 5 1 1 5596
0 5598 7 1 2 32565 5597
0 5599 5 1 1 5598
0 5600 7 1 2 24049 5599
0 5601 5 1 1 5600
0 5602 7 1 2 5591 5601
0 5603 5 1 1 5602
0 5604 7 1 2 25051 5603
0 5605 5 1 1 5604
0 5606 7 2 2 24520 25052
0 5607 5 2 1 32569
0 5608 7 1 2 31533 32571
0 5609 5 18 1 5608
0 5610 7 2 2 21903 24374
0 5611 7 2 2 24050 32591
0 5612 7 1 2 27578 32593
0 5613 5 1 1 5612
0 5614 7 1 2 27849 5613
0 5615 5 1 1 5614
0 5616 7 1 2 27173 5615
0 5617 5 1 1 5616
0 5618 7 6 2 22014 24375
0 5619 7 3 2 28067 32595
0 5620 7 1 2 28215 32601
0 5621 5 1 1 5620
0 5622 7 1 2 4524 5621
0 5623 7 1 2 5617 5622
0 5624 5 1 1 5623
0 5625 7 1 2 32573 5624
0 5626 5 1 1 5625
0 5627 7 1 2 5605 5626
0 5628 7 1 2 5582 5627
0 5629 5 1 1 5628
0 5630 7 1 2 5565 5629
0 5631 5 1 1 5630
0 5632 7 1 2 5561 5631
0 5633 5 1 1 5632
0 5634 7 1 2 28791 5633
0 5635 5 1 1 5634
0 5636 7 1 2 5533 5635
0 5637 7 1 2 5388 5636
0 5638 7 1 2 5224 5637
0 5639 5 1 1 5638
0 5640 7 1 2 28526 5639
0 5641 5 1 1 5640
0 5642 7 9 2 25573 30918
0 5643 7 1 2 26107 32604
0 5644 5 2 1 5643
0 5645 7 9 2 23633 25910
0 5646 7 3 2 23939 29778
0 5647 5 11 1 32624
0 5648 7 2 2 32615 32627
0 5649 5 1 1 32638
0 5650 7 1 2 32613 5649
0 5651 5 1 1 5650
0 5652 7 1 2 26061 5651
0 5653 5 1 1 5652
0 5654 7 7 2 23634 32628
0 5655 7 1 2 27687 32640
0 5656 5 1 1 5655
0 5657 7 1 2 5653 5656
0 5658 5 1 1 5657
0 5659 7 1 2 25663 5658
0 5660 5 1 1 5659
0 5661 7 2 2 25574 26001
0 5662 5 1 1 32647
0 5663 7 1 2 5660 5662
0 5664 5 2 1 5663
0 5665 7 1 2 32522 32649
0 5666 5 1 1 5665
0 5667 7 1 2 28021 31024
0 5668 5 1 1 5667
0 5669 7 1 2 27667 5668
0 5670 5 1 1 5669
0 5671 7 1 2 23814 5670
0 5672 5 1 1 5671
0 5673 7 3 2 21805 26153
0 5674 5 1 1 32651
0 5675 7 1 2 28022 32652
0 5676 5 1 1 5675
0 5677 7 1 2 27670 5676
0 5678 7 1 2 5672 5677
0 5679 5 1 1 5678
0 5680 7 1 2 23940 5679
0 5681 5 1 1 5680
0 5682 7 2 2 22379 23001
0 5683 7 1 2 27820 32654
0 5684 7 1 2 29189 5683
0 5685 5 1 1 5684
0 5686 7 1 2 5681 5685
0 5687 5 1 1 5686
0 5688 7 1 2 22641 5687
0 5689 5 1 1 5688
0 5690 7 1 2 21806 31991
0 5691 5 1 1 5690
0 5692 7 2 2 27404 32147
0 5693 7 1 2 26505 32656
0 5694 5 1 1 5693
0 5695 7 1 2 5691 5694
0 5696 5 1 1 5695
0 5697 7 1 2 30268 5696
0 5698 5 1 1 5697
0 5699 7 1 2 28023 29538
0 5700 5 1 1 5699
0 5701 7 1 2 5698 5700
0 5702 5 1 1 5701
0 5703 7 1 2 24597 5702
0 5704 5 1 1 5703
0 5705 7 1 2 27603 31025
0 5706 5 1 1 5705
0 5707 7 1 2 27630 5706
0 5708 5 1 1 5707
0 5709 7 1 2 23815 5708
0 5710 5 1 1 5709
0 5711 7 1 2 27604 32653
0 5712 5 1 1 5711
0 5713 7 1 2 27633 5712
0 5714 7 1 2 5710 5713
0 5715 5 1 1 5714
0 5716 7 1 2 23941 5715
0 5717 5 1 1 5716
0 5718 7 1 2 22642 30492
0 5719 7 1 2 5717 5718
0 5720 5 1 1 5719
0 5721 7 1 2 27440 27605
0 5722 5 1 1 5721
0 5723 7 1 2 26332 28095
0 5724 5 1 1 5723
0 5725 7 1 2 5722 5724
0 5726 5 1 1 5725
0 5727 7 1 2 30269 5726
0 5728 5 1 1 5727
0 5729 7 1 2 27606 29539
0 5730 5 1 1 5729
0 5731 7 1 2 24598 5730
0 5732 7 1 2 5728 5731
0 5733 5 1 1 5732
0 5734 7 1 2 25911 5733
0 5735 7 1 2 5720 5734
0 5736 5 1 1 5735
0 5737 7 1 2 5704 5736
0 5738 7 1 2 5689 5737
0 5739 7 1 2 5666 5738
0 5740 5 1 1 5739
0 5741 7 4 2 24521 30449
0 5742 7 1 2 26839 32658
0 5743 5 1 1 5742
0 5744 7 1 2 26845 29082
0 5745 5 1 1 5744
0 5746 7 1 2 5743 5745
0 5747 5 1 1 5746
0 5748 7 1 2 28527 5747
0 5749 7 1 2 5740 5748
0 5750 5 1 1 5749
0 5751 7 1 2 22015 23002
0 5752 5 2 1 5751
0 5753 7 1 2 21904 31026
0 5754 5 1 1 5753
0 5755 7 1 2 32662 5754
0 5756 5 1 1 5755
0 5757 7 1 2 23816 5756
0 5758 5 1 1 5757
0 5759 7 1 2 28196 28207
0 5760 5 2 1 5759
0 5761 7 1 2 32220 32664
0 5762 7 1 2 5758 5761
0 5763 5 3 1 5762
0 5764 7 1 2 26405 32666
0 5765 5 1 1 5764
0 5766 7 1 2 22016 28229
0 5767 5 9 1 5766
0 5768 7 1 2 26627 32291
0 5769 7 1 2 32669 5768
0 5770 5 1 1 5769
0 5771 7 1 2 5765 5770
0 5772 5 2 1 5771
0 5773 7 1 2 24376 32678
0 5774 5 1 1 5773
0 5775 7 3 2 23635 32667
0 5776 7 2 2 25880 32680
0 5777 5 1 1 32683
0 5778 7 1 2 5774 5777
0 5779 5 2 1 5778
0 5780 7 1 2 32574 32685
0 5781 5 1 1 5780
0 5782 7 3 2 22380 26464
0 5783 5 2 1 32687
0 5784 7 1 2 24469 26628
0 5785 5 1 1 5784
0 5786 7 1 2 26419 5785
0 5787 5 4 1 5786
0 5788 7 1 2 24377 32692
0 5789 5 1 1 5788
0 5790 7 1 2 32690 5789
0 5791 5 4 1 5790
0 5792 7 4 2 23817 32208
0 5793 7 2 2 29387 32700
0 5794 5 2 1 32704
0 5795 7 1 2 32696 32705
0 5796 5 1 1 5795
0 5797 7 3 2 27441 31651
0 5798 5 1 1 32708
0 5799 7 1 2 27321 32709
0 5800 5 1 1 5799
0 5801 7 1 2 25912 29787
0 5802 7 1 2 29405 5801
0 5803 5 1 1 5802
0 5804 7 1 2 5800 5803
0 5805 5 1 1 5804
0 5806 7 1 2 32305 5805
0 5807 5 1 1 5806
0 5808 7 1 2 5796 5807
0 5809 7 1 2 5781 5808
0 5810 5 1 1 5809
0 5811 7 1 2 26062 5810
0 5812 5 1 1 5811
0 5813 7 4 2 24051 29004
0 5814 5 1 1 32711
0 5815 7 2 2 29788 32712
0 5816 5 2 1 32715
0 5817 7 2 2 3054 5674
0 5818 5 19 1 32719
0 5819 7 1 2 32721 32575
0 5820 5 1 1 5819
0 5821 7 1 2 32717 5820
0 5822 5 1 1 5821
0 5823 7 1 2 21905 5822
0 5824 5 1 1 5823
0 5825 7 1 2 21906 29789
0 5826 5 2 1 5825
0 5827 7 1 2 22017 32740
0 5828 5 1 1 5827
0 5829 7 1 2 23942 28425
0 5830 5 1 1 5829
0 5831 7 1 2 5828 5830
0 5832 5 1 1 5831
0 5833 7 1 2 32576 5832
0 5834 5 1 1 5833
0 5835 7 1 2 32706 5834
0 5836 7 1 2 5824 5835
0 5837 5 3 1 5836
0 5838 7 1 2 27700 32742
0 5839 5 1 1 5838
0 5840 7 1 2 5812 5839
0 5841 5 1 1 5840
0 5842 7 1 2 25664 5841
0 5843 5 1 1 5842
0 5844 7 1 2 30919 32577
0 5845 5 1 1 5844
0 5846 7 2 2 21907 29893
0 5847 5 1 1 32745
0 5848 7 1 2 27442 32746
0 5849 5 2 1 5848
0 5850 7 1 2 29005 32306
0 5851 5 2 1 5850
0 5852 7 5 2 22018 29111
0 5853 5 1 1 32751
0 5854 7 2 2 23943 32752
0 5855 5 2 1 32756
0 5856 7 1 2 32749 32758
0 5857 7 2 2 32747 5856
0 5858 5 3 1 32760
0 5859 7 1 2 5845 32761
0 5860 5 3 1 5859
0 5861 7 1 2 28117 32765
0 5862 5 1 1 5861
0 5863 7 4 2 23090 28106
0 5864 5 1 1 32768
0 5865 7 1 2 29754 29493
0 5866 5 1 1 5865
0 5867 7 1 2 24052 30643
0 5868 7 1 2 5866 5867
0 5869 5 1 1 5868
0 5870 7 1 2 32769 5869
0 5871 5 1 1 5870
0 5872 7 1 2 5862 5871
0 5873 5 1 1 5872
0 5874 7 1 2 23732 5873
0 5875 5 1 1 5874
0 5876 7 1 2 5843 5875
0 5877 5 1 1 5876
0 5878 7 2 2 30496 29883
0 5879 5 1 1 32772
0 5880 7 1 2 22643 26846
0 5881 5 1 1 5880
0 5882 7 1 2 5879 5881
0 5883 5 1 1 5882
0 5884 7 1 2 28528 5883
0 5885 7 1 2 5877 5884
0 5886 5 1 1 5885
0 5887 7 1 2 5750 5886
0 5888 7 1 2 5641 5887
0 5889 7 1 2 1057 28333
0 5890 5 1 1 5889
0 5891 7 1 2 32322 5890
0 5892 5 1 1 5891
0 5893 7 11 2 22190 25233
0 5894 7 1 2 22906 23202
0 5895 7 1 2 32396 5894
0 5896 7 1 2 32774 5895
0 5897 7 4 2 25386 29252
0 5898 7 2 2 22381 31955
0 5899 7 1 2 32785 32789
0 5900 7 1 2 5896 5899
0 5901 5 1 1 5900
0 5902 7 1 2 5892 5901
0 5903 5 1 1 5902
0 5904 7 1 2 24522 5903
0 5905 5 1 1 5904
0 5906 7 1 2 22907 26898
0 5907 7 1 2 28099 5906
0 5908 7 1 2 31931 5907
0 5909 5 1 1 5908
0 5910 7 1 2 5905 5909
0 5911 5 1 1 5910
0 5912 7 1 2 23944 5911
0 5913 5 1 1 5912
0 5914 7 3 2 25053 27961
0 5915 5 1 1 32791
0 5916 7 1 2 23203 3103
0 5917 5 1 1 5916
0 5918 7 1 2 24599 326
0 5919 7 1 2 5917 5918
0 5920 5 1 1 5919
0 5921 7 1 2 5915 5920
0 5922 5 1 1 5921
0 5923 7 1 2 26787 28251
0 5924 7 1 2 29379 5923
0 5925 7 1 2 5922 5924
0 5926 5 1 1 5925
0 5927 7 1 2 5913 5926
0 5928 5 1 1 5927
0 5929 7 1 2 23003 5928
0 5930 5 1 1 5929
0 5931 7 2 2 28481 31927
0 5932 7 2 2 23280 27133
0 5933 7 1 2 26201 32796
0 5934 7 1 2 32794 5933
0 5935 5 1 1 5934
0 5936 7 1 2 22908 27502
0 5937 7 1 2 31928 5936
0 5938 5 1 1 5937
0 5939 7 2 2 26764 27134
0 5940 7 1 2 26629 30241
0 5941 7 1 2 32798 5940
0 5942 5 1 1 5941
0 5943 7 1 2 5938 5942
0 5944 5 1 1 5943
0 5945 7 1 2 22382 5944
0 5946 5 1 1 5945
0 5947 7 1 2 26765 25875
0 5948 7 1 2 30242 5947
0 5949 7 1 2 32428 5948
0 5950 5 1 1 5949
0 5951 7 1 2 5946 5950
0 5952 5 1 1 5951
0 5953 7 1 2 29995 32323
0 5954 7 1 2 5952 5953
0 5955 5 1 1 5954
0 5956 7 1 2 5935 5955
0 5957 5 1 1 5956
0 5958 7 1 2 28792 5957
0 5959 5 1 1 5958
0 5960 7 2 2 28407 28482
0 5961 7 1 2 28290 32800
0 5962 5 1 1 5961
0 5963 7 4 2 23516 31579
0 5964 7 1 2 26917 29656
0 5965 7 1 2 32802 5964
0 5966 5 1 1 5965
0 5967 7 1 2 5962 5966
0 5968 5 1 1 5967
0 5969 7 1 2 28381 31855
0 5970 7 1 2 5968 5969
0 5971 5 1 1 5970
0 5972 7 1 2 5959 5971
0 5973 7 1 2 5930 5972
0 5974 5 1 1 5973
0 5975 7 1 2 24053 5974
0 5976 5 1 1 5975
0 5977 7 2 2 25463 28483
0 5978 7 4 2 27135 32806
0 5979 5 1 1 32808
0 5980 7 1 2 25748 32043
0 5981 5 1 1 5980
0 5982 7 1 2 4385 5981
0 5983 5 1 1 5982
0 5984 7 1 2 32809 5983
0 5985 5 1 1 5984
0 5986 7 2 2 22856 25387
0 5987 7 1 2 26766 32812
0 5988 7 1 2 32803 5987
0 5989 5 1 1 5988
0 5990 7 1 2 5985 5989
0 5991 5 1 1 5990
0 5992 7 1 2 30869 5991
0 5993 5 1 1 5992
0 5994 7 1 2 30021 32801
0 5995 5 1 1 5994
0 5996 7 1 2 5993 5995
0 5997 5 1 1 5996
0 5998 7 1 2 22313 5997
0 5999 5 1 1 5998
0 6000 7 2 2 27136 28705
0 6001 7 1 2 32814 32795
0 6002 5 1 1 6001
0 6003 7 1 2 5999 6002
0 6004 5 1 1 6003
0 6005 7 1 2 29448 6004
0 6006 5 1 1 6005
0 6007 7 1 2 26767 28360
0 6008 7 1 2 29202 6007
0 6009 7 1 2 32804 6008
0 6010 5 1 1 6009
0 6011 7 1 2 6006 6010
0 6012 5 1 1 6011
0 6013 7 2 2 22909 23281
0 6014 7 1 2 22383 29591
0 6015 7 1 2 32816 6014
0 6016 7 1 2 6012 6015
0 6017 5 1 1 6016
0 6018 7 1 2 5976 6017
0 6019 5 1 1 6018
0 6020 7 1 2 23733 6019
0 6021 5 1 1 6020
0 6022 7 2 2 27300 27838
0 6023 5 1 1 32818
0 6024 7 1 2 32324 32819
0 6025 5 2 1 6024
0 6026 7 3 2 26614 32348
0 6027 7 2 2 29303 32822
0 6028 5 1 1 32825
0 6029 7 1 2 24470 32826
0 6030 5 1 1 6029
0 6031 7 1 2 32820 6030
0 6032 5 1 1 6031
0 6033 7 1 2 23945 6032
0 6034 5 1 1 6033
0 6035 7 7 2 23734 32325
0 6036 7 3 2 22910 32827
0 6037 7 2 2 29182 32834
0 6038 7 1 2 27301 32837
0 6039 5 1 1 6038
0 6040 7 1 2 6034 6039
0 6041 5 1 1 6040
0 6042 7 1 2 23818 6041
0 6043 5 1 1 6042
0 6044 7 2 2 28197 29866
0 6045 7 2 2 29592 32839
0 6046 7 7 2 27772 32326
0 6047 5 2 1 32843
0 6048 7 1 2 32841 32844
0 6049 5 1 1 6048
0 6050 7 1 2 6043 6049
0 6051 5 2 1 6050
0 6052 7 1 2 31998 32852
0 6053 5 1 1 6052
0 6054 7 1 2 26490 32823
0 6055 5 1 1 6054
0 6056 7 1 2 32850 6055
0 6057 5 3 1 6056
0 6058 7 1 2 23819 32854
0 6059 5 1 1 6058
0 6060 7 1 2 32821 6059
0 6061 5 1 1 6060
0 6062 7 1 2 24523 6061
0 6063 5 1 1 6062
0 6064 7 1 2 27210 32845
0 6065 5 1 1 6064
0 6066 7 1 2 6063 6065
0 6067 5 1 1 6066
0 6068 7 1 2 23946 6067
0 6069 5 1 1 6068
0 6070 7 1 2 29810 32846
0 6071 5 1 1 6070
0 6072 7 1 2 6069 6071
0 6073 5 1 1 6072
0 6074 7 2 2 24798 31906
0 6075 5 1 1 32857
0 6076 7 1 2 6073 32858
0 6077 5 1 1 6076
0 6078 7 1 2 6053 6077
0 6079 5 1 1 6078
0 6080 7 1 2 25575 6079
0 6081 5 1 1 6080
0 6082 7 2 2 27377 32327
0 6083 7 1 2 32025 32859
0 6084 5 1 1 6083
0 6085 7 1 2 4493 6075
0 6086 5 1 1 6085
0 6087 7 1 2 27590 6086
0 6088 7 1 2 32437 6087
0 6089 5 1 1 6088
0 6090 7 1 2 6084 6089
0 6091 5 1 1 6090
0 6092 7 1 2 29449 6091
0 6093 5 1 1 6092
0 6094 7 1 2 29740 32016
0 6095 7 1 2 31871 6094
0 6096 7 1 2 32328 6095
0 6097 5 1 1 6096
0 6098 7 1 2 6093 6097
0 6099 5 1 1 6098
0 6100 7 1 2 25913 29593
0 6101 7 1 2 6099 6100
0 6102 5 1 1 6101
0 6103 7 1 2 32851 6028
0 6104 5 1 1 6103
0 6105 7 1 2 27503 6104
0 6106 5 1 1 6105
0 6107 7 1 2 30572 32847
0 6108 5 1 1 6107
0 6109 7 1 2 27570 29239
0 6110 7 1 2 32354 6109
0 6111 5 1 1 6110
0 6112 7 1 2 6108 6111
0 6113 7 1 2 6106 6112
0 6114 5 1 1 6113
0 6115 7 1 2 23947 6114
0 6116 5 1 1 6115
0 6117 7 2 2 23004 31582
0 6118 5 1 1 32861
0 6119 7 1 2 32848 32862
0 6120 5 1 1 6119
0 6121 7 1 2 27504 32838
0 6122 5 1 1 6121
0 6123 7 1 2 6120 6122
0 6124 7 1 2 6116 6123
0 6125 5 1 1 6124
0 6126 7 1 2 28927 31964
0 6127 7 1 2 6125 6126
0 6128 5 1 1 6127
0 6129 7 1 2 6102 6128
0 6130 7 1 2 6081 6129
0 6131 5 1 1 6130
0 6132 7 1 2 24054 6131
0 6133 5 1 1 6132
0 6134 7 3 2 22911 27922
0 6135 7 2 2 29663 29836
0 6136 5 1 1 32866
0 6137 7 1 2 32863 32867
0 6138 7 1 2 32007 6137
0 6139 7 1 2 32828 6138
0 6140 5 1 1 6139
0 6141 7 1 2 23517 6140
0 6142 7 1 2 6133 6141
0 6143 5 1 1 6142
0 6144 7 1 2 23948 29827
0 6145 5 1 1 6144
0 6146 7 1 2 29815 6145
0 6147 5 5 1 6146
0 6148 7 2 2 31318 32868
0 6149 7 1 2 26063 27839
0 6150 5 1 1 6149
0 6151 7 1 2 4775 6150
0 6152 5 1 1 6151
0 6153 7 1 2 32873 6152
0 6154 5 1 1 6153
0 6155 7 1 2 31027 32701
0 6156 5 1 1 6155
0 6157 7 1 2 22019 32269
0 6158 5 2 1 6157
0 6159 7 2 2 21807 32875
0 6160 5 1 1 32877
0 6161 7 1 2 24055 28473
0 6162 5 2 1 6161
0 6163 7 1 2 32878 32879
0 6164 5 1 1 6163
0 6165 7 1 2 6156 6164
0 6166 5 2 1 6165
0 6167 7 2 2 22529 23282
0 6168 7 1 2 25786 32883
0 6169 7 1 2 25778 6168
0 6170 7 1 2 32881 6169
0 6171 5 1 1 6170
0 6172 7 1 2 6154 6171
0 6173 5 1 1 6172
0 6174 7 1 2 28141 6173
0 6175 5 1 1 6174
0 6176 7 3 2 25388 23735
0 6177 7 1 2 31301 32885
0 6178 7 1 2 32035 6177
0 6179 7 1 2 32869 6178
0 6180 5 1 1 6179
0 6181 7 1 2 6175 6180
0 6182 5 1 1 6181
0 6183 7 1 2 26263 6182
0 6184 5 1 1 6183
0 6185 7 2 2 23736 32870
0 6186 7 1 2 25914 32056
0 6187 5 1 1 6186
0 6188 7 1 2 27072 32161
0 6189 5 1 1 6188
0 6190 7 1 2 6187 6189
0 6191 5 1 1 6190
0 6192 7 1 2 24056 26693
0 6193 7 1 2 6191 6192
0 6194 7 1 2 32888 6193
0 6195 5 1 1 6194
0 6196 7 1 2 6184 6195
0 6197 5 1 1 6196
0 6198 7 1 2 25576 6197
0 6199 5 1 1 6198
0 6200 7 1 2 30007 32057
0 6201 7 1 2 32849 6200
0 6202 5 1 1 6201
0 6203 7 2 2 23428 31818
0 6204 7 1 2 25749 32890
0 6205 7 1 2 32438 6204
0 6206 5 1 1 6205
0 6207 7 1 2 26108 29741
0 6208 7 1 2 32339 6207
0 6209 7 1 2 32040 6208
0 6210 5 1 1 6209
0 6211 7 1 2 6206 6210
0 6212 5 1 1 6211
0 6213 7 1 2 25665 29450
0 6214 7 1 2 6212 6213
0 6215 5 1 1 6214
0 6216 7 1 2 6202 6215
0 6217 5 1 1 6216
0 6218 7 1 2 23636 31182
0 6219 7 1 2 6217 6218
0 6220 5 1 1 6219
0 6221 7 1 2 25464 6220
0 6222 7 1 2 6199 6221
0 6223 5 1 1 6222
0 6224 7 1 2 23091 6223
0 6225 7 1 2 6143 6224
0 6226 5 1 1 6225
0 6227 7 1 2 6021 6226
0 6228 5 1 1 6227
0 6229 7 1 2 25323 6228
0 6230 5 1 1 6229
0 6231 7 1 2 31343 31283
0 6232 7 2 2 31732 6231
0 6233 5 1 1 32892
0 6234 7 3 2 24684 23283
0 6235 7 1 2 25465 32284
0 6236 7 2 2 32894 6235
0 6237 7 1 2 32265 32897
0 6238 5 1 1 6237
0 6239 7 1 2 6233 6238
0 6240 5 1 1 6239
0 6241 7 1 2 21808 6240
0 6242 5 1 1 6241
0 6243 7 1 2 22467 32893
0 6244 5 1 1 6243
0 6245 7 4 2 23949 31031
0 6246 5 1 1 32899
0 6247 7 1 2 32900 32898
0 6248 5 1 1 6247
0 6249 7 1 2 6244 6248
0 6250 7 1 2 6242 6249
0 6251 5 1 1 6250
0 6252 7 1 2 25324 6251
0 6253 5 1 1 6252
0 6254 7 3 2 24057 22745
0 6255 7 1 2 26840 32903
0 6256 7 1 2 28216 6255
0 6257 5 1 1 6256
0 6258 7 1 2 6253 6257
0 6259 5 1 1 6258
0 6260 7 1 2 24197 6259
0 6261 5 1 1 6260
0 6262 7 12 2 24685 23360
0 6263 5 1 1 32906
0 6264 7 2 2 28291 32907
0 6265 5 1 1 32918
0 6266 7 1 2 26788 31164
0 6267 5 1 1 6266
0 6268 7 1 2 6265 6267
0 6269 5 10 1 6268
0 6270 7 6 2 23284 31288
0 6271 7 2 2 28217 32930
0 6272 5 1 1 32936
0 6273 7 1 2 32920 32937
0 6274 5 1 1 6273
0 6275 7 1 2 6261 6274
0 6276 5 1 1 6275
0 6277 7 1 2 26630 6276
0 6278 5 1 1 6277
0 6279 7 2 2 22912 31289
0 6280 7 3 2 31856 32498
0 6281 7 3 2 32921 32940
0 6282 7 1 2 32938 32943
0 6283 5 1 1 6282
0 6284 7 1 2 6278 6283
0 6285 5 1 1 6284
0 6286 7 1 2 24378 6285
0 6287 5 1 1 6286
0 6288 7 2 2 25881 31290
0 6289 7 1 2 32944 32946
0 6290 5 1 1 6289
0 6291 7 1 2 6287 6290
0 6292 5 1 1 6291
0 6293 7 1 2 26064 6292
0 6294 5 1 1 6293
0 6295 7 12 2 24686 25325
0 6296 5 1 1 32948
0 6297 7 1 2 31255 6296
0 6298 5 37 1 6297
0 6299 7 3 2 22020 25577
0 6300 7 2 2 29344 32997
0 6301 7 2 2 27573 31713
0 6302 7 1 2 30405 33002
0 6303 7 1 2 33000 6302
0 6304 5 1 1 6303
0 6305 7 9 2 24198 23285
0 6306 7 2 2 33004 32285
0 6307 7 1 2 25466 33013
0 6308 7 1 2 32499 6307
0 6309 7 1 2 32616 6308
0 6310 5 1 1 6309
0 6311 7 1 2 6304 6310
0 6312 5 1 1 6311
0 6313 7 1 2 26065 6312
0 6314 5 1 1 6313
0 6315 7 2 2 23637 32500
0 6316 7 4 2 24849 25467
0 6317 7 2 2 27981 33017
0 6318 7 1 2 33014 33021
0 6319 7 1 2 33015 6318
0 6320 5 1 1 6319
0 6321 7 1 2 6314 6320
0 6322 5 1 1 6321
0 6323 7 1 2 32960 6322
0 6324 5 1 1 6323
0 6325 7 1 2 27688 31291
0 6326 7 1 2 32945 6325
0 6327 5 1 1 6326
0 6328 7 1 2 6324 6327
0 6329 7 1 2 6294 6328
0 6330 5 1 1 6329
0 6331 7 1 2 32578 6330
0 6332 5 1 1 6331
0 6333 7 11 2 22191 23286
0 6334 7 9 2 23638 31819
0 6335 7 1 2 24471 29905
0 6336 7 3 2 31481 6335
0 6337 5 1 1 33043
0 6338 7 1 2 33034 33044
0 6339 5 1 1 6338
0 6340 7 3 2 24058 28736
0 6341 5 1 1 33046
0 6342 7 2 2 33035 33047
0 6343 5 1 1 33049
0 6344 7 1 2 22021 29006
0 6345 5 5 1 6344
0 6346 7 1 2 23005 31446
0 6347 7 2 2 33051 6346
0 6348 7 1 2 26066 32697
0 6349 5 1 1 6348
0 6350 7 1 2 653 6349
0 6351 5 2 1 6350
0 6352 7 1 2 33056 33058
0 6353 5 1 1 6352
0 6354 7 1 2 6343 6353
0 6355 5 1 1 6354
0 6356 7 1 2 23950 6355
0 6357 5 1 1 6356
0 6358 7 1 2 6339 6357
0 6359 5 1 1 6358
0 6360 7 1 2 23820 6359
0 6361 5 1 1 6360
0 6362 7 1 2 30888 33050
0 6363 5 1 1 6362
0 6364 7 1 2 6361 6363
0 6365 5 1 1 6364
0 6366 7 1 2 33023 6365
0 6367 5 1 1 6366
0 6368 7 2 2 25787 29695
0 6369 7 1 2 28741 28904
0 6370 7 1 2 33060 6369
0 6371 5 1 1 6370
0 6372 7 1 2 28230 29007
0 6373 5 2 1 6372
0 6374 7 1 2 29980 33062
0 6375 5 5 1 6374
0 6376 7 1 2 33036 33064
0 6377 5 1 1 6376
0 6378 7 1 2 6371 6377
0 6379 5 1 1 6378
0 6380 7 1 2 31811 6379
0 6381 5 1 1 6380
0 6382 7 1 2 6367 6381
0 6383 5 1 1 6382
0 6384 7 1 2 32922 6383
0 6385 5 1 1 6384
0 6386 7 2 2 25468 26829
0 6387 7 3 2 32961 33037
0 6388 5 1 1 33071
0 6389 7 1 2 28417 33048
0 6390 7 1 2 33072 6389
0 6391 5 1 1 6390
0 6392 7 2 2 24472 31242
0 6393 5 1 1 33074
0 6394 7 3 2 26109 27898
0 6395 7 1 2 33075 33076
0 6396 5 1 1 6395
0 6397 7 1 2 6388 6396
0 6398 5 1 1 6397
0 6399 7 2 2 23821 33057
0 6400 7 1 2 6398 33079
0 6401 5 1 1 6400
0 6402 7 1 2 6391 6401
0 6403 5 1 1 6402
0 6404 7 1 2 23951 6403
0 6405 5 1 1 6404
0 6406 7 1 2 23822 33045
0 6407 7 1 2 33073 6406
0 6408 5 1 1 6407
0 6409 7 1 2 6405 6408
0 6410 5 1 1 6409
0 6411 7 1 2 33069 6410
0 6412 5 1 1 6411
0 6413 7 1 2 31724 31947
0 6414 7 1 2 32596 6413
0 6415 7 2 2 25054 26922
0 6416 7 2 2 25234 29428
0 6417 7 1 2 26615 29721
0 6418 7 1 2 33083 6417
0 6419 7 1 2 33081 6418
0 6420 7 1 2 6414 6419
0 6421 5 1 1 6420
0 6422 7 1 2 6412 6421
0 6423 5 1 1 6422
0 6424 7 1 2 24199 6423
0 6425 5 1 1 6424
0 6426 7 1 2 26406 2072
0 6427 5 1 1 6426
0 6428 7 1 2 25578 30941
0 6429 5 1 1 6428
0 6430 7 1 2 22530 26468
0 6431 7 1 2 6429 6430
0 6432 5 1 1 6431
0 6433 7 2 2 22913 28756
0 6434 5 1 1 33085
0 6435 7 3 2 26631 29388
0 6436 5 1 1 33087
0 6437 7 4 2 24941 23639
0 6438 7 1 2 22914 33090
0 6439 5 1 1 6438
0 6440 7 1 2 6436 6439
0 6441 5 1 1 6440
0 6442 7 1 2 22468 6441
0 6443 5 1 1 6442
0 6444 7 1 2 6434 6443
0 6445 7 1 2 6432 6444
0 6446 5 1 1 6445
0 6447 7 1 2 21809 6446
0 6448 5 1 1 6447
0 6449 7 1 2 6427 6448
0 6450 5 1 1 6449
0 6451 7 1 2 24379 6450
0 6452 5 1 1 6451
0 6453 7 1 2 30035 30050
0 6454 5 2 1 6453
0 6455 7 2 2 26465 33094
0 6456 7 1 2 22384 33096
0 6457 5 1 1 6456
0 6458 7 1 2 6452 6457
0 6459 5 2 1 6458
0 6460 7 1 2 26067 33098
0 6461 5 1 1 6460
0 6462 7 2 2 27982 33097
0 6463 5 1 1 33100
0 6464 7 1 2 6461 6463
0 6465 5 1 1 6464
0 6466 7 1 2 21908 6465
0 6467 5 1 1 6466
0 6468 7 2 2 29406 31054
0 6469 7 1 2 31820 33102
0 6470 5 1 1 6469
0 6471 7 1 2 6467 6470
0 6472 5 1 1 6471
0 6473 7 5 2 22022 22192
0 6474 7 2 2 32962 33104
0 6475 7 1 2 30406 33109
0 6476 7 1 2 6472 6475
0 6477 5 1 1 6476
0 6478 7 1 2 6425 6477
0 6479 7 1 2 6385 6478
0 6480 7 1 2 6332 6479
0 6481 5 1 1 6480
0 6482 7 1 2 25666 6481
0 6483 5 1 1 6482
0 6484 7 2 2 26491 29240
0 6485 7 1 2 32560 33111
0 6486 5 1 1 6485
0 6487 7 1 2 6023 6486
0 6488 5 1 1 6487
0 6489 7 1 2 23092 6488
0 6490 5 1 1 6489
0 6491 7 1 2 27773 29837
0 6492 5 1 1 6491
0 6493 7 1 2 6490 6492
0 6494 5 1 1 6493
0 6495 7 1 2 23952 6494
0 6496 5 1 1 6495
0 6497 7 1 2 24473 29187
0 6498 5 1 1 6497
0 6499 7 1 2 6496 6498
0 6500 5 1 1 6499
0 6501 7 1 2 23823 6500
0 6502 5 1 1 6501
0 6503 7 1 2 29170 32266
0 6504 5 1 1 6503
0 6505 7 1 2 23824 27731
0 6506 7 1 2 32579 6505
0 6507 5 1 1 6506
0 6508 7 1 2 27794 6507
0 6509 5 1 1 6508
0 6510 7 1 2 28198 6509
0 6511 5 1 1 6510
0 6512 7 1 2 27302 32580
0 6513 5 1 1 6512
0 6514 7 1 2 22531 29742
0 6515 5 1 1 6514
0 6516 7 1 2 6513 6515
0 6517 5 1 1 6516
0 6518 7 1 2 24380 29152
0 6519 7 1 2 6517 6518
0 6520 5 1 1 6519
0 6521 7 1 2 23093 27840
0 6522 5 1 1 6521
0 6523 7 1 2 22532 29790
0 6524 5 1 1 6523
0 6525 7 1 2 27774 6524
0 6526 5 1 1 6525
0 6527 7 1 2 6522 6526
0 6528 7 1 2 6520 6527
0 6529 7 1 2 6511 6528
0 6530 5 1 1 6529
0 6531 7 1 2 24059 6530
0 6532 5 1 1 6531
0 6533 7 1 2 6504 6532
0 6534 7 1 2 6502 6533
0 6535 5 2 1 6534
0 6536 7 1 2 33005 32475
0 6537 7 1 2 33113 6536
0 6538 5 1 1 6537
0 6539 7 1 2 22469 29083
0 6540 5 1 1 6539
0 6541 7 1 2 31275 6540
0 6542 5 1 1 6541
0 6543 7 1 2 21909 6542
0 6544 5 1 1 6543
0 6545 7 2 2 24942 29008
0 6546 5 2 1 33115
0 6547 7 1 2 1934 33117
0 6548 5 1 1 6547
0 6549 7 1 2 22023 6548
0 6550 5 1 1 6549
0 6551 7 1 2 6544 6550
0 6552 5 1 1 6551
0 6553 7 1 2 21810 6552
0 6554 5 1 1 6553
0 6555 7 1 2 28474 28977
0 6556 5 1 1 6555
0 6557 7 1 2 22024 28205
0 6558 7 1 2 6556 6557
0 6559 5 1 1 6558
0 6560 7 1 2 6554 6559
0 6561 5 2 1 6560
0 6562 7 1 2 30243 32775
0 6563 7 1 2 32125 6562
0 6564 7 1 2 33119 6563
0 6565 5 1 1 6564
0 6566 7 1 2 6538 6565
0 6567 5 1 1 6566
0 6568 7 1 2 25579 6567
0 6569 5 1 1 6568
0 6570 7 5 2 22025 27775
0 6571 5 1 1 33121
0 6572 7 2 2 22026 29304
0 6573 7 1 2 27579 33126
0 6574 5 1 1 6573
0 6575 7 1 2 32566 6574
0 6576 5 1 1 6575
0 6577 7 1 2 21910 6576
0 6578 5 1 1 6577
0 6579 7 1 2 6571 6578
0 6580 5 1 1 6579
0 6581 7 1 2 27174 6580
0 6582 5 1 1 6581
0 6583 7 1 2 24060 27505
0 6584 5 3 1 6583
0 6585 7 1 2 29840 33128
0 6586 5 1 1 6585
0 6587 7 1 2 23953 6586
0 6588 5 1 1 6587
0 6589 7 1 2 27841 5569
0 6590 7 1 2 6588 6589
0 6591 5 1 1 6590
0 6592 7 1 2 6582 6591
0 6593 5 1 1 6592
0 6594 7 1 2 25055 6593
0 6595 5 1 1 6594
0 6596 7 1 2 30790 32003
0 6597 5 1 1 6596
0 6598 7 1 2 29345 29706
0 6599 5 2 1 6598
0 6600 7 3 2 29959 31652
0 6601 5 1 1 33133
0 6602 7 1 2 33131 6601
0 6603 5 1 1 6602
0 6604 7 1 2 32602 6603
0 6605 5 1 1 6604
0 6606 7 1 2 6597 6605
0 6607 7 1 2 6595 6606
0 6608 5 2 1 6607
0 6609 7 1 2 30820 32776
0 6610 7 1 2 33136 6609
0 6611 5 1 1 6610
0 6612 7 1 2 6569 6611
0 6613 5 1 1 6612
0 6614 7 1 2 32963 6613
0 6615 5 1 1 6614
0 6616 7 1 2 30258 31284
0 6617 7 1 2 33120 6616
0 6618 5 1 1 6617
0 6619 7 1 2 25056 2030
0 6620 5 1 1 6619
0 6621 7 1 2 22533 32501
0 6622 5 1 1 6621
0 6623 7 1 2 28612 32572
0 6624 7 1 2 6622 6623
0 6625 5 1 1 6624
0 6626 7 1 2 24061 6625
0 6627 7 1 2 6620 6626
0 6628 5 1 1 6627
0 6629 7 2 2 22027 28978
0 6630 5 4 1 33138
0 6631 7 1 2 33139 32625
0 6632 5 1 1 6631
0 6633 7 1 2 6628 6632
0 6634 5 1 1 6633
0 6635 7 1 2 30292 32895
0 6636 7 1 2 6634 6635
0 6637 5 1 1 6636
0 6638 7 1 2 6618 6637
0 6639 5 1 1 6638
0 6640 7 1 2 25326 6639
0 6641 5 1 1 6640
0 6642 7 3 2 22028 24687
0 6643 7 1 2 25801 33144
0 6644 7 1 2 30293 6643
0 6645 7 1 2 33065 6644
0 6646 5 1 1 6645
0 6647 7 1 2 6641 6646
0 6648 5 1 1 6647
0 6649 7 1 2 24200 6648
0 6650 5 1 1 6649
0 6651 7 1 2 24062 28218
0 6652 5 1 1 6651
0 6653 7 1 2 21811 32880
0 6654 5 1 1 6653
0 6655 7 5 2 32876 6654
0 6656 5 6 1 33147
0 6657 7 1 2 29112 33148
0 6658 5 1 1 6657
0 6659 7 2 2 6652 6658
0 6660 5 1 1 33158
0 6661 7 1 2 31165 33024
0 6662 7 1 2 30259 6661
0 6663 7 1 2 6660 6662
0 6664 5 1 1 6663
0 6665 7 1 2 6650 6664
0 6666 5 1 1 6665
0 6667 7 1 2 25915 6666
0 6668 5 1 1 6667
0 6669 7 1 2 31166 30862
0 6670 5 1 1 6669
0 6671 7 5 2 23429 32908
0 6672 7 1 2 28670 33160
0 6673 5 1 1 6672
0 6674 7 1 2 6670 6673
0 6675 5 5 1 6674
0 6676 7 9 2 24201 25235
0 6677 7 1 2 33170 33137
0 6678 5 1 1 6677
0 6679 7 1 2 33025 33114
0 6680 5 1 1 6679
0 6681 7 1 2 6678 6680
0 6682 5 1 1 6681
0 6683 7 1 2 33165 6682
0 6684 5 1 1 6683
0 6685 7 1 2 6668 6684
0 6686 7 1 2 6615 6685
0 6687 5 1 1 6686
0 6688 7 1 2 28793 6687
0 6689 5 1 1 6688
0 6690 7 3 2 22193 31243
0 6691 5 3 1 33179
0 6692 7 2 2 28529 31222
0 6693 5 1 1 33185
0 6694 7 1 2 33182 6693
0 6695 5 1 1 6694
0 6696 7 1 2 26789 6695
0 6697 5 1 1 6696
0 6698 7 2 2 28142 26833
0 6699 5 1 1 33187
0 6700 7 1 2 29755 33188
0 6701 5 1 1 6700
0 6702 7 1 2 6697 6701
0 6703 5 1 1 6702
0 6704 7 1 2 31188 6703
0 6705 5 1 1 6704
0 6706 7 2 2 22470 32949
0 6707 5 1 1 33189
0 6708 7 1 2 31256 6707
0 6709 5 2 1 6708
0 6710 7 1 2 22194 33191
0 6711 5 1 1 6710
0 6712 7 2 2 24202 31167
0 6713 5 1 1 33193
0 6714 7 1 2 22471 33194
0 6715 5 1 1 6714
0 6716 7 1 2 6711 6715
0 6717 5 1 1 6716
0 6718 7 1 2 26790 6717
0 6719 5 1 1 6718
0 6720 7 1 2 29884 31162
0 6721 5 1 1 6720
0 6722 7 1 2 6719 6721
0 6723 5 1 1 6722
0 6724 7 1 2 21812 6723
0 6725 5 1 1 6724
0 6726 7 1 2 23518 26571
0 6727 7 1 2 31727 6726
0 6728 5 1 1 6727
0 6729 7 1 2 6725 6728
0 6730 5 1 1 6729
0 6731 7 1 2 24943 6730
0 6732 5 1 1 6731
0 6733 7 1 2 24203 33145
0 6734 7 1 2 29885 6733
0 6735 5 1 1 6734
0 6736 7 1 2 6732 6735
0 6737 5 1 1 6736
0 6738 7 1 2 29494 6737
0 6739 5 1 1 6738
0 6740 7 1 2 6705 6739
0 6741 5 1 1 6740
0 6742 7 1 2 28107 6741
0 6743 5 1 1 6742
0 6744 7 1 2 22029 30843
0 6745 5 2 1 6744
0 6746 7 1 2 29657 33195
0 6747 5 1 1 6746
0 6748 7 3 2 22195 32950
0 6749 5 1 1 33197
0 6750 7 1 2 6749 33183
0 6751 7 1 2 6713 6750
0 6752 5 7 1 6751
0 6753 7 1 2 26791 33200
0 6754 5 1 1 6753
0 6755 7 1 2 6754 6699
0 6756 5 2 1 6755
0 6757 7 1 2 28118 33207
0 6758 7 1 2 6747 6757
0 6759 5 1 1 6758
0 6760 7 1 2 6743 6759
0 6761 5 1 1 6760
0 6762 7 1 2 25057 6761
0 6763 5 1 1 6762
0 6764 7 1 2 31664 31771
0 6765 7 1 2 33208 6764
0 6766 5 1 1 6765
0 6767 7 1 2 25236 6766
0 6768 7 1 2 6763 6767
0 6769 5 1 1 6768
0 6770 7 1 2 29122 32226
0 6771 5 1 1 6770
0 6772 7 1 2 27378 31438
0 6773 5 1 1 6772
0 6774 7 1 2 6771 6773
0 6775 5 3 1 6774
0 6776 7 2 2 22196 32923
0 6777 5 1 1 33212
0 6778 7 5 2 24204 32964
0 6779 5 1 1 33214
0 6780 7 2 2 28292 33215
0 6781 5 1 1 33219
0 6782 7 1 2 6777 6781
0 6783 5 3 1 6782
0 6784 7 1 2 25580 33221
0 6785 7 2 2 33209 6784
0 6786 7 1 2 25916 33224
0 6787 5 1 1 6786
0 6788 7 8 2 22746 23094
0 6789 5 1 1 33226
0 6790 7 2 2 26842 33227
0 6791 5 1 1 33234
0 6792 7 4 2 24688 23006
0 6793 7 1 2 23825 33236
0 6794 7 1 2 29886 6793
0 6795 5 1 1 6794
0 6796 7 1 2 6791 6795
0 6797 5 1 1 6796
0 6798 7 1 2 22197 6797
0 6799 5 1 1 6798
0 6800 7 1 2 29779 33220
0 6801 5 1 1 6800
0 6802 7 1 2 6799 6801
0 6803 5 1 1 6802
0 6804 7 1 2 31458 6803
0 6805 5 1 1 6804
0 6806 7 2 2 22198 32909
0 6807 5 1 1 33240
0 6808 7 1 2 6779 6807
0 6809 5 8 1 6808
0 6810 7 1 2 31447 6136
0 6811 5 1 1 6810
0 6812 7 1 2 33242 6811
0 6813 5 1 1 6812
0 6814 7 7 2 23954 24205
0 6815 7 2 2 25327 33250
0 6816 7 1 2 29764 33237
0 6817 7 1 2 33257 6816
0 6818 5 1 1 6817
0 6819 7 1 2 6813 6818
0 6820 5 1 1 6819
0 6821 7 1 2 28293 6820
0 6822 5 1 1 6821
0 6823 7 1 2 6805 6822
0 6824 5 1 1 6823
0 6825 7 1 2 26424 6824
0 6826 5 1 1 6825
0 6827 7 1 2 6787 6826
0 6828 5 1 1 6827
0 6829 7 1 2 25848 6828
0 6830 5 1 1 6829
0 6831 7 1 2 25971 33225
0 6832 5 1 1 6831
0 6833 7 1 2 23287 6832
0 6834 7 1 2 6830 6833
0 6835 7 1 2 22534 28193
0 6836 5 5 1 6835
0 6837 7 3 2 23826 28119
0 6838 5 1 1 33264
0 6839 7 1 2 33265 33222
0 6840 5 1 1 6839
0 6841 7 1 2 26202 28945
0 6842 7 1 2 33243 6841
0 6843 5 1 1 6842
0 6844 7 1 2 6840 6843
0 6845 5 1 1 6844
0 6846 7 1 2 24063 6845
0 6847 5 1 1 6846
0 6848 7 3 2 26792 27712
0 6849 7 1 2 28247 28958
0 6850 7 1 2 33228 6849
0 6851 7 2 2 33267 6850
0 6852 5 1 1 33270
0 6853 7 1 2 23827 33271
0 6854 5 1 1 6853
0 6855 7 1 2 6847 6854
0 6856 5 1 1 6855
0 6857 7 1 2 33259 6856
0 6858 5 1 1 6857
0 6859 7 4 2 24064 28120
0 6860 5 1 1 33272
0 6861 7 2 2 33273 33223
0 6862 5 1 1 33276
0 6863 7 1 2 6862 6852
0 6864 5 1 1 6863
0 6865 7 1 2 27303 6864
0 6866 5 1 1 6865
0 6867 7 5 2 23095 23430
0 6868 7 1 2 27137 28959
0 6869 7 1 2 33278 6868
0 6870 7 1 2 28279 28688
0 6871 7 1 2 6869 6870
0 6872 5 1 1 6871
0 6873 7 1 2 6866 6872
0 6874 5 1 1 6873
0 6875 7 1 2 29594 6874
0 6876 5 1 1 6875
0 6877 7 1 2 6858 6876
0 6878 7 1 2 6834 6877
0 6879 5 1 1 6878
0 6880 7 1 2 23737 6879
0 6881 7 1 2 6769 6880
0 6882 5 1 1 6881
0 6883 7 1 2 6689 6882
0 6884 7 1 2 6483 6883
0 6885 5 1 1 6884
0 6886 7 1 2 30144 6885
0 6887 5 1 1 6886
0 6888 7 1 2 6230 6887
0 6889 7 1 2 5888 6888
0 6890 7 1 2 4931 6889
0 6891 5 1 1 6890
0 6892 7 1 2 25698 6891
0 6893 5 1 1 6892
0 6894 7 53 2 22243 22787
0 6895 5 1 1 33283
0 6896 7 1 2 33284 32084
0 6897 5 1 1 6896
0 6898 7 55 2 24256 24731
0 6899 5 1 1 33336
0 6900 7 5 2 22915 28794
0 6901 7 2 2 33337 33391
0 6902 5 1 1 33396
0 6903 7 1 2 6897 6902
0 6904 5 1 1 6903
0 6905 7 1 2 22385 6904
0 6906 5 1 1 6905
0 6907 7 8 2 22244 22314
0 6908 7 12 2 22788 33398
0 6909 7 2 2 33406 31966
0 6910 5 2 1 33418
0 6911 7 1 2 6906 33420
0 6912 5 7 1 6911
0 6913 7 6 2 23519 23738
0 6914 7 2 2 33422 33429
0 6915 7 3 2 25328 28530
0 6916 5 1 1 33437
0 6917 7 1 2 29009 33438
0 6918 5 1 1 6917
0 6919 7 1 2 22535 33180
0 6920 5 1 1 6919
0 6921 7 1 2 6918 6920
0 6922 5 1 1 6921
0 6923 7 1 2 33435 6922
0 6924 5 1 1 6923
0 6925 7 1 2 23361 27039
0 6926 7 1 2 30206 30771
0 6927 7 1 2 6925 6926
0 6928 7 5 2 24732 24799
0 6929 7 4 2 25788 33440
0 6930 7 11 2 22199 24257
0 6931 7 2 2 31687 33449
0 6932 7 1 2 33445 33460
0 6933 7 1 2 6927 6932
0 6934 5 1 1 6933
0 6935 7 1 2 6924 6934
0 6936 5 1 1 6935
0 6937 7 1 2 22644 6936
0 6938 5 1 1 6937
0 6939 7 5 2 27776 29213
0 6940 5 2 1 33462
0 6941 7 3 2 25469 27574
0 6942 7 1 2 33469 32581
0 6943 7 1 2 32072 6942
0 6944 5 1 1 6943
0 6945 7 1 2 33467 6944
0 6946 5 1 1 6945
0 6947 7 1 2 22645 6946
0 6948 5 1 1 6947
0 6949 7 1 2 27777 29084
0 6950 7 1 2 32182 6949
0 6951 5 1 1 6950
0 6952 7 1 2 6948 6951
0 6953 5 1 1 6952
0 6954 7 1 2 24322 6953
0 6955 5 1 1 6954
0 6956 7 8 2 22916 23520
0 6957 7 2 2 24800 33472
0 6958 5 2 1 33480
0 6959 7 1 2 22857 33470
0 6960 5 1 1 6959
0 6961 7 1 2 33482 6960
0 6962 5 1 1 6961
0 6963 7 1 2 22386 6962
0 6964 5 1 1 6963
0 6965 7 1 2 32173 31967
0 6966 5 1 1 6965
0 6967 7 1 2 6964 6966
0 6968 5 1 1 6967
0 6969 7 1 2 29085 6968
0 6970 5 1 1 6969
0 6971 7 1 2 28436 33481
0 6972 5 1 1 6971
0 6973 7 1 2 6970 6972
0 6974 5 1 1 6973
0 6975 7 1 2 28497 6974
0 6976 5 1 1 6975
0 6977 7 1 2 6955 6976
0 6978 5 1 1 6977
0 6979 7 1 2 33338 6978
0 6980 5 1 1 6979
0 6981 7 4 2 23739 33285
0 6982 7 1 2 29086 30690
0 6983 5 1 1 6982
0 6984 7 1 2 5496 6983
0 6985 5 1 1 6984
0 6986 7 1 2 25917 6985
0 6987 5 1 1 6986
0 6988 7 1 2 24600 29113
0 6989 5 4 1 6988
0 6990 7 2 2 23521 33488
0 6991 7 1 2 25972 33492
0 6992 5 1 1 6991
0 6993 7 1 2 6987 6992
0 6994 5 1 1 6993
0 6995 7 1 2 33484 6994
0 6996 5 1 1 6995
0 6997 7 1 2 6980 6996
0 6998 5 1 1 6997
0 6999 7 1 2 33181 6998
0 7000 5 1 1 6999
0 7001 7 3 2 25058 25470
0 7002 7 2 2 30566 33494
0 7003 7 7 2 24258 22315
0 7004 7 6 2 24733 22858
0 7005 7 5 2 33499 33506
0 7006 5 1 1 33512
0 7007 7 3 2 28795 33286
0 7008 5 1 1 33517
0 7009 7 1 2 7006 7008
0 7010 5 17 1 7009
0 7011 7 2 2 25918 33520
0 7012 5 2 1 33537
0 7013 7 2 2 25973 33339
0 7014 5 2 1 33541
0 7015 7 1 2 33539 33543
0 7016 5 4 1 7015
0 7017 7 1 2 33497 33545
0 7018 5 1 1 7017
0 7019 7 1 2 33423 33493
0 7020 5 1 1 7019
0 7021 7 1 2 7018 7020
0 7022 5 1 1 7021
0 7023 7 1 2 23740 33439
0 7024 7 1 2 7022 7023
0 7025 5 1 1 7024
0 7026 7 1 2 7000 7025
0 7027 5 1 1 7026
0 7028 7 1 2 21911 7027
0 7029 5 1 1 7028
0 7030 7 1 2 6938 7029
0 7031 5 1 1 7030
0 7032 7 1 2 23204 7031
0 7033 5 1 1 7032
0 7034 7 1 2 27058 33186
0 7035 5 1 1 7034
0 7036 7 1 2 33184 6916
0 7037 5 1 1 7036
0 7038 7 1 2 23096 29495
0 7039 7 1 2 7037 7038
0 7040 5 1 1 7039
0 7041 7 1 2 7035 7040
0 7042 5 1 1 7041
0 7043 7 1 2 23741 28561
0 7044 7 1 2 7042 7043
0 7045 7 1 2 33424 7044
0 7046 5 1 1 7045
0 7047 7 1 2 7033 7046
0 7048 5 1 1 7047
0 7049 7 1 2 25581 7048
0 7050 5 1 1 7049
0 7051 7 1 2 30521 31141
0 7052 5 1 1 7051
0 7053 7 1 2 24944 32466
0 7054 5 1 1 7053
0 7055 7 1 2 7052 7054
0 7056 5 1 1 7055
0 7057 7 1 2 23205 7056
0 7058 5 1 1 7057
0 7059 7 1 2 22859 23097
0 7060 7 3 2 29362 7059
0 7061 7 1 2 30122 33549
0 7062 5 1 1 7061
0 7063 7 1 2 7058 7062
0 7064 5 1 1 7063
0 7065 7 1 2 33287 7064
0 7066 5 1 1 7065
0 7067 7 3 2 22316 24734
0 7068 7 3 2 24259 33552
0 7069 7 2 2 29564 33555
0 7070 7 1 2 30809 32187
0 7071 7 1 2 33558 7070
0 7072 5 1 1 7071
0 7073 7 14 2 25471 33521
0 7074 7 2 2 30609 33560
0 7075 5 1 1 33574
0 7076 7 2 2 27233 32194
0 7077 5 1 1 33576
0 7078 7 1 2 33407 33577
0 7079 5 1 1 7078
0 7080 7 1 2 7075 7079
0 7081 5 2 1 7080
0 7082 7 1 2 29496 33578
0 7083 5 1 1 7082
0 7084 7 1 2 7072 7083
0 7085 7 1 2 7066 7084
0 7086 5 1 1 7085
0 7087 7 1 2 33201 32065
0 7088 7 1 2 7086 7087
0 7089 5 1 1 7088
0 7090 7 1 2 7050 7089
0 7091 5 1 1 7090
0 7092 7 1 2 25237 7091
0 7093 5 1 1 7092
0 7094 7 5 2 24260 22387
0 7095 7 3 2 24735 33473
0 7096 7 2 2 33580 33585
0 7097 5 1 1 33588
0 7098 7 5 2 25582 33589
0 7099 5 1 1 33590
0 7100 7 9 2 25472 33288
0 7101 7 1 2 26219 26482
0 7102 5 1 1 7101
0 7103 7 1 2 33595 7102
0 7104 7 1 2 26363 7103
0 7105 5 1 1 7104
0 7106 7 1 2 7099 7105
0 7107 5 1 1 7106
0 7108 7 1 2 28796 7107
0 7109 5 1 1 7108
0 7110 7 3 2 24736 33581
0 7111 7 2 2 22917 28658
0 7112 5 1 1 33607
0 7113 7 3 2 33604 33608
0 7114 5 2 1 33609
0 7115 7 5 2 22789 23522
0 7116 7 12 2 22245 33614
0 7117 5 3 1 33619
0 7118 7 2 2 33340 32174
0 7119 5 1 1 33634
0 7120 7 1 2 33631 7119
0 7121 5 5 1 7120
0 7122 7 1 2 28121 33636
0 7123 5 1 1 7122
0 7124 7 1 2 33612 7123
0 7125 7 1 2 7109 7124
0 7126 5 1 1 7125
0 7127 7 1 2 29565 7126
0 7128 5 1 1 7127
0 7129 7 2 2 28949 33289
0 7130 7 3 2 29260 33641
0 7131 7 1 2 28727 29497
0 7132 7 1 2 33643 7131
0 7133 5 1 1 7132
0 7134 7 1 2 7128 7133
0 7135 5 1 1 7134
0 7136 7 2 2 23742 27018
0 7137 7 1 2 26694 33646
0 7138 7 1 2 33202 7137
0 7139 7 1 2 7135 7138
0 7140 5 1 1 7139
0 7141 7 1 2 7093 7140
0 7142 5 1 1 7141
0 7143 7 1 2 23431 7142
0 7144 5 1 1 7143
0 7145 7 1 2 25238 33579
0 7146 5 1 1 7145
0 7147 7 6 2 22790 22860
0 7148 7 10 2 33399 33648
0 7149 7 1 2 28880 30711
0 7150 7 1 2 33654 7149
0 7151 5 1 1 7150
0 7152 7 1 2 7146 7151
0 7153 5 1 1 7152
0 7154 7 1 2 29498 7153
0 7155 5 1 1 7154
0 7156 7 1 2 33561 32373
0 7157 5 1 1 7156
0 7158 7 3 2 23523 30610
0 7159 7 1 2 30755 33655
0 7160 7 1 2 33664 7159
0 7161 5 1 1 7160
0 7162 7 1 2 7157 7161
0 7163 7 1 2 7155 7162
0 7164 5 1 1 7163
0 7165 7 1 2 23640 7164
0 7166 5 1 1 7165
0 7167 7 1 2 33341 32447
0 7168 5 1 1 7167
0 7169 7 3 2 24323 33290
0 7170 5 1 1 33667
0 7171 7 3 2 33668 31912
0 7172 5 2 1 33670
0 7173 7 1 2 7168 33673
0 7174 5 5 1 7173
0 7175 7 2 2 33675 32368
0 7176 7 1 2 26473 30436
0 7177 7 1 2 33680 7176
0 7178 5 1 1 7177
0 7179 7 1 2 26203 7178
0 7180 7 1 2 7166 7179
0 7181 5 1 1 7180
0 7182 7 1 2 30736 33291
0 7183 5 1 1 7182
0 7184 7 4 2 24737 33500
0 7185 7 4 2 30663 33682
0 7186 5 1 1 33686
0 7187 7 1 2 7183 7186
0 7188 5 6 1 7187
0 7189 7 5 2 21912 30567
0 7190 5 1 1 33696
0 7191 7 1 2 30531 33697
0 7192 7 1 2 32369 7191
0 7193 7 1 2 33690 7192
0 7194 5 1 1 7193
0 7195 7 1 2 26220 7194
0 7196 5 1 1 7195
0 7197 7 4 2 23362 23743
0 7198 7 1 2 26129 33701
0 7199 7 1 2 28186 7198
0 7200 7 1 2 7196 7199
0 7201 7 1 2 7181 7200
0 7202 5 1 1 7201
0 7203 7 1 2 7144 7202
0 7204 5 1 1 7203
0 7205 7 1 2 22030 7204
0 7206 5 1 1 7205
0 7207 7 2 2 25849 29263
0 7208 5 1 1 33705
0 7209 7 1 2 27059 27899
0 7210 5 1 1 7209
0 7211 7 1 2 7208 7210
0 7212 5 1 1 7211
0 7213 7 1 2 33292 7212
0 7214 5 1 1 7213
0 7215 7 6 2 25583 33342
0 7216 7 3 2 28797 33707
0 7217 7 1 2 27060 33713
0 7218 5 1 1 7217
0 7219 7 1 2 7214 7218
0 7220 5 1 1 7219
0 7221 7 1 2 25164 7220
0 7222 5 1 1 7221
0 7223 7 5 2 22246 33649
0 7224 7 1 2 28013 30108
0 7225 7 1 2 33716 7224
0 7226 5 1 1 7225
0 7227 7 1 2 7222 7226
0 7228 5 1 1 7227
0 7229 7 1 2 24945 7228
0 7230 5 1 1 7229
0 7231 7 2 2 28798 33343
0 7232 5 1 1 33721
0 7233 7 8 2 26068 33293
0 7234 5 1 1 33723
0 7235 7 1 2 7232 7234
0 7236 5 13 1 7235
0 7237 7 7 2 25584 33731
0 7238 7 2 2 23206 27019
0 7239 7 1 2 33744 33751
0 7240 5 1 1 7239
0 7241 7 1 2 7230 7240
0 7242 5 1 1 7241
0 7243 7 1 2 22536 7242
0 7244 5 1 1 7243
0 7245 7 1 2 31112 33745
0 7246 5 1 1 7245
0 7247 7 1 2 7244 7246
0 7248 5 1 1 7247
0 7249 7 1 2 30972 7248
0 7250 5 1 1 7249
0 7251 7 2 2 26848 30806
0 7252 5 1 1 33753
0 7253 7 1 2 33746 33754
0 7254 5 1 1 7253
0 7255 7 1 2 7250 7254
0 7256 5 1 1 7255
0 7257 7 1 2 28531 7256
0 7258 5 1 1 7257
0 7259 7 2 2 30080 33400
0 7260 7 2 2 22791 23363
0 7261 7 4 2 22537 25239
0 7262 7 1 2 33757 33759
0 7263 7 1 2 33755 7262
0 7264 7 1 2 28345 7263
0 7265 7 1 2 30624 7264
0 7266 5 1 1 7265
0 7267 7 1 2 7258 7266
0 7268 5 1 1 7267
0 7269 7 1 2 21913 7268
0 7270 5 1 1 7269
0 7271 7 1 2 23007 30980
0 7272 5 1 1 7271
0 7273 7 1 2 31528 31207
0 7274 7 2 2 7272 7273
0 7275 5 1 1 33763
0 7276 7 1 2 28532 33747
0 7277 7 1 2 33764 7276
0 7278 5 1 1 7277
0 7279 7 1 2 7270 7278
0 7280 5 1 1 7279
0 7281 7 1 2 22918 7280
0 7282 5 1 1 7281
0 7283 7 2 2 24850 33656
0 7284 7 4 2 22646 29058
0 7285 5 3 1 33767
0 7286 7 1 2 31393 33771
0 7287 5 1 1 7286
0 7288 7 1 2 30973 7287
0 7289 5 1 1 7288
0 7290 7 1 2 7252 7289
0 7291 5 1 1 7290
0 7292 7 1 2 21914 7291
0 7293 5 1 1 7292
0 7294 7 1 2 7275 7293
0 7295 5 1 1 7294
0 7296 7 1 2 25585 28533
0 7297 7 2 2 7295 7296
0 7298 7 1 2 33765 33774
0 7299 5 1 1 7298
0 7300 7 1 2 7282 7299
0 7301 5 1 1 7300
0 7302 7 1 2 22388 7301
0 7303 5 1 1 7302
0 7304 7 1 2 33419 33775
0 7305 5 1 1 7304
0 7306 7 1 2 7303 7305
0 7307 5 1 1 7306
0 7308 7 1 2 33430 7307
0 7309 5 1 1 7308
0 7310 7 1 2 7206 7309
0 7311 5 1 1 7310
0 7312 7 1 2 27175 7311
0 7313 5 1 1 7312
0 7314 7 1 2 29071 31061
0 7315 5 3 1 7314
0 7316 7 2 2 31568 31292
0 7317 5 1 1 33779
0 7318 7 2 2 25699 26069
0 7319 7 1 2 25882 32629
0 7320 7 1 2 32924 7319
0 7321 7 1 2 33781 7320
0 7322 5 1 1 7321
0 7323 7 3 2 25473 32085
0 7324 7 8 2 24689 28912
0 7325 7 3 2 23828 30889
0 7326 5 11 1 33794
0 7327 7 2 2 33786 33797
0 7328 7 1 2 33783 33808
0 7329 5 1 1 7328
0 7330 7 6 2 25389 31168
0 7331 7 1 2 30522 30920
0 7332 5 1 1 7331
0 7333 7 2 2 25850 32630
0 7334 7 1 2 23524 33816
0 7335 5 1 1 7334
0 7336 7 1 2 7332 7335
0 7337 5 1 1 7336
0 7338 7 1 2 24851 7337
0 7339 5 1 1 7338
0 7340 7 2 2 26070 33474
0 7341 5 1 1 33818
0 7342 7 1 2 32631 33819
0 7343 5 1 1 7342
0 7344 7 1 2 7339 7343
0 7345 5 1 1 7344
0 7346 7 1 2 33810 7345
0 7347 5 1 1 7346
0 7348 7 1 2 7329 7347
0 7349 5 1 1 7348
0 7350 7 1 2 24381 25700
0 7351 7 1 2 7349 7350
0 7352 5 1 1 7351
0 7353 7 1 2 7322 7352
0 7354 5 1 1 7353
0 7355 7 1 2 33780 7354
0 7356 5 1 1 7355
0 7357 7 6 2 23432 33294
0 7358 7 1 2 28503 33820
0 7359 5 1 1 7358
0 7360 7 6 2 25390 30921
0 7361 7 1 2 25701 33826
0 7362 5 1 1 7361
0 7363 7 1 2 7359 7362
0 7364 5 1 1 7363
0 7365 7 1 2 22031 7364
0 7366 5 1 1 7365
0 7367 7 3 2 22472 22792
0 7368 7 2 2 22247 33832
0 7369 7 1 2 24946 32163
0 7370 7 1 2 33835 7369
0 7371 5 1 1 7370
0 7372 7 1 2 7366 7371
0 7373 5 1 1 7372
0 7374 7 1 2 30824 7373
0 7375 5 1 1 7374
0 7376 7 2 2 26849 33798
0 7377 7 2 2 29918 33837
0 7378 5 1 1 33839
0 7379 7 1 2 33295 33840
0 7380 5 1 1 7379
0 7381 7 1 2 7375 7380
0 7382 5 1 1 7381
0 7383 7 1 2 28799 7382
0 7384 5 1 1 7383
0 7385 7 1 2 26856 30779
0 7386 7 1 2 33152 7385
0 7387 5 1 1 7386
0 7388 7 1 2 7378 7387
0 7389 5 1 1 7388
0 7390 7 1 2 33513 7389
0 7391 5 1 1 7390
0 7392 7 1 2 7384 7391
0 7393 5 1 1 7392
0 7394 7 1 2 25474 7393
0 7395 5 1 1 7394
0 7396 7 2 2 25702 33153
0 7397 7 1 2 25851 30780
0 7398 7 1 2 29880 7397
0 7399 7 1 2 33841 7398
0 7400 5 1 1 7399
0 7401 7 1 2 7395 7400
0 7402 5 1 1 7401
0 7403 7 1 2 24852 7402
0 7404 5 1 1 7403
0 7405 7 3 2 22793 26793
0 7406 5 2 1 33843
0 7407 7 3 2 24738 28294
0 7408 5 1 1 33848
0 7409 7 1 2 33846 7408
0 7410 5 11 1 7409
0 7411 7 1 2 24261 33851
0 7412 5 1 1 7411
0 7413 7 2 2 25691 26794
0 7414 5 1 1 33862
0 7415 7 1 2 7412 7414
0 7416 5 5 1 7415
0 7417 7 1 2 22032 30825
0 7418 7 1 2 33864 7417
0 7419 5 1 1 7418
0 7420 7 9 2 24739 25475
0 7421 7 5 2 24065 24262
0 7422 7 3 2 33869 33878
0 7423 5 1 1 33883
0 7424 7 1 2 26572 31569
0 7425 7 1 2 33884 7424
0 7426 5 1 1 7425
0 7427 7 1 2 7419 7426
0 7428 5 1 1 7427
0 7429 7 1 2 32632 7428
0 7430 5 1 1 7429
0 7431 7 1 2 24066 31523
0 7432 5 2 1 7431
0 7433 7 3 2 22473 33886
0 7434 7 1 2 30826 33888
0 7435 7 1 2 33865 7434
0 7436 5 1 1 7435
0 7437 7 1 2 7430 7436
0 7438 5 2 1 7437
0 7439 7 1 2 26506 33891
0 7440 5 1 1 7439
0 7441 7 1 2 7404 7440
0 7442 5 1 1 7441
0 7443 7 1 2 24382 7442
0 7444 5 1 1 7443
0 7445 7 1 2 26071 25883
0 7446 7 1 2 33892 7445
0 7447 5 1 1 7446
0 7448 7 1 2 22747 7447
0 7449 7 1 2 7444 7448
0 7450 5 1 1 7449
0 7451 7 2 2 26015 29919
0 7452 5 1 1 33893
0 7453 7 1 2 25802 31131
0 7454 5 1 1 7453
0 7455 7 1 2 7452 7454
0 7456 5 1 1 7455
0 7457 7 3 2 22794 25476
0 7458 7 4 2 22248 24383
0 7459 7 1 2 24853 33898
0 7460 7 4 2 33895 7459
0 7461 5 1 1 33902
0 7462 7 1 2 33827 33903
0 7463 5 1 1 7462
0 7464 7 4 2 25703 25919
0 7465 7 3 2 32476 33906
0 7466 7 1 2 33910 33799
0 7467 5 1 1 7466
0 7468 7 1 2 7463 7467
0 7469 5 1 1 7468
0 7470 7 1 2 28800 7469
0 7471 5 1 1 7470
0 7472 7 21 2 25477 33344
0 7473 7 1 2 31821 33913
0 7474 7 1 2 33828 7473
0 7475 5 1 1 7474
0 7476 7 1 2 7471 7475
0 7477 5 1 1 7476
0 7478 7 1 2 7456 7477
0 7479 5 1 1 7478
0 7480 7 1 2 33022 33842
0 7481 5 1 1 7480
0 7482 7 2 2 22033 32633
0 7483 5 1 1 33934
0 7484 7 1 2 29031 33935
0 7485 5 1 1 7484
0 7486 7 1 2 32448 33889
0 7487 5 1 1 7486
0 7488 7 1 2 7485 7487
0 7489 5 1 1 7488
0 7490 7 1 2 33907 7489
0 7491 5 1 1 7490
0 7492 7 1 2 7481 7491
0 7493 5 1 1 7492
0 7494 7 7 2 25240 23433
0 7495 7 1 2 31490 33936
0 7496 7 1 2 7493 7495
0 7497 5 1 1 7496
0 7498 7 1 2 24690 7497
0 7499 7 1 2 7479 7498
0 7500 5 1 1 7499
0 7501 7 1 2 24206 7500
0 7502 7 1 2 7450 7501
0 7503 5 1 1 7502
0 7504 7 1 2 7356 7503
0 7505 5 1 1 7504
0 7506 7 1 2 23641 7505
0 7507 5 1 1 7506
0 7508 7 3 2 27879 32634
0 7509 5 1 1 33943
0 7510 7 9 2 22795 24854
0 7511 7 2 2 23434 33946
0 7512 7 1 2 33944 33955
0 7513 5 1 1 7512
0 7514 7 3 2 22796 22919
0 7515 7 3 2 30280 33957
0 7516 5 1 1 33960
0 7517 7 22 2 24740 25391
0 7518 5 1 1 33963
0 7519 7 1 2 26632 33964
0 7520 7 1 2 32722 7519
0 7521 5 1 1 7520
0 7522 7 1 2 7516 7521
0 7523 5 1 1 7522
0 7524 7 1 2 21915 7523
0 7525 5 1 1 7524
0 7526 7 1 2 29791 33961
0 7527 5 1 1 7526
0 7528 7 5 2 22474 24741
0 7529 7 3 2 21813 33985
0 7530 7 3 2 24855 25392
0 7531 7 2 2 26474 33993
0 7532 7 1 2 23955 33996
0 7533 7 1 2 33990 7532
0 7534 5 1 1 7533
0 7535 7 1 2 7527 7534
0 7536 7 1 2 7525 7535
0 7537 5 1 1 7536
0 7538 7 1 2 26072 7537
0 7539 5 1 1 7538
0 7540 7 1 2 7513 7539
0 7541 5 1 1 7540
0 7542 7 1 2 24263 7541
0 7543 5 1 1 7542
0 7544 7 4 2 23642 32086
0 7545 7 9 2 24742 23435
0 7546 5 2 1 34002
0 7547 7 2 2 22249 34003
0 7548 5 1 1 34013
0 7549 7 1 2 34014 32635
0 7550 7 1 2 33998 7549
0 7551 5 1 1 7550
0 7552 7 1 2 7543 7551
0 7553 5 1 1 7552
0 7554 7 1 2 24067 7553
0 7555 5 1 1 7554
0 7556 7 4 2 23956 23436
0 7557 7 1 2 25704 34015
0 7558 7 1 2 32723 7557
0 7559 7 1 2 33999 7558
0 7560 5 1 1 7559
0 7561 7 1 2 25478 7560
0 7562 7 1 2 7555 7561
0 7563 5 1 1 7562
0 7564 7 6 2 23288 27976
0 7565 7 4 2 24264 28801
0 7566 7 2 2 6246 6160
0 7567 5 3 1 34029
0 7568 7 1 2 24068 30894
0 7569 5 1 1 7568
0 7570 7 3 2 34030 7569
0 7571 5 6 1 34034
0 7572 7 8 2 24743 22920
0 7573 7 1 2 28928 34043
0 7574 7 1 2 34037 7573
0 7575 5 1 1 7574
0 7576 7 1 2 24069 33956
0 7577 7 1 2 32605 7576
0 7578 5 1 1 7577
0 7579 7 1 2 7575 7578
0 7580 5 1 1 7579
0 7581 7 1 2 34025 7580
0 7582 5 1 1 7581
0 7583 7 3 2 25393 33296
0 7584 5 1 1 34051
0 7585 7 1 2 34000 34038
0 7586 5 1 1 7585
0 7587 7 4 2 24070 24324
0 7588 7 2 2 24801 34054
0 7589 7 1 2 26633 34058
0 7590 7 1 2 30922 7589
0 7591 5 1 1 7590
0 7592 7 1 2 7586 7591
0 7593 5 1 1 7592
0 7594 7 1 2 34052 7593
0 7595 5 1 1 7594
0 7596 7 1 2 23525 7595
0 7597 7 1 2 7582 7596
0 7598 5 1 1 7597
0 7599 7 1 2 34019 7598
0 7600 7 1 2 7563 7599
0 7601 5 1 1 7600
0 7602 7 1 2 22250 24856
0 7603 7 7 2 33896 7602
0 7604 5 1 1 34060
0 7605 7 8 2 33475 33345
0 7606 5 3 1 34067
0 7607 7 1 2 7604 34075
0 7608 5 8 1 7607
0 7609 7 1 2 28802 34078
0 7610 5 2 1 7609
0 7611 7 1 2 33346 33784
0 7612 5 1 1 7611
0 7613 7 1 2 34086 7612
0 7614 5 1 1 7613
0 7615 7 2 2 23437 7614
0 7616 5 1 1 34088
0 7617 7 1 2 28504 34089
0 7618 5 1 1 7617
0 7619 7 1 2 24802 30212
0 7620 5 1 1 7619
0 7621 7 1 2 30505 30629
0 7622 7 1 2 7620 7621
0 7623 5 1 1 7622
0 7624 7 1 2 7341 7623
0 7625 5 1 1 7624
0 7626 7 1 2 27176 7625
0 7627 5 1 1 7626
0 7628 7 1 2 23526 30895
0 7629 7 1 2 32087 7628
0 7630 5 1 1 7629
0 7631 7 1 2 28574 30506
0 7632 7 1 2 30852 7631
0 7633 5 1 1 7632
0 7634 7 1 2 7630 7633
0 7635 7 1 2 7627 7634
0 7636 5 1 1 7635
0 7637 7 1 2 22251 33965
0 7638 7 1 2 7636 7637
0 7639 5 1 1 7638
0 7640 7 1 2 7618 7639
0 7641 5 1 1 7640
0 7642 7 1 2 22034 7641
0 7643 5 1 1 7642
0 7644 7 1 2 32088 33863
0 7645 5 1 1 7644
0 7646 7 1 2 7616 7645
0 7647 5 1 1 7646
0 7648 7 1 2 29977 7647
0 7649 5 1 1 7648
0 7650 7 1 2 7643 7649
0 7651 5 1 1 7650
0 7652 7 1 2 31684 32468
0 7653 7 1 2 7651 7652
0 7654 5 1 1 7653
0 7655 7 1 2 7601 7654
0 7656 5 1 1 7655
0 7657 7 1 2 24384 7656
0 7658 5 1 1 7657
0 7659 7 5 2 23643 25884
0 7660 7 2 2 24803 26795
0 7661 7 2 2 33556 34095
0 7662 5 1 1 34097
0 7663 7 18 2 22797 23438
0 7664 5 4 1 34099
0 7665 7 6 2 24265 25479
0 7666 7 2 2 34100 34121
0 7667 5 1 1 34127
0 7668 7 2 2 22252 33852
0 7669 5 2 1 34129
0 7670 7 1 2 7667 34131
0 7671 5 2 1 7670
0 7672 7 1 2 24804 34133
0 7673 5 1 1 7672
0 7674 7 12 2 23527 33347
0 7675 7 1 2 34135 32813
0 7676 5 1 1 7675
0 7677 7 1 2 7673 7676
0 7678 5 1 1 7677
0 7679 7 1 2 24325 7678
0 7680 5 1 1 7679
0 7681 7 1 2 7662 7680
0 7682 5 1 1 7681
0 7683 7 1 2 34020 34039
0 7684 7 1 2 7682 7683
0 7685 5 1 1 7684
0 7686 7 2 2 23439 32449
0 7687 7 1 2 24266 34147
0 7688 5 1 1 7687
0 7689 7 3 2 22253 24326
0 7690 7 1 2 34096 34149
0 7691 5 1 1 7690
0 7692 7 1 2 7688 7691
0 7693 5 1 1 7692
0 7694 7 4 2 22647 24744
0 7695 7 2 2 34152 32777
0 7696 7 1 2 33154 34156
0 7697 7 1 2 7693 7696
0 7698 5 1 1 7697
0 7699 7 1 2 7685 7698
0 7700 5 1 1 7699
0 7701 7 1 2 34090 7700
0 7702 5 1 1 7701
0 7703 7 1 2 7658 7702
0 7704 5 1 1 7703
0 7705 7 1 2 32965 7704
0 7706 5 1 1 7705
0 7707 7 1 2 25329 31913
0 7708 7 2 2 31894 7707
0 7709 5 1 1 34158
0 7710 7 4 2 25330 32477
0 7711 7 1 2 34160 31939
0 7712 5 1 1 7711
0 7713 7 1 2 24805 33213
0 7714 5 1 1 7713
0 7715 7 1 2 7712 7714
0 7716 5 1 1 7715
0 7717 7 1 2 24327 7716
0 7718 5 1 1 7717
0 7719 7 1 2 7709 7718
0 7720 5 1 1 7719
0 7721 7 1 2 25920 7720
0 7722 5 1 1 7721
0 7723 7 3 2 31806 31958
0 7724 7 1 2 32925 34164
0 7725 5 1 1 7724
0 7726 7 1 2 7722 7725
0 7727 5 1 1 7726
0 7728 7 1 2 23957 23644
0 7729 7 1 2 7727 7728
0 7730 5 1 1 7729
0 7731 7 5 2 24857 25331
0 7732 7 1 2 24385 34167
0 7733 7 1 2 34055 7732
0 7734 7 2 2 28073 30299
0 7735 7 1 2 28143 34172
0 7736 7 1 2 7733 7735
0 7737 5 1 1 7736
0 7738 7 1 2 7730 7737
0 7739 5 1 1 7738
0 7740 7 1 2 25705 7739
0 7741 5 1 1 7740
0 7742 7 11 2 24267 24328
0 7743 7 9 2 24745 34174
0 7744 7 5 2 26496 34185
0 7745 5 1 1 34194
0 7746 7 1 2 24858 33522
0 7747 5 1 1 7746
0 7748 7 1 2 7745 7747
0 7749 5 1 1 7748
0 7750 7 1 2 24386 7749
0 7751 5 1 1 7750
0 7752 7 4 2 24268 27648
0 7753 7 4 2 24746 24859
0 7754 7 4 2 24806 34203
0 7755 7 5 2 34199 34207
0 7756 5 1 1 34211
0 7757 7 1 2 7751 7756
0 7758 5 4 1 7757
0 7759 7 4 2 23645 34216
0 7760 7 2 2 26834 31900
0 7761 7 1 2 33251 34224
0 7762 7 1 2 34220 7761
0 7763 5 1 1 7762
0 7764 7 1 2 7741 7763
0 7765 5 1 1 7764
0 7766 7 1 2 31570 7765
0 7767 5 1 1 7766
0 7768 7 1 2 31693 31718
0 7769 7 3 2 25241 33450
0 7770 7 4 2 25332 27029
0 7771 7 1 2 34226 34229
0 7772 7 1 2 33446 7771
0 7773 7 1 2 7768 7772
0 7774 5 1 1 7773
0 7775 7 1 2 7767 7774
0 7776 5 1 1 7775
0 7777 7 1 2 32724 7776
0 7778 5 1 1 7777
0 7779 7 5 2 25586 26110
0 7780 7 2 2 30781 31372
0 7781 5 1 1 34238
0 7782 7 1 2 7781 7317
0 7783 5 3 1 7782
0 7784 7 1 2 31914 33811
0 7785 5 1 1 7784
0 7786 7 1 2 30630 33161
0 7787 5 1 1 7786
0 7788 7 1 2 7785 7787
0 7789 5 1 1 7788
0 7790 7 1 2 24329 7789
0 7791 5 1 1 7790
0 7792 7 1 2 32441 33787
0 7793 5 1 1 7792
0 7794 7 1 2 7791 7793
0 7795 5 3 1 7794
0 7796 7 1 2 30847 34243
0 7797 5 1 1 7796
0 7798 7 1 2 1948 4377
0 7799 5 1 1 7798
0 7800 7 1 2 974 1750
0 7801 7 2 2 7799 7800
0 7802 7 1 2 24330 34246
0 7803 5 1 1 7802
0 7804 7 1 2 28617 33788
0 7805 5 1 1 7804
0 7806 7 1 2 7803 7805
0 7807 5 1 1 7806
0 7808 7 1 2 23528 30909
0 7809 7 1 2 7807 7808
0 7810 5 1 1 7809
0 7811 7 1 2 7797 7810
0 7812 5 1 1 7811
0 7813 7 1 2 34240 7812
0 7814 5 1 1 7813
0 7815 7 1 2 28517 30923
0 7816 5 1 1 7815
0 7817 7 1 2 28511 30910
0 7818 5 1 1 7817
0 7819 7 1 2 7816 7818
0 7820 5 1 1 7819
0 7821 7 1 2 23364 7820
0 7822 5 1 1 7821
0 7823 7 1 2 28415 31157
0 7824 7 1 2 33258 7823
0 7825 5 1 1 7824
0 7826 7 1 2 7822 7825
0 7827 5 1 1 7826
0 7828 7 2 2 28295 26073
0 7829 7 2 2 23289 29920
0 7830 7 1 2 34248 34250
0 7831 7 1 2 7827 7830
0 7832 5 1 1 7831
0 7833 7 1 2 7814 7832
0 7834 5 1 1 7833
0 7835 7 1 2 25706 7834
0 7836 5 1 1 7835
0 7837 7 3 2 24691 31223
0 7838 5 1 1 34252
0 7839 7 3 2 23958 22475
0 7840 7 2 2 21814 34255
0 7841 7 1 2 34253 34258
0 7842 5 1 1 7841
0 7843 7 2 2 27506 31244
0 7844 5 1 1 34260
0 7845 7 1 2 21916 34261
0 7846 5 1 1 7845
0 7847 7 1 2 7842 7846
0 7848 5 1 1 7847
0 7849 7 3 2 22648 34186
0 7850 7 8 2 22200 33937
0 7851 7 2 2 22035 28575
0 7852 7 1 2 34265 34273
0 7853 7 1 2 34262 7852
0 7854 7 1 2 7848 7853
0 7855 5 1 1 7854
0 7856 7 1 2 7836 7855
0 7857 5 1 1 7856
0 7858 7 1 2 34233 7857
0 7859 5 1 1 7858
0 7860 7 1 2 7778 7859
0 7861 7 1 2 7706 7860
0 7862 7 1 2 7507 7861
0 7863 5 1 1 7862
0 7864 7 1 2 25667 7863
0 7865 5 1 1 7864
0 7866 7 4 2 24692 26573
0 7867 5 1 1 34275
0 7868 7 6 2 22748 26857
0 7869 5 3 1 34279
0 7870 7 1 2 7867 34285
0 7871 5 22 1 7870
0 7872 7 8 2 23290 31228
0 7873 7 3 2 30300 33485
0 7874 5 2 1 34318
0 7875 7 1 2 32670 34319
0 7876 5 1 1 7875
0 7877 7 2 2 25668 34040
0 7878 7 1 2 23646 34136
0 7879 7 1 2 34323 7878
0 7880 5 1 1 7879
0 7881 7 2 2 7876 7880
0 7882 5 1 1 34325
0 7883 7 1 2 34310 7882
0 7884 5 1 1 7883
0 7885 7 3 2 24207 22649
0 7886 7 2 2 25242 34327
0 7887 7 2 2 24269 33986
0 7888 7 1 2 30097 34332
0 7889 5 1 1 7888
0 7890 7 1 2 34321 7889
0 7891 5 1 1 7890
0 7892 7 1 2 33887 7891
0 7893 5 1 1 7892
0 7894 7 3 2 22036 33348
0 7895 7 1 2 30098 33800
0 7896 7 1 2 34334 7895
0 7897 5 1 1 7896
0 7898 7 7 2 25480 23744
0 7899 7 1 2 21917 26475
0 7900 7 1 2 34337 7899
0 7901 7 1 2 33836 7900
0 7902 5 1 1 7901
0 7903 7 1 2 7897 7902
0 7904 7 2 2 7893 7903
0 7905 5 1 1 34344
0 7906 7 1 2 34330 7905
0 7907 5 1 1 7906
0 7908 7 1 2 7884 7907
0 7909 5 1 1 7908
0 7910 7 1 2 28803 7909
0 7911 5 1 1 7910
0 7912 7 11 2 24270 33870
0 7913 5 1 1 34346
0 7914 7 1 2 33632 7913
0 7915 5 16 1 7914
0 7916 7 1 2 34357 34311
0 7917 7 1 2 34041 7916
0 7918 5 1 1 7917
0 7919 7 6 2 24208 22254
0 7920 7 8 2 22650 22798
0 7921 7 4 2 25243 23529
0 7922 7 3 2 34379 34387
0 7923 7 1 2 34373 34391
0 7924 7 1 2 33155 7923
0 7925 5 1 1 7924
0 7926 7 1 2 7918 7925
0 7927 5 1 1 7926
0 7928 7 1 2 27607 7927
0 7929 5 1 1 7928
0 7930 7 1 2 34312 32671
0 7931 5 1 1 7930
0 7932 7 3 2 25244 32292
0 7933 7 1 2 34328 34394
0 7934 5 1 1 7933
0 7935 7 1 2 7931 7934
0 7936 5 3 1 7935
0 7937 7 1 2 33914 34397
0 7938 5 1 1 7937
0 7939 7 24 2 23530 33297
0 7940 5 2 1 34400
0 7941 7 1 2 27857 34401
0 7942 7 1 2 34313 7941
0 7943 5 1 1 7942
0 7944 7 1 2 7938 7943
0 7945 5 1 1 7944
0 7946 7 1 2 27622 7945
0 7947 5 1 1 7946
0 7948 7 1 2 7929 7947
0 7949 7 1 2 7911 7948
0 7950 5 1 1 7949
0 7951 7 1 2 25921 7950
0 7952 5 1 1 7951
0 7953 7 8 2 28641 33298
0 7954 5 2 1 34426
0 7955 7 2 2 27778 32502
0 7956 5 1 1 34436
0 7957 7 1 2 26111 34324
0 7958 5 1 1 7957
0 7959 7 1 2 7956 7958
0 7960 5 1 1 7959
0 7961 7 1 2 34427 7960
0 7962 5 1 1 7961
0 7963 7 8 2 28671 33349
0 7964 5 1 1 34438
0 7965 7 1 2 27779 27858
0 7966 7 1 2 34439 7965
0 7967 5 1 1 7966
0 7968 7 1 2 7962 7967
0 7969 5 1 1 7968
0 7970 7 1 2 28804 7969
0 7971 5 1 1 7970
0 7972 7 2 2 29724 33299
0 7973 5 2 1 34446
0 7974 7 4 2 23959 24271
0 7975 7 2 2 33871 34450
0 7976 5 1 1 34454
0 7977 7 1 2 34448 7976
0 7978 5 1 1 7977
0 7979 7 1 2 27507 7978
0 7980 5 1 1 7979
0 7981 7 2 2 23008 29351
0 7982 5 1 1 34456
0 7983 7 1 2 33915 34457
0 7984 5 1 1 7983
0 7985 7 1 2 7980 7984
0 7986 5 1 1 7985
0 7987 7 1 2 27661 7986
0 7988 5 1 1 7987
0 7989 7 1 2 34347 34042
0 7990 5 1 1 7989
0 7991 7 1 2 33620 34031
0 7992 5 1 1 7991
0 7993 7 1 2 7990 7992
0 7994 5 1 1 7993
0 7995 7 1 2 27732 7994
0 7996 5 1 1 7995
0 7997 7 7 2 33582 34044
0 7998 7 1 2 34458 34338
0 7999 7 1 2 32503 7998
0 8000 5 1 1 7999
0 8001 7 1 2 7996 8000
0 8002 5 1 1 8001
0 8003 7 1 2 27713 8002
0 8004 5 1 1 8003
0 8005 7 1 2 7988 8004
0 8006 7 1 2 7971 8005
0 8007 5 1 1 8006
0 8008 7 1 2 34314 8007
0 8009 5 1 1 8008
0 8010 7 2 2 27995 34187
0 8011 7 3 2 25481 34465
0 8012 7 1 2 21918 31032
0 8013 5 1 1 8012
0 8014 7 1 2 32665 8013
0 8015 5 4 1 8014
0 8016 7 1 2 34467 34470
0 8017 5 2 1 8016
0 8018 7 1 2 27900 30853
0 8019 5 1 1 8018
0 8020 7 1 2 27714 30896
0 8021 5 1 1 8020
0 8022 7 1 2 8019 8021
0 8023 5 1 1 8022
0 8024 7 1 2 33300 8023
0 8025 5 1 1 8024
0 8026 7 1 2 30854 33714
0 8027 5 1 1 8026
0 8028 7 1 2 8025 8027
0 8029 5 1 1 8028
0 8030 7 1 2 23531 8029
0 8031 5 1 1 8030
0 8032 7 1 2 34474 8031
0 8033 5 1 1 8032
0 8034 7 1 2 27733 8033
0 8035 5 1 1 8034
0 8036 7 6 2 24272 22921
0 8037 7 9 2 22389 24747
0 8038 7 2 2 26074 34482
0 8039 7 2 2 34476 34491
0 8040 5 1 1 34493
0 8041 7 1 2 31151 34494
0 8042 5 1 1 8041
0 8043 7 1 2 8035 8042
0 8044 5 1 1 8043
0 8045 7 1 2 34241 8044
0 8046 5 1 1 8045
0 8047 7 1 2 24807 28728
0 8048 7 1 2 31775 33171
0 8049 7 1 2 8047 8048
0 8050 7 1 2 30316 8049
0 8051 7 1 2 34263 8050
0 8052 5 1 1 8051
0 8053 7 1 2 30207 34242
0 8054 7 1 2 33748 8053
0 8055 5 1 1 8054
0 8056 7 1 2 22255 34380
0 8057 7 1 2 27880 8056
0 8058 7 1 2 31812 8057
0 8059 5 1 1 8058
0 8060 7 1 2 8055 8059
0 8061 5 1 1 8060
0 8062 7 1 2 23532 27734
0 8063 7 1 2 8061 8062
0 8064 5 1 1 8063
0 8065 7 1 2 8052 8064
0 8066 5 1 1 8065
0 8067 7 1 2 27177 8066
0 8068 5 1 1 8067
0 8069 7 2 2 22476 27985
0 8070 7 4 2 27674 33650
0 8071 7 1 2 29429 34374
0 8072 7 1 2 30787 8071
0 8073 7 1 2 34497 8072
0 8074 7 1 2 34495 8073
0 8075 5 1 1 8074
0 8076 7 1 2 8068 8075
0 8077 7 1 2 8046 8076
0 8078 7 1 2 8009 8077
0 8079 7 1 2 7952 8078
0 8080 5 1 1 8079
0 8081 7 1 2 34288 8080
0 8082 5 1 1 8081
0 8083 7 2 2 33301 33006
0 8084 7 1 2 29921 34501
0 8085 5 1 1 8084
0 8086 7 1 2 25707 31685
0 8087 7 1 2 34395 8086
0 8088 5 1 1 8087
0 8089 7 1 2 8085 8088
0 8090 5 1 1 8089
0 8091 7 1 2 24808 8090
0 8092 5 1 1 8091
0 8093 7 9 2 24209 24273
0 8094 7 2 2 24071 34503
0 8095 7 3 2 24601 22861
0 8096 7 2 2 24748 23291
0 8097 7 2 2 34514 34517
0 8098 7 1 2 34512 34519
0 8099 5 1 1 8098
0 8100 7 1 2 8092 8099
0 8101 5 1 1 8100
0 8102 7 1 2 24331 8101
0 8103 5 1 1 8102
0 8104 7 2 2 33007 32397
0 8105 7 1 2 33441 33879
0 8106 7 1 2 34521 8105
0 8107 5 1 1 8106
0 8108 7 1 2 8103 8107
0 8109 5 1 1 8108
0 8110 7 1 2 22390 33476
0 8111 7 1 2 8109 8110
0 8112 5 1 1 8111
0 8113 7 1 2 32293 34157
0 8114 5 2 1 8113
0 8115 7 2 2 22799 23292
0 8116 7 3 2 27977 34525
0 8117 7 1 2 24072 34527
0 8118 5 1 1 8117
0 8119 7 1 2 34523 8118
0 8120 5 1 1 8119
0 8121 7 1 2 30737 8120
0 8122 5 1 1 8121
0 8123 7 1 2 30523 34528
0 8124 7 1 2 28219 8123
0 8125 5 1 1 8124
0 8126 7 1 2 8122 8125
0 8127 5 1 1 8126
0 8128 7 1 2 22256 8127
0 8129 5 1 1 8128
0 8130 7 1 2 25852 33451
0 8131 7 1 2 34392 8130
0 8132 7 1 2 32294 8131
0 8133 5 1 1 8132
0 8134 7 1 2 8129 8133
0 8135 5 1 1 8134
0 8136 7 1 2 25922 8135
0 8137 5 1 1 8136
0 8138 7 1 2 25394 8137
0 8139 7 1 2 8112 8138
0 8140 5 1 1 8139
0 8141 7 3 2 25482 25982
0 8142 7 1 2 32672 34529
0 8143 5 1 1 8142
0 8144 7 1 2 34524 8143
0 8145 5 1 1 8144
0 8146 7 1 2 34530 8145
0 8147 5 1 1 8146
0 8148 7 2 2 22391 34021
0 8149 7 7 2 24332 22800
0 8150 7 3 2 23533 34535
0 8151 7 1 2 28258 34542
0 8152 7 1 2 32504 8151
0 8153 7 1 2 34533 8152
0 8154 5 1 1 8153
0 8155 7 1 2 8147 8154
0 8156 5 1 1 8155
0 8157 7 1 2 24274 8156
0 8158 5 1 1 8157
0 8159 7 1 2 23440 8158
0 8160 5 1 1 8159
0 8161 7 1 2 27405 8160
0 8162 7 1 2 8140 8161
0 8163 5 1 1 8162
0 8164 7 1 2 34045 34339
0 8165 7 2 2 34534 8164
0 8166 7 1 2 32673 34545
0 8167 5 1 1 8166
0 8168 7 2 2 26112 33105
0 8169 7 2 2 32517 34547
0 8170 7 1 2 34549 34393
0 8171 5 1 1 8170
0 8172 7 1 2 8167 8171
0 8173 5 1 1 8172
0 8174 7 1 2 26075 8173
0 8175 5 1 1 8174
0 8176 7 2 2 34381 33106
0 8177 7 4 2 25245 25483
0 8178 7 1 2 27821 34553
0 8179 7 1 2 34551 8178
0 8180 5 1 1 8179
0 8181 7 8 2 24073 24210
0 8182 7 1 2 23534 34557
0 8183 7 1 2 34518 8182
0 8184 7 1 2 29773 8183
0 8185 7 1 2 30855 8184
0 8186 5 1 1 8185
0 8187 7 1 2 8180 8186
0 8188 5 1 1 8187
0 8189 7 1 2 24387 8188
0 8190 5 1 1 8189
0 8191 7 1 2 24388 29288
0 8192 7 1 2 30285 34204
0 8193 7 1 2 8191 8192
0 8194 7 1 2 34022 8193
0 8195 5 1 1 8194
0 8196 7 1 2 32200 34554
0 8197 7 1 2 34382 8196
0 8198 7 1 2 32126 8197
0 8199 5 1 1 8198
0 8200 7 1 2 8195 8199
0 8201 5 1 1 8200
0 8202 7 1 2 29625 8201
0 8203 5 1 1 8202
0 8204 7 2 2 25246 28437
0 8205 7 1 2 33107 34340
0 8206 7 1 2 33947 8205
0 8207 7 1 2 34565 8206
0 8208 5 1 1 8207
0 8209 7 1 2 8203 8208
0 8210 7 1 2 8190 8209
0 8211 5 1 1 8210
0 8212 7 1 2 28805 8211
0 8213 5 1 1 8212
0 8214 7 1 2 25484 28267
0 8215 7 1 2 34520 8214
0 8216 7 1 2 32127 8215
0 8217 7 1 2 32674 8216
0 8218 5 1 1 8217
0 8219 7 1 2 25587 8218
0 8220 7 1 2 8213 8219
0 8221 7 1 2 8175 8220
0 8222 5 1 1 8221
0 8223 7 3 2 24275 25395
0 8224 5 1 1 34567
0 8225 7 2 2 22257 23441
0 8226 5 1 1 34570
0 8227 7 1 2 8224 8226
0 8228 5 2 1 8227
0 8229 7 1 2 32505 34546
0 8230 5 1 1 8229
0 8231 7 2 2 25669 31714
0 8232 7 1 2 30788 33948
0 8233 7 1 2 34574 8232
0 8234 7 1 2 33156 8233
0 8235 5 1 1 8234
0 8236 7 1 2 8230 8235
0 8237 5 1 1 8236
0 8238 7 1 2 25853 8237
0 8239 5 1 1 8238
0 8240 7 1 2 30286 34383
0 8241 7 1 2 32778 8240
0 8242 7 1 2 31816 8241
0 8243 7 1 2 33157 8242
0 8244 5 1 1 8243
0 8245 7 1 2 23647 8244
0 8246 7 1 2 8239 8245
0 8247 5 1 1 8246
0 8248 7 1 2 34572 8247
0 8249 7 1 2 8222 8248
0 8250 5 1 1 8249
0 8251 7 1 2 1042 28806
0 8252 7 2 2 34117 7518
0 8253 5 16 1 34576
0 8254 7 1 2 462 1291
0 8255 5 1 1 8254
0 8256 7 1 2 34577 8255
0 8257 7 4 2 8251 8256
0 8258 5 1 1 34594
0 8259 7 3 2 22258 24602
0 8260 7 1 2 33008 34598
0 8261 7 1 2 34437 8260
0 8262 5 1 1 8261
0 8263 7 1 2 30782 33452
0 8264 7 1 2 32603 8263
0 8265 7 1 2 30924 8264
0 8266 5 1 1 8265
0 8267 7 1 2 8262 8266
0 8268 5 1 1 8267
0 8269 7 1 2 34595 8268
0 8270 5 1 1 8269
0 8271 7 1 2 30401 34153
0 8272 7 1 2 34150 8271
0 8273 7 1 2 34550 8272
0 8274 5 1 1 8273
0 8275 7 1 2 22392 23745
0 8276 7 1 2 25689 8275
0 8277 7 1 2 32154 8276
0 8278 7 1 2 34522 8277
0 8279 7 1 2 32506 8278
0 8280 5 1 1 8279
0 8281 7 1 2 8274 8280
0 8282 5 1 1 8281
0 8283 7 1 2 28693 8282
0 8284 5 1 1 8283
0 8285 7 1 2 8270 8284
0 8286 7 1 2 8250 8285
0 8287 7 1 2 8163 8286
0 8288 5 1 1 8287
0 8289 7 1 2 32966 8288
0 8290 5 1 1 8289
0 8291 7 2 2 28706 33812
0 8292 5 1 1 34601
0 8293 7 1 2 22317 34247
0 8294 5 1 1 8293
0 8295 7 1 2 8292 8294
0 8296 5 3 1 8295
0 8297 7 1 2 25923 34603
0 8298 5 1 1 8297
0 8299 7 1 2 25974 33789
0 8300 5 1 1 8299
0 8301 7 1 2 8298 8300
0 8302 5 2 1 8301
0 8303 7 1 2 25588 34606
0 8304 7 1 2 34398 8303
0 8305 5 1 1 8304
0 8306 7 1 2 26338 34315
0 8307 7 1 2 32507 8306
0 8308 7 1 2 34604 8307
0 8309 5 1 1 8308
0 8310 7 1 2 8305 8309
0 8311 5 1 1 8310
0 8312 7 1 2 25485 8311
0 8313 5 1 1 8312
0 8314 7 2 2 25983 33813
0 8315 7 1 2 34608 34399
0 8316 5 1 1 8315
0 8317 7 2 2 27928 31229
0 8318 7 1 2 23442 28271
0 8319 7 1 2 34610 8318
0 8320 7 1 2 32508 8319
0 8321 7 1 2 33392 8320
0 8322 5 1 1 8321
0 8323 7 1 2 8316 8322
0 8324 5 1 1 8323
0 8325 7 1 2 28672 8324
0 8326 5 1 1 8325
0 8327 7 1 2 8313 8326
0 8328 5 1 1 8327
0 8329 7 1 2 25708 8328
0 8330 5 1 1 8329
0 8331 7 2 2 28220 26016
0 8332 7 1 2 24603 34612
0 8333 5 1 1 8332
0 8334 7 1 2 31491 34396
0 8335 5 1 1 8334
0 8336 7 1 2 8333 8335
0 8337 5 1 1 8336
0 8338 7 1 2 24693 8337
0 8339 5 1 1 8338
0 8340 7 2 2 22749 27859
0 8341 7 2 2 24604 27929
0 8342 7 1 2 34614 34616
0 8343 5 1 1 8342
0 8344 7 1 2 8339 8343
0 8345 5 1 1 8344
0 8346 7 1 2 24211 8345
0 8347 5 1 1 8346
0 8348 7 1 2 24074 24694
0 8349 7 1 2 34611 8348
0 8350 5 1 1 8349
0 8351 7 1 2 8347 8350
0 8352 5 1 1 8351
0 8353 7 1 2 25396 8352
0 8354 5 1 1 8353
0 8355 7 1 2 31169 34016
0 8356 7 1 2 34316 8355
0 8357 5 1 1 8356
0 8358 7 1 2 8354 8357
0 8359 5 1 1 8358
0 8360 7 2 2 28673 33425
0 8361 7 1 2 8359 34618
0 8362 5 1 1 8361
0 8363 7 1 2 8330 8362
0 8364 5 1 1 8363
0 8365 7 1 2 23746 8364
0 8366 5 1 1 8365
0 8367 7 1 2 8290 8366
0 8368 7 1 2 8082 8367
0 8369 7 1 2 7865 8368
0 8370 5 1 1 8369
0 8371 7 1 2 33776 8370
0 8372 5 1 1 8371
0 8373 7 1 2 28047 32209
0 8374 7 1 2 26031 8373
0 8375 5 1 1 8374
0 8376 7 2 2 24947 26278
0 8377 5 1 1 34620
0 8378 7 1 2 26321 8377
0 8379 5 1 1 8378
0 8380 7 1 2 22477 32307
0 8381 7 1 2 8379 8380
0 8382 5 1 1 8381
0 8383 7 1 2 8375 8382
0 8384 5 1 1 8383
0 8385 7 1 2 21815 8384
0 8386 5 1 1 8385
0 8387 7 2 2 26017 27328
0 8388 7 1 2 30141 34622
0 8389 5 1 1 8388
0 8390 7 1 2 24474 34621
0 8391 5 1 1 8390
0 8392 7 1 2 8389 8391
0 8393 5 1 1 8392
0 8394 7 1 2 23829 8393
0 8395 5 1 1 8394
0 8396 7 1 2 26316 27379
0 8397 5 1 1 8396
0 8398 7 1 2 8395 8397
0 8399 5 1 1 8398
0 8400 7 1 2 23960 8399
0 8401 5 1 1 8400
0 8402 7 1 2 25803 30432
0 8403 5 1 1 8402
0 8404 7 1 2 8401 8403
0 8405 5 1 1 8404
0 8406 7 1 2 22037 8405
0 8407 5 1 1 8406
0 8408 7 1 2 8386 8407
0 8409 5 1 1 8408
0 8410 7 1 2 22538 8409
0 8411 5 1 1 8410
0 8412 7 1 2 30273 32534
0 8413 7 1 2 26317 8412
0 8414 7 1 2 31410 8413
0 8415 5 1 1 8414
0 8416 7 1 2 8411 8415
0 8417 5 1 1 8416
0 8418 7 1 2 23098 8417
0 8419 5 1 1 8418
0 8420 7 1 2 22651 26028
0 8421 5 2 1 8420
0 8422 7 1 2 24524 30129
0 8423 5 1 1 8422
0 8424 7 1 2 34624 8423
0 8425 5 1 1 8424
0 8426 7 1 2 29499 31310
0 8427 7 1 2 30877 8426
0 8428 7 1 2 8425 8427
0 8429 5 1 1 8428
0 8430 7 1 2 8419 8429
0 8431 5 1 1 8430
0 8432 7 1 2 27735 8431
0 8433 5 1 1 8432
0 8434 7 3 2 30064 32329
0 8435 7 1 2 31304 34626
0 8436 5 1 1 8435
0 8437 7 1 2 25247 30347
0 8438 5 1 1 8437
0 8439 7 2 2 22539 25817
0 8440 7 2 2 21919 34629
0 8441 7 1 2 30222 34631
0 8442 5 1 1 8441
0 8443 7 1 2 8438 8442
0 8444 5 3 1 8443
0 8445 7 1 2 23365 31311
0 8446 7 1 2 34633 8445
0 8447 5 1 1 8446
0 8448 7 1 2 8436 8447
0 8449 5 3 1 8448
0 8450 7 1 2 27780 34636
0 8451 5 1 1 8450
0 8452 7 1 2 8433 8451
0 8453 5 1 1 8452
0 8454 7 1 2 26076 8453
0 8455 5 1 1 8454
0 8456 7 1 2 32123 34637
0 8457 5 1 1 8456
0 8458 7 1 2 8455 8457
0 8459 5 1 1 8458
0 8460 7 1 2 33350 8459
0 8461 5 1 1 8460
0 8462 7 1 2 33518 32128
0 8463 7 1 2 34638 8462
0 8464 5 1 1 8463
0 8465 7 1 2 8461 8464
0 8466 5 1 1 8465
0 8467 7 1 2 22750 8466
0 8468 5 1 1 8467
0 8469 7 1 2 33540 8040
0 8470 5 3 1 8469
0 8471 7 2 2 22038 23747
0 8472 7 1 2 27443 32951
0 8473 7 1 2 34642 8472
0 8474 7 1 2 34639 8473
0 8475 7 1 2 34634 8474
0 8476 5 1 1 8475
0 8477 7 1 2 25486 8476
0 8478 7 1 2 8468 8477
0 8479 5 1 1 8478
0 8480 7 1 2 23099 32853
0 8481 5 1 1 8480
0 8482 7 1 2 29997 32330
0 8483 5 1 1 8482
0 8484 7 1 2 28484 32797
0 8485 5 1 1 8484
0 8486 7 1 2 8483 8485
0 8487 5 1 1 8486
0 8488 7 1 2 27781 8487
0 8489 5 1 1 8488
0 8490 7 1 2 8481 8489
0 8491 5 1 1 8490
0 8492 7 1 2 24075 8491
0 8493 5 1 1 8492
0 8494 7 2 2 23748 28485
0 8495 7 4 2 24525 22922
0 8496 7 1 2 23293 34646
0 8497 7 1 2 29376 8496
0 8498 7 1 2 34644 8497
0 8499 5 1 1 8498
0 8500 7 1 2 8493 8499
0 8501 5 1 1 8500
0 8502 7 1 2 25333 8501
0 8503 5 1 1 8502
0 8504 7 1 2 30611 31574
0 8505 5 2 1 8504
0 8506 7 2 2 23207 32455
0 8507 5 1 1 34652
0 8508 7 1 2 25059 34653
0 8509 5 1 1 8508
0 8510 7 1 2 34650 8509
0 8511 5 1 1 8510
0 8512 7 1 2 25248 8511
0 8513 5 1 1 8512
0 8514 7 2 2 23294 32456
0 8515 7 1 2 28507 34654
0 8516 5 1 1 8515
0 8517 7 1 2 8513 8516
0 8518 5 1 1 8517
0 8519 7 1 2 24948 8518
0 8520 5 1 1 8519
0 8521 7 1 2 31067 33760
0 8522 5 1 1 8521
0 8523 7 1 2 8520 8522
0 8524 5 1 1 8523
0 8525 7 1 2 22039 8524
0 8526 5 1 1 8525
0 8527 7 1 2 25249 31074
0 8528 5 1 1 8527
0 8529 7 2 2 8526 8528
0 8530 5 1 1 34656
0 8531 7 1 2 23366 27842
0 8532 7 1 2 8530 8531
0 8533 5 1 1 8532
0 8534 7 1 2 8503 8533
0 8535 5 1 1 8534
0 8536 7 1 2 22751 8535
0 8537 5 1 1 8536
0 8538 7 1 2 29066 32142
0 8539 5 1 1 8538
0 8540 7 1 2 29932 29500
0 8541 7 1 2 8539 8540
0 8542 5 1 1 8541
0 8543 7 1 2 31336 32251
0 8544 5 1 1 8543
0 8545 7 1 2 27444 33768
0 8546 5 1 1 8545
0 8547 7 1 2 8544 8546
0 8548 7 1 2 8542 8547
0 8549 5 1 1 8548
0 8550 7 1 2 24949 8549
0 8551 5 1 1 8550
0 8552 7 1 2 27445 28602
0 8553 5 1 1 8552
0 8554 7 3 2 24950 29765
0 8555 7 1 2 30612 34658
0 8556 5 1 1 8555
0 8557 7 1 2 8553 8556
0 8558 5 1 1 8557
0 8559 7 1 2 31189 8558
0 8560 5 1 1 8559
0 8561 7 7 2 24076 25060
0 8562 7 1 2 26305 34661
0 8563 5 1 1 8562
0 8564 7 1 2 22040 31068
0 8565 5 1 1 8564
0 8566 7 1 2 8563 8565
0 8567 5 1 1 8566
0 8568 7 1 2 22540 8567
0 8569 5 1 1 8568
0 8570 7 1 2 8560 8569
0 8571 7 1 2 8551 8570
0 8572 5 3 1 8571
0 8573 7 1 2 25250 34668
0 8574 5 1 1 8573
0 8575 7 3 2 26884 31495
0 8576 7 1 2 32461 34671
0 8577 5 1 1 8576
0 8578 7 1 2 8574 8577
0 8579 5 2 1 8578
0 8580 7 1 2 27843 32952
0 8581 7 1 2 34674 8580
0 8582 5 1 1 8581
0 8583 7 1 2 8537 8582
0 8584 5 1 1 8583
0 8585 7 1 2 33732 8584
0 8586 5 1 1 8585
0 8587 7 1 2 23367 34657
0 8588 5 1 1 8587
0 8589 7 1 2 25334 34675
0 8590 5 1 1 8589
0 8591 7 1 2 24695 8590
0 8592 5 1 1 8591
0 8593 7 2 2 29140 31433
0 8594 5 2 1 34676
0 8595 7 1 2 29059 31183
0 8596 5 2 1 8595
0 8597 7 1 2 32413 34680
0 8598 5 1 1 8597
0 8599 7 1 2 24475 8598
0 8600 5 1 1 8599
0 8601 7 1 2 34678 8600
0 8602 5 2 1 8601
0 8603 7 1 2 23295 34682
0 8604 5 1 1 8603
0 8605 7 1 2 29595 30551
0 8606 5 1 1 8605
0 8607 7 1 2 2023 8606
0 8608 5 1 1 8607
0 8609 7 1 2 30468 8608
0 8610 5 1 1 8609
0 8611 7 1 2 8604 8610
0 8612 5 1 1 8611
0 8613 7 1 2 23830 8612
0 8614 5 1 1 8613
0 8615 7 1 2 31101 32383
0 8616 5 1 1 8615
0 8617 7 1 2 31170 8616
0 8618 7 1 2 8614 8617
0 8619 5 1 1 8618
0 8620 7 1 2 33657 32129
0 8621 7 1 2 8619 8620
0 8622 7 1 2 8592 8621
0 8623 7 1 2 8588 8622
0 8624 5 1 1 8623
0 8625 7 1 2 23535 8624
0 8626 7 1 2 8586 8625
0 8627 5 1 1 8626
0 8628 7 1 2 23443 8627
0 8629 7 1 2 8479 8628
0 8630 5 1 1 8629
0 8631 7 1 2 30469 30065
0 8632 5 1 1 8631
0 8633 7 1 2 27508 29289
0 8634 5 3 1 8633
0 8635 7 1 2 24526 33149
0 8636 5 1 1 8635
0 8637 7 1 2 34684 8636
0 8638 5 1 1 8637
0 8639 7 1 2 25165 8638
0 8640 5 1 1 8639
0 8641 7 1 2 28428 31459
0 8642 5 2 1 8641
0 8643 7 1 2 29296 34687
0 8644 5 1 1 8643
0 8645 7 1 2 25166 8644
0 8646 5 1 1 8645
0 8647 7 1 2 29501 32106
0 8648 5 2 1 8647
0 8649 7 1 2 8646 34689
0 8650 5 1 1 8649
0 8651 7 1 2 23100 8650
0 8652 5 1 1 8651
0 8653 7 1 2 29352 31058
0 8654 5 2 1 8653
0 8655 7 1 2 29353 32423
0 8656 5 1 1 8655
0 8657 7 1 2 34691 8656
0 8658 7 1 2 8652 8657
0 8659 7 1 2 8640 8658
0 8660 5 1 1 8659
0 8661 7 1 2 24605 8660
0 8662 5 1 1 8661
0 8663 7 2 2 29060 30274
0 8664 7 1 2 22541 30897
0 8665 5 1 1 8664
0 8666 7 1 2 34693 8665
0 8667 5 1 1 8666
0 8668 7 1 2 34625 8667
0 8669 5 1 1 8668
0 8670 7 1 2 27509 8669
0 8671 5 1 1 8670
0 8672 7 1 2 27267 29451
0 8673 5 2 1 8672
0 8674 7 1 2 30117 34695
0 8675 5 1 1 8674
0 8676 7 1 2 30109 29596
0 8677 5 1 1 8676
0 8678 7 1 2 28554 8677
0 8679 5 1 1 8678
0 8680 7 1 2 8675 8679
0 8681 5 1 1 8680
0 8682 7 1 2 8671 8681
0 8683 5 1 1 8682
0 8684 7 1 2 24077 8683
0 8685 5 1 1 8684
0 8686 7 1 2 28892 31001
0 8687 5 1 1 8686
0 8688 7 4 2 23961 22652
0 8689 7 1 2 23208 34697
0 8690 7 1 2 8687 8689
0 8691 5 3 1 8690
0 8692 7 1 2 8685 34701
0 8693 7 1 2 8662 8692
0 8694 5 1 1 8693
0 8695 7 1 2 23296 8694
0 8696 5 1 1 8695
0 8697 7 1 2 8632 8696
0 8698 5 1 1 8697
0 8699 7 1 2 34068 8698
0 8700 5 1 1 8699
0 8701 7 2 2 25487 34627
0 8702 7 3 2 24078 22259
0 8703 7 1 2 33949 34706
0 8704 7 1 2 34704 8703
0 8705 5 1 1 8704
0 8706 7 1 2 8700 8705
0 8707 5 1 1 8706
0 8708 7 1 2 22393 8707
0 8709 5 1 1 8708
0 8710 7 1 2 24389 33958
0 8711 7 1 2 34707 8710
0 8712 7 1 2 34705 8711
0 8713 5 1 1 8712
0 8714 7 1 2 8709 8713
0 8715 5 1 1 8714
0 8716 7 1 2 23749 8715
0 8717 5 1 1 8716
0 8718 7 1 2 24079 34137
0 8719 7 3 2 29780 30961
0 8720 7 1 2 34709 33112
0 8721 7 1 2 8718 8720
0 8722 7 1 2 32349 8721
0 8723 5 1 1 8722
0 8724 7 1 2 8717 8723
0 8725 5 1 1 8724
0 8726 7 1 2 28807 8725
0 8727 5 1 1 8726
0 8728 7 3 2 26002 33916
0 8729 7 1 2 34712 34628
0 8730 5 1 1 8729
0 8731 7 1 2 27329 31085
0 8732 5 1 1 8731
0 8733 7 1 2 2201 8732
0 8734 5 1 1 8733
0 8735 7 1 2 23209 8734
0 8736 5 1 1 8735
0 8737 7 1 2 26695 31421
0 8738 5 1 1 8737
0 8739 7 1 2 22653 27864
0 8740 5 1 1 8739
0 8741 7 1 2 26696 8740
0 8742 5 1 1 8741
0 8743 7 2 2 29781 30420
0 8744 5 1 1 34715
0 8745 7 1 2 8742 8744
0 8746 5 1 1 8745
0 8747 7 1 2 23101 8746
0 8748 5 1 1 8747
0 8749 7 1 2 8738 8748
0 8750 7 1 2 8736 8749
0 8751 5 1 1 8750
0 8752 7 1 2 26003 8751
0 8753 5 1 1 8752
0 8754 7 1 2 26077 32855
0 8755 5 1 1 8754
0 8756 7 1 2 25965 32829
0 8757 5 1 1 8756
0 8758 7 1 2 8755 8757
0 8759 5 1 1 8758
0 8760 7 1 2 23831 8759
0 8761 5 1 1 8760
0 8762 7 1 2 27304 25984
0 8763 7 1 2 32830 8762
0 8764 5 1 1 8763
0 8765 7 1 2 8761 8764
0 8766 5 2 1 8765
0 8767 7 1 2 28979 34717
0 8768 5 1 1 8767
0 8769 7 1 2 8753 8768
0 8770 5 1 1 8769
0 8771 7 1 2 23962 8770
0 8772 5 1 1 8771
0 8773 7 1 2 28980 34716
0 8774 5 1 1 8773
0 8775 7 1 2 25167 31125
0 8776 5 1 1 8775
0 8777 7 1 2 27342 29087
0 8778 5 1 1 8777
0 8779 7 1 2 22654 8778
0 8780 5 1 1 8779
0 8781 7 1 2 8776 8780
0 8782 5 1 1 8781
0 8783 7 1 2 23009 31104
0 8784 5 1 1 8783
0 8785 7 1 2 26306 8784
0 8786 5 1 1 8785
0 8787 7 1 2 23297 8786
0 8788 7 1 2 8782 8787
0 8789 5 1 1 8788
0 8790 7 1 2 8774 8789
0 8791 5 1 1 8790
0 8792 7 1 2 26004 8791
0 8793 5 1 1 8792
0 8794 7 1 2 8772 8793
0 8795 5 1 1 8794
0 8796 7 1 2 34402 8795
0 8797 5 1 1 8796
0 8798 7 1 2 8730 8797
0 8799 5 1 1 8798
0 8800 7 1 2 24080 8799
0 8801 5 1 1 8800
0 8802 7 1 2 25168 29452
0 8803 7 1 2 27380 8802
0 8804 5 1 1 8803
0 8805 7 1 2 34690 8804
0 8806 5 1 1 8805
0 8807 7 1 2 23102 8806
0 8808 5 1 1 8807
0 8809 7 1 2 23963 31059
0 8810 5 1 1 8809
0 8811 7 1 2 31062 34696
0 8812 5 1 1 8811
0 8813 7 1 2 27138 8812
0 8814 5 1 1 8813
0 8815 7 1 2 8810 8814
0 8816 7 1 2 8808 8815
0 8817 5 1 1 8816
0 8818 7 1 2 24606 8817
0 8819 5 1 1 8818
0 8820 7 1 2 34702 8819
0 8821 5 1 1 8820
0 8822 7 8 2 22260 23536
0 8823 7 1 2 34719 34526
0 8824 7 1 2 26005 8823
0 8825 7 1 2 8821 8824
0 8826 5 1 1 8825
0 8827 7 1 2 8801 8826
0 8828 7 1 2 8727 8827
0 8829 5 1 1 8828
0 8830 7 1 2 34276 8829
0 8831 5 1 1 8830
0 8832 7 1 2 22201 8831
0 8833 7 1 2 8630 8832
0 8834 5 1 1 8833
0 8835 7 3 2 29766 5189
0 8836 5 6 1 34727
0 8837 7 1 2 29128 34728
0 8838 5 1 1 8837
0 8839 7 1 2 27247 8838
0 8840 5 1 1 8839
0 8841 7 1 2 30110 31675
0 8842 5 1 1 8841
0 8843 7 1 2 8840 8842
0 8844 5 1 1 8843
0 8845 7 1 2 31245 8844
0 8846 5 1 1 8845
0 8847 7 2 2 30118 3020
0 8848 5 1 1 34736
0 8849 7 1 2 28597 29910
0 8850 5 1 1 8849
0 8851 7 1 2 34737 8850
0 8852 5 1 1 8851
0 8853 7 1 2 31246 8852
0 8854 5 1 1 8853
0 8855 7 2 2 24476 32953
0 8856 5 1 1 34738
0 8857 7 2 2 29782 34739
0 8858 7 1 2 29061 34740
0 8859 5 1 1 8858
0 8860 7 1 2 8854 8859
0 8861 5 1 1 8860
0 8862 7 1 2 29597 8861
0 8863 5 1 1 8862
0 8864 7 1 2 8846 8863
0 8865 5 1 1 8864
0 8866 7 1 2 23298 33436
0 8867 7 1 2 8865 8866
0 8868 5 1 1 8867
0 8869 7 1 2 32860 34713
0 8870 5 1 1 8869
0 8871 7 1 2 34403 34718
0 8872 5 1 1 8871
0 8873 7 1 2 8870 8872
0 8874 5 1 1 8873
0 8875 7 1 2 23103 8874
0 8876 5 1 1 8875
0 8877 7 1 2 34138 32856
0 8878 5 1 1 8877
0 8879 7 4 2 25924 33596
0 8880 5 1 1 34742
0 8881 7 1 2 34743 32831
0 8882 5 1 1 8881
0 8883 7 1 2 8878 8882
0 8884 5 1 1 8883
0 8885 7 1 2 32273 8884
0 8886 5 1 1 8885
0 8887 7 1 2 7097 8880
0 8888 5 2 1 8887
0 8889 7 1 2 27221 30555
0 8890 5 1 1 8889
0 8891 7 1 2 34746 8890
0 8892 7 1 2 32832 8891
0 8893 5 1 1 8892
0 8894 7 1 2 8886 8893
0 8895 5 1 1 8894
0 8896 7 1 2 28808 8895
0 8897 5 1 1 8896
0 8898 7 2 2 25985 34358
0 8899 7 1 2 27211 32833
0 8900 7 1 2 34748 8899
0 8901 5 1 1 8900
0 8902 7 1 2 8897 8901
0 8903 7 1 2 8876 8902
0 8904 5 1 1 8903
0 8905 7 1 2 29453 8904
0 8906 5 1 1 8905
0 8907 7 1 2 26899 34404
0 8908 5 1 1 8907
0 8909 7 1 2 33917 32331
0 8910 5 1 1 8909
0 8911 7 1 2 8908 8910
0 8912 5 1 1 8911
0 8913 7 1 2 25986 8912
0 8914 5 1 1 8913
0 8915 7 1 2 34744 32332
0 8916 5 1 1 8915
0 8917 7 3 2 24607 34483
0 8918 7 2 2 24276 34750
0 8919 7 1 2 30172 33477
0 8920 7 1 2 34753 8919
0 8921 5 1 1 8920
0 8922 7 1 2 8916 8921
0 8923 5 1 1 8922
0 8924 7 1 2 28809 8923
0 8925 5 1 1 8924
0 8926 7 1 2 8914 8925
0 8927 5 1 1 8926
0 8928 7 2 2 28883 29783
0 8929 7 1 2 23750 34755
0 8930 7 1 2 8927 8929
0 8931 5 1 1 8930
0 8932 7 1 2 8906 8931
0 8933 5 1 1 8932
0 8934 7 1 2 29598 32967
0 8935 7 1 2 8933 8934
0 8936 5 1 1 8935
0 8937 7 1 2 8868 8936
0 8938 5 1 1 8937
0 8939 7 1 2 24081 8938
0 8940 5 1 1 8939
0 8941 7 2 2 30497 33229
0 8942 5 1 1 34757
0 8943 7 7 2 24696 25251
0 8944 7 1 2 34759 32301
0 8945 5 1 1 8944
0 8946 7 1 2 8942 8945
0 8947 5 1 1 8946
0 8948 7 1 2 29502 8947
0 8949 5 1 1 8948
0 8950 7 2 2 25061 31752
0 8951 7 1 2 31344 34766
0 8952 7 1 2 32370 8951
0 8953 5 1 1 8952
0 8954 7 1 2 8949 8953
0 8955 5 1 1 8954
0 8956 7 1 2 27446 8955
0 8957 5 1 1 8956
0 8958 7 4 2 22752 23299
0 8959 7 4 2 29454 34730
0 8960 5 1 1 34772
0 8961 7 1 2 25169 34773
0 8962 5 1 1 8961
0 8963 7 1 2 34692 8962
0 8964 5 1 1 8963
0 8965 7 1 2 24608 8964
0 8966 5 1 1 8965
0 8967 7 1 2 34703 8966
0 8968 5 1 1 8967
0 8969 7 1 2 34768 8968
0 8970 5 1 1 8969
0 8971 7 1 2 8957 8970
0 8972 5 2 1 8971
0 8973 7 1 2 34069 34776
0 8974 5 1 1 8973
0 8975 7 3 2 26875 34635
0 8976 7 3 2 22261 33950
0 8977 7 2 2 31312 34781
0 8978 7 1 2 34778 34784
0 8979 5 1 1 8978
0 8980 7 1 2 8974 8979
0 8981 5 1 1 8980
0 8982 7 1 2 22394 8981
0 8983 5 1 1 8982
0 8984 7 3 2 22923 33302
0 8985 7 1 2 27447 32597
0 8986 7 2 2 34786 8985
0 8987 7 1 2 34779 34789
0 8988 5 1 1 8987
0 8989 7 1 2 8983 8988
0 8990 5 1 1 8989
0 8991 7 1 2 28810 8990
0 8992 5 1 1 8991
0 8993 7 4 2 24277 27448
0 8994 7 3 2 22041 24749
0 8995 7 2 2 34791 34795
0 8996 7 1 2 34780 34798
0 8997 5 1 1 8996
0 8998 7 1 2 33621 34777
0 8999 5 1 1 8998
0 9000 7 1 2 8997 8999
0 9001 5 1 1 9000
0 9002 7 1 2 25987 9001
0 9003 5 1 1 9002
0 9004 7 1 2 8992 9003
0 9005 5 1 1 9004
0 9006 7 1 2 33702 9005
0 9007 5 1 1 9006
0 9008 7 1 2 8940 9007
0 9009 5 1 1 9008
0 9010 7 1 2 25397 9009
0 9011 5 1 1 9010
0 9012 7 3 2 25488 30348
0 9013 7 1 2 34785 34800
0 9014 5 1 1 9013
0 9015 7 1 2 34070 34669
0 9016 5 1 1 9015
0 9017 7 1 2 9014 9016
0 9018 5 1 1 9017
0 9019 7 1 2 22395 9018
0 9020 5 1 1 9019
0 9021 7 1 2 34790 34801
0 9022 5 1 1 9021
0 9023 7 1 2 9020 9022
0 9024 5 1 1 9023
0 9025 7 1 2 25252 9024
0 9026 5 1 1 9025
0 9027 7 1 2 30716 34459
0 9028 5 1 1 9027
0 9029 7 1 2 22542 34745
0 9030 5 1 1 9029
0 9031 7 1 2 9028 9030
0 9032 5 1 1 9031
0 9033 7 1 2 29960 9032
0 9034 5 1 1 9033
0 9035 7 2 2 22543 31411
0 9036 5 1 1 34803
0 9037 7 1 2 31511 34071
0 9038 7 1 2 34804 9037
0 9039 5 1 1 9038
0 9040 7 1 2 9034 9039
0 9041 5 1 1 9040
0 9042 7 1 2 34672 9041
0 9043 5 1 1 9042
0 9044 7 1 2 9026 9043
0 9045 5 1 1 9044
0 9046 7 1 2 28811 9045
0 9047 5 1 1 9046
0 9048 7 1 2 34799 34802
0 9049 5 1 1 9048
0 9050 7 1 2 33622 34670
0 9051 5 1 1 9050
0 9052 7 1 2 9049 9051
0 9053 5 1 1 9052
0 9054 7 1 2 25253 9053
0 9055 5 1 1 9054
0 9056 7 2 2 30717 33303
0 9057 7 1 2 29966 9036
0 9058 5 2 1 9057
0 9059 7 1 2 34805 34807
0 9060 5 1 1 9059
0 9061 7 2 2 22544 27449
0 9062 7 3 2 21920 24278
0 9063 7 2 2 33872 34811
0 9064 5 1 1 34814
0 9065 7 1 2 34809 34815
0 9066 5 1 1 9065
0 9067 7 1 2 9060 9066
0 9068 5 1 1 9067
0 9069 7 1 2 34673 9068
0 9070 5 1 1 9069
0 9071 7 1 2 9055 9070
0 9072 5 1 1 9071
0 9073 7 1 2 25988 9072
0 9074 5 1 1 9073
0 9075 7 1 2 9047 9074
0 9076 5 1 1 9075
0 9077 7 1 2 23751 34280
0 9078 7 1 2 9076 9077
0 9079 5 1 1 9078
0 9080 7 1 2 24212 9079
0 9081 7 1 2 9011 9080
0 9082 5 1 1 9081
0 9083 7 1 2 25589 9082
0 9084 7 1 2 8834 9083
0 9085 5 1 1 9084
0 9086 7 1 2 34405 33099
0 9087 5 1 1 9086
0 9088 7 1 2 34348 32617
0 9089 7 1 2 33095 9088
0 9090 5 1 1 9089
0 9091 7 1 2 9087 9090
0 9092 5 1 1 9091
0 9093 7 1 2 26078 9092
0 9094 5 1 1 9093
0 9095 7 1 2 34359 33101
0 9096 5 1 1 9095
0 9097 7 1 2 9094 9096
0 9098 5 1 1 9097
0 9099 7 1 2 21921 9098
0 9100 5 1 1 9099
0 9101 7 3 2 31822 34360
0 9102 7 1 2 34816 33103
0 9103 5 1 1 9102
0 9104 7 1 2 9100 9103
0 9105 5 1 1 9104
0 9106 7 1 2 34266 9105
0 9107 5 1 1 9106
0 9108 7 4 2 23104 25398
0 9109 7 2 2 23537 34819
0 9110 7 1 2 29784 29455
0 9111 7 1 2 34823 9110
0 9112 7 1 2 34502 9111
0 9113 7 1 2 33059 9112
0 9114 5 1 1 9113
0 9115 7 1 2 9107 9114
0 9116 5 1 1 9115
0 9117 7 1 2 22042 9116
0 9118 5 1 1 9117
0 9119 7 7 2 25399 33009
0 9120 7 2 2 28447 28981
0 9121 7 1 2 34825 34832
0 9122 7 1 2 32693 9121
0 9123 5 1 1 9122
0 9124 7 2 2 25590 30772
0 9125 7 1 2 29961 34267
0 9126 7 1 2 34834 9125
0 9127 5 1 1 9126
0 9128 7 1 2 9123 9127
0 9129 5 1 1 9128
0 9130 7 1 2 23010 9129
0 9131 5 1 1 9130
0 9132 7 2 2 26634 29696
0 9133 7 1 2 31529 34836
0 9134 5 2 1 9133
0 9135 7 2 2 23648 33066
0 9136 7 1 2 22924 34840
0 9137 5 1 1 9136
0 9138 7 1 2 34838 9137
0 9139 5 2 1 9138
0 9140 7 1 2 34268 34842
0 9141 5 1 1 9140
0 9142 7 1 2 9131 9141
0 9143 5 1 1 9142
0 9144 7 1 2 24390 9143
0 9145 5 1 1 9144
0 9146 7 17 2 24213 25400
0 9147 7 2 2 34844 32472
0 9148 5 1 1 34861
0 9149 7 1 2 33795 34862
0 9150 5 1 1 9149
0 9151 7 2 2 23444 33067
0 9152 7 1 2 32779 34863
0 9153 5 1 1 9152
0 9154 7 1 2 9150 9153
0 9155 5 1 1 9154
0 9156 7 1 2 34091 9155
0 9157 5 1 1 9156
0 9158 7 1 2 9145 9157
0 9159 5 1 1 9158
0 9160 7 1 2 22043 9159
0 9161 5 1 1 9160
0 9162 7 5 2 31043 34558
0 9163 7 1 2 3101 30844
0 9164 5 2 1 9163
0 9165 7 1 2 25062 34870
0 9166 5 1 1 9165
0 9167 7 1 2 1283 9166
0 9168 5 4 1 9167
0 9169 7 1 2 32618 34872
0 9170 5 1 1 9169
0 9171 7 1 2 31550 33088
0 9172 5 1 1 9171
0 9173 7 1 2 9170 9172
0 9174 5 2 1 9173
0 9175 7 1 2 34865 34876
0 9176 5 1 1 9175
0 9177 7 1 2 9161 9176
0 9178 5 1 1 9177
0 9179 7 1 2 34139 9178
0 9180 5 1 1 9179
0 9181 7 1 2 34555 33821
0 9182 7 1 2 34548 9181
0 9183 7 1 2 34841 9182
0 9184 5 1 1 9183
0 9185 7 1 2 9180 9184
0 9186 5 1 1 9185
0 9187 7 1 2 28812 9186
0 9188 5 1 1 9187
0 9189 7 1 2 33038 34873
0 9190 5 1 1 9189
0 9191 7 4 2 27212 30198
0 9192 5 1 1 34878
0 9193 7 1 2 34879 33077
0 9194 5 1 1 9193
0 9195 7 1 2 9190 9194
0 9196 5 1 1 9195
0 9197 7 1 2 33623 34866
0 9198 7 1 2 9196 9197
0 9199 5 1 1 9198
0 9200 7 1 2 9188 9199
0 9201 7 1 2 9118 9200
0 9202 5 1 1 9201
0 9203 7 1 2 32968 9202
0 9204 5 1 1 9203
0 9205 7 2 2 33026 34833
0 9206 7 1 2 32694 34882
0 9207 5 1 1 9206
0 9208 7 1 2 25254 31624
0 9209 7 1 2 34835 9208
0 9210 5 1 1 9209
0 9211 7 1 2 9207 9210
0 9212 5 1 1 9211
0 9213 7 1 2 23011 9212
0 9214 5 1 1 9213
0 9215 7 1 2 33172 34843
0 9216 5 1 1 9215
0 9217 7 1 2 9214 9216
0 9218 5 1 1 9217
0 9219 7 1 2 24391 9218
0 9220 5 1 1 9219
0 9221 7 2 2 33173 33068
0 9222 5 1 1 34884
0 9223 7 1 2 23012 34883
0 9224 5 1 1 9223
0 9225 7 1 2 9222 9224
0 9226 5 1 1 9225
0 9227 7 1 2 34092 9226
0 9228 5 1 1 9227
0 9229 7 1 2 9220 9228
0 9230 5 1 1 9229
0 9231 7 1 2 22044 9230
0 9232 5 1 1 9231
0 9233 7 1 2 32931 34877
0 9234 5 1 1 9233
0 9235 7 1 2 9232 9234
0 9236 5 2 1 9235
0 9237 7 1 2 26079 34886
0 9238 5 1 1 9237
0 9239 7 1 2 29894 32210
0 9240 5 1 1 9239
0 9241 7 1 2 6341 9240
0 9242 5 1 1 9241
0 9243 7 1 2 24527 9242
0 9244 5 1 1 9243
0 9245 7 2 2 24082 27305
0 9246 7 1 2 29906 30955
0 9247 7 1 2 34888 9246
0 9248 5 1 1 9247
0 9249 7 1 2 9244 9248
0 9250 5 1 1 9249
0 9251 7 1 2 23832 9250
0 9252 5 1 1 9251
0 9253 7 1 2 32267 34662
0 9254 5 1 1 9253
0 9255 7 1 2 9252 9254
0 9256 5 3 1 9255
0 9257 7 1 2 33027 34890
0 9258 5 1 1 9257
0 9259 7 1 2 22045 34885
0 9260 5 1 1 9259
0 9261 7 1 2 9258 9260
0 9262 5 1 1 9261
0 9263 7 1 2 27701 9262
0 9264 5 1 1 9263
0 9265 7 1 2 9238 9264
0 9266 5 1 1 9265
0 9267 7 1 2 34406 9266
0 9268 5 1 1 9267
0 9269 7 5 2 22202 33351
0 9270 7 1 2 34893 32388
0 9271 7 1 2 31823 9270
0 9272 7 1 2 34891 9271
0 9273 5 1 1 9272
0 9274 7 1 2 9268 9273
0 9275 5 1 1 9274
0 9276 7 1 2 34289 9275
0 9277 5 1 1 9276
0 9278 7 1 2 34140 34887
0 9279 5 1 1 9278
0 9280 7 2 2 26113 33897
0 9281 7 10 2 22203 22262
0 9282 7 1 2 31857 34900
0 9283 7 1 2 34898 9282
0 9284 7 1 2 34892 9283
0 9285 5 1 1 9284
0 9286 7 1 2 9279 9285
0 9287 5 1 1 9286
0 9288 7 1 2 34290 9287
0 9289 5 1 1 9288
0 9290 7 1 2 34760 33134
0 9291 5 1 1 9290
0 9292 7 4 2 23833 29456
0 9293 7 1 2 29895 34769
0 9294 7 1 2 34910 9293
0 9295 5 1 1 9294
0 9296 7 1 2 9291 9295
0 9297 5 1 1 9296
0 9298 7 1 2 22046 9297
0 9299 5 1 1 9298
0 9300 7 1 2 23300 32904
0 9301 7 1 2 34874 9300
0 9302 5 1 1 9301
0 9303 7 1 2 9299 9302
0 9304 5 1 1 9303
0 9305 7 1 2 23368 9304
0 9306 5 1 1 9305
0 9307 7 1 2 25335 29664
0 9308 7 1 2 32896 9307
0 9309 7 1 2 33080 9308
0 9310 5 1 1 9309
0 9311 7 1 2 9306 9310
0 9312 5 1 1 9311
0 9313 7 1 2 25401 9312
0 9314 5 1 1 9313
0 9315 7 4 2 22047 25336
0 9316 7 1 2 31285 34914
0 9317 7 1 2 34864 9316
0 9318 5 1 1 9317
0 9319 7 1 2 9314 9318
0 9320 5 2 1 9319
0 9321 7 1 2 23649 34375
0 9322 7 1 2 34899 9321
0 9323 7 1 2 34918 9322
0 9324 5 1 1 9323
0 9325 7 1 2 9289 9324
0 9326 5 1 1 9325
0 9327 7 1 2 28813 9326
0 9328 5 1 1 9327
0 9329 7 2 2 28576 32725
0 9330 5 1 1 34920
0 9331 7 1 2 34188 34921
0 9332 5 1 1 9331
0 9333 7 23 2 23538 33733
0 9334 5 1 1 34922
0 9335 7 1 2 27381 34923
0 9336 5 1 1 9335
0 9337 7 1 2 9332 9336
0 9338 5 1 1 9337
0 9339 7 1 2 23964 9338
0 9340 5 1 1 9339
0 9341 7 1 2 27213 34924
0 9342 5 1 1 9341
0 9343 7 1 2 9340 9342
0 9344 5 1 1 9343
0 9345 7 1 2 25591 9344
0 9346 5 1 1 9345
0 9347 7 7 2 25854 34407
0 9348 7 1 2 34945 33016
0 9349 5 1 1 9348
0 9350 7 1 2 9346 9349
0 9351 5 1 1 9350
0 9352 7 1 2 26114 9351
0 9353 5 1 1 9352
0 9354 7 3 2 23650 26130
0 9355 7 1 2 32509 34952
0 9356 7 1 2 34925 9355
0 9357 5 1 1 9356
0 9358 7 1 2 9353 9357
0 9359 5 1 1 9358
0 9360 7 1 2 26221 34867
0 9361 7 1 2 9359 9360
0 9362 5 1 1 9361
0 9363 7 2 2 31345 30834
0 9364 7 1 2 27030 33003
0 9365 7 1 2 34955 9364
0 9366 7 1 2 34926 9365
0 9367 5 1 1 9366
0 9368 7 1 2 9362 9367
0 9369 5 1 1 9368
0 9370 7 1 2 32969 9369
0 9371 5 1 1 9370
0 9372 7 2 2 33676 32941
0 9373 7 1 2 32939 34957
0 9374 5 1 1 9373
0 9375 7 1 2 31813 32029
0 9376 5 1 1 9375
0 9377 7 1 2 6272 9376
0 9378 5 1 1 9377
0 9379 7 1 2 23539 33722
0 9380 5 1 1 9379
0 9381 7 1 2 33674 9380
0 9382 5 1 1 9381
0 9383 7 1 2 9378 9382
0 9384 5 1 1 9383
0 9385 7 1 2 28471 31814
0 9386 5 1 1 9385
0 9387 7 1 2 32268 32932
0 9388 5 1 1 9387
0 9389 7 1 2 9386 9388
0 9390 5 1 1 9389
0 9391 7 1 2 21816 9390
0 9392 5 1 1 9391
0 9393 7 1 2 32901 32933
0 9394 5 1 1 9393
0 9395 7 1 2 9392 9394
0 9396 5 1 1 9395
0 9397 7 1 2 29032 33352
0 9398 7 1 2 9396 9397
0 9399 5 1 1 9398
0 9400 7 1 2 9384 9399
0 9401 5 1 1 9400
0 9402 7 1 2 25592 9401
0 9403 5 1 1 9402
0 9404 7 1 2 31293 32942
0 9405 7 1 2 33691 9404
0 9406 5 1 1 9405
0 9407 7 1 2 9403 9406
0 9408 5 1 1 9407
0 9409 7 1 2 24860 9408
0 9410 5 1 1 9409
0 9411 7 1 2 9374 9410
0 9412 5 1 1 9411
0 9413 7 1 2 24392 9412
0 9414 5 1 1 9413
0 9415 7 1 2 32947 34958
0 9416 5 1 1 9415
0 9417 7 1 2 9414 9416
0 9418 5 1 1 9417
0 9419 7 1 2 34291 9418
0 9420 5 1 1 9419
0 9421 7 1 2 24951 23369
0 9422 7 1 2 34956 9421
0 9423 5 1 1 9422
0 9424 7 1 2 24083 34613
0 9425 5 1 1 9424
0 9426 7 1 2 9423 9425
0 9427 5 1 1 9426
0 9428 7 1 2 24697 9427
0 9429 5 1 1 9428
0 9430 7 1 2 27930 32905
0 9431 7 1 2 32510 9430
0 9432 5 1 1 9431
0 9433 7 1 2 9429 9432
0 9434 5 1 1 9433
0 9435 7 1 2 34845 34221
0 9436 7 1 2 9434 9435
0 9437 5 1 1 9436
0 9438 7 4 2 24698 24750
0 9439 7 1 2 25771 30756
0 9440 7 1 2 34959 9439
0 9441 7 2 2 34175 32133
0 9442 7 1 2 34963 34230
0 9443 7 1 2 9440 9442
0 9444 7 1 2 31838 9443
0 9445 5 1 1 9444
0 9446 7 1 2 9437 9445
0 9447 5 1 1 9446
0 9448 7 1 2 25489 9447
0 9449 5 1 1 9448
0 9450 7 1 2 9420 9449
0 9451 7 1 2 9371 9450
0 9452 5 1 1 9451
0 9453 7 1 2 32582 9452
0 9454 5 1 1 9453
0 9455 7 1 2 24214 33039
0 9456 7 1 2 34919 9455
0 9457 5 1 1 9456
0 9458 7 1 2 29760 31688
0 9459 7 1 2 30939 33938
0 9460 7 1 2 9458 9459
0 9461 7 1 2 26141 9460
0 9462 7 1 2 31839 9461
0 9463 5 1 1 9462
0 9464 7 1 2 9457 9463
0 9465 5 1 1 9464
0 9466 7 1 2 33918 9465
0 9467 5 1 1 9466
0 9468 7 1 2 25670 9467
0 9469 7 1 2 9454 9468
0 9470 7 1 2 9328 9469
0 9471 7 1 2 9277 9470
0 9472 7 1 2 9204 9471
0 9473 5 1 1 9472
0 9474 7 3 2 24084 27554
0 9475 5 1 1 34965
0 9476 7 1 2 30275 34966
0 9477 5 1 1 9476
0 9478 7 2 2 27139 29599
0 9479 7 1 2 26425 34968
0 9480 5 1 1 9479
0 9481 7 1 2 9477 9480
0 9482 5 1 1 9481
0 9483 7 1 2 23105 9482
0 9484 5 1 1 9483
0 9485 7 3 2 24085 22396
0 9486 7 2 2 26407 34970
0 9487 5 1 1 34973
0 9488 7 1 2 23965 34974
0 9489 5 1 1 9488
0 9490 7 3 2 23966 26154
0 9491 7 2 2 23834 27555
0 9492 5 1 1 34978
0 9493 7 1 2 34975 34979
0 9494 5 1 1 9493
0 9495 7 1 2 9487 9494
0 9496 5 1 1 9495
0 9497 7 1 2 29114 9496
0 9498 5 1 1 9497
0 9499 7 1 2 9489 9498
0 9500 7 1 2 9484 9499
0 9501 5 1 1 9500
0 9502 7 1 2 33523 9501
0 9503 5 1 1 9502
0 9504 7 1 2 30276 31439
0 9505 5 1 1 9504
0 9506 7 1 2 29123 29743
0 9507 5 1 1 9506
0 9508 7 1 2 9505 9507
0 9509 5 1 1 9508
0 9510 7 1 2 25975 33708
0 9511 7 1 2 9509 9510
0 9512 5 1 1 9511
0 9513 7 1 2 9503 9512
0 9514 5 1 1 9513
0 9515 7 1 2 25490 9514
0 9516 5 1 1 9515
0 9517 7 1 2 22048 29129
0 9518 5 3 1 9517
0 9519 7 1 2 26243 34980
0 9520 5 1 1 9519
0 9521 7 1 2 30440 34967
0 9522 5 1 1 9521
0 9523 7 1 2 9520 9522
0 9524 5 1 1 9523
0 9525 7 1 2 33597 9524
0 9526 5 1 1 9525
0 9527 7 2 2 30890 34460
0 9528 7 2 2 23106 28674
0 9529 7 1 2 34983 34985
0 9530 5 1 1 9529
0 9531 7 1 2 9526 9530
0 9532 5 1 1 9531
0 9533 7 1 2 28814 9532
0 9534 5 1 1 9533
0 9535 7 2 2 26941 33353
0 9536 7 1 2 34987 34981
0 9537 5 1 1 9536
0 9538 7 1 2 31641 33624
0 9539 5 1 1 9538
0 9540 7 1 2 9537 9539
0 9541 5 1 1 9540
0 9542 7 1 2 28108 9541
0 9543 5 1 1 9542
0 9544 7 2 2 30962 33304
0 9545 7 1 2 29725 34989
0 9546 5 1 1 9545
0 9547 7 1 2 7423 9546
0 9548 5 1 1 9547
0 9549 7 1 2 30441 9548
0 9550 7 1 2 28122 9549
0 9551 5 1 1 9550
0 9552 7 1 2 9543 9551
0 9553 7 1 2 9534 9552
0 9554 5 1 1 9553
0 9555 7 1 2 27510 9554
0 9556 5 1 1 9555
0 9557 7 3 2 22925 33644
0 9558 5 3 1 34991
0 9559 7 1 2 31440 34992
0 9560 5 1 1 9559
0 9561 7 1 2 32205 33546
0 9562 5 1 1 9561
0 9563 7 1 2 29178 33645
0 9564 5 1 1 9563
0 9565 7 1 2 9562 9564
0 9566 5 2 1 9565
0 9567 7 2 2 23967 30573
0 9568 5 1 1 34999
0 9569 7 1 2 9568 6118
0 9570 5 1 1 9569
0 9571 7 1 2 34997 9570
0 9572 5 1 1 9571
0 9573 7 1 2 9560 9572
0 9574 7 1 2 9556 9573
0 9575 7 1 2 9516 9574
0 9576 5 1 1 9575
0 9577 7 1 2 26850 9576
0 9578 5 1 1 9577
0 9579 7 2 2 25491 32998
0 9580 7 1 2 33547 35001
0 9581 5 1 1 9580
0 9582 7 1 2 25063 34993
0 9583 5 1 1 9582
0 9584 7 1 2 9581 9583
0 9585 5 1 1 9584
0 9586 7 1 2 27178 9585
0 9587 5 1 1 9586
0 9588 7 5 2 22926 25064
0 9589 7 5 2 23651 33524
0 9590 7 3 2 25492 35008
0 9591 7 2 2 35003 35013
0 9592 7 1 2 32149 35016
0 9593 5 1 1 9592
0 9594 7 1 2 9587 9593
0 9595 5 1 1 9594
0 9596 7 1 2 24952 9595
0 9597 5 2 1 9596
0 9598 7 1 2 27680 33642
0 9599 5 1 1 9598
0 9600 7 1 2 33421 9599
0 9601 5 1 1 9600
0 9602 7 1 2 28675 9601
0 9603 5 1 1 9602
0 9604 7 2 2 22318 33354
0 9605 5 1 1 35020
0 9606 7 1 2 7170 9605
0 9607 5 6 1 9606
0 9608 7 1 2 28694 35022
0 9609 5 1 1 9608
0 9610 7 1 2 28707 34440
0 9611 5 1 1 9610
0 9612 7 1 2 24809 28642
0 9613 7 1 2 33408 9612
0 9614 5 1 1 9613
0 9615 7 1 2 9611 9614
0 9616 7 1 2 9609 9615
0 9617 5 1 1 9616
0 9618 7 1 2 26204 9617
0 9619 5 1 1 9618
0 9620 7 1 2 9603 9619
0 9621 5 1 1 9620
0 9622 7 1 2 31496 9621
0 9623 5 1 1 9622
0 9624 7 1 2 35018 9623
0 9625 5 1 1 9624
0 9626 7 1 2 29503 9625
0 9627 5 1 1 9626
0 9628 7 3 2 30301 31356
0 9629 7 1 2 35028 33548
0 9630 5 1 1 9629
0 9631 7 4 2 22478 25593
0 9632 5 1 1 35031
0 9633 7 1 2 26222 9632
0 9634 5 1 1 9633
0 9635 7 1 2 21817 9634
0 9636 7 1 2 26364 9635
0 9637 5 1 1 9636
0 9638 7 1 2 32138 9637
0 9639 5 2 1 9638
0 9640 7 1 2 33525 35035
0 9641 5 1 1 9640
0 9642 7 5 2 21818 25594
0 9643 7 2 2 34200 35037
0 9644 7 1 2 30648 34046
0 9645 7 1 2 35042 9644
0 9646 5 1 1 9645
0 9647 7 1 2 9641 9646
0 9648 5 1 1 9647
0 9649 7 1 2 25493 9648
0 9650 5 1 1 9649
0 9651 7 1 2 34994 9650
0 9652 5 1 1 9651
0 9653 7 1 2 31190 9652
0 9654 5 1 1 9653
0 9655 7 1 2 30838 35002
0 9656 7 1 2 34640 9655
0 9657 5 1 1 9656
0 9658 7 1 2 9654 9657
0 9659 5 1 1 9658
0 9660 7 1 2 25065 9659
0 9661 5 1 1 9660
0 9662 7 1 2 9630 9661
0 9663 7 1 2 9627 9662
0 9664 5 1 1 9663
0 9665 7 1 2 30974 9664
0 9666 5 1 1 9665
0 9667 7 1 2 9578 9666
0 9668 5 1 1 9667
0 9669 7 1 2 28534 9668
0 9670 5 1 1 9669
0 9671 7 1 2 29785 33562
0 9672 5 1 1 9671
0 9673 7 1 2 33305 33550
0 9674 5 1 1 9673
0 9675 7 1 2 9672 9674
0 9676 5 1 1 9675
0 9677 7 1 2 31460 9676
0 9678 5 1 1 9677
0 9679 7 1 2 22479 32276
0 9680 5 1 1 9679
0 9681 7 1 2 23013 29124
0 9682 7 1 2 9680 9681
0 9683 5 1 1 9682
0 9684 7 1 2 31448 9683
0 9685 5 1 1 9684
0 9686 7 1 2 33563 9685
0 9687 5 1 1 9686
0 9688 7 1 2 9678 9687
0 9689 5 1 1 9688
0 9690 7 1 2 23652 9689
0 9691 5 1 1 9690
0 9692 7 1 2 34468 33210
0 9693 5 1 1 9692
0 9694 7 1 2 9691 9693
0 9695 5 1 1 9694
0 9696 7 1 2 26205 9695
0 9697 5 1 1 9696
0 9698 7 1 2 27306 34998
0 9699 5 1 1 9698
0 9700 7 1 2 28884 32864
0 9701 7 1 2 35014 9700
0 9702 5 1 1 9701
0 9703 7 1 2 9699 9702
0 9704 5 1 1 9703
0 9705 7 1 2 29600 9704
0 9706 5 1 1 9705
0 9707 7 2 2 29264 32865
0 9708 5 1 1 35044
0 9709 7 1 2 34946 35045
0 9710 5 2 1 9709
0 9711 7 3 2 24086 25494
0 9712 7 1 2 26430 9492
0 9713 5 2 1 9712
0 9714 7 1 2 33526 35051
0 9715 5 1 1 9714
0 9716 7 2 2 23835 24279
0 9717 7 1 2 34484 35053
0 9718 7 1 2 28101 9717
0 9719 5 1 1 9718
0 9720 7 1 2 9715 9719
0 9721 5 1 1 9720
0 9722 7 1 2 35048 9721
0 9723 5 1 1 9722
0 9724 7 1 2 35046 9723
0 9725 5 1 1 9724
0 9726 7 1 2 33260 9725
0 9727 5 1 1 9726
0 9728 7 1 2 30302 33538
0 9729 7 1 2 33211 9728
0 9730 5 1 1 9729
0 9731 7 1 2 9727 9730
0 9732 7 1 2 9706 9731
0 9733 7 1 2 9697 9732
0 9734 5 1 1 9733
0 9735 7 1 2 26018 9734
0 9736 5 1 1 9735
0 9737 7 3 2 22049 22397
0 9738 7 1 2 35055 35017
0 9739 5 1 1 9738
0 9740 7 1 2 35019 9739
0 9741 5 1 1 9740
0 9742 7 1 2 29504 9741
0 9743 5 1 1 9742
0 9744 7 1 2 25855 35036
0 9745 5 1 1 9744
0 9746 7 3 2 26206 27901
0 9747 7 1 2 27450 35058
0 9748 5 1 1 9747
0 9749 7 1 2 9745 9748
0 9750 5 1 1 9749
0 9751 7 1 2 33919 9750
0 9752 5 1 1 9751
0 9753 7 1 2 34995 9752
0 9754 5 1 1 9753
0 9755 7 1 2 31191 9754
0 9756 5 1 1 9755
0 9757 7 2 2 21922 34361
0 9758 5 1 1 35061
0 9759 7 1 2 29626 33920
0 9760 5 1 1 9759
0 9761 7 1 2 9758 9760
0 9762 5 1 1 9761
0 9763 7 1 2 31772 9762
0 9764 5 1 1 9763
0 9765 7 1 2 9756 9764
0 9766 5 1 1 9765
0 9767 7 1 2 25066 9766
0 9768 5 1 1 9767
0 9769 7 1 2 29403 33052
0 9770 5 1 1 9769
0 9771 7 1 2 21923 9770
0 9772 5 1 1 9771
0 9773 7 1 2 27343 31497
0 9774 5 1 1 9773
0 9775 7 1 2 9772 9774
0 9776 5 1 1 9775
0 9777 7 1 2 27556 9776
0 9778 5 1 1 9777
0 9779 7 4 2 25067 31192
0 9780 7 1 2 26339 29756
0 9781 7 1 2 35063 9780
0 9782 5 1 1 9781
0 9783 7 1 2 9778 9782
0 9784 5 1 1 9783
0 9785 7 1 2 33598 9784
0 9786 5 1 1 9785
0 9787 7 1 2 30592 31346
0 9788 7 1 2 34461 9787
0 9789 5 1 1 9788
0 9790 7 1 2 9786 9789
0 9791 5 1 1 9790
0 9792 7 1 2 28815 9791
0 9793 5 1 1 9792
0 9794 7 4 2 25595 34531
0 9795 7 1 2 29566 34335
0 9796 7 1 2 35067 9795
0 9797 5 1 1 9796
0 9798 7 1 2 9793 9797
0 9799 7 1 2 9768 9798
0 9800 7 1 2 9743 9799
0 9801 5 1 1 9800
0 9802 7 1 2 25804 9801
0 9803 5 1 1 9802
0 9804 7 1 2 9736 9803
0 9805 5 1 1 9804
0 9806 7 1 2 28346 9805
0 9807 5 1 1 9806
0 9808 7 1 2 24087 32741
0 9809 5 1 1 9808
0 9810 7 1 2 29088 9809
0 9811 5 1 1 9810
0 9812 7 1 2 28191 7483
0 9813 7 1 2 9811 9812
0 9814 5 1 1 9813
0 9815 7 1 2 28187 31482
0 9816 5 1 1 9815
0 9817 7 1 2 31637 31477
0 9818 5 1 1 9817
0 9819 7 1 2 9816 9818
0 9820 5 1 1 9819
0 9821 7 1 2 23014 9820
0 9822 5 1 1 9821
0 9823 7 2 2 28174 34559
0 9824 5 1 1 35071
0 9825 7 11 2 23445 26768
0 9826 5 1 1 35073
0 9827 7 1 2 28885 35074
0 9828 5 1 1 9827
0 9829 7 1 2 9824 9828
0 9830 5 1 1 9829
0 9831 7 1 2 21819 30898
0 9832 5 1 1 9831
0 9833 7 1 2 29601 9832
0 9834 7 1 2 9830 9833
0 9835 5 1 1 9834
0 9836 7 1 2 1773 29942
0 9837 7 1 2 35072 9836
0 9838 5 1 1 9837
0 9839 7 1 2 9835 9838
0 9840 7 1 2 9822 9839
0 9841 7 1 2 9814 9840
0 9842 5 1 1 9841
0 9843 7 1 2 26019 9842
0 9844 5 1 1 9843
0 9845 7 1 2 28188 31269
0 9846 5 1 1 9845
0 9847 7 1 2 29089 35075
0 9848 5 1 1 9847
0 9849 7 1 2 9846 9848
0 9850 5 1 1 9849
0 9851 7 1 2 21924 9850
0 9852 5 1 1 9851
0 9853 7 6 2 25402 25750
0 9854 7 1 2 35084 33116
0 9855 5 1 1 9854
0 9856 7 1 2 25068 35076
0 9857 5 1 1 9856
0 9858 7 1 2 9855 9857
0 9859 5 1 1 9858
0 9860 7 1 2 22050 9859
0 9861 5 1 1 9860
0 9862 7 1 2 9852 9861
0 9863 5 1 1 9862
0 9864 7 1 2 27179 9863
0 9865 5 1 1 9864
0 9866 7 2 2 31626 31880
0 9867 5 1 1 35090
0 9868 7 3 2 21820 31158
0 9869 7 2 2 34846 35092
0 9870 5 1 1 35095
0 9871 7 1 2 9867 9870
0 9872 5 1 1 9871
0 9873 7 1 2 31193 9872
0 9874 5 1 1 9873
0 9875 7 1 2 27367 29505
0 9876 5 2 1 9875
0 9877 7 1 2 3989 35097
0 9878 5 1 1 9877
0 9879 7 1 2 35077 9878
0 9880 5 1 1 9879
0 9881 7 1 2 9874 9880
0 9882 5 1 1 9881
0 9883 7 1 2 25069 9882
0 9884 5 1 1 9883
0 9885 7 1 2 25403 31753
0 9886 7 1 2 31748 9885
0 9887 5 1 1 9886
0 9888 7 1 2 9884 9887
0 9889 7 1 2 9865 9888
0 9890 5 1 1 9889
0 9891 7 1 2 25805 9890
0 9892 5 1 1 9891
0 9893 7 1 2 9844 9892
0 9894 5 1 1 9893
0 9895 7 1 2 34619 9894
0 9896 5 1 1 9895
0 9897 7 1 2 23752 9896
0 9898 7 1 2 9807 9897
0 9899 7 1 2 9670 9898
0 9900 5 1 1 9899
0 9901 7 1 2 30145 9900
0 9902 7 1 2 9473 9901
0 9903 5 1 1 9902
0 9904 7 3 2 24215 31428
0 9905 7 1 2 31119 35099
0 9906 5 1 1 9905
0 9907 7 5 2 23836 29290
0 9908 7 1 2 22204 24528
0 9909 7 1 2 28886 9908
0 9910 7 1 2 35102 9909
0 9911 5 1 1 9910
0 9912 7 1 2 9906 9911
0 9913 5 1 1 9912
0 9914 7 1 2 34292 9913
0 9915 5 1 1 9914
0 9916 7 1 2 31120 32164
0 9917 7 1 2 33110 9916
0 9918 5 1 1 9917
0 9919 7 7 2 24529 22753
0 9920 7 2 2 31441 35107
0 9921 7 2 2 24216 26574
0 9922 7 1 2 31378 35116
0 9923 7 1 2 35114 9922
0 9924 5 1 1 9923
0 9925 7 1 2 9918 9924
0 9926 7 1 2 9915 9925
0 9927 5 1 1 9926
0 9928 7 1 2 26697 9927
0 9929 5 1 1 9928
0 9930 7 2 2 23446 33203
0 9931 5 1 1 35118
0 9932 7 4 2 31142 31848
0 9933 7 2 2 30173 35120
0 9934 7 1 2 35119 35124
0 9935 5 1 1 9934
0 9936 7 1 2 9929 9935
0 9937 5 1 1 9936
0 9938 7 1 2 34362 32089
0 9939 5 1 1 9938
0 9940 7 1 2 34087 9939
0 9941 5 2 1 9940
0 9942 7 1 2 9937 35126
0 9943 5 1 1 9942
0 9944 7 4 2 22801 34376
0 9945 7 3 2 24699 35128
0 9946 5 1 1 35132
0 9947 7 1 2 32090 35133
0 9948 5 1 1 9947
0 9949 7 1 2 25751 33397
0 9950 5 1 1 9949
0 9951 7 1 2 9948 9950
0 9952 5 1 1 9951
0 9953 7 1 2 23370 35125
0 9954 5 1 1 9953
0 9955 7 1 2 26020 29069
0 9956 7 1 2 29669 9955
0 9957 5 1 1 9956
0 9958 7 1 2 9954 9957
0 9959 5 1 1 9958
0 9960 7 1 2 26796 9959
0 9961 7 1 2 9952 9960
0 9962 5 1 1 9961
0 9963 7 1 2 9943 9962
0 9964 5 1 1 9963
0 9965 7 1 2 24953 9964
0 9966 5 1 1 9965
0 9967 7 7 2 28982 29291
0 9968 7 3 2 32954 34847
0 9969 7 2 2 23837 30421
0 9970 5 1 1 35145
0 9971 7 1 2 32435 9970
0 9972 5 2 1 9971
0 9973 7 1 2 34408 35147
0 9974 5 1 1 9973
0 9975 7 2 2 27140 33921
0 9976 7 1 2 32432 35149
0 9977 5 1 1 9976
0 9978 7 1 2 9974 9977
0 9979 5 1 1 9978
0 9980 7 1 2 32091 9979
0 9981 5 1 1 9980
0 9982 7 1 2 34072 35146
0 9983 5 1 1 9982
0 9984 7 1 2 27180 34076
0 9985 5 1 1 9984
0 9986 7 1 2 34079 9985
0 9987 7 1 2 32433 9986
0 9988 5 1 1 9987
0 9989 7 1 2 9983 9988
0 9990 5 1 1 9989
0 9991 7 1 2 28816 9990
0 9992 5 1 1 9991
0 9993 7 1 2 9981 9992
0 9994 5 1 1 9993
0 9995 7 1 2 35142 9994
0 9996 5 1 1 9995
0 9997 7 1 2 22205 34293
0 9998 5 2 1 9997
0 9999 7 1 2 22754 35117
0 10000 5 1 1 9999
0 10001 7 1 2 35151 10000
0 10002 5 5 1 10001
0 10003 7 1 2 35153 35127
0 10004 7 1 2 35148 10003
0 10005 5 1 1 10004
0 10006 7 1 2 9996 10005
0 10007 5 1 1 10006
0 10008 7 1 2 35135 10007
0 10009 5 1 1 10008
0 10010 7 1 2 9966 10009
0 10011 5 1 1 10010
0 10012 7 1 2 27548 10011
0 10013 5 1 1 10012
0 10014 7 1 2 22862 32175
0 10015 7 2 2 33683 10014
0 10016 5 1 1 35158
0 10017 7 1 2 30691 33306
0 10018 5 1 1 10017
0 10019 7 1 2 10016 10018
0 10020 5 2 1 10019
0 10021 7 1 2 30613 35160
0 10022 5 1 1 10021
0 10023 7 1 2 30791 30810
0 10024 7 1 2 33527 10023
0 10025 5 1 1 10024
0 10026 7 1 2 10022 10025
0 10027 5 1 1 10026
0 10028 7 1 2 25255 10027
0 10029 5 1 1 10028
0 10030 7 1 2 29860 30883
0 10031 7 1 2 33564 10030
0 10032 5 1 1 10031
0 10033 7 1 2 10029 10032
0 10034 5 1 1 10033
0 10035 7 1 2 22051 10034
0 10036 5 1 1 10035
0 10037 7 1 2 25256 27451
0 10038 7 1 2 33409 10037
0 10039 7 1 2 32198 10038
0 10040 5 1 1 10039
0 10041 7 1 2 10036 10040
0 10042 5 1 1 10041
0 10043 7 1 2 29506 10042
0 10044 5 1 1 10043
0 10045 7 4 2 27452 31194
0 10046 5 1 1 35162
0 10047 7 2 2 30614 35163
0 10048 5 1 1 35166
0 10049 7 1 2 26969 31357
0 10050 5 1 1 10049
0 10051 7 1 2 10048 10050
0 10052 5 1 1 10051
0 10053 7 1 2 25257 10052
0 10054 5 1 1 10053
0 10055 7 1 2 31565 31705
0 10056 5 1 1 10055
0 10057 7 1 2 10054 10056
0 10058 5 1 1 10057
0 10059 7 1 2 35161 10058
0 10060 5 1 1 10059
0 10061 7 1 2 31347 33761
0 10062 7 1 2 33575 10061
0 10063 5 1 1 10062
0 10064 7 1 2 10060 10063
0 10065 7 1 2 10044 10064
0 10066 5 1 1 10065
0 10067 7 1 2 27822 10066
0 10068 5 2 1 10067
0 10069 7 1 2 28068 29542
0 10070 7 2 2 30581 10069
0 10071 7 1 2 33681 35170
0 10072 5 1 1 10071
0 10073 7 1 2 35168 10072
0 10074 5 1 1 10073
0 10075 7 1 2 31627 10074
0 10076 5 1 1 10075
0 10077 7 1 2 31580 31461
0 10078 5 1 1 10077
0 10079 7 1 2 34681 10078
0 10080 5 1 1 10079
0 10081 7 1 2 29214 10080
0 10082 5 1 1 10081
0 10083 7 1 2 28577 34677
0 10084 5 1 1 10083
0 10085 7 1 2 10082 10084
0 10086 5 1 1 10085
0 10087 7 1 2 23301 10086
0 10088 5 1 1 10087
0 10089 7 1 2 31642 32404
0 10090 5 1 1 10089
0 10091 7 1 2 29457 32401
0 10092 5 1 1 10091
0 10093 7 1 2 10090 10092
0 10094 5 1 1 10093
0 10095 7 1 2 30470 10094
0 10096 5 1 1 10095
0 10097 7 1 2 10088 10096
0 10098 5 1 1 10097
0 10099 7 1 2 22319 10098
0 10100 5 1 1 10099
0 10101 7 1 2 22863 26942
0 10102 7 1 2 29136 10101
0 10103 7 2 2 32333 10102
0 10104 7 1 2 34056 35172
0 10105 5 1 1 10104
0 10106 7 1 2 10100 10105
0 10107 5 1 1 10106
0 10108 7 1 2 33307 10107
0 10109 5 1 1 10108
0 10110 7 2 2 24088 22320
0 10111 7 1 2 33355 35174
0 10112 7 1 2 35173 10111
0 10113 5 1 1 10112
0 10114 7 1 2 10109 10113
0 10115 5 1 1 10114
0 10116 7 1 2 27823 10115
0 10117 5 2 1 10116
0 10118 7 2 2 35136 32824
0 10119 7 1 2 34927 35178
0 10120 5 1 1 10119
0 10121 7 1 2 35176 10120
0 10122 5 1 1 10121
0 10123 7 1 2 27511 10122
0 10124 5 1 1 10123
0 10125 7 2 2 22321 33651
0 10126 7 1 2 34720 35180
0 10127 7 2 2 32022 10126
0 10128 5 1 1 35182
0 10129 7 1 2 33528 32807
0 10130 5 1 1 10129
0 10131 7 1 2 10128 10130
0 10132 5 1 1 10131
0 10133 7 1 2 30024 10132
0 10134 5 1 1 10133
0 10135 7 1 2 31594 34947
0 10136 5 1 1 10135
0 10137 7 1 2 10134 10136
0 10138 5 1 1 10137
0 10139 7 1 2 23302 10138
0 10140 5 1 1 10139
0 10141 7 2 2 22864 29458
0 10142 7 2 2 24609 22802
0 10143 7 1 2 33401 35186
0 10144 7 1 2 34388 10143
0 10145 7 1 2 35184 10144
0 10146 7 1 2 30452 10145
0 10147 5 1 1 10146
0 10148 7 1 2 10140 10147
0 10149 5 1 1 10148
0 10150 7 1 2 27824 10149
0 10151 5 2 1 10150
0 10152 7 3 2 23753 32817
0 10153 7 1 2 24810 5979
0 10154 5 1 1 10153
0 10155 7 2 2 7190 32805
0 10156 5 1 1 35193
0 10157 7 1 2 22865 10156
0 10158 5 1 1 10157
0 10159 7 1 2 22322 10158
0 10160 7 1 2 10154 10159
0 10161 5 1 1 10160
0 10162 7 1 2 28708 32810
0 10163 5 1 1 10162
0 10164 7 1 2 10161 10163
0 10165 5 1 1 10164
0 10166 7 1 2 33308 10165
0 10167 5 1 1 10166
0 10168 7 1 2 22866 33557
0 10169 7 1 2 32811 10168
0 10170 5 1 1 10169
0 10171 7 1 2 10167 10170
0 10172 5 1 1 10171
0 10173 7 1 2 35190 10172
0 10174 5 1 1 10173
0 10175 7 3 2 25856 32835
0 10176 7 1 2 30574 35195
0 10177 5 1 1 10176
0 10178 7 1 2 29241 32358
0 10179 7 1 2 32355 10178
0 10180 5 1 1 10179
0 10181 7 1 2 10177 10180
0 10182 5 1 1 10181
0 10183 7 1 2 34409 10182
0 10184 5 1 1 10183
0 10185 7 1 2 31583 33687
0 10186 7 1 2 32836 10185
0 10187 5 1 1 10186
0 10188 7 1 2 10184 10187
0 10189 5 1 1 10188
0 10190 7 1 2 23968 10189
0 10191 5 1 1 10190
0 10192 7 2 2 34341 32334
0 10193 7 2 2 34787 35198
0 10194 5 1 1 35200
0 10195 7 1 2 31589 35201
0 10196 5 1 1 10195
0 10197 7 2 2 23540 34205
0 10198 7 1 2 24530 34451
0 10199 7 1 2 35202 10198
0 10200 7 2 2 32356 10199
0 10201 5 1 1 35204
0 10202 7 1 2 34969 35205
0 10203 5 1 1 10202
0 10204 7 1 2 10196 10203
0 10205 5 1 1 10204
0 10206 7 1 2 28817 10205
0 10207 5 1 1 10206
0 10208 7 1 2 24531 33922
0 10209 5 1 1 10208
0 10210 7 1 2 34449 10209
0 10211 5 1 1 10210
0 10212 7 1 2 27141 10211
0 10213 5 1 1 10212
0 10214 7 1 2 29838 34410
0 10215 5 1 1 10214
0 10216 7 1 2 10213 10215
0 10217 5 1 1 10216
0 10218 7 1 2 35196 10217
0 10219 5 2 1 10218
0 10220 7 1 2 10207 35206
0 10221 7 1 2 10191 10220
0 10222 5 1 1 10221
0 10223 7 1 2 23107 10222
0 10224 5 1 1 10223
0 10225 7 1 2 10174 10224
0 10226 5 1 1 10225
0 10227 7 1 2 24089 10226
0 10228 5 1 1 10227
0 10229 7 1 2 35188 10228
0 10230 7 1 2 10124 10229
0 10231 5 1 1 10230
0 10232 7 1 2 34848 10231
0 10233 5 1 1 10232
0 10234 7 1 2 10076 10233
0 10235 5 1 1 10234
0 10236 7 1 2 32970 10235
0 10237 5 1 1 10236
0 10238 7 1 2 25857 26988
0 10239 7 6 2 24700 23210
0 10240 7 3 2 24090 22927
0 10241 7 1 2 35208 35214
0 10242 7 1 2 10238 10241
0 10243 7 1 2 26843 33486
0 10244 7 1 2 10242 10243
0 10245 7 1 2 31592 10244
0 10246 5 1 1 10245
0 10247 7 9 2 24532 29292
0 10248 5 1 1 35217
0 10249 7 2 2 35218 34820
0 10250 7 1 2 31247 32439
0 10251 5 1 1 10250
0 10252 7 1 2 32340 34741
0 10253 5 1 1 10252
0 10254 7 1 2 10251 10253
0 10255 5 1 1 10254
0 10256 7 1 2 35226 10255
0 10257 5 1 1 10256
0 10258 7 1 2 27234 29858
0 10259 7 1 2 31689 10258
0 10260 7 1 2 31429 30975
0 10261 7 1 2 10259 10260
0 10262 5 1 1 10261
0 10263 7 1 2 10257 10262
0 10264 5 1 1 10263
0 10265 7 6 2 26080 33356
0 10266 7 1 2 25671 33018
0 10267 7 1 2 35228 10266
0 10268 7 1 2 10264 10267
0 10269 5 1 1 10268
0 10270 7 1 2 10246 10269
0 10271 5 1 1 10270
0 10272 7 1 2 24217 10271
0 10273 5 1 1 10272
0 10274 7 1 2 33677 35179
0 10275 5 1 1 10274
0 10276 7 1 2 35177 10275
0 10277 5 1 1 10276
0 10278 7 1 2 27512 10277
0 10279 5 1 1 10278
0 10280 7 1 2 30575 34411
0 10281 5 1 1 10280
0 10282 7 1 2 31584 33923
0 10283 5 1 1 10282
0 10284 7 1 2 10281 10283
0 10285 5 1 1 10284
0 10286 7 1 2 35197 10285
0 10287 5 1 1 10286
0 10288 7 1 2 24333 25779
0 10289 7 1 2 31081 10288
0 10290 7 1 2 34363 32352
0 10291 7 1 2 10289 10290
0 10292 5 1 1 10291
0 10293 7 1 2 10287 10292
0 10294 5 1 1 10293
0 10295 7 1 2 23969 10294
0 10296 5 1 1 10295
0 10297 7 1 2 35207 10296
0 10298 5 1 1 10297
0 10299 7 1 2 23108 10298
0 10300 5 1 1 10299
0 10301 7 1 2 10194 10201
0 10302 5 1 1 10301
0 10303 7 1 2 31643 10302
0 10304 5 1 1 10303
0 10305 7 1 2 28159 34788
0 10306 7 1 2 34645 10305
0 10307 5 1 1 10306
0 10308 7 1 2 10304 10307
0 10309 5 1 1 10308
0 10310 7 1 2 27142 10309
0 10311 5 1 1 10310
0 10312 7 1 2 34647 34990
0 10313 7 1 2 35199 10312
0 10314 5 1 1 10313
0 10315 7 1 2 10311 10314
0 10316 5 1 1 10315
0 10317 7 1 2 28818 10316
0 10318 5 1 1 10317
0 10319 7 1 2 33309 35194
0 10320 5 1 1 10319
0 10321 7 1 2 28486 35150
0 10322 5 1 1 10321
0 10323 7 1 2 10320 10322
0 10324 5 1 1 10323
0 10325 7 1 2 25858 35191
0 10326 7 1 2 10324 10325
0 10327 5 1 1 10326
0 10328 7 1 2 10318 10327
0 10329 7 1 2 10300 10328
0 10330 5 1 1 10329
0 10331 7 1 2 24091 10330
0 10332 5 1 1 10331
0 10333 7 1 2 22206 35189
0 10334 7 1 2 10332 10333
0 10335 7 1 2 10279 10334
0 10336 5 1 1 10335
0 10337 7 1 2 34928 32371
0 10338 5 1 1 10337
0 10339 7 4 2 24811 25170
0 10340 7 1 2 28160 35234
0 10341 7 1 2 34264 10340
0 10342 5 1 1 10341
0 10343 7 1 2 10338 10342
0 10344 5 1 1 10343
0 10345 7 1 2 35171 10344
0 10346 5 1 1 10345
0 10347 7 1 2 24218 10346
0 10348 7 1 2 35169 10347
0 10349 5 1 1 10348
0 10350 7 1 2 34294 10349
0 10351 7 1 2 10336 10350
0 10352 5 1 1 10351
0 10353 7 1 2 10273 10352
0 10354 7 1 2 10237 10353
0 10355 5 1 1 10354
0 10356 7 1 2 22398 10355
0 10357 5 1 1 10356
0 10358 7 1 2 10013 10357
0 10359 5 1 1 10358
0 10360 7 1 2 23653 10359
0 10361 5 1 1 10360
0 10362 7 1 2 32514 35015
0 10363 5 1 1 10362
0 10364 7 2 2 22655 32112
0 10365 7 1 2 33671 35238
0 10366 5 1 1 10365
0 10367 7 1 2 29162 35239
0 10368 5 1 1 10367
0 10369 7 2 2 24610 32295
0 10370 5 1 1 35240
0 10371 7 1 2 22656 32675
0 10372 5 1 1 10371
0 10373 7 1 2 10370 10372
0 10374 5 3 1 10373
0 10375 7 1 2 29033 35242
0 10376 5 1 1 10375
0 10377 7 1 2 10368 10376
0 10378 5 1 1 10377
0 10379 7 1 2 33357 10378
0 10380 5 1 1 10379
0 10381 7 1 2 10366 10380
0 10382 5 1 1 10381
0 10383 7 1 2 25596 10382
0 10384 5 1 1 10383
0 10385 7 1 2 10363 10384
0 10386 5 1 1 10385
0 10387 7 1 2 27782 10386
0 10388 5 1 1 10387
0 10389 7 1 2 22657 34326
0 10390 5 1 1 10389
0 10391 7 1 2 24611 34345
0 10392 5 1 1 10391
0 10393 7 1 2 28819 10392
0 10394 7 1 2 10390 10393
0 10395 5 1 1 10394
0 10396 7 2 2 34721 34384
0 10397 7 1 2 35245 32113
0 10398 5 1 1 10397
0 10399 7 1 2 34349 35243
0 10400 5 1 1 10399
0 10401 7 1 2 10398 10400
0 10402 5 1 1 10401
0 10403 7 1 2 27623 10402
0 10404 5 1 1 10403
0 10405 7 1 2 22658 34035
0 10406 5 1 1 10405
0 10407 7 1 2 24612 33150
0 10408 5 1 1 10407
0 10409 7 1 2 27608 34364
0 10410 7 1 2 10408 10409
0 10411 7 1 2 10406 10410
0 10412 5 1 1 10411
0 10413 7 1 2 10404 10412
0 10414 7 1 2 10395 10413
0 10415 5 1 1 10414
0 10416 7 1 2 25925 10415
0 10417 5 1 1 10416
0 10418 7 1 2 30925 34412
0 10419 5 1 1 10418
0 10420 7 1 2 32176 34452
0 10421 7 1 2 33991 10420
0 10422 5 1 1 10421
0 10423 7 1 2 10419 10422
0 10424 5 1 1 10423
0 10425 7 1 2 27902 10424
0 10426 5 1 1 10425
0 10427 7 1 2 34365 33945
0 10428 5 1 1 10427
0 10429 7 1 2 34428 32636
0 10430 5 1 1 10429
0 10431 7 1 2 30926 34441
0 10432 5 1 1 10431
0 10433 7 1 2 10430 10432
0 10434 5 1 1 10433
0 10435 7 1 2 28820 10434
0 10436 5 1 1 10435
0 10437 7 1 2 10428 10436
0 10438 7 1 2 10426 10437
0 10439 5 1 1 10438
0 10440 7 1 2 32523 10439
0 10441 5 1 1 10440
0 10442 7 3 2 27881 33625
0 10443 5 1 1 35247
0 10444 7 3 2 28868 33310
0 10445 5 1 1 35250
0 10446 7 1 2 27871 35021
0 10447 5 1 1 10446
0 10448 7 1 2 10445 10447
0 10449 5 1 1 10448
0 10450 7 1 2 25495 10449
0 10451 5 1 1 10450
0 10452 7 1 2 10443 10451
0 10453 5 1 1 10452
0 10454 7 1 2 34698 10453
0 10455 5 1 1 10454
0 10456 7 1 2 34350 32524
0 10457 7 1 2 32000 10456
0 10458 5 1 1 10457
0 10459 7 1 2 10455 10458
0 10460 5 1 1 10459
0 10461 7 1 2 32726 10460
0 10462 5 1 1 10461
0 10463 7 2 2 24613 33890
0 10464 5 1 1 35253
0 10465 7 1 2 23654 35254
0 10466 7 1 2 33692 10465
0 10467 5 1 1 10466
0 10468 7 1 2 10462 10467
0 10469 7 1 2 10441 10468
0 10470 5 1 1 10469
0 10471 7 1 2 27736 10470
0 10472 5 1 1 10471
0 10473 7 1 2 10417 10472
0 10474 7 1 2 10388 10473
0 10475 5 1 1 10474
0 10476 7 2 2 25404 31618
0 10477 7 1 2 35255 32473
0 10478 5 1 1 10477
0 10479 7 1 2 30976 34630
0 10480 5 1 1 10479
0 10481 7 1 2 10478 10480
0 10482 5 1 1 10481
0 10483 7 1 2 10475 10482
0 10484 5 1 1 10483
0 10485 7 1 2 28578 32882
0 10486 5 1 1 10485
0 10487 7 1 2 22052 29215
0 10488 7 1 2 28221 10487
0 10489 5 1 1 10488
0 10490 7 1 2 10486 10489
0 10491 5 1 1 10490
0 10492 7 1 2 24334 10491
0 10493 5 1 1 10492
0 10494 7 2 2 22053 22323
0 10495 7 2 2 28222 31915
0 10496 7 1 2 35257 35259
0 10497 5 1 1 10496
0 10498 7 1 2 10493 10497
0 10499 5 1 1 10498
0 10500 7 1 2 33358 10499
0 10501 5 1 1 10500
0 10502 7 2 2 22054 33311
0 10503 7 1 2 24335 35261
0 10504 7 1 2 35260 10503
0 10505 5 1 1 10504
0 10506 7 1 2 10501 10505
0 10507 5 1 1 10506
0 10508 7 1 2 25597 10507
0 10509 5 1 1 10508
0 10510 7 1 2 33693 32681
0 10511 5 1 1 10510
0 10512 7 1 2 26115 10511
0 10513 7 1 2 10509 10512
0 10514 5 1 1 10513
0 10515 7 1 2 33678 32682
0 10516 5 1 1 10515
0 10517 7 1 2 26131 10516
0 10518 5 1 1 10517
0 10519 7 1 2 25672 26223
0 10520 7 1 2 10518 10519
0 10521 7 1 2 10514 10520
0 10522 5 1 1 10521
0 10523 7 1 2 23970 34714
0 10524 5 1 1 10523
0 10525 7 1 2 24861 30287
0 10526 7 2 2 32594 10525
0 10527 7 1 2 33724 35263
0 10528 5 1 1 10527
0 10529 7 1 2 10524 10528
0 10530 5 1 1 10529
0 10531 7 1 2 26476 10530
0 10532 5 1 1 10531
0 10533 7 1 2 23754 33610
0 10534 5 1 1 10533
0 10535 7 2 2 25496 33487
0 10536 7 1 2 27557 30208
0 10537 5 1 1 10536
0 10538 7 1 2 26431 10537
0 10539 5 1 1 10538
0 10540 7 1 2 35265 10539
0 10541 5 1 1 10540
0 10542 7 1 2 24954 33709
0 10543 7 1 2 35264 10542
0 10544 5 1 1 10543
0 10545 7 1 2 10541 10544
0 10546 5 1 1 10545
0 10547 7 1 2 28821 10546
0 10548 5 1 1 10547
0 10549 7 1 2 10534 10548
0 10550 7 1 2 10532 10549
0 10551 5 1 1 10550
0 10552 7 1 2 27181 10551
0 10553 5 1 1 10552
0 10554 7 1 2 27558 30856
0 10555 5 1 1 10554
0 10556 7 1 2 21925 26426
0 10557 5 1 1 10556
0 10558 7 1 2 10555 10557
0 10559 5 1 1 10558
0 10560 7 1 2 33599 10559
0 10561 5 1 1 10560
0 10562 7 1 2 21926 33591
0 10563 5 1 1 10562
0 10564 7 1 2 10561 10563
0 10565 5 1 1 10564
0 10566 7 1 2 28822 10565
0 10567 5 1 1 10566
0 10568 7 1 2 27453 34424
0 10569 5 1 1 10568
0 10570 7 1 2 35062 10569
0 10571 5 1 1 10570
0 10572 7 1 2 24751 26943
0 10573 7 1 2 34792 10572
0 10574 5 1 1 10573
0 10575 7 1 2 10571 10574
0 10576 5 1 1 10575
0 10577 7 1 2 28123 10576
0 10578 5 1 1 10577
0 10579 7 1 2 33633 9064
0 10580 5 1 1 10579
0 10581 7 1 2 28109 10580
0 10582 5 1 1 10581
0 10583 7 1 2 10578 10582
0 10584 7 1 2 10567 10583
0 10585 5 1 1 10584
0 10586 7 1 2 23755 10585
0 10587 5 1 1 10586
0 10588 7 1 2 10553 10587
0 10589 7 1 2 10522 10588
0 10590 5 1 1 10589
0 10591 7 1 2 32583 10590
0 10592 5 1 1 10591
0 10593 7 3 2 25673 32308
0 10594 7 1 2 24393 32131
0 10595 5 1 1 10594
0 10596 7 1 2 32691 10595
0 10597 5 1 1 10596
0 10598 7 1 2 35267 10597
0 10599 5 1 1 10598
0 10600 7 4 2 24533 25598
0 10601 7 1 2 35270 32102
0 10602 5 1 1 10601
0 10603 7 1 2 10599 10602
0 10604 5 1 1 10603
0 10605 7 1 2 21821 10604
0 10606 5 1 1 10605
0 10607 7 1 2 32619 35268
0 10608 5 1 1 10607
0 10609 7 1 2 22480 29183
0 10610 7 1 2 27654 10609
0 10611 5 1 1 10610
0 10612 7 1 2 10608 10611
0 10613 5 1 1 10612
0 10614 7 1 2 24955 10613
0 10615 5 1 1 10614
0 10616 7 1 2 10606 10615
0 10617 5 1 1 10616
0 10618 7 1 2 34141 10617
0 10619 5 1 1 10618
0 10620 7 1 2 27844 28607
0 10621 5 1 1 10620
0 10622 7 1 2 32564 10621
0 10623 5 1 1 10622
0 10624 7 1 2 33600 10623
0 10625 5 1 1 10624
0 10626 7 2 2 23541 25926
0 10627 7 1 2 33359 32211
0 10628 7 1 2 32557 10627
0 10629 7 1 2 35274 10628
0 10630 5 1 1 10629
0 10631 7 1 2 10625 10630
0 10632 5 1 1 10631
0 10633 7 1 2 23655 10632
0 10634 5 1 1 10633
0 10635 7 1 2 34442 32212
0 10636 7 1 2 27745 10635
0 10637 5 1 1 10636
0 10638 7 1 2 10634 10637
0 10639 5 1 1 10638
0 10640 7 1 2 23838 10639
0 10641 5 1 1 10640
0 10642 7 1 2 21927 27559
0 10643 5 1 1 10642
0 10644 7 1 2 22545 26340
0 10645 5 1 1 10644
0 10646 7 1 2 10643 10645
0 10647 5 1 1 10646
0 10648 7 1 2 23756 10647
0 10649 5 1 1 10648
0 10650 7 1 2 24862 27591
0 10651 7 1 2 29792 32592
0 10652 7 1 2 10650 10651
0 10653 5 1 1 10652
0 10654 7 1 2 10649 10653
0 10655 5 1 1 10654
0 10656 7 1 2 33312 35049
0 10657 7 1 2 10655 10656
0 10658 5 1 1 10657
0 10659 7 1 2 10641 10658
0 10660 7 1 2 10619 10659
0 10661 5 1 1 10660
0 10662 7 1 2 25070 10661
0 10663 5 1 1 10662
0 10664 7 1 2 34429 32551
0 10665 5 1 1 10664
0 10666 7 1 2 34443 32753
0 10667 5 1 1 10666
0 10668 7 1 2 10665 10667
0 10669 5 1 1 10668
0 10670 7 1 2 27783 10669
0 10671 5 1 1 10670
0 10672 7 1 2 29896 35032
0 10673 7 1 2 35266 10672
0 10674 5 1 1 10673
0 10675 7 4 2 24092 22546
0 10676 5 1 1 35276
0 10677 7 1 2 33360 35277
0 10678 7 1 2 30099 10677
0 10679 5 1 1 10678
0 10680 7 1 2 10674 10679
0 10681 5 1 1 10680
0 10682 7 1 2 21822 10681
0 10683 5 1 1 10682
0 10684 7 1 2 27806 34142
0 10685 5 1 1 10684
0 10686 7 1 2 34322 10685
0 10687 5 1 1 10686
0 10688 7 1 2 35278 10687
0 10689 5 1 1 10688
0 10690 7 1 2 10683 10689
0 10691 5 1 1 10690
0 10692 7 1 2 21928 10691
0 10693 5 1 1 10692
0 10694 7 1 2 32757 34320
0 10695 5 1 1 10694
0 10696 7 1 2 10693 10695
0 10697 5 1 1 10696
0 10698 7 1 2 25927 10697
0 10699 5 1 1 10698
0 10700 7 1 2 34333 34986
0 10701 5 1 1 10700
0 10702 7 1 2 34434 10701
0 10703 5 1 1 10702
0 10704 7 1 2 21823 10703
0 10705 5 1 1 10704
0 10706 7 1 2 33601 33091
0 10707 5 1 1 10706
0 10708 7 1 2 10705 10707
0 10709 5 1 1 10708
0 10710 7 2 2 22547 27737
0 10711 5 1 1 35280
0 10712 7 2 2 32309 35281
0 10713 7 1 2 10709 35282
0 10714 5 1 1 10713
0 10715 7 1 2 10699 10714
0 10716 7 1 2 10671 10715
0 10717 7 1 2 10663 10716
0 10718 5 1 1 10717
0 10719 7 1 2 28823 10718
0 10720 5 1 1 10719
0 10721 7 1 2 25928 27609
0 10722 5 1 1 10721
0 10723 7 1 2 810 10722
0 10724 5 1 1 10723
0 10725 7 1 2 32310 10724
0 10726 5 1 1 10725
0 10727 7 1 2 29037 32648
0 10728 5 1 1 10727
0 10729 7 1 2 10726 10728
0 10730 5 1 1 10729
0 10731 7 1 2 29793 10730
0 10732 5 1 1 10731
0 10733 7 2 2 25929 35038
0 10734 5 1 1 35284
0 10735 7 1 2 31094 35285
0 10736 5 1 1 10735
0 10737 7 1 2 26341 28492
0 10738 5 1 1 10737
0 10739 7 1 2 10736 10738
0 10740 5 1 1 10739
0 10741 7 1 2 25859 10740
0 10742 5 1 1 10741
0 10743 7 2 2 21824 26507
0 10744 7 1 2 31512 35271
0 10745 7 1 2 35286 10744
0 10746 5 1 1 10745
0 10747 7 1 2 10742 10746
0 10748 5 1 1 10747
0 10749 7 1 2 23757 10748
0 10750 5 1 1 10749
0 10751 7 2 2 27996 28006
0 10752 7 1 2 33061 35288
0 10753 5 1 1 10752
0 10754 7 1 2 26355 10753
0 10755 5 1 1 10754
0 10756 7 1 2 24093 10755
0 10757 5 1 1 10756
0 10758 7 1 2 10750 10757
0 10759 7 1 2 10732 10758
0 10760 5 1 1 10759
0 10761 7 1 2 34413 10760
0 10762 5 1 1 10761
0 10763 7 3 2 28377 33684
0 10764 7 3 2 22928 28643
0 10765 7 1 2 31808 35293
0 10766 7 1 2 35290 10765
0 10767 5 1 1 10766
0 10768 7 1 2 33899 32213
0 10769 7 1 2 34543 10768
0 10770 7 1 2 35289 10769
0 10771 5 1 1 10770
0 10772 7 1 2 10767 10771
0 10773 5 1 1 10772
0 10774 7 1 2 24477 10773
0 10775 5 1 1 10774
0 10776 7 1 2 34817 32562
0 10777 5 1 1 10776
0 10778 7 1 2 33410 33463
0 10779 5 1 1 10778
0 10780 7 1 2 10777 10779
0 10781 5 1 1 10780
0 10782 7 1 2 23656 10781
0 10783 5 1 1 10782
0 10784 7 1 2 10775 10783
0 10785 5 1 1 10784
0 10786 7 1 2 23839 10785
0 10787 5 1 1 10786
0 10788 7 1 2 27610 29794
0 10789 5 1 1 10788
0 10790 7 1 2 27631 10789
0 10791 5 1 1 10790
0 10792 7 1 2 25930 10791
0 10793 5 1 1 10792
0 10794 7 1 2 28024 29795
0 10795 5 1 1 10794
0 10796 7 1 2 27668 10795
0 10797 7 1 2 10793 10796
0 10798 5 1 1 10797
0 10799 7 1 2 21929 10798
0 10800 5 1 1 10799
0 10801 7 1 2 22548 26353
0 10802 5 1 1 10801
0 10803 7 1 2 10800 10802
0 10804 5 1 1 10803
0 10805 7 1 2 33885 10804
0 10806 5 1 1 10805
0 10807 7 1 2 10787 10806
0 10808 7 1 2 10762 10807
0 10809 5 1 1 10808
0 10810 7 1 2 25071 10809
0 10811 5 1 1 10810
0 10812 7 2 2 27882 29757
0 10813 5 1 1 35296
0 10814 7 1 2 28081 29715
0 10815 5 1 1 10814
0 10816 7 1 2 10813 10815
0 10817 5 1 1 10816
0 10818 7 1 2 23109 10817
0 10819 5 1 1 10818
0 10820 7 3 2 22549 27903
0 10821 5 1 1 35298
0 10822 7 1 2 24094 35299
0 10823 5 1 1 10822
0 10824 7 1 2 10819 10823
0 10825 5 1 1 10824
0 10826 7 1 2 21930 10825
0 10827 5 1 1 10826
0 10828 7 1 2 24534 27513
0 10829 5 2 1 10828
0 10830 7 1 2 24956 35301
0 10831 7 1 2 33706 10830
0 10832 5 1 1 10831
0 10833 7 1 2 10827 10832
0 10834 5 1 1 10833
0 10835 7 1 2 33924 10834
0 10836 5 1 1 10835
0 10837 7 3 2 23971 27904
0 10838 5 1 1 35303
0 10839 7 1 2 27890 10838
0 10840 5 1 1 10839
0 10841 7 1 2 33925 10840
0 10842 5 1 1 10841
0 10843 7 1 2 28684 33669
0 10844 5 1 1 10843
0 10845 7 1 2 10842 10844
0 10846 5 1 1 10845
0 10847 7 1 2 29115 10846
0 10848 5 1 1 10847
0 10849 7 1 2 29266 33411
0 10850 5 1 1 10849
0 10851 7 1 2 10848 10850
0 10852 5 1 1 10851
0 10853 7 1 2 22055 10852
0 10854 5 1 1 10853
0 10855 7 2 2 23110 33658
0 10856 7 1 2 29253 35306
0 10857 7 1 2 30845 10856
0 10858 5 1 1 10857
0 10859 7 1 2 10854 10858
0 10860 7 1 2 10836 10859
0 10861 5 1 1 10860
0 10862 7 1 2 27784 10861
0 10863 5 1 1 10862
0 10864 7 2 2 29796 34366
0 10865 7 1 2 27715 35308
0 10866 5 1 1 10865
0 10867 7 1 2 22263 28742
0 10868 7 1 2 30653 10867
0 10869 7 1 2 34544 10868
0 10870 5 1 1 10869
0 10871 7 1 2 10866 10870
0 10872 5 1 1 10871
0 10873 7 1 2 35283 10872
0 10874 5 1 1 10873
0 10875 7 1 2 31195 34982
0 10876 5 1 1 10875
0 10877 7 1 2 32748 10876
0 10878 5 1 1 10877
0 10879 7 1 2 33926 10878
0 10880 5 1 1 10879
0 10881 7 1 2 33626 32754
0 10882 5 1 1 10881
0 10883 7 1 2 10880 10882
0 10884 5 1 1 10883
0 10885 7 1 2 27624 10884
0 10886 5 1 1 10885
0 10887 7 3 2 22550 24812
0 10888 7 1 2 24336 23657
0 10889 7 1 2 35310 10888
0 10890 7 1 2 35269 10889
0 10891 7 1 2 35309 10890
0 10892 5 1 1 10891
0 10893 7 1 2 10886 10892
0 10894 5 1 1 10893
0 10895 7 1 2 25931 10894
0 10896 5 1 1 10895
0 10897 7 1 2 10874 10896
0 10898 7 1 2 10863 10897
0 10899 7 1 2 10811 10898
0 10900 7 1 2 10720 10899
0 10901 7 1 2 10592 10900
0 10902 5 1 1 10901
0 10903 7 1 2 31208 10902
0 10904 5 1 1 10903
0 10905 7 1 2 10484 10904
0 10906 5 1 1 10905
0 10907 7 1 2 28535 10906
0 10908 5 1 1 10907
0 10909 7 1 2 28240 30878
0 10910 5 1 1 10909
0 10911 7 1 2 28983 30352
0 10912 5 1 1 10911
0 10913 7 1 2 10910 10912
0 10914 5 1 1 10913
0 10915 7 3 2 24280 22755
0 10916 7 2 2 22207 35313
0 10917 5 1 1 35316
0 10918 7 3 2 22264 24701
0 10919 7 1 2 24219 35318
0 10920 5 1 1 10919
0 10921 7 1 2 10917 10920
0 10922 5 4 1 10921
0 10923 7 1 2 34596 32532
0 10924 5 1 1 10923
0 10925 7 1 2 28296 33507
0 10926 5 1 1 10925
0 10927 7 9 2 22803 25405
0 10928 5 2 1 35325
0 10929 7 1 2 30631 35326
0 10930 5 1 1 10929
0 10931 7 1 2 10926 10930
0 10932 5 1 1 10931
0 10933 7 1 2 22324 10932
0 10934 5 1 1 10933
0 10935 7 1 2 30733 35327
0 10936 5 1 1 10935
0 10937 7 1 2 10934 10936
0 10938 5 2 1 10937
0 10939 7 1 2 25932 35336
0 10940 5 1 1 10939
0 10941 7 1 2 25976 33853
0 10942 5 1 1 10941
0 10943 7 1 2 10940 10942
0 10944 5 1 1 10943
0 10945 7 4 2 25599 10944
0 10946 7 1 2 23972 35338
0 10947 5 1 1 10946
0 10948 7 2 2 28310 28026
0 10949 7 2 2 25860 34485
0 10950 7 1 2 35342 35344
0 10951 5 1 1 10950
0 10952 7 1 2 10947 10951
0 10953 5 1 1 10952
0 10954 7 1 2 27514 10953
0 10955 5 1 1 10954
0 10956 7 1 2 22056 7982
0 10957 5 1 1 10956
0 10958 7 1 2 35339 10957
0 10959 5 1 1 10958
0 10960 7 3 2 23973 22325
0 10961 7 1 2 34486 35346
0 10962 7 1 2 28315 10961
0 10963 5 1 1 10962
0 10964 7 1 2 10959 10963
0 10965 7 1 2 10955 10964
0 10966 5 1 1 10965
0 10967 7 1 2 22659 10966
0 10968 5 1 1 10967
0 10969 7 1 2 35340 35241
0 10970 5 1 1 10969
0 10971 7 1 2 23758 10970
0 10972 7 1 2 10968 10971
0 10973 5 1 1 10972
0 10974 7 1 2 33854 32639
0 10975 5 1 1 10974
0 10976 7 1 2 27515 33844
0 10977 5 1 1 10976
0 10978 7 2 2 28297 32727
0 10979 7 1 2 24752 35349
0 10980 5 1 1 10979
0 10981 7 1 2 10977 10980
0 10982 5 1 1 10981
0 10983 7 1 2 21931 10982
0 10984 5 1 1 10983
0 10985 7 1 2 28298 33987
0 10986 5 1 1 10985
0 10987 7 1 2 33847 10986
0 10988 5 1 1 10987
0 10989 7 1 2 30209 10988
0 10990 5 1 1 10989
0 10991 7 1 2 22481 28361
0 10992 7 1 2 33615 10991
0 10993 5 1 1 10992
0 10994 7 1 2 10990 10993
0 10995 5 1 1 10994
0 10996 7 1 2 21825 10995
0 10997 5 1 1 10996
0 10998 7 1 2 23974 33833
0 10999 7 1 2 31733 10998
0 11000 5 1 1 10999
0 11001 7 1 2 10997 11000
0 11002 7 1 2 10984 11001
0 11003 5 1 1 11002
0 11004 7 1 2 27322 11003
0 11005 5 1 1 11004
0 11006 7 1 2 10975 11005
0 11007 5 1 1 11006
0 11008 7 1 2 24813 11007
0 11009 5 1 1 11008
0 11010 7 2 2 25933 34004
0 11011 7 1 2 30511 33801
0 11012 7 1 2 35351 11011
0 11013 5 1 1 11012
0 11014 7 1 2 24337 11013
0 11015 7 1 2 11009 11014
0 11016 5 1 1 11015
0 11017 7 2 2 22867 33019
0 11018 5 1 1 35353
0 11019 7 1 2 11018 33483
0 11020 5 1 1 11019
0 11021 7 1 2 34005 11020
0 11022 5 1 1 11021
0 11023 7 3 2 22804 27681
0 11024 7 1 2 26797 35355
0 11025 5 1 1 11024
0 11026 7 1 2 11022 11025
0 11027 5 1 1 11026
0 11028 7 1 2 24394 11027
0 11029 5 1 1 11028
0 11030 7 2 2 22399 33442
0 11031 7 2 2 23542 32074
0 11032 7 1 2 35358 35360
0 11033 5 1 1 11032
0 11034 7 1 2 11029 11033
0 11035 5 1 1 11034
0 11036 7 1 2 32641 11035
0 11037 5 1 1 11036
0 11038 7 1 2 22326 11037
0 11039 5 1 1 11038
0 11040 7 1 2 32525 11039
0 11041 7 1 2 11016 11040
0 11042 5 1 1 11041
0 11043 7 1 2 27689 33855
0 11044 5 1 1 11043
0 11045 7 1 2 32450 34006
0 11046 5 1 1 11045
0 11047 7 1 2 25406 31916
0 11048 7 1 2 34536 11047
0 11049 5 1 1 11048
0 11050 7 1 2 11046 11049
0 11051 5 1 1 11050
0 11052 7 1 2 25934 11051
0 11053 5 1 1 11052
0 11054 7 1 2 11044 11053
0 11055 5 1 1 11054
0 11056 7 3 2 23975 32728
0 11057 5 1 1 35362
0 11058 7 1 2 22660 35363
0 11059 5 1 1 11058
0 11060 7 1 2 10464 11059
0 11061 5 2 1 11060
0 11062 7 1 2 23658 35365
0 11063 7 1 2 11055 11062
0 11064 5 1 1 11063
0 11065 7 1 2 25674 11064
0 11066 7 1 2 11042 11065
0 11067 5 1 1 11066
0 11068 7 1 2 10973 11067
0 11069 5 1 1 11068
0 11070 7 1 2 10924 11069
0 11071 5 1 1 11070
0 11072 7 1 2 35321 11071
0 11073 5 1 1 11072
0 11074 7 2 2 24281 24702
0 11075 7 4 2 28390 35367
0 11076 7 2 2 35369 32409
0 11077 7 1 2 34471 35373
0 11078 5 1 1 11077
0 11079 7 3 2 22756 24814
0 11080 7 3 2 22208 34151
0 11081 7 3 2 35375 35378
0 11082 5 1 1 35381
0 11083 7 1 2 25752 34026
0 11084 5 1 1 11083
0 11085 7 1 2 11082 11084
0 11086 5 4 1 11085
0 11087 7 1 2 32606 35384
0 11088 5 1 1 11087
0 11089 7 9 2 22757 34901
0 11090 7 6 2 25861 35388
0 11091 7 1 2 32642 35397
0 11092 5 1 1 11091
0 11093 7 1 2 11088 11092
0 11094 5 1 1 11093
0 11095 7 1 2 23543 11094
0 11096 5 1 1 11095
0 11097 7 1 2 11078 11096
0 11098 5 1 1 11097
0 11099 7 1 2 26116 11098
0 11100 5 1 1 11099
0 11101 7 1 2 26132 29254
0 11102 7 2 2 33802 11101
0 11103 7 1 2 35403 35385
0 11104 5 1 1 11103
0 11105 7 1 2 11100 11104
0 11106 5 1 1 11105
0 11107 7 1 2 26224 32526
0 11108 7 1 2 11106 11107
0 11109 5 1 1 11108
0 11110 7 1 2 25935 35386
0 11111 5 1 1 11110
0 11112 7 1 2 26117 35398
0 11113 5 1 1 11112
0 11114 7 1 2 11111 11113
0 11115 5 1 1 11114
0 11116 7 1 2 29255 35366
0 11117 7 1 2 11115 11116
0 11118 5 1 1 11117
0 11119 7 1 2 11109 11118
0 11120 5 1 1 11119
0 11121 7 1 2 25675 11120
0 11122 5 1 1 11121
0 11123 7 1 2 28824 35389
0 11124 5 1 1 11123
0 11125 7 1 2 33501 31940
0 11126 5 1 1 11125
0 11127 7 1 2 11124 11126
0 11128 5 6 1 11127
0 11129 7 1 2 25936 35405
0 11130 5 1 1 11129
0 11131 7 3 2 22400 26497
0 11132 7 1 2 35370 35411
0 11133 5 1 1 11132
0 11134 7 1 2 11130 11133
0 11135 5 1 1 11134
0 11136 7 1 2 25600 11135
0 11137 7 1 2 35244 11136
0 11138 5 1 1 11137
0 11139 7 1 2 26342 32515
0 11140 7 1 2 35406 11139
0 11141 5 1 1 11140
0 11142 7 1 2 11138 11141
0 11143 5 1 1 11142
0 11144 7 1 2 34342 11143
0 11145 5 1 1 11144
0 11146 7 1 2 11122 11145
0 11147 5 1 1 11146
0 11148 7 1 2 34578 11147
0 11149 5 1 1 11148
0 11150 7 5 2 23544 27406
0 11151 7 2 2 28337 35414
0 11152 7 2 2 24703 34504
0 11153 7 2 2 34487 35421
0 11154 7 2 2 35419 35423
0 11155 5 1 1 35425
0 11156 7 3 2 26769 33900
0 11157 7 4 2 25676 28644
0 11158 7 1 2 34101 33803
0 11159 5 1 1 11158
0 11160 7 1 2 24753 33829
0 11161 5 1 1 11160
0 11162 7 1 2 11159 11161
0 11163 5 1 1 11162
0 11164 7 2 2 35430 11163
0 11165 7 2 2 24863 35434
0 11166 7 1 2 35427 35436
0 11167 5 1 1 11166
0 11168 7 1 2 11155 11167
0 11169 5 1 1 11168
0 11170 7 1 2 28825 11169
0 11171 5 1 1 11170
0 11172 7 1 2 34488 35382
0 11173 7 1 2 35420 11172
0 11174 5 2 1 11173
0 11175 7 3 2 24282 25753
0 11176 7 2 2 27983 35440
0 11177 7 1 2 35443 35437
0 11178 5 1 1 11177
0 11179 7 1 2 35438 11178
0 11180 7 1 2 11171 11179
0 11181 5 1 1 11180
0 11182 7 1 2 32527 11181
0 11183 5 1 1 11182
0 11184 7 4 2 26081 35441
0 11185 7 1 2 35435 35445
0 11186 5 1 1 11185
0 11187 7 2 2 22209 33402
0 11188 7 1 2 27407 33508
0 11189 7 1 2 31602 11188
0 11190 7 2 2 35449 11189
0 11191 5 2 1 35451
0 11192 7 1 2 11186 35453
0 11193 5 1 1 11192
0 11194 7 1 2 32528 11193
0 11195 5 1 1 11194
0 11196 7 2 2 32729 35431
0 11197 7 1 2 35446 35455
0 11198 5 1 1 11197
0 11199 7 1 2 35415 35399
0 11200 5 1 1 11199
0 11201 7 1 2 11198 11200
0 11202 5 1 1 11201
0 11203 7 1 2 34102 11202
0 11204 5 1 1 11203
0 11205 7 1 2 27382 35452
0 11206 5 1 1 11205
0 11207 7 1 2 11204 11206
0 11208 5 1 1 11207
0 11209 7 1 2 23976 11208
0 11210 5 1 1 11209
0 11211 7 1 2 23840 33966
0 11212 5 1 1 11211
0 11213 7 1 2 34118 11212
0 11214 5 2 1 11213
0 11215 7 2 2 23841 22805
0 11216 5 1 1 35459
0 11217 7 1 2 22482 11216
0 11218 5 1 1 11217
0 11219 7 1 2 26370 33431
0 11220 7 1 2 11218 11219
0 11221 7 2 2 35457 11220
0 11222 7 1 2 35400 35461
0 11223 5 1 1 11222
0 11224 7 1 2 11210 11223
0 11225 5 1 1 11224
0 11226 7 1 2 22661 11225
0 11227 5 1 1 11226
0 11228 7 1 2 11195 11227
0 11229 5 1 1 11228
0 11230 7 1 2 25937 11229
0 11231 5 1 1 11230
0 11232 7 2 2 24864 35456
0 11233 7 1 2 35463 35428
0 11234 5 1 1 11233
0 11235 7 2 2 28272 34505
0 11236 7 1 2 27825 28676
0 11237 7 1 2 35465 11236
0 11238 5 1 1 11237
0 11239 7 1 2 11234 11238
0 11240 5 1 1 11239
0 11241 7 1 2 34103 11240
0 11242 5 1 1 11241
0 11243 7 1 2 26798 27383
0 11244 7 2 2 27655 11243
0 11245 7 1 2 35467 35424
0 11246 5 1 1 11245
0 11247 7 1 2 11242 11246
0 11248 5 1 1 11247
0 11249 7 1 2 23977 11248
0 11250 5 1 1 11249
0 11251 7 2 2 22929 35462
0 11252 7 1 2 35469 35466
0 11253 5 1 1 11252
0 11254 7 1 2 22662 11253
0 11255 7 1 2 11250 11254
0 11256 5 1 1 11255
0 11257 7 1 2 27182 35426
0 11258 5 1 1 11257
0 11259 7 3 2 26118 34430
0 11260 5 1 1 35471
0 11261 7 1 2 31728 32098
0 11262 7 2 2 35472 11261
0 11263 7 1 2 21826 35474
0 11264 5 1 1 11263
0 11265 7 1 2 11258 11264
0 11266 5 1 1 11265
0 11267 7 1 2 30270 11266
0 11268 5 1 1 11267
0 11269 7 1 2 22057 35475
0 11270 5 1 1 11269
0 11271 7 1 2 24614 11270
0 11272 7 1 2 11268 11271
0 11273 5 1 1 11272
0 11274 7 1 2 28826 11273
0 11275 7 1 2 11256 11274
0 11276 5 1 1 11275
0 11277 7 1 2 35464 35444
0 11278 5 1 1 11277
0 11279 7 1 2 26207 35416
0 11280 7 1 2 35383 11279
0 11281 5 1 1 11280
0 11282 7 1 2 11278 11281
0 11283 5 1 1 11282
0 11284 7 1 2 34104 11283
0 11285 5 1 1 11284
0 11286 7 4 2 22758 24754
0 11287 7 2 2 24815 35476
0 11288 7 1 2 27649 34902
0 11289 7 1 2 35480 11288
0 11290 7 1 2 35468 11289
0 11291 5 1 1 11290
0 11292 7 1 2 11285 11291
0 11293 5 1 1 11292
0 11294 7 1 2 23978 11293
0 11295 5 1 1 11294
0 11296 7 1 2 27652 35390
0 11297 7 1 2 35470 11296
0 11298 5 1 1 11297
0 11299 7 1 2 11295 11298
0 11300 5 1 1 11299
0 11301 7 1 2 22663 11300
0 11302 5 1 1 11301
0 11303 7 3 2 25497 34105
0 11304 7 1 2 27592 30649
0 11305 7 1 2 35482 11304
0 11306 7 2 2 35371 11305
0 11307 5 1 1 35485
0 11308 7 1 2 35454 11307
0 11309 5 1 1 11308
0 11310 7 1 2 25938 11309
0 11311 5 1 1 11310
0 11312 7 1 2 28299 27593
0 11313 7 2 2 35356 11312
0 11314 7 1 2 33502 32079
0 11315 7 1 2 35487 11314
0 11316 5 1 1 11315
0 11317 7 1 2 35439 11316
0 11318 7 1 2 11311 11317
0 11319 5 1 1 11318
0 11320 7 1 2 21827 11319
0 11321 5 1 1 11320
0 11322 7 3 2 22483 22868
0 11323 5 1 1 35489
0 11324 7 1 2 25692 35490
0 11325 7 1 2 25939 11324
0 11326 7 1 2 35417 11325
0 11327 7 1 2 31872 11326
0 11328 5 1 1 11327
0 11329 7 2 2 24755 26498
0 11330 7 1 2 31603 35492
0 11331 7 1 2 35379 32657
0 11332 7 1 2 11330 11331
0 11333 5 1 1 11332
0 11334 7 1 2 11328 11333
0 11335 7 1 2 11321 11334
0 11336 5 1 1 11335
0 11337 7 1 2 30271 11336
0 11338 5 1 1 11337
0 11339 7 1 2 22058 25940
0 11340 7 1 2 35486 11339
0 11341 5 1 1 11340
0 11342 7 2 2 22327 34506
0 11343 7 1 2 32134 33146
0 11344 7 1 2 35494 11343
0 11345 7 1 2 35488 11344
0 11346 5 1 1 11345
0 11347 7 1 2 11341 11346
0 11348 7 1 2 11338 11347
0 11349 5 1 1 11348
0 11350 7 1 2 24615 11349
0 11351 5 1 1 11350
0 11352 7 1 2 11302 11351
0 11353 7 1 2 11276 11352
0 11354 7 1 2 11231 11353
0 11355 7 1 2 11183 11354
0 11356 7 1 2 11149 11355
0 11357 7 1 2 11073 11356
0 11358 5 1 1 11357
0 11359 7 1 2 10914 11358
0 11360 5 1 1 11359
0 11361 7 2 2 22265 34579
0 11362 5 1 1 35496
0 11363 7 2 2 24283 35328
0 11364 5 1 1 35498
0 11365 7 1 2 11362 11364
0 11366 5 6 1 11365
0 11367 7 1 2 26770 35500
0 11368 5 1 1 11367
0 11369 7 1 2 33313 35085
0 11370 5 1 1 11369
0 11371 7 1 2 11368 11370
0 11372 5 1 1 11371
0 11373 7 1 2 27682 11372
0 11374 7 1 2 32743 11373
0 11375 5 1 1 11374
0 11376 7 2 2 24284 34580
0 11377 5 1 1 35506
0 11378 7 1 2 11377 7548
0 11379 5 2 1 11378
0 11380 7 1 2 25754 35508
0 11381 5 1 1 11380
0 11382 7 1 2 26598 34894
0 11383 5 1 1 11382
0 11384 7 1 2 11381 11383
0 11385 5 2 1 11384
0 11386 7 1 2 21932 32716
0 11387 5 1 1 11386
0 11388 7 1 2 32707 11387
0 11389 5 3 1 11388
0 11390 7 1 2 26499 35512
0 11391 7 1 2 35510 11390
0 11392 5 1 1 11391
0 11393 7 1 2 11375 11392
0 11394 5 1 1 11393
0 11395 7 1 2 22328 11394
0 11396 5 1 1 11395
0 11397 7 2 2 34903 35376
0 11398 5 1 1 35515
0 11399 7 1 2 24285 31941
0 11400 5 1 1 11399
0 11401 7 1 2 11398 11400
0 11402 5 1 1 11401
0 11403 7 1 2 34581 11402
0 11404 5 1 1 11403
0 11405 7 1 2 22806 4383
0 11406 5 1 1 11405
0 11407 7 1 2 24756 4645
0 11408 5 1 1 11407
0 11409 7 2 2 11406 11408
0 11410 7 1 2 35517 35322
0 11411 5 1 1 11410
0 11412 7 1 2 11404 11411
0 11413 5 1 1 11412
0 11414 7 1 2 25969 35513
0 11415 7 1 2 11413 11414
0 11416 5 1 1 11415
0 11417 7 1 2 11396 11416
0 11418 5 1 1 11417
0 11419 7 1 2 24395 11418
0 11420 5 1 1 11419
0 11421 7 1 2 34582 35387
0 11422 5 1 1 11421
0 11423 7 1 2 28775 35334
0 11424 5 1 1 11423
0 11425 7 1 2 26099 34011
0 11426 5 1 1 11425
0 11427 7 3 2 11424 11426
0 11428 7 1 2 35519 35323
0 11429 5 1 1 11428
0 11430 7 1 2 11422 11429
0 11431 5 2 1 11430
0 11432 7 1 2 25885 35514
0 11433 7 1 2 35522 11432
0 11434 5 1 1 11433
0 11435 7 1 2 11420 11434
0 11436 5 1 1 11435
0 11437 7 1 2 23659 11436
0 11438 5 1 1 11437
0 11439 7 4 2 22807 24816
0 11440 7 4 2 22266 35524
0 11441 7 1 2 28347 35528
0 11442 5 1 1 11441
0 11443 7 1 2 25709 31951
0 11444 5 1 1 11443
0 11445 7 1 2 11442 11444
0 11446 5 1 1 11445
0 11447 7 1 2 32584 11446
0 11448 5 1 1 11447
0 11449 7 1 2 33509 33279
0 11450 7 1 2 33461 11449
0 11451 5 1 1 11450
0 11452 7 2 2 25710 25755
0 11453 5 1 1 35532
0 11454 7 1 2 31530 32044
0 11455 7 1 2 35533 11454
0 11456 5 1 1 11455
0 11457 7 1 2 11451 11456
0 11458 7 1 2 11448 11457
0 11459 5 1 1 11458
0 11460 7 1 2 24338 11459
0 11461 5 1 1 11460
0 11462 7 2 2 26771 33361
0 11463 5 1 1 35534
0 11464 7 1 2 11463 11453
0 11465 5 2 1 11464
0 11466 7 1 2 22551 28618
0 11467 7 1 2 33280 11466
0 11468 7 1 2 35536 11467
0 11469 5 1 1 11468
0 11470 7 1 2 11461 11469
0 11471 5 1 1 11470
0 11472 7 1 2 32686 11471
0 11473 5 1 1 11472
0 11474 7 1 2 22059 34880
0 11475 5 1 1 11474
0 11476 7 2 2 31653 32311
0 11477 7 1 2 27454 35538
0 11478 5 1 1 11477
0 11479 7 2 2 11475 11478
0 11480 5 3 1 35540
0 11481 7 1 2 34234 35542
0 11482 7 1 2 35523 11481
0 11483 5 1 1 11482
0 11484 7 1 2 11473 11483
0 11485 7 1 2 11438 11484
0 11486 5 1 1 11485
0 11487 7 1 2 23545 11486
0 11488 5 1 1 11487
0 11489 7 2 2 24478 28579
0 11490 5 1 1 35545
0 11491 7 1 2 35546 32702
0 11492 5 1 1 11491
0 11493 7 1 2 22484 28580
0 11494 5 1 1 11493
0 11495 7 1 2 29228 11494
0 11496 5 2 1 11495
0 11497 7 1 2 23842 11323
0 11498 5 1 1 11497
0 11499 7 1 2 32312 11498
0 11500 7 1 2 35547 11499
0 11501 5 1 1 11500
0 11502 7 1 2 11492 11501
0 11503 5 1 1 11502
0 11504 7 1 2 24957 11503
0 11505 5 1 1 11504
0 11506 7 3 2 23843 29216
0 11507 5 1 1 35549
0 11508 7 1 2 28199 35550
0 11509 5 1 1 11508
0 11510 7 4 2 27183 27516
0 11511 7 1 2 35552 32405
0 11512 5 1 1 11511
0 11513 7 1 2 1866 11512
0 11514 5 1 1 11513
0 11515 7 1 2 23979 11514
0 11516 5 1 1 11515
0 11517 7 1 2 11509 11516
0 11518 5 1 1 11517
0 11519 7 1 2 22060 11518
0 11520 5 1 1 11519
0 11521 7 1 2 11505 11520
0 11522 5 1 1 11521
0 11523 7 1 2 26635 11522
0 11524 5 1 1 11523
0 11525 7 4 2 27872 33478
0 11526 7 1 2 35556 32668
0 11527 5 1 1 11526
0 11528 7 1 2 11524 11527
0 11529 5 1 1 11528
0 11530 7 1 2 24339 11529
0 11531 5 1 1 11530
0 11532 7 1 2 32442 32679
0 11533 5 1 1 11532
0 11534 7 1 2 11531 11533
0 11535 5 1 1 11534
0 11536 7 1 2 24396 11535
0 11537 5 1 1 11536
0 11538 7 1 2 29163 32684
0 11539 5 1 1 11538
0 11540 7 1 2 11537 11539
0 11541 5 1 1 11540
0 11542 7 1 2 32570 35511
0 11543 5 1 1 11542
0 11544 7 2 2 24220 33362
0 11545 7 1 2 31754 34821
0 11546 7 1 2 35560 11545
0 11547 5 1 1 11546
0 11548 7 1 2 11543 11547
0 11549 5 1 1 11548
0 11550 7 1 2 11541 11549
0 11551 5 1 1 11550
0 11552 7 1 2 31824 35537
0 11553 5 1 1 11552
0 11554 7 1 2 28827 33951
0 11555 7 1 2 35429 11554
0 11556 5 1 1 11555
0 11557 7 1 2 11553 11556
0 11558 5 1 1 11557
0 11559 7 1 2 32744 11558
0 11560 5 1 1 11559
0 11561 7 1 2 23447 11560
0 11562 5 1 1 11561
0 11563 7 1 2 29627 32585
0 11564 5 1 1 11563
0 11565 7 1 2 5798 11564
0 11566 5 1 1 11565
0 11567 7 1 2 32313 11566
0 11568 5 1 1 11567
0 11569 7 1 2 28223 32586
0 11570 5 1 1 11569
0 11571 7 1 2 9192 11570
0 11572 5 1 1 11571
0 11573 7 1 2 22061 11572
0 11574 5 1 1 11573
0 11575 7 1 2 11568 11574
0 11576 5 1 1 11575
0 11577 7 1 2 25756 34212
0 11578 5 1 1 11577
0 11579 7 1 2 25711 26772
0 11580 5 1 1 11579
0 11581 7 1 2 9946 11580
0 11582 5 1 1 11581
0 11583 7 1 2 28828 11582
0 11584 5 1 1 11583
0 11585 7 1 2 25757 33514
0 11586 5 1 1 11585
0 11587 7 1 2 24865 11586
0 11588 7 1 2 11584 11587
0 11589 5 1 1 11588
0 11590 7 1 2 24757 35447
0 11591 5 1 1 11590
0 11592 7 1 2 22930 11591
0 11593 5 1 1 11592
0 11594 7 1 2 24397 11593
0 11595 7 1 2 11589 11594
0 11596 5 1 1 11595
0 11597 7 1 2 11578 11596
0 11598 5 1 1 11597
0 11599 7 1 2 11576 11598
0 11600 5 1 1 11599
0 11601 7 1 2 25407 11600
0 11602 5 1 1 11601
0 11603 7 1 2 28645 11602
0 11604 7 1 2 11562 11603
0 11605 5 1 1 11604
0 11606 7 1 2 25677 11605
0 11607 7 1 2 11551 11606
0 11608 7 1 2 11488 11607
0 11609 5 1 1 11608
0 11610 7 2 2 28829 34007
0 11611 7 1 2 28613 10676
0 11612 5 2 1 11611
0 11613 7 1 2 25072 35564
0 11614 5 1 1 11613
0 11615 7 1 2 32548 11614
0 11616 5 2 1 11615
0 11617 7 1 2 35562 35566
0 11618 5 1 1 11617
0 11619 7 2 2 25408 32762
0 11620 7 1 2 24817 34537
0 11621 7 1 2 35568 11620
0 11622 5 1 1 11621
0 11623 7 1 2 11618 11622
0 11624 5 1 1 11623
0 11625 7 1 2 22931 11624
0 11626 5 1 1 11625
0 11627 7 1 2 25862 33952
0 11628 7 1 2 35569 11627
0 11629 5 1 1 11628
0 11630 7 1 2 11626 11629
0 11631 5 1 1 11630
0 11632 7 1 2 25601 11631
0 11633 5 1 1 11632
0 11634 7 2 2 25073 29546
0 11635 5 1 1 35570
0 11636 7 1 2 29293 30998
0 11637 5 1 1 11636
0 11638 7 2 2 23111 11637
0 11639 5 1 1 35572
0 11640 7 1 2 11635 11639
0 11641 5 1 1 11640
0 11642 7 3 2 22329 22808
0 11643 7 1 2 28343 35574
0 11644 7 1 2 11641 11643
0 11645 5 1 1 11644
0 11646 7 1 2 11633 11645
0 11647 5 1 1 11646
0 11648 7 1 2 22401 11647
0 11649 5 1 1 11648
0 11650 7 3 2 22402 22809
0 11651 7 1 2 28338 35577
0 11652 7 1 2 27883 11651
0 11653 5 2 1 11652
0 11654 7 2 2 25989 33830
0 11655 7 1 2 22810 35582
0 11656 5 1 1 11655
0 11657 7 1 2 22932 31383
0 11658 7 3 2 31971 11657
0 11659 7 1 2 34489 35584
0 11660 5 1 1 11659
0 11661 7 1 2 11656 11660
0 11662 5 1 1 11661
0 11663 7 1 2 25602 11662
0 11664 5 1 1 11663
0 11665 7 1 2 35580 11664
0 11666 5 1 1 11665
0 11667 7 1 2 32587 11666
0 11668 5 1 1 11667
0 11669 7 1 2 25603 28339
0 11670 7 1 2 34498 11669
0 11671 7 1 2 32763 11670
0 11672 5 1 1 11671
0 11673 7 1 2 23546 11672
0 11674 7 1 2 11668 11673
0 11675 7 1 2 11649 11674
0 11676 5 1 1 11675
0 11677 7 1 2 28776 34012
0 11678 5 1 1 11677
0 11679 7 1 2 25872 35335
0 11680 5 1 1 11679
0 11681 7 5 2 11678 11680
0 11682 7 1 2 26343 35567
0 11683 5 1 1 11682
0 11684 7 5 2 28463 26427
0 11685 5 1 1 35592
0 11686 7 1 2 27560 30927
0 11687 5 1 1 11686
0 11688 7 1 2 11685 11687
0 11689 5 1 1 11688
0 11690 7 1 2 32588 11689
0 11691 5 1 1 11690
0 11692 7 1 2 27561 32764
0 11693 5 1 1 11692
0 11694 7 1 2 11691 11693
0 11695 7 1 2 11683 11694
0 11696 5 1 1 11695
0 11697 7 1 2 35587 11696
0 11698 5 1 1 11697
0 11699 7 2 2 34492 32155
0 11700 5 1 1 35597
0 11701 7 1 2 25604 35598
0 11702 7 1 2 32766 11701
0 11703 5 1 1 11702
0 11704 7 1 2 25498 11703
0 11705 7 1 2 11698 11704
0 11706 5 1 1 11705
0 11707 7 1 2 35324 11706
0 11708 7 1 2 11676 11707
0 11709 5 1 1 11708
0 11710 7 2 2 29256 35401
0 11711 5 2 1 35599
0 11712 7 2 2 24221 34176
0 11713 7 1 2 29716 35603
0 11714 7 1 2 35093 11713
0 11715 5 2 1 11714
0 11716 7 1 2 32062 35407
0 11717 5 1 1 11716
0 11718 7 1 2 35605 11717
0 11719 5 1 1 11718
0 11720 7 1 2 25499 11719
0 11721 5 1 1 11720
0 11722 7 1 2 35601 11721
0 11723 5 1 1 11722
0 11724 7 1 2 29507 11723
0 11725 5 1 1 11724
0 11726 7 2 2 33252 34177
0 11727 7 3 2 22552 28581
0 11728 5 2 1 35609
0 11729 7 2 2 24704 25605
0 11730 7 1 2 35610 35614
0 11731 7 1 2 35607 11730
0 11732 5 1 1 11731
0 11733 7 1 2 35602 11732
0 11734 5 1 1 11733
0 11735 7 1 2 27184 11734
0 11736 5 1 1 11735
0 11737 7 2 2 25500 27455
0 11738 5 1 1 35616
0 11739 7 3 2 23660 35408
0 11740 5 3 1 35618
0 11741 7 1 2 35617 35619
0 11742 5 1 1 11741
0 11743 7 1 2 11736 11742
0 11744 5 1 1 11743
0 11745 7 1 2 24958 11744
0 11746 5 1 1 11745
0 11747 7 1 2 30539 35391
0 11748 7 1 2 33129 11747
0 11749 5 1 1 11748
0 11750 7 1 2 25501 31196
0 11751 7 1 2 35409 11750
0 11752 5 1 1 11751
0 11753 7 1 2 11749 11752
0 11754 5 1 1 11753
0 11755 7 1 2 23661 11754
0 11756 5 1 1 11755
0 11757 7 1 2 27517 29567
0 11758 5 2 1 11757
0 11759 7 1 2 35624 32221
0 11760 5 1 1 11759
0 11761 7 1 2 35374 11760
0 11762 5 1 1 11761
0 11763 7 1 2 23112 11762
0 11764 7 1 2 11756 11763
0 11765 7 1 2 11746 11764
0 11766 7 1 2 11725 11765
0 11767 5 1 1 11766
0 11768 7 3 2 25606 27518
0 11769 7 1 2 35626 35448
0 11770 5 1 1 11769
0 11771 7 1 2 35621 11770
0 11772 5 1 1 11771
0 11773 7 1 2 21933 11772
0 11774 5 1 1 11773
0 11775 7 1 2 26477 27065
0 11776 7 1 2 35608 11775
0 11777 5 1 1 11776
0 11778 7 1 2 35622 11777
0 11779 5 1 1 11778
0 11780 7 1 2 27185 11779
0 11781 5 1 1 11780
0 11782 7 1 2 35606 11781
0 11783 7 1 2 11774 11782
0 11784 5 1 1 11783
0 11785 7 1 2 24535 11784
0 11786 5 1 1 11785
0 11787 7 1 2 24705 34560
0 11788 7 1 2 34812 11787
0 11789 7 2 2 27905 11788
0 11790 5 1 1 35629
0 11791 7 1 2 35620 35565
0 11792 5 1 1 11791
0 11793 7 1 2 11790 11792
0 11794 7 1 2 11786 11793
0 11795 5 1 1 11794
0 11796 7 1 2 25502 11795
0 11797 5 1 1 11796
0 11798 7 6 2 29568 31313
0 11799 5 2 1 35631
0 11800 7 1 2 35637 35600
0 11801 5 1 1 11800
0 11802 7 1 2 25074 11801
0 11803 7 1 2 11797 11802
0 11804 5 1 1 11803
0 11805 7 1 2 11767 11804
0 11806 5 1 1 11805
0 11807 7 1 2 35304 35422
0 11808 5 1 1 11807
0 11809 7 1 2 35623 11808
0 11810 5 1 1 11809
0 11811 7 1 2 32535 11810
0 11812 5 1 1 11811
0 11813 7 1 2 22553 35630
0 11814 5 1 1 11813
0 11815 7 1 2 11812 11814
0 11816 5 1 1 11815
0 11817 7 1 2 25503 11816
0 11818 5 1 1 11817
0 11819 7 1 2 26208 11818
0 11820 7 1 2 11806 11819
0 11821 5 1 1 11820
0 11822 7 1 2 30303 35410
0 11823 7 1 2 32767 11822
0 11824 5 1 1 11823
0 11825 7 1 2 26225 11824
0 11826 5 1 1 11825
0 11827 7 1 2 26133 34583
0 11828 7 1 2 11826 11827
0 11829 7 1 2 11821 11828
0 11830 5 1 1 11829
0 11831 7 1 2 28362 33992
0 11832 5 1 1 11831
0 11833 7 1 2 29758 34106
0 11834 5 1 1 11833
0 11835 7 1 2 11832 11834
0 11836 5 1 1 11835
0 11837 7 1 2 23113 11836
0 11838 5 1 1 11837
0 11839 7 1 2 33967 32713
0 11840 5 1 1 11839
0 11841 7 1 2 11838 11840
0 11842 5 1 1 11841
0 11843 7 1 2 21934 11842
0 11844 5 1 1 11843
0 11845 7 1 2 29981 33968
0 11846 7 1 2 30905 11845
0 11847 5 1 1 11846
0 11848 7 1 2 34119 11847
0 11849 5 1 1 11848
0 11850 7 1 2 31384 32589
0 11851 7 1 2 11849 11850
0 11852 5 1 1 11851
0 11853 7 1 2 23980 33969
0 11854 5 1 1 11853
0 11855 7 1 2 34120 11854
0 11856 5 1 1 11855
0 11857 7 1 2 32755 11856
0 11858 5 1 1 11857
0 11859 7 1 2 28558 34659
0 11860 5 2 1 11859
0 11861 7 1 2 22554 29907
0 11862 7 1 2 31504 11861
0 11863 5 1 1 11862
0 11864 7 1 2 35639 11863
0 11865 5 1 1 11864
0 11866 7 1 2 34107 11865
0 11867 5 1 1 11866
0 11868 7 1 2 11858 11867
0 11869 7 1 2 11852 11868
0 11870 7 1 2 11844 11869
0 11871 5 1 1 11870
0 11872 7 1 2 35392 32092
0 11873 5 1 1 11872
0 11874 7 1 2 33393 35442
0 11875 5 1 1 11874
0 11876 7 1 2 11873 11875
0 11877 5 1 1 11876
0 11878 7 1 2 22403 11877
0 11879 5 1 1 11878
0 11880 7 1 2 25876 35402
0 11881 5 1 1 11880
0 11882 7 1 2 11879 11881
0 11883 5 1 1 11882
0 11884 7 1 2 28677 11883
0 11885 7 1 2 11871 11884
0 11886 5 1 1 11885
0 11887 7 1 2 23759 11886
0 11888 7 1 2 11830 11887
0 11889 7 1 2 11709 11888
0 11890 5 1 1 11889
0 11891 7 1 2 26325 11890
0 11892 7 1 2 11609 11891
0 11893 5 1 1 11892
0 11894 7 1 2 11360 11893
0 11895 7 1 2 10908 11894
0 11896 7 1 2 10361 11895
0 11897 7 1 2 9903 11896
0 11898 7 1 2 9085 11897
0 11899 7 1 2 8372 11898
0 11900 7 1 2 7313 11899
0 11901 7 1 2 6893 11900
0 11902 5 1 1 11901
0 11903 7 1 2 252 26681
0 11904 7 1 2 11902 11903
0 11905 5 1 1 11904
0 11906 7 1 2 25075 34032
0 11907 5 1 1 11906
0 11908 7 1 2 3561 11907
0 11909 5 1 1 11908
0 11910 7 1 2 22555 11909
0 11911 5 2 1 11910
0 11912 7 1 2 25076 31403
0 11913 5 1 1 11912
0 11914 7 2 2 35641 11913
0 11915 5 2 1 35643
0 11916 7 1 2 30174 35645
0 11917 5 1 1 11916
0 11918 7 1 2 29978 31386
0 11919 5 1 1 11918
0 11920 7 1 2 11917 11919
0 11921 5 1 1 11920
0 11922 7 1 2 24616 11921
0 11923 5 1 1 11922
0 11924 7 1 2 27456 29148
0 11925 5 1 1 11924
0 11926 7 1 2 30460 11925
0 11927 5 2 1 11926
0 11928 7 1 2 24959 35647
0 11929 5 1 1 11928
0 11930 7 1 2 30442 11929
0 11931 5 1 1 11930
0 11932 7 1 2 24617 11931
0 11933 5 1 1 11932
0 11934 7 1 2 23981 29908
0 11935 5 1 1 11934
0 11936 7 1 2 5847 11935
0 11937 5 1 1 11936
0 11938 7 1 2 22664 26389
0 11939 7 1 2 11937 11938
0 11940 5 1 1 11939
0 11941 7 1 2 25171 11940
0 11942 7 1 2 11933 11941
0 11943 5 1 1 11942
0 11944 7 1 2 29016 29702
0 11945 5 1 1 11944
0 11946 7 1 2 29116 31408
0 11947 5 1 1 11946
0 11948 7 1 2 33489 11947
0 11949 7 1 2 11945 11948
0 11950 5 1 1 11949
0 11951 7 1 2 23211 11950
0 11952 5 1 1 11951
0 11953 7 1 2 23303 11952
0 11954 7 1 2 11943 11953
0 11955 5 1 1 11954
0 11956 7 1 2 30153 31389
0 11957 5 1 1 11956
0 11958 7 1 2 26885 30199
0 11959 5 1 1 11958
0 11960 7 1 2 11957 11959
0 11961 5 1 1 11960
0 11962 7 1 2 24536 11961
0 11963 5 1 1 11962
0 11964 7 6 2 23982 29389
0 11965 5 1 1 35649
0 11966 7 1 2 30187 35650
0 11967 5 1 1 11966
0 11968 7 1 2 11963 11967
0 11969 7 1 2 11955 11968
0 11970 5 1 1 11969
0 11971 7 1 2 22062 11970
0 11972 5 1 1 11971
0 11973 7 1 2 21828 29665
0 11974 5 1 1 11973
0 11975 7 2 2 30899 11974
0 11976 7 1 2 32104 35655
0 11977 5 1 1 11976
0 11978 7 1 2 23212 29697
0 11979 5 1 1 11978
0 11980 7 1 2 11977 11979
0 11981 5 1 1 11980
0 11982 7 1 2 29090 30223
0 11983 7 1 2 11981 11982
0 11984 5 1 1 11983
0 11985 7 1 2 11972 11984
0 11986 7 1 2 11923 11985
0 11987 5 1 1 11986
0 11988 7 1 2 22759 11987
0 11989 5 1 1 11988
0 11990 7 2 2 26307 35632
0 11991 7 1 2 30320 32167
0 11992 7 1 2 35657 11991
0 11993 5 1 1 11992
0 11994 7 1 2 11989 11993
0 11995 5 1 1 11994
0 11996 7 1 2 23371 11995
0 11997 5 1 1 11996
0 11998 7 1 2 28085 32170
0 11999 7 1 2 35633 11998
0 12000 5 1 1 11999
0 12001 7 1 2 11997 12000
0 12002 5 1 1 12001
0 12003 7 1 2 25678 32620
0 12004 7 1 2 12002 12003
0 12005 5 1 1 12004
0 12006 7 1 2 25337 29673
0 12007 5 1 1 12006
0 12008 7 1 2 30765 31647
0 12009 5 1 1 12008
0 12010 7 1 2 30443 12009
0 12011 5 5 1 12010
0 12012 7 1 2 23372 31277
0 12013 7 1 2 35659 12012
0 12014 5 1 1 12013
0 12015 7 1 2 12007 12014
0 12016 5 1 1 12015
0 12017 7 1 2 26731 35615
0 12018 7 1 2 27845 12017
0 12019 7 1 2 12016 12018
0 12020 5 1 1 12019
0 12021 7 1 2 12005 12020
0 12022 5 1 1 12021
0 12023 7 1 2 23448 12022
0 12024 5 1 1 12023
0 12025 7 2 2 27408 27972
0 12026 7 2 2 26437 30091
0 12027 7 4 2 24706 22933
0 12028 7 1 2 35668 35103
0 12029 7 1 2 35666 12028
0 12030 7 1 2 35664 12029
0 12031 5 1 1 12030
0 12032 7 1 2 12024 12031
0 12033 5 1 1 12032
0 12034 7 1 2 33363 12033
0 12035 5 1 1 12034
0 12036 7 1 2 27850 10711
0 12037 5 1 1 12036
0 12038 7 1 2 28761 12037
0 12039 5 1 1 12038
0 12040 7 1 2 25941 30532
0 12041 5 1 1 12040
0 12042 7 1 2 4814 12041
0 12043 5 1 1 12042
0 12044 7 2 2 23760 12043
0 12045 7 1 2 22556 35672
0 12046 5 1 1 12045
0 12047 7 1 2 12039 12046
0 12048 5 1 1 12047
0 12049 7 1 2 29962 12048
0 12050 5 1 1 12049
0 12051 7 1 2 30568 35004
0 12052 7 1 2 28041 12051
0 12053 7 1 2 31412 12052
0 12054 5 1 1 12053
0 12055 7 1 2 12050 12054
0 12056 5 1 1 12055
0 12057 7 1 2 22063 31711
0 12058 7 1 2 30235 12057
0 12059 7 1 2 34053 12058
0 12060 7 1 2 12056 12059
0 12061 5 1 1 12060
0 12062 7 1 2 12035 12061
0 12063 5 1 1 12062
0 12064 7 1 2 23547 12063
0 12065 5 1 1 12064
0 12066 7 2 2 24758 29874
0 12067 7 1 2 35314 35674
0 12068 5 1 1 12067
0 12069 7 2 2 34571 33758
0 12070 7 1 2 24707 35676
0 12071 5 1 1 12070
0 12072 7 1 2 12068 12071
0 12073 5 2 1 12072
0 12074 7 1 2 35673 35678
0 12075 5 1 1 12074
0 12076 7 4 2 23373 27594
0 12077 7 4 2 26119 33314
0 12078 7 3 2 25077 23449
0 12079 7 1 2 35688 32168
0 12080 7 1 2 35684 12079
0 12081 7 1 2 35680 12080
0 12082 5 1 1 12081
0 12083 7 1 2 12075 12082
0 12084 5 1 1 12083
0 12085 7 1 2 29650 12084
0 12086 5 1 1 12085
0 12087 7 1 2 22404 28757
0 12088 7 1 2 28731 12087
0 12089 7 1 2 35679 12088
0 12090 7 1 2 34808 12089
0 12091 5 1 1 12090
0 12092 7 1 2 12086 12091
0 12093 5 1 1 12092
0 12094 7 4 2 25172 34556
0 12095 7 1 2 31132 35691
0 12096 7 1 2 12093 12095
0 12097 5 1 1 12096
0 12098 7 1 2 22210 12097
0 12099 7 1 2 12065 12098
0 12100 5 1 1 12099
0 12101 7 4 2 23761 33592
0 12102 7 2 2 26732 30066
0 12103 7 1 2 24095 35699
0 12104 5 1 1 12103
0 12105 7 3 2 23304 30349
0 12106 7 1 2 31314 35701
0 12107 5 1 1 12106
0 12108 7 1 2 12104 12107
0 12109 5 3 1 12108
0 12110 7 1 2 35695 35704
0 12111 5 1 1 12110
0 12112 7 1 2 24096 29703
0 12113 5 2 1 12112
0 12114 7 1 2 30418 35707
0 12115 5 1 1 12114
0 12116 7 1 2 23213 31413
0 12117 5 1 1 12116
0 12118 7 2 2 28494 12117
0 12119 5 1 1 35709
0 12120 7 1 2 24097 35710
0 12121 5 1 1 12120
0 12122 7 1 2 25258 32256
0 12123 7 1 2 12121 12122
0 12124 7 1 2 33196 12123
0 12125 5 1 1 12124
0 12126 7 1 2 12115 12125
0 12127 5 1 1 12126
0 12128 7 1 2 23114 12127
0 12129 5 1 1 12128
0 12130 7 2 2 23214 28429
0 12131 7 1 2 29294 30321
0 12132 7 1 2 35711 12131
0 12133 5 1 1 12132
0 12134 7 1 2 12129 12133
0 12135 5 1 1 12134
0 12136 7 1 2 24537 12135
0 12137 5 1 1 12136
0 12138 7 1 2 29797 30465
0 12139 5 1 1 12138
0 12140 7 1 2 30444 12139
0 12141 5 2 1 12140
0 12142 7 2 2 26698 35713
0 12143 5 1 1 35715
0 12144 7 3 2 24479 22557
0 12145 5 1 1 35717
0 12146 7 1 2 23115 35718
0 12147 5 1 1 12146
0 12148 7 1 2 11965 12147
0 12149 5 1 1 12148
0 12150 7 1 2 23844 12149
0 12151 5 1 1 12150
0 12152 7 2 2 23983 29010
0 12153 7 1 2 30042 35720
0 12154 5 1 1 12153
0 12155 7 2 2 12151 12154
0 12156 5 1 1 35722
0 12157 7 1 2 30175 12156
0 12158 5 1 1 12157
0 12159 7 1 2 12143 12158
0 12160 5 1 1 12159
0 12161 7 1 2 24098 12160
0 12162 5 1 1 12161
0 12163 7 1 2 26706 31010
0 12164 7 1 2 32730 12163
0 12165 5 1 1 12164
0 12166 7 1 2 12162 12165
0 12167 7 1 2 12137 12166
0 12168 5 1 1 12167
0 12169 7 1 2 22665 12168
0 12170 5 1 1 12169
0 12171 7 1 2 24480 35651
0 12172 5 1 1 12171
0 12173 7 1 2 31021 12172
0 12174 5 1 1 12173
0 12175 7 1 2 23845 12174
0 12176 5 1 1 12175
0 12177 7 1 2 29530 3551
0 12178 5 2 1 12177
0 12179 7 1 2 28984 35724
0 12180 5 1 1 12179
0 12181 7 1 2 12176 12180
0 12182 5 1 1 12181
0 12183 7 1 2 24099 12182
0 12184 5 1 1 12183
0 12185 7 1 2 30061 32214
0 12186 5 1 1 12185
0 12187 7 1 2 12184 12186
0 12188 5 1 1 12187
0 12189 7 1 2 25173 12188
0 12190 5 1 1 12189
0 12191 7 1 2 23846 29011
0 12192 7 1 2 30942 12191
0 12193 7 1 2 29943 12192
0 12194 5 1 1 12193
0 12195 7 1 2 30040 30557
0 12196 5 1 1 12195
0 12197 7 1 2 35721 12196
0 12198 5 1 1 12197
0 12199 7 1 2 29043 12198
0 12200 7 2 2 12194 12199
0 12201 5 2 1 35726
0 12202 7 1 2 22064 35727
0 12203 5 1 1 12202
0 12204 7 2 2 29534 35625
0 12205 5 2 1 35730
0 12206 7 1 2 25078 35731
0 12207 5 1 1 12206
0 12208 7 1 2 1805 12207
0 12209 5 2 1 12208
0 12210 7 1 2 24100 35734
0 12211 5 1 1 12210
0 12212 7 1 2 23215 12211
0 12213 7 1 2 12203 12212
0 12214 5 1 1 12213
0 12215 7 1 2 12190 12214
0 12216 5 1 1 12215
0 12217 7 1 2 26989 12216
0 12218 5 1 1 12217
0 12219 7 1 2 12170 12218
0 12220 5 1 1 12219
0 12221 7 1 2 27595 33904
0 12222 7 1 2 12220 12221
0 12223 5 1 1 12222
0 12224 7 1 2 12111 12223
0 12225 5 1 1 12224
0 12226 7 1 2 24708 12225
0 12227 5 1 1 12226
0 12228 7 1 2 29185 33432
0 12229 7 2 2 33710 12228
0 12230 7 1 2 32114 35736
0 12231 5 1 1 12230
0 12232 7 2 2 29173 33315
0 12233 7 2 2 29305 35432
0 12234 7 1 2 35738 35740
0 12235 5 1 1 12234
0 12236 7 1 2 29117 35696
0 12237 5 1 1 12236
0 12238 7 1 2 12235 12237
0 12239 5 1 1 12238
0 12240 7 1 2 30841 12239
0 12241 5 1 1 12240
0 12242 7 1 2 12231 12241
0 12243 5 1 1 12242
0 12244 7 1 2 31331 34770
0 12245 7 1 2 12243 12244
0 12246 5 1 1 12245
0 12247 7 1 2 12227 12246
0 12248 5 1 1 12247
0 12249 7 1 2 23374 12248
0 12250 5 1 1 12249
0 12251 7 1 2 30058 35697
0 12252 5 1 1 12251
0 12253 7 1 2 34782 34756
0 12254 7 1 2 35741 12253
0 12255 5 1 1 12254
0 12256 7 1 2 12252 12255
0 12257 5 1 1 12256
0 12258 7 1 2 23984 12257
0 12259 5 1 1 12258
0 12260 7 1 2 29744 35737
0 12261 5 1 1 12260
0 12262 7 1 2 12259 12261
0 12263 5 1 1 12262
0 12264 7 1 2 35209 33894
0 12265 7 1 2 12263 12264
0 12266 5 1 1 12265
0 12267 7 1 2 12250 12266
0 12268 5 1 1 12267
0 12269 7 1 2 25409 12268
0 12270 5 1 1 12269
0 12271 7 1 2 31072 32241
0 12272 5 1 1 12271
0 12273 7 1 2 23216 35660
0 12274 5 1 1 12273
0 12275 7 1 2 34651 12274
0 12276 5 1 1 12275
0 12277 7 1 2 31270 12276
0 12278 5 1 1 12277
0 12279 7 1 2 12272 12278
0 12280 5 1 1 12279
0 12281 7 1 2 23305 12280
0 12282 5 2 1 12281
0 12283 7 7 2 24101 25174
0 12284 5 1 1 35744
0 12285 7 1 2 30461 35745
0 12286 5 1 1 12285
0 12287 7 1 2 32414 12286
0 12288 5 1 1 12287
0 12289 7 1 2 24481 12288
0 12290 5 1 1 12289
0 12291 7 1 2 12290 34679
0 12292 5 1 1 12291
0 12293 7 1 2 23847 12292
0 12294 5 1 1 12293
0 12295 7 1 2 31102 35746
0 12296 5 2 1 12295
0 12297 7 1 2 12294 35751
0 12298 5 1 1 12297
0 12299 7 1 2 25259 12298
0 12300 5 1 1 12299
0 12301 7 1 2 35742 12300
0 12302 5 1 1 12301
0 12303 7 1 2 25338 12302
0 12304 5 1 1 12303
0 12305 7 2 2 25825 32457
0 12306 7 1 2 31278 35753
0 12307 5 1 1 12306
0 12308 7 1 2 12304 12307
0 12309 5 1 1 12308
0 12310 7 1 2 12309 35698
0 12311 5 1 1 12310
0 12312 7 2 2 25679 27360
0 12313 7 5 2 23116 25260
0 12314 7 1 2 25339 27365
0 12315 7 1 2 35757 12314
0 12316 7 1 2 29310 34061
0 12317 7 1 2 12315 12316
0 12318 7 1 2 35755 12317
0 12319 5 1 1 12318
0 12320 7 1 2 12311 12319
0 12321 5 1 1 12320
0 12322 7 1 2 22760 12321
0 12323 5 1 1 12322
0 12324 7 1 2 26450 33988
0 12325 7 1 2 34477 35056
0 12326 7 1 2 12324 12325
0 12327 7 1 2 29434 31367
0 12328 7 1 2 35418 12327
0 12329 7 1 2 12326 12328
0 12330 5 1 1 12329
0 12331 7 1 2 12323 12330
0 12332 5 1 1 12331
0 12333 7 1 2 23450 12332
0 12334 5 1 1 12333
0 12335 7 1 2 24222 12334
0 12336 7 1 2 12270 12335
0 12337 5 1 1 12336
0 12338 7 1 2 22141 12337
0 12339 7 1 2 12100 12338
0 12340 5 1 1 12339
0 12341 7 3 2 27409 32478
0 12342 7 2 2 26329 35762
0 12343 7 2 2 22934 35765
0 12344 7 2 2 33583 35477
0 12345 7 3 2 30025 31294
0 12346 7 1 2 35769 35771
0 12347 7 1 2 35767 12346
0 12348 5 1 1 12347
0 12349 7 1 2 12340 12348
0 12350 5 1 1 12349
0 12351 7 1 2 28830 12350
0 12352 5 1 1 12351
0 12353 7 2 2 22142 25680
0 12354 7 3 2 23662 33316
0 12355 7 2 2 27690 35776
0 12356 7 1 2 27519 35779
0 12357 5 1 1 12356
0 12358 7 1 2 27143 34235
0 12359 5 1 1 12358
0 12360 7 2 2 25942 27520
0 12361 7 1 2 23663 35781
0 12362 5 1 1 12361
0 12363 7 1 2 12359 12362
0 12364 5 1 1 12363
0 12365 7 1 2 33734 12364
0 12366 5 1 1 12365
0 12367 7 1 2 12357 12366
0 12368 5 1 1 12367
0 12369 7 2 2 23015 12368
0 12370 7 3 2 30783 31628
0 12371 7 1 2 25175 35785
0 12372 5 2 1 12371
0 12373 7 7 2 25410 27962
0 12374 7 1 2 27978 35790
0 12375 5 2 1 12374
0 12376 7 1 2 35788 35797
0 12377 5 1 1 12376
0 12378 7 1 2 35783 12377
0 12379 5 1 1 12378
0 12380 7 2 2 25943 33735
0 12381 5 1 1 35799
0 12382 7 3 2 22267 27675
0 12383 7 3 2 35357 35801
0 12384 5 2 1 35804
0 12385 7 1 2 12381 35807
0 12386 5 5 1 12385
0 12387 7 2 2 23451 32780
0 12388 7 1 2 30123 35814
0 12389 5 1 1 12388
0 12390 7 1 2 35798 12389
0 12391 5 1 1 12390
0 12392 7 1 2 29197 12391
0 12393 7 1 2 35809 12392
0 12394 5 1 1 12393
0 12395 7 1 2 12379 12394
0 12396 5 1 1 12395
0 12397 7 1 2 23548 12396
0 12398 5 1 1 12397
0 12399 7 2 2 27350 34217
0 12400 7 1 2 22211 26733
0 12401 7 1 2 27332 12400
0 12402 7 1 2 28311 12401
0 12403 7 1 2 35816 12402
0 12404 5 1 1 12403
0 12405 7 1 2 12398 12404
0 12406 5 1 1 12405
0 12407 7 1 2 35137 12406
0 12408 5 1 1 12407
0 12409 7 2 2 26734 34080
0 12410 7 1 2 34329 35818
0 12411 5 1 1 12410
0 12412 7 3 2 23217 28161
0 12413 7 1 2 34904 33953
0 12414 7 1 2 35820 12413
0 12415 5 1 1 12414
0 12416 7 1 2 12411 12415
0 12417 5 1 1 12416
0 12418 7 1 2 24398 12417
0 12419 5 1 1 12418
0 12420 7 1 2 25176 34507
0 12421 7 1 2 35203 12420
0 12422 7 1 2 34566 12421
0 12423 5 1 1 12422
0 12424 7 1 2 12419 12423
0 12425 5 1 1 12424
0 12426 7 1 2 28831 12425
0 12427 5 1 1 12426
0 12428 7 5 2 26308 33174
0 12429 5 2 1 35823
0 12430 7 1 2 35824 34367
0 12431 5 1 1 12430
0 12432 7 1 2 35821 34895
0 12433 5 1 1 12432
0 12434 7 1 2 12431 12433
0 12435 5 1 1 12434
0 12436 7 1 2 31825 12435
0 12437 5 1 1 12436
0 12438 7 1 2 12427 12437
0 12439 5 1 1 12438
0 12440 7 3 2 31849 33698
0 12441 7 2 2 28758 35830
0 12442 7 1 2 23452 35833
0 12443 7 1 2 12439 12442
0 12444 5 1 1 12443
0 12445 7 1 2 12408 12444
0 12446 5 1 1 12445
0 12447 7 1 2 35774 12446
0 12448 5 1 1 12447
0 12449 7 1 2 23848 34683
0 12450 5 1 1 12449
0 12451 7 1 2 35752 12450
0 12452 5 1 1 12451
0 12453 7 1 2 25261 12452
0 12454 5 1 1 12453
0 12455 7 1 2 35743 12454
0 12456 5 3 1 12455
0 12457 7 1 2 22212 35835
0 12458 5 1 1 12457
0 12459 7 2 2 35661 34239
0 12460 5 1 1 35838
0 12461 7 1 2 30124 35839
0 12462 5 1 1 12461
0 12463 7 1 2 12458 12462
0 12464 5 1 1 12463
0 12465 7 1 2 23453 12464
0 12466 5 1 1 12465
0 12467 7 1 2 26264 34868
0 12468 7 1 2 30012 12467
0 12469 5 1 1 12468
0 12470 7 1 2 12466 12469
0 12471 5 1 1 12470
0 12472 7 1 2 22143 12471
0 12473 5 1 1 12472
0 12474 7 2 2 28881 34269
0 12475 5 1 1 35840
0 12476 7 1 2 25177 35841
0 12477 5 1 1 12476
0 12478 7 1 2 26396 26292
0 12479 5 2 1 12478
0 12480 7 1 2 34826 35842
0 12481 5 1 1 12480
0 12482 7 1 2 12477 12481
0 12483 5 1 1 12482
0 12484 7 1 2 29674 12483
0 12485 5 1 1 12484
0 12486 7 1 2 12473 12485
0 12487 5 1 1 12486
0 12488 7 1 2 33565 12487
0 12489 5 1 1 12488
0 12490 7 1 2 21829 30704
0 12491 5 1 1 12490
0 12492 7 1 2 31745 12491
0 12493 5 1 1 12492
0 12494 7 1 2 29508 12493
0 12495 5 1 1 12494
0 12496 7 1 2 23117 35164
0 12497 5 1 1 12496
0 12498 7 1 2 12495 12497
0 12499 5 1 1 12498
0 12500 7 1 2 23306 12499
0 12501 5 2 1 12500
0 12502 7 1 2 29824 2972
0 12503 5 1 1 12502
0 12504 7 1 2 5032 12503
0 12505 5 1 1 12504
0 12506 7 1 2 25262 12505
0 12507 5 1 1 12506
0 12508 7 1 2 35844 12507
0 12509 5 1 1 12508
0 12510 7 1 2 22213 12509
0 12511 5 1 1 12510
0 12512 7 1 2 12460 12511
0 12513 5 1 1 12512
0 12514 7 1 2 22144 12513
0 12515 5 1 1 12514
0 12516 7 2 2 24102 29811
0 12517 7 1 2 27020 32781
0 12518 7 1 2 35846 12517
0 12519 5 1 1 12518
0 12520 7 1 2 12515 12519
0 12521 5 1 1 12520
0 12522 7 1 2 23454 12521
0 12523 5 1 1 12522
0 12524 7 1 2 30986 31449
0 12525 5 1 1 12524
0 12526 7 1 2 22145 12525
0 12527 5 1 1 12526
0 12528 7 1 2 30200 32259
0 12529 5 1 1 12528
0 12530 7 1 2 12527 12529
0 12531 5 1 1 12530
0 12532 7 1 2 34270 12531
0 12533 5 1 1 12532
0 12534 7 3 2 24223 31044
0 12535 7 1 2 31507 35848
0 12536 5 1 1 12535
0 12537 7 1 2 12533 12536
0 12538 5 1 1 12537
0 12539 7 1 2 29828 12538
0 12540 5 1 1 12539
0 12541 7 9 2 24161 24224
0 12542 7 2 2 31045 35851
0 12543 7 1 2 35860 35847
0 12544 5 1 1 12543
0 12545 7 1 2 25178 12544
0 12546 7 1 2 12540 12545
0 12547 7 1 2 12523 12546
0 12548 5 1 1 12547
0 12549 7 11 2 22146 22214
0 12550 7 2 2 23455 35862
0 12551 7 1 2 22666 31453
0 12552 5 1 1 12551
0 12553 7 1 2 29933 29615
0 12554 7 1 2 35165 12553
0 12555 5 1 1 12554
0 12556 7 1 2 12552 12555
0 12557 5 1 1 12556
0 12558 7 1 2 23307 12557
0 12559 5 2 1 12558
0 12560 7 2 2 1908 31425
0 12561 5 1 1 35877
0 12562 7 1 2 25263 35878
0 12563 5 1 1 12562
0 12564 7 1 2 29934 30766
0 12565 5 1 1 12564
0 12566 7 1 2 23308 31707
0 12567 7 1 2 12565 12566
0 12568 5 1 1 12567
0 12569 7 1 2 25079 12568
0 12570 7 1 2 12563 12569
0 12571 5 1 1 12570
0 12572 7 1 2 35875 12571
0 12573 5 2 1 12572
0 12574 7 1 2 35873 35879
0 12575 5 1 1 12574
0 12576 7 1 2 29675 35758
0 12577 5 1 1 12576
0 12578 7 1 2 23309 27061
0 12579 5 1 1 12578
0 12580 7 1 2 12577 12579
0 12581 5 1 1 12580
0 12582 7 1 2 24162 12581
0 12583 5 1 1 12582
0 12584 7 2 2 27144 31462
0 12585 5 1 1 35881
0 12586 7 1 2 31197 12585
0 12587 5 1 1 12586
0 12588 7 1 2 28769 12587
0 12589 5 1 1 12588
0 12590 7 1 2 31590 34663
0 12591 5 1 1 12590
0 12592 7 1 2 12589 12591
0 12593 5 1 1 12592
0 12594 7 1 2 31571 12593
0 12595 5 1 1 12594
0 12596 7 1 2 12583 12595
0 12597 5 1 1 12596
0 12598 7 1 2 23016 12597
0 12599 5 1 1 12598
0 12600 7 1 2 28985 30872
0 12601 5 1 1 12600
0 12602 7 1 2 24163 23118
0 12603 5 1 1 12602
0 12604 7 1 2 27521 12603
0 12605 7 1 2 30462 12604
0 12606 5 1 1 12605
0 12607 7 1 2 12601 12606
0 12608 5 1 1 12607
0 12609 7 1 2 34251 12608
0 12610 5 1 1 12609
0 12611 7 1 2 12599 12610
0 12612 5 2 1 12611
0 12613 7 1 2 34849 35883
0 12614 5 1 1 12613
0 12615 7 1 2 23218 12614
0 12616 7 1 2 12575 12615
0 12617 5 1 1 12616
0 12618 7 1 2 34948 12617
0 12619 7 1 2 12548 12618
0 12620 5 1 1 12619
0 12621 7 1 2 12489 12620
0 12622 5 1 1 12621
0 12623 7 1 2 23664 12622
0 12624 5 1 1 12623
0 12625 7 1 2 25264 35235
0 12626 7 2 2 34189 12625
0 12627 7 1 2 31629 35885
0 12628 5 1 1 12627
0 12629 7 3 2 33970 34508
0 12630 7 1 2 26082 30498
0 12631 7 1 2 35887 12630
0 12632 5 1 1 12631
0 12633 7 1 2 12628 12632
0 12634 5 1 1 12633
0 12635 7 1 2 30070 12634
0 12636 5 1 1 12635
0 12637 7 1 2 23017 29150
0 12638 5 1 1 12637
0 12639 7 1 2 31587 31644
0 12640 5 1 1 12639
0 12641 7 1 2 28092 12640
0 12642 7 1 2 12638 12641
0 12643 5 1 1 12642
0 12644 7 1 2 25179 12643
0 12645 5 1 1 12644
0 12646 7 1 2 26981 27145
0 12647 5 1 1 12646
0 12648 7 1 2 12645 12647
0 12649 5 1 1 12648
0 12650 7 1 2 34929 35815
0 12651 7 1 2 12649 12650
0 12652 5 1 1 12651
0 12653 7 1 2 12636 12652
0 12654 5 1 1 12653
0 12655 7 1 2 24103 12654
0 12656 5 1 1 12655
0 12657 7 2 2 30718 33736
0 12658 7 1 2 35167 35890
0 12659 5 1 1 12658
0 12660 7 1 2 23219 34660
0 12661 5 1 1 12660
0 12662 7 1 2 30597 12661
0 12663 5 1 1 12662
0 12664 7 1 2 34930 12663
0 12665 5 1 1 12664
0 12666 7 2 2 25504 33443
0 12667 7 2 2 24286 22485
0 12668 7 1 2 21830 24340
0 12669 7 1 2 35894 12668
0 12670 7 2 2 35892 12669
0 12671 7 1 2 26970 35896
0 12672 5 1 1 12671
0 12673 7 1 2 12665 12672
0 12674 5 1 1 12673
0 12675 7 1 2 29569 12674
0 12676 5 1 1 12675
0 12677 7 2 2 30338 33364
0 12678 7 1 2 30799 35898
0 12679 5 1 1 12678
0 12680 7 1 2 30598 32143
0 12681 5 1 1 12680
0 12682 7 1 2 35891 12681
0 12683 5 1 1 12682
0 12684 7 1 2 12679 12683
0 12685 5 1 1 12684
0 12686 7 1 2 29509 12685
0 12687 5 1 1 12686
0 12688 7 1 2 12676 12687
0 12689 5 1 1 12688
0 12690 7 1 2 22065 12689
0 12691 5 1 1 12690
0 12692 7 1 2 12659 12691
0 12693 5 1 1 12692
0 12694 7 1 2 23310 12693
0 12695 5 1 1 12694
0 12696 7 1 2 31089 34931
0 12697 5 1 1 12696
0 12698 7 1 2 12695 12697
0 12699 5 1 1 12698
0 12700 7 1 2 22215 12699
0 12701 5 1 1 12700
0 12702 7 1 2 24960 33672
0 12703 5 1 1 12702
0 12704 7 1 2 28832 30719
0 12705 5 1 1 12704
0 12706 7 1 2 26083 33495
0 12707 5 1 1 12706
0 12708 7 1 2 12705 12707
0 12709 5 1 1 12708
0 12710 7 1 2 33365 12709
0 12711 5 1 1 12710
0 12712 7 1 2 12703 12711
0 12713 5 1 1 12712
0 12714 7 1 2 31749 31547
0 12715 7 2 2 34810 12714
0 12716 7 1 2 12713 35900
0 12717 5 1 1 12716
0 12718 7 1 2 12701 12717
0 12719 5 1 1 12718
0 12720 7 1 2 23456 12719
0 12721 5 1 1 12720
0 12722 7 1 2 12656 12721
0 12723 5 1 1 12722
0 12724 7 1 2 26607 12723
0 12725 5 1 1 12724
0 12726 7 1 2 12624 12725
0 12727 5 1 1 12726
0 12728 7 1 2 26209 12727
0 12729 5 1 1 12728
0 12730 7 4 2 22869 30720
0 12731 5 2 1 35902
0 12732 7 1 2 25080 28582
0 12733 5 1 1 12732
0 12734 7 1 2 35906 12733
0 12735 5 1 1 12734
0 12736 7 1 2 22330 12735
0 12737 5 1 1 12736
0 12738 7 1 2 28709 33496
0 12739 5 1 1 12738
0 12740 7 1 2 12737 12739
0 12741 5 1 1 12740
0 12742 7 1 2 35901 12741
0 12743 5 1 1 12742
0 12744 7 1 2 30524 35705
0 12745 5 1 1 12744
0 12746 7 1 2 30540 35836
0 12747 5 1 1 12746
0 12748 7 1 2 12745 12747
0 12749 5 1 1 12748
0 12750 7 1 2 22216 12749
0 12751 5 1 1 12750
0 12752 7 1 2 12743 12751
0 12753 5 1 1 12752
0 12754 7 1 2 23457 12753
0 12755 5 1 1 12754
0 12756 7 3 2 26265 30067
0 12757 7 2 2 35908 34869
0 12758 5 1 1 35911
0 12759 7 1 2 30525 35912
0 12760 5 1 1 12759
0 12761 7 1 2 12755 12760
0 12762 5 1 1 12761
0 12763 7 1 2 33317 12762
0 12764 5 1 1 12763
0 12765 7 1 2 34331 34632
0 12766 5 2 1 12765
0 12767 7 1 2 22217 35702
0 12768 5 1 1 12767
0 12769 7 1 2 35913 12768
0 12770 5 2 1 12769
0 12771 7 1 2 31315 35915
0 12772 5 1 1 12771
0 12773 7 1 2 31295 35700
0 12774 5 1 1 12773
0 12775 7 1 2 12772 12774
0 12776 5 1 1 12775
0 12777 7 1 2 23458 12776
0 12778 5 1 1 12777
0 12779 7 1 2 12758 12778
0 12780 5 1 1 12779
0 12781 7 1 2 33688 12780
0 12782 5 1 1 12781
0 12783 7 1 2 12764 12782
0 12784 5 1 1 12783
0 12785 7 1 2 22147 27562
0 12786 7 1 2 12784 12785
0 12787 5 1 1 12786
0 12788 7 1 2 12729 12787
0 12789 5 1 1 12788
0 12790 7 1 2 23762 12789
0 12791 5 1 1 12790
0 12792 7 1 2 12448 12791
0 12793 5 1 1 12792
0 12794 7 1 2 32971 12793
0 12795 5 1 1 12794
0 12796 7 4 2 22218 22558
0 12797 7 1 2 31498 33939
0 12798 7 1 2 35917 12797
0 12799 5 1 1 12798
0 12800 7 1 2 9148 12799
0 12801 5 1 1 12800
0 12802 7 1 2 27457 12801
0 12803 5 1 1 12802
0 12804 7 1 2 35849 32714
0 12805 5 1 1 12804
0 12806 7 1 2 12803 12805
0 12807 5 1 1 12806
0 12808 7 1 2 21935 12807
0 12809 5 1 1 12808
0 12810 7 1 2 22066 28464
0 12811 5 2 1 12810
0 12812 7 1 2 29091 35921
0 12813 5 1 1 12812
0 12814 7 1 2 33140 12813
0 12815 5 1 1 12814
0 12816 7 1 2 34827 12815
0 12817 5 1 1 12816
0 12818 7 1 2 12809 12817
0 12819 5 1 1 12818
0 12820 7 1 2 24961 12819
0 12821 5 1 1 12820
0 12822 7 1 2 29711 35759
0 12823 5 2 1 12822
0 12824 7 1 2 27146 35923
0 12825 5 1 1 12824
0 12826 7 2 2 22559 27007
0 12827 5 1 1 35925
0 12828 7 1 2 27186 12827
0 12829 5 1 1 12828
0 12830 7 1 2 30904 12829
0 12831 7 1 2 12825 12830
0 12832 5 1 1 12831
0 12833 7 1 2 30445 2533
0 12834 5 1 1 12833
0 12835 7 1 2 30427 31648
0 12836 7 1 2 12834 12835
0 12837 5 1 1 12836
0 12838 7 1 2 12832 12837
0 12839 5 1 1 12838
0 12840 7 1 2 34850 12839
0 12841 5 1 1 12840
0 12842 7 1 2 12821 12841
0 12843 5 1 1 12842
0 12844 7 1 2 32910 12843
0 12845 5 1 1 12844
0 12846 7 2 2 31171 31261
0 12847 5 1 1 35927
0 12848 7 1 2 27522 33175
0 12849 7 1 2 35138 12848
0 12850 7 1 2 35928 12849
0 12851 5 1 1 12850
0 12852 7 1 2 12845 12851
0 12853 5 1 1 12852
0 12854 7 1 2 27738 12853
0 12855 5 1 1 12854
0 12856 7 1 2 22067 28732
0 12857 7 5 2 23375 28273
0 12858 7 1 2 34271 35929
0 12859 7 1 2 12856 12858
0 12860 7 1 2 35662 12859
0 12861 5 1 1 12860
0 12862 7 1 2 12855 12861
0 12863 5 1 1 12862
0 12864 7 1 2 33515 12863
0 12865 5 1 1 12864
0 12866 7 2 2 32886 35663
0 12867 7 2 2 22405 22761
0 12868 7 2 2 33725 35936
0 12869 7 1 2 28729 34915
0 12870 7 1 2 32782 12869
0 12871 7 1 2 35938 12870
0 12872 7 1 2 35934 12871
0 12873 5 1 1 12872
0 12874 7 1 2 12865 12873
0 12875 5 1 1 12874
0 12876 7 1 2 25180 12875
0 12877 5 1 1 12876
0 12878 7 1 2 31585 31414
0 12879 5 1 1 12878
0 12880 7 1 2 3039 12879
0 12881 5 1 1 12880
0 12882 7 1 2 23119 12881
0 12883 5 1 1 12882
0 12884 7 1 2 27523 30576
0 12885 5 1 1 12884
0 12886 7 1 2 29841 12885
0 12887 5 2 1 12886
0 12888 7 2 2 25081 35940
0 12889 5 1 1 35942
0 12890 7 1 2 23985 35943
0 12891 5 1 1 12890
0 12892 7 1 2 12883 12891
0 12893 5 1 1 12892
0 12894 7 1 2 24104 12893
0 12895 5 1 1 12894
0 12896 7 1 2 28986 32215
0 12897 7 1 2 27351 12896
0 12898 5 1 1 12897
0 12899 7 1 2 12895 12898
0 12900 5 1 1 12899
0 12901 7 1 2 28017 34960
0 12902 7 1 2 30993 35495
0 12903 7 1 2 12901 12902
0 12904 7 1 2 12900 12903
0 12905 5 1 1 12904
0 12906 7 1 2 12877 12905
0 12907 5 1 1 12906
0 12908 7 1 2 22667 12907
0 12909 5 1 1 12908
0 12910 7 3 2 24618 25411
0 12911 7 1 2 23220 29570
0 12912 5 1 1 12911
0 12913 7 1 2 5299 12912
0 12914 5 1 1 12913
0 12915 7 1 2 27458 12914
0 12916 5 1 1 12915
0 12917 7 2 2 21936 24538
0 12918 7 1 2 28598 35947
0 12919 5 1 1 12918
0 12920 7 1 2 12916 12919
0 12921 5 1 1 12920
0 12922 7 1 2 34761 12921
0 12923 5 1 1 12922
0 12924 7 2 2 27352 31790
0 12925 7 1 2 29459 35949
0 12926 5 1 1 12925
0 12927 7 1 2 12923 12926
0 12928 5 1 1 12927
0 12929 7 1 2 23376 12928
0 12930 5 1 1 12929
0 12931 7 1 2 24709 26032
0 12932 7 1 2 30026 12931
0 12933 5 1 1 12932
0 12934 7 1 2 12930 12933
0 12935 5 1 1 12934
0 12936 7 1 2 35944 12935
0 12937 5 1 1 12936
0 12938 7 1 2 28459 35108
0 12939 7 1 2 31226 12938
0 12940 5 1 1 12939
0 12941 7 1 2 12937 12940
0 12942 5 1 1 12941
0 12943 7 1 2 23120 12942
0 12944 5 1 1 12943
0 12945 7 1 2 23221 35732
0 12946 5 1 1 12945
0 12947 7 1 2 28495 12946
0 12948 5 1 1 12947
0 12949 7 2 2 26575 34762
0 12950 7 1 2 27062 35951
0 12951 7 1 2 12948 12950
0 12952 5 1 1 12951
0 12953 7 1 2 12944 12952
0 12954 5 1 1 12953
0 12955 7 1 2 24105 12954
0 12956 5 1 1 12955
0 12957 7 2 2 34911 32237
0 12958 5 1 1 35953
0 12959 7 1 2 23222 35728
0 12960 5 1 1 12959
0 12961 7 1 2 12958 12960
0 12962 5 1 1 12961
0 12963 7 1 2 32519 35952
0 12964 7 1 2 12962 12963
0 12965 5 1 1 12964
0 12966 7 1 2 12956 12965
0 12967 5 1 1 12966
0 12968 7 3 2 24225 22870
0 12969 7 1 2 33366 35955
0 12970 7 1 2 30509 12969
0 12971 7 1 2 12967 12970
0 12972 5 1 1 12971
0 12973 7 1 2 12909 12972
0 12974 5 1 1 12973
0 12975 7 1 2 23665 12974
0 12976 5 1 1 12975
0 12977 7 4 2 24399 22762
0 12978 7 1 2 29875 35958
0 12979 7 1 2 33766 12978
0 12980 5 1 1 12979
0 12981 7 1 2 35229 32156
0 12982 7 1 2 35930 12981
0 12983 5 1 1 12982
0 12984 7 1 2 12980 12983
0 12985 5 1 1 12984
0 12986 7 1 2 29543 33647
0 12987 7 1 2 12985 12986
0 12988 5 1 1 12987
0 12989 7 2 2 25789 33880
0 12990 7 2 2 28913 35962
0 12991 7 2 2 33444 35964
0 12992 7 1 2 29769 33230
0 12993 7 1 2 35966 12992
0 12994 7 1 2 32282 12993
0 12995 5 1 1 12994
0 12996 7 1 2 12988 12995
0 12997 5 1 1 12996
0 12998 7 1 2 22560 12997
0 12999 5 1 1 12998
0 13000 7 1 2 27801 28890
0 13001 5 1 1 13000
0 13002 7 1 2 25082 32720
0 13003 5 1 1 13002
0 13004 7 1 2 24619 29767
0 13005 7 1 2 13003 13004
0 13006 5 1 1 13005
0 13007 7 1 2 13001 13006
0 13008 5 1 1 13007
0 13009 7 1 2 23986 13008
0 13010 5 1 1 13009
0 13011 7 1 2 30154 29897
0 13012 5 1 1 13011
0 13013 7 1 2 13010 13012
0 13014 5 1 1 13013
0 13015 7 1 2 28069 35109
0 13016 7 1 2 35967 13015
0 13017 7 1 2 13014 13016
0 13018 5 1 1 13017
0 13019 7 1 2 12999 13018
0 13020 5 1 1 13019
0 13021 7 1 2 25181 13020
0 13022 5 1 1 13021
0 13023 7 1 2 25083 31379
0 13024 5 1 1 13023
0 13025 7 1 2 29044 13024
0 13026 5 1 1 13025
0 13027 7 2 2 23377 32099
0 13028 7 2 2 22668 35968
0 13029 7 1 2 22763 23223
0 13030 7 1 2 26616 13029
0 13031 7 1 2 33881 13030
0 13032 7 1 2 33447 13031
0 13033 7 1 2 35970 13032
0 13034 7 1 2 13026 13033
0 13035 5 1 1 13034
0 13036 7 1 2 13022 13035
0 13037 5 1 1 13036
0 13038 7 1 2 25607 32783
0 13039 7 1 2 13037 13038
0 13040 5 1 1 13039
0 13041 7 1 2 12976 13040
0 13042 5 1 1 13041
0 13043 7 1 2 25505 13042
0 13044 5 1 1 13043
0 13045 7 4 2 22331 28929
0 13046 7 1 2 29986 35972
0 13047 7 2 2 25084 33510
0 13048 7 1 2 31415 34227
0 13049 7 1 2 35976 13048
0 13050 7 1 2 13046 13049
0 13051 5 1 1 13050
0 13052 7 1 2 28391 26830
0 13053 7 1 2 28743 13052
0 13054 7 1 2 31575 35529
0 13055 7 1 2 13053 13054
0 13056 5 1 1 13055
0 13057 7 1 2 13051 13056
0 13058 5 1 1 13057
0 13059 7 1 2 24962 13058
0 13060 5 1 1 13059
0 13061 7 2 2 23121 33010
0 13062 7 1 2 33822 35978
0 13063 5 1 1 13062
0 13064 7 1 2 30322 33971
0 13065 7 1 2 35895 13064
0 13066 7 1 2 31737 13065
0 13067 5 1 1 13066
0 13068 7 1 2 13063 13067
0 13069 5 1 1 13068
0 13070 7 1 2 21937 35300
0 13071 7 1 2 13069 13070
0 13072 5 1 1 13071
0 13073 7 1 2 13060 13072
0 13074 5 1 1 13073
0 13075 7 1 2 22068 13074
0 13076 5 1 1 13075
0 13077 7 1 2 25265 31486
0 13078 5 1 1 13077
0 13079 7 1 2 30569 30696
0 13080 7 1 2 29698 13079
0 13081 5 1 1 13080
0 13082 7 1 2 13078 13081
0 13083 5 1 1 13082
0 13084 7 1 2 28392 27031
0 13085 7 1 2 35530 13084
0 13086 7 1 2 13083 13085
0 13087 5 1 1 13086
0 13088 7 1 2 13076 13087
0 13089 5 1 1 13088
0 13090 7 1 2 27785 13089
0 13091 5 1 1 13090
0 13092 7 1 2 28002 33553
0 13093 7 1 2 32188 34568
0 13094 7 1 2 33762 13093
0 13095 7 1 2 13092 13094
0 13096 7 1 2 31840 34496
0 13097 7 1 2 13095 13096
0 13098 5 1 1 13097
0 13099 7 1 2 13091 13098
0 13100 5 1 1 13099
0 13101 7 1 2 25340 13100
0 13102 5 1 1 13101
0 13103 7 1 2 27021 35000
0 13104 5 1 1 13103
0 13105 7 1 2 21938 29911
0 13106 7 1 2 33490 13105
0 13107 5 1 1 13106
0 13108 7 1 2 13104 13107
0 13109 5 1 1 13108
0 13110 7 1 2 22069 13109
0 13111 5 1 1 13110
0 13112 7 1 2 27524 29092
0 13113 5 1 1 13112
0 13114 7 1 2 31746 13113
0 13115 5 1 1 13114
0 13116 7 1 2 34699 13115
0 13117 5 1 1 13116
0 13118 7 2 2 22070 29093
0 13119 5 1 1 35980
0 13120 7 1 2 29704 13119
0 13121 5 1 1 13120
0 13122 7 1 2 24620 31483
0 13123 7 1 2 13121 13122
0 13124 5 1 1 13123
0 13125 7 1 2 13117 13124
0 13126 5 1 1 13125
0 13127 7 1 2 24963 13126
0 13128 5 1 1 13127
0 13129 7 1 2 29390 29987
0 13130 7 1 2 31397 13129
0 13131 5 1 1 13130
0 13132 7 1 2 13128 13131
0 13133 7 1 2 13111 13132
0 13134 5 1 1 13133
0 13135 7 1 2 31859 34165
0 13136 7 1 2 13134 13135
0 13137 5 1 1 13136
0 13138 7 1 2 27022 31271
0 13139 7 1 2 33176 13138
0 13140 7 1 2 27662 13139
0 13141 7 1 2 32458 13140
0 13142 5 1 1 13141
0 13143 7 1 2 13137 13142
0 13144 5 1 1 13143
0 13145 7 1 2 35677 13144
0 13146 5 1 1 13145
0 13147 7 1 2 13102 13146
0 13148 5 1 1 13147
0 13149 7 1 2 25182 13148
0 13150 5 1 1 13149
0 13151 7 3 2 23224 33318
0 13152 7 3 2 28393 25967
0 13153 7 1 2 27656 31224
0 13154 7 2 2 35985 13153
0 13155 5 1 1 35988
0 13156 7 1 2 31416 35989
0 13157 5 1 1 13156
0 13158 7 1 2 29699 35681
0 13159 7 1 2 34166 13158
0 13160 5 1 1 13159
0 13161 7 1 2 13157 13160
0 13162 5 1 1 13161
0 13163 7 1 2 33491 13162
0 13164 5 1 1 13163
0 13165 7 2 2 31804 31959
0 13166 7 2 2 35682 35990
0 13167 7 1 2 30773 35992
0 13168 5 2 1 13167
0 13169 7 1 2 27410 28960
0 13170 7 1 2 30900 13169
0 13171 7 1 2 35986 13170
0 13172 5 1 1 13171
0 13173 7 1 2 35994 13172
0 13174 5 1 1 13173
0 13175 7 1 2 29988 13174
0 13176 5 1 1 13175
0 13177 7 1 2 13164 13176
0 13178 5 1 1 13177
0 13179 7 1 2 22071 13178
0 13180 5 1 1 13179
0 13181 7 1 2 13155 35995
0 13182 5 1 1 13181
0 13183 7 1 2 30084 13182
0 13184 5 1 1 13183
0 13185 7 1 2 13180 13184
0 13186 5 1 1 13185
0 13187 7 1 2 23459 13186
0 13188 5 1 1 13187
0 13189 7 1 2 23763 29922
0 13190 7 1 2 29761 34851
0 13191 7 1 2 13189 13190
0 13192 7 1 2 25977 13191
0 13193 7 1 2 29949 13192
0 13194 5 1 1 13193
0 13195 7 1 2 13188 13194
0 13196 5 1 1 13195
0 13197 7 1 2 23311 13196
0 13198 5 1 1 13197
0 13199 7 1 2 22561 34033
0 13200 5 1 1 13199
0 13201 7 1 2 22072 32626
0 13202 5 1 1 13201
0 13203 7 1 2 13200 13202
0 13204 5 1 1 13203
0 13205 7 1 2 29770 35993
0 13206 7 1 2 13204 13205
0 13207 5 1 1 13206
0 13208 7 2 2 24226 25341
0 13209 7 1 2 31809 35996
0 13210 7 1 2 31463 13209
0 13211 7 2 2 22406 26461
0 13212 7 1 2 35998 32359
0 13213 7 1 2 13210 13212
0 13214 5 1 1 13213
0 13215 7 1 2 13207 13214
0 13216 5 1 1 13215
0 13217 7 1 2 25085 13216
0 13218 5 1 1 13217
0 13219 7 2 2 23122 23378
0 13220 7 1 2 30155 31960
0 13221 7 1 2 36000 13220
0 13222 7 1 2 27683 27596
0 13223 7 1 2 33127 13222
0 13224 7 1 2 13221 13223
0 13225 5 1 1 13224
0 13226 7 1 2 13218 13225
0 13227 5 1 1 13226
0 13228 7 1 2 33940 13227
0 13229 5 1 1 13228
0 13230 7 1 2 13198 13229
0 13231 5 1 1 13230
0 13232 7 1 2 35982 13231
0 13233 5 1 1 13232
0 13234 7 1 2 13150 13233
0 13235 5 1 1 13234
0 13236 7 1 2 22764 13235
0 13237 5 1 1 13236
0 13238 7 1 2 27691 27597
0 13239 7 2 2 31248 33028
0 13240 7 1 2 31417 36002
0 13241 7 1 2 13238 13240
0 13242 7 1 2 30136 13241
0 13243 5 1 1 13242
0 13244 7 1 2 24818 31881
0 13245 7 1 2 30353 13244
0 13246 7 1 2 32068 13245
0 13247 5 1 1 13246
0 13248 7 1 2 27891 4190
0 13249 5 2 1 13248
0 13250 7 1 2 26318 28512
0 13251 7 1 2 36004 13250
0 13252 5 1 1 13251
0 13253 7 1 2 13247 13252
0 13254 5 1 1 13253
0 13255 7 1 2 27846 29963
0 13256 7 1 2 13254 13255
0 13257 5 1 1 13256
0 13258 7 1 2 13243 13257
0 13259 5 1 1 13258
0 13260 7 1 2 33823 13259
0 13261 5 1 1 13260
0 13262 7 1 2 28490 27054
0 13263 7 1 2 28877 34478
0 13264 7 1 2 13262 13263
0 13265 7 1 2 26773 28037
0 13266 7 1 2 31364 13265
0 13267 7 1 2 35345 13266
0 13268 7 1 2 13264 13267
0 13269 5 1 1 13268
0 13270 7 1 2 13261 13269
0 13271 5 1 1 13270
0 13272 7 1 2 22073 13271
0 13273 5 1 1 13272
0 13274 7 1 2 30281 31619
0 13275 7 1 2 29774 13274
0 13276 7 1 2 31302 33659
0 13277 7 1 2 32568 13276
0 13278 7 1 2 13275 13277
0 13279 5 1 1 13278
0 13280 7 1 2 13273 13279
0 13281 5 1 1 13280
0 13282 7 1 2 29012 13281
0 13283 5 1 1 13282
0 13284 7 5 2 22811 35319
0 13285 7 1 2 27986 35991
0 13286 7 1 2 30357 13285
0 13287 5 1 1 13286
0 13288 7 1 2 29372 35825
0 13289 7 1 2 35059 13288
0 13290 5 1 1 13289
0 13291 7 1 2 13287 13290
0 13292 5 1 1 13291
0 13293 7 1 2 23460 13292
0 13294 5 1 1 13293
0 13295 7 1 2 28394 27936
0 13296 7 1 2 35412 31877
0 13297 7 1 2 13295 13296
0 13298 5 1 1 13297
0 13299 7 1 2 13294 13298
0 13300 5 1 1 13299
0 13301 7 1 2 21939 13300
0 13302 5 1 1 13301
0 13303 7 2 2 33703 36005
0 13304 7 1 2 27389 35786
0 13305 7 1 2 36011 13304
0 13306 5 1 1 13305
0 13307 7 1 2 13302 13306
0 13308 5 1 1 13307
0 13309 7 1 2 29094 13308
0 13310 5 1 1 13309
0 13311 7 1 2 26576 29510
0 13312 7 1 2 35987 13311
0 13313 7 1 2 35192 13312
0 13314 7 1 2 30657 13313
0 13315 5 1 1 13314
0 13316 7 1 2 13310 13315
0 13317 5 1 1 13316
0 13318 7 1 2 27459 13317
0 13319 5 1 1 13318
0 13320 7 1 2 28248 26735
0 13321 7 1 2 27023 29571
0 13322 7 1 2 32157 13321
0 13323 7 1 2 13320 13322
0 13324 7 1 2 36012 13323
0 13325 5 1 1 13324
0 13326 7 1 2 13319 13325
0 13327 5 1 1 13326
0 13328 7 1 2 22074 13327
0 13329 5 1 1 13328
0 13330 7 1 2 22219 30027
0 13331 7 1 2 26869 13330
0 13332 5 1 1 13331
0 13333 7 1 2 27214 31645
0 13334 5 1 1 13333
0 13335 7 1 2 8960 13334
0 13336 5 1 1 13335
0 13337 7 1 2 26286 34852
0 13338 7 1 2 13336 13337
0 13339 5 1 1 13338
0 13340 7 1 2 13332 13339
0 13341 5 1 1 13340
0 13342 7 1 2 24106 27663
0 13343 7 1 2 13341 13342
0 13344 5 1 1 13343
0 13345 7 1 2 13329 13344
0 13346 5 1 1 13345
0 13347 7 1 2 36006 13346
0 13348 5 1 1 13347
0 13349 7 1 2 13283 13348
0 13350 7 1 2 13237 13349
0 13351 5 1 1 13350
0 13352 7 1 2 23549 13351
0 13353 5 1 1 13352
0 13354 7 1 2 29898 34828
0 13355 5 1 1 13354
0 13356 7 1 2 12475 13355
0 13357 5 1 1 13356
0 13358 7 1 2 29511 13357
0 13359 5 1 1 13358
0 13360 7 1 2 35787 33699
0 13361 5 1 1 13360
0 13362 7 1 2 13359 13361
0 13363 5 1 1 13362
0 13364 7 1 2 27460 13363
0 13365 5 1 1 13364
0 13366 7 2 2 29989 32201
0 13367 7 2 2 26381 33941
0 13368 7 1 2 36013 36015
0 13369 5 1 1 13368
0 13370 7 1 2 13365 13369
0 13371 5 1 1 13370
0 13372 7 1 2 22075 13371
0 13373 5 1 1 13372
0 13374 7 1 2 30402 34561
0 13375 7 1 2 30068 13374
0 13376 5 1 1 13375
0 13377 7 1 2 13373 13376
0 13378 5 1 1 13377
0 13379 7 1 2 25183 13378
0 13380 5 1 1 13379
0 13381 7 1 2 31373 31338
0 13382 5 1 1 13381
0 13383 7 1 2 29676 31230
0 13384 5 1 1 13383
0 13385 7 1 2 13382 13384
0 13386 5 1 1 13385
0 13387 7 1 2 35791 13386
0 13388 5 1 1 13387
0 13389 7 1 2 13380 13388
0 13390 5 1 1 13389
0 13391 7 1 2 24710 13390
0 13392 5 1 1 13391
0 13393 7 2 2 29923 35792
0 13394 7 1 2 29950 36017
0 13395 5 1 1 13394
0 13396 7 1 2 23461 31133
0 13397 7 1 2 31846 13396
0 13398 7 1 2 32459 13397
0 13399 5 1 1 13398
0 13400 7 1 2 13395 13399
0 13401 5 1 1 13400
0 13402 7 1 2 28518 13401
0 13403 5 1 1 13402
0 13404 7 1 2 13392 13403
0 13405 5 1 1 13404
0 13406 7 1 2 34414 13405
0 13407 5 1 1 13406
0 13408 7 2 2 33873 35689
0 13409 7 2 2 26309 34763
0 13410 5 2 1 36021
0 13411 7 1 2 33453 36022
0 13412 7 1 2 36019 13411
0 13413 7 1 2 35634 13412
0 13414 5 1 1 13413
0 13415 7 1 2 13407 13414
0 13416 5 1 1 13415
0 13417 7 1 2 27625 13416
0 13418 5 1 1 13417
0 13419 7 3 2 29572 31499
0 13420 5 1 1 36025
0 13421 7 1 2 22076 35648
0 13422 5 1 1 13421
0 13423 7 1 2 27461 30437
0 13424 5 1 1 13423
0 13425 7 1 2 13422 13424
0 13426 5 1 1 13425
0 13427 7 1 2 24964 13426
0 13428 5 1 1 13427
0 13429 7 1 2 13420 13428
0 13430 5 1 1 13429
0 13431 7 1 2 27248 13430
0 13432 5 1 1 13431
0 13433 7 1 2 26971 35635
0 13434 5 1 1 13433
0 13435 7 1 2 30901 34694
0 13436 5 1 1 13435
0 13437 7 1 2 8507 13436
0 13438 5 1 1 13437
0 13439 7 1 2 22077 13438
0 13440 5 1 1 13439
0 13441 7 2 2 31464 10046
0 13442 5 1 1 36028
0 13443 7 1 2 23225 36029
0 13444 5 1 1 13443
0 13445 7 2 2 22562 28200
0 13446 5 1 1 36030
0 13447 7 1 2 36031 35656
0 13448 5 1 1 13447
0 13449 7 1 2 30577 32216
0 13450 5 1 1 13449
0 13451 7 1 2 25184 13450
0 13452 7 1 2 13448 13451
0 13453 5 1 1 13452
0 13454 7 1 2 25086 13453
0 13455 7 1 2 13444 13454
0 13456 5 1 1 13455
0 13457 7 1 2 13440 13456
0 13458 5 1 1 13457
0 13459 7 1 2 22669 13458
0 13460 5 1 1 13459
0 13461 7 1 2 13434 13460
0 13462 7 1 2 13432 13461
0 13463 5 1 1 13462
0 13464 7 1 2 31630 33627
0 13465 7 1 2 13463 13464
0 13466 5 1 1 13465
0 13467 7 3 2 25506 27353
0 13468 7 1 2 29144 31332
0 13469 7 1 2 35888 13468
0 13470 7 1 2 36032 13469
0 13471 5 1 1 13470
0 13472 7 1 2 13466 13471
0 13473 5 1 1 13472
0 13474 7 1 2 22765 13473
0 13475 5 1 1 13474
0 13476 7 1 2 29798 32314
0 13477 5 3 1 13476
0 13478 7 1 2 23123 36035
0 13479 5 2 1 13478
0 13480 7 1 2 36036 34036
0 13481 5 1 1 13480
0 13482 7 2 2 36038 13481
0 13483 7 1 2 22563 36040
0 13484 5 1 1 13483
0 13485 7 1 2 28627 32536
0 13486 5 2 1 13485
0 13487 7 1 2 28426 28987
0 13488 5 3 1 13487
0 13489 7 1 2 29799 34664
0 13490 5 1 1 13489
0 13491 7 1 2 36044 13490
0 13492 5 3 1 13491
0 13493 7 1 2 21940 36047
0 13494 5 3 1 13493
0 13495 7 1 2 36042 36050
0 13496 7 1 2 13484 13495
0 13497 5 1 1 13496
0 13498 7 2 2 33874 34509
0 13499 7 1 2 28175 26310
0 13500 7 1 2 36053 13499
0 13501 7 1 2 13497 13500
0 13502 5 1 1 13501
0 13503 7 1 2 23312 13502
0 13504 7 1 2 13475 13503
0 13505 5 1 1 13504
0 13506 7 1 2 27288 32253
0 13507 7 1 2 35918 13506
0 13508 7 1 2 32165 13507
0 13509 7 1 2 34368 13508
0 13510 5 1 1 13509
0 13511 7 2 2 33253 33882
0 13512 7 2 2 24759 23226
0 13513 7 1 2 30244 36057
0 13514 7 1 2 36055 13513
0 13515 7 1 2 35941 13514
0 13516 5 1 1 13515
0 13517 7 1 2 13510 13516
0 13518 5 1 1 13517
0 13519 7 1 2 22670 13518
0 13520 5 1 1 13519
0 13521 7 1 2 24107 35733
0 13522 5 1 1 13521
0 13523 7 1 2 30989 32217
0 13524 5 1 1 13523
0 13525 7 1 2 13522 13524
0 13526 5 1 1 13525
0 13527 7 1 2 23227 13526
0 13528 5 1 1 13527
0 13529 7 1 2 27268 29670
0 13530 5 1 1 13529
0 13531 7 1 2 13528 13530
0 13532 5 1 1 13531
0 13533 7 1 2 35945 36054
0 13534 7 1 2 13532 13533
0 13535 5 1 1 13534
0 13536 7 1 2 13520 13535
0 13537 5 1 1 13536
0 13538 7 1 2 25087 13537
0 13539 5 1 1 13538
0 13540 7 1 2 28500 35747
0 13541 5 1 1 13540
0 13542 7 1 2 22078 30906
0 13543 5 1 1 13542
0 13544 7 1 2 23228 29297
0 13545 7 1 2 13543 13544
0 13546 5 1 1 13545
0 13547 7 1 2 13541 13546
0 13548 5 1 1 13547
0 13549 7 1 2 22671 13548
0 13550 5 1 1 13549
0 13551 7 1 2 28599 32315
0 13552 5 1 1 13551
0 13553 7 1 2 23229 31316
0 13554 5 1 1 13553
0 13555 7 1 2 13552 13554
0 13556 5 1 1 13555
0 13557 7 1 2 24621 13556
0 13558 5 1 1 13557
0 13559 7 1 2 35922 33130
0 13560 7 1 2 8848 13559
0 13561 5 1 1 13560
0 13562 7 1 2 13558 13561
0 13563 7 1 2 13550 13562
0 13564 5 1 1 13563
0 13565 7 1 2 24539 13564
0 13566 5 1 1 13565
0 13567 7 1 2 29354 32529
0 13568 5 1 1 13567
0 13569 7 1 2 29924 29700
0 13570 5 1 1 13569
0 13571 7 1 2 13568 13570
0 13572 5 1 1 13571
0 13573 7 1 2 32425 13572
0 13574 5 1 1 13573
0 13575 7 1 2 13566 13574
0 13576 5 1 1 13575
0 13577 7 1 2 29409 35889
0 13578 7 1 2 13576 13577
0 13579 5 1 1 13578
0 13580 7 1 2 13539 13579
0 13581 5 1 1 13580
0 13582 7 1 2 24711 13581
0 13583 5 1 1 13582
0 13584 7 1 2 28448 29391
0 13585 5 3 1 13584
0 13586 7 1 2 31022 36059
0 13587 5 5 1 13586
0 13588 7 2 2 22079 36062
0 13589 5 1 1 36067
0 13590 7 1 2 35644 13589
0 13591 5 1 1 13590
0 13592 7 3 2 28168 34415
0 13593 7 1 2 26266 36069
0 13594 7 1 2 13591 13593
0 13595 5 1 1 13594
0 13596 7 1 2 25266 13595
0 13597 7 1 2 13583 13596
0 13598 5 1 1 13597
0 13599 7 1 2 27611 13598
0 13600 7 1 2 13505 13599
0 13601 5 1 1 13600
0 13602 7 1 2 23379 13601
0 13603 7 1 2 13418 13602
0 13604 5 1 1 13603
0 13605 7 1 2 31121 33367
0 13606 7 1 2 31841 13605
0 13607 7 1 2 32013 13606
0 13608 5 1 1 13607
0 13609 7 2 2 33403 34108
0 13610 7 2 2 35956 36072
0 13611 7 1 2 27411 36074
0 13612 7 1 2 31487 13611
0 13613 5 1 1 13612
0 13614 7 1 2 13608 13613
0 13615 5 1 1 13614
0 13616 7 1 2 25267 13615
0 13617 5 1 1 13616
0 13618 7 1 2 24965 13442
0 13619 5 1 1 13618
0 13620 7 1 2 31708 13619
0 13621 5 1 1 13620
0 13622 7 1 2 32017 35979
0 13623 7 1 2 36073 13622
0 13624 7 1 2 13621 13623
0 13625 5 1 1 13624
0 13626 7 1 2 13617 13625
0 13627 5 1 1 13626
0 13628 7 1 2 25185 13627
0 13629 5 1 1 13628
0 13630 7 2 2 25268 35882
0 13631 5 1 1 36076
0 13632 7 1 2 22080 34655
0 13633 5 1 1 13632
0 13634 7 1 2 13631 13633
0 13635 5 1 1 13634
0 13636 7 1 2 25088 13635
0 13637 5 1 1 13636
0 13638 7 1 2 35876 13637
0 13639 5 1 1 13638
0 13640 7 1 2 24966 13639
0 13641 5 1 1 13640
0 13642 7 1 2 13641 5093
0 13643 5 1 1 13642
0 13644 7 1 2 30396 36075
0 13645 7 1 2 13643 13644
0 13646 5 1 1 13645
0 13647 7 1 2 13629 13646
0 13648 5 1 1 13647
0 13649 7 1 2 22766 13648
0 13650 5 1 1 13649
0 13651 7 2 2 22220 27963
0 13652 5 1 1 36078
0 13653 7 1 2 27809 36079
0 13654 5 1 1 13653
0 13655 7 1 2 27626 35826
0 13656 5 1 1 13655
0 13657 7 1 2 13654 13656
0 13658 5 1 1 13657
0 13659 7 1 2 35121 13658
0 13660 5 1 1 13659
0 13661 7 1 2 22871 25186
0 13662 7 1 2 23764 13661
0 13663 7 1 2 32784 13662
0 13664 7 3 2 29295 35272
0 13665 7 1 2 29248 36080
0 13666 7 1 2 13663 13665
0 13667 5 1 1 13666
0 13668 7 1 2 13660 13667
0 13669 5 1 1 13668
0 13670 7 1 2 23462 13669
0 13671 5 1 1 13670
0 13672 7 1 2 25863 34853
0 13673 7 1 2 30430 13672
0 13674 7 1 2 30477 13673
0 13675 5 1 1 13674
0 13676 7 1 2 13671 13675
0 13677 5 1 1 13676
0 13678 7 1 2 36007 13677
0 13679 5 1 1 13678
0 13680 7 1 2 23550 13679
0 13681 7 1 2 13650 13680
0 13682 5 1 1 13681
0 13683 7 3 2 25187 31286
0 13684 7 3 2 24540 24760
0 13685 7 1 2 26084 36086
0 13686 7 1 2 33281 13685
0 13687 7 1 2 36056 13686
0 13688 7 1 2 35756 13687
0 13689 5 1 1 13688
0 13690 7 1 2 33756 34552
0 13691 7 1 2 35935 13690
0 13692 5 1 1 13691
0 13693 7 1 2 13689 13692
0 13694 5 1 1 13693
0 13695 7 1 2 36083 13694
0 13696 5 1 1 13695
0 13697 7 2 2 23124 35230
0 13698 7 1 2 31785 32558
0 13699 7 3 2 31046 35210
0 13700 5 2 1 36091
0 13701 7 2 2 28449 34562
0 13702 7 1 2 36092 36096
0 13703 7 1 2 13698 13702
0 13704 7 1 2 36089 13703
0 13705 5 1 1 13704
0 13706 7 1 2 13696 13705
0 13707 5 1 1 13706
0 13708 7 1 2 23666 13707
0 13709 5 1 1 13708
0 13710 7 1 2 25089 36084
0 13711 7 1 2 33726 31878
0 13712 7 1 2 13710 13711
0 13713 7 1 2 31843 13712
0 13714 5 1 1 13713
0 13715 7 1 2 25507 13714
0 13716 7 1 2 13709 13715
0 13717 5 1 1 13716
0 13718 7 1 2 13682 13717
0 13719 5 1 1 13718
0 13720 7 1 2 25342 13719
0 13721 5 1 1 13720
0 13722 7 1 2 25944 13721
0 13723 7 1 2 13604 13722
0 13724 5 1 1 13723
0 13725 7 1 2 13353 13724
0 13726 7 1 2 13044 13725
0 13727 5 1 1 13726
0 13728 7 1 2 22148 13727
0 13729 5 1 1 13728
0 13730 7 1 2 31238 35828
0 13731 5 1 1 13730
0 13732 7 1 2 35784 13731
0 13733 5 1 1 13732
0 13734 7 1 2 30125 33177
0 13735 5 1 1 13734
0 13736 7 1 2 31239 13735
0 13737 5 1 1 13736
0 13738 7 1 2 29198 13737
0 13739 7 1 2 35810 13738
0 13740 5 1 1 13739
0 13741 7 1 2 13733 13740
0 13742 5 1 1 13741
0 13743 7 1 2 23551 13742
0 13744 5 1 1 13743
0 13745 7 1 2 28646 31235
0 13746 7 1 2 35817 13745
0 13747 5 1 1 13746
0 13748 7 1 2 13744 13747
0 13749 5 1 1 13748
0 13750 7 1 2 35139 13749
0 13751 5 1 1 13750
0 13752 7 1 2 25945 34190
0 13753 5 1 1 13752
0 13754 7 1 2 22332 35685
0 13755 5 1 1 13754
0 13756 7 1 2 13753 13755
0 13757 5 1 1 13756
0 13758 7 1 2 30632 13757
0 13759 5 1 1 13758
0 13760 7 1 2 25892 2610
0 13761 5 1 1 13760
0 13762 7 1 2 26134 4317
0 13763 5 1 1 13762
0 13764 7 1 2 35023 13763
0 13765 7 1 2 13761 13764
0 13766 5 1 1 13765
0 13767 7 1 2 13759 13766
0 13768 5 1 1 13767
0 13769 7 1 2 33092 32884
0 13770 7 1 2 32230 13769
0 13771 7 1 2 35100 13770
0 13772 7 1 2 13768 13771
0 13773 5 1 1 13772
0 13774 7 1 2 13751 13773
0 13775 5 1 1 13774
0 13776 7 1 2 35775 13775
0 13777 5 1 1 13776
0 13778 7 1 2 31296 35909
0 13779 5 1 1 13778
0 13780 7 2 2 21831 31374
0 13781 7 1 2 31765 36098
0 13782 5 1 1 13781
0 13783 7 1 2 13779 13782
0 13784 5 1 1 13783
0 13785 7 1 2 28583 13784
0 13786 5 1 1 13785
0 13787 7 2 2 23552 30013
0 13788 7 2 2 31297 36100
0 13789 7 1 2 23230 34515
0 13790 7 1 2 36102 13789
0 13791 5 1 1 13790
0 13792 7 1 2 13786 13791
0 13793 5 1 1 13792
0 13794 7 1 2 24341 13793
0 13795 5 1 1 13794
0 13796 7 2 2 28076 36101
0 13797 7 1 2 31298 32398
0 13798 7 1 2 36104 13797
0 13799 5 1 1 13798
0 13800 7 1 2 13795 13799
0 13801 5 1 1 13800
0 13802 7 1 2 33368 13801
0 13803 5 1 1 13802
0 13804 7 2 2 34905 34538
0 13805 7 1 2 29925 36106
0 13806 7 1 2 36105 13805
0 13807 5 1 1 13806
0 13808 7 1 2 13803 13807
0 13809 5 1 1 13808
0 13810 7 1 2 23313 13809
0 13811 5 1 1 13810
0 13812 7 1 2 34563 35886
0 13813 7 1 2 30071 13812
0 13814 5 1 1 13813
0 13815 7 1 2 13811 13814
0 13816 5 1 1 13815
0 13817 7 1 2 26608 13816
0 13818 5 1 1 13817
0 13819 7 1 2 24227 35837
0 13820 5 1 1 13819
0 13821 7 1 2 26267 32934
0 13822 7 1 2 30014 13821
0 13823 5 1 1 13822
0 13824 7 1 2 13820 13823
0 13825 5 1 1 13824
0 13826 7 1 2 22149 13825
0 13827 5 1 1 13826
0 13828 7 1 2 33029 35843
0 13829 5 1 1 13828
0 13830 7 1 2 26382 35827
0 13831 5 1 1 13830
0 13832 7 1 2 13829 13831
0 13833 5 1 1 13832
0 13834 7 1 2 29677 13833
0 13835 5 1 1 13834
0 13836 7 1 2 13827 13835
0 13837 5 1 1 13836
0 13838 7 1 2 33566 13837
0 13839 5 1 1 13838
0 13840 7 1 2 22221 35884
0 13841 5 1 1 13840
0 13842 7 1 2 26949 35880
0 13843 5 1 1 13842
0 13844 7 1 2 23231 13843
0 13845 7 1 2 13841 13844
0 13846 5 1 1 13845
0 13847 7 1 2 29017 33151
0 13848 5 1 1 13847
0 13849 7 1 2 28224 31451
0 13850 5 1 1 13849
0 13851 7 1 2 2411 13850
0 13852 7 1 2 13848 13851
0 13853 5 1 1 13852
0 13854 7 1 2 25269 13853
0 13855 5 1 1 13854
0 13856 7 1 2 35845 13855
0 13857 5 1 1 13856
0 13858 7 1 2 22150 13857
0 13859 5 1 1 13858
0 13860 7 1 2 27024 32874
0 13861 5 1 1 13860
0 13862 7 1 2 13859 13861
0 13863 5 1 1 13862
0 13864 7 1 2 24228 13863
0 13865 5 1 1 13864
0 13866 7 3 2 24164 22222
0 13867 7 1 2 30428 36108
0 13868 7 1 2 32871 13867
0 13869 5 1 1 13868
0 13870 7 1 2 25188 13869
0 13871 7 1 2 13865 13870
0 13872 5 1 1 13871
0 13873 7 1 2 34949 13872
0 13874 7 1 2 13846 13873
0 13875 5 1 1 13874
0 13876 7 1 2 13839 13875
0 13877 5 1 1 13876
0 13878 7 1 2 23667 13877
0 13879 5 1 1 13878
0 13880 7 1 2 26210 13879
0 13881 7 1 2 13818 13880
0 13882 5 1 1 13881
0 13883 7 3 2 23765 26135
0 13884 7 1 2 24229 35706
0 13885 5 1 1 13884
0 13886 7 1 2 35910 32935
0 13887 5 1 1 13886
0 13888 7 1 2 13885 13887
0 13889 5 1 1 13888
0 13890 7 1 2 33567 13889
0 13891 5 1 1 13890
0 13892 7 2 2 33319 32399
0 13893 7 1 2 22872 27964
0 13894 7 1 2 36114 13893
0 13895 7 1 2 36103 13894
0 13896 5 1 1 13895
0 13897 7 1 2 13891 13896
0 13898 5 1 1 13897
0 13899 7 1 2 26609 13898
0 13900 5 1 1 13899
0 13901 7 1 2 26226 13900
0 13902 5 1 1 13901
0 13903 7 1 2 36111 13902
0 13904 7 1 2 13882 13903
0 13905 5 1 1 13904
0 13906 7 1 2 13777 13905
0 13907 5 1 1 13906
0 13908 7 1 2 34295 13907
0 13909 5 1 1 13908
0 13910 7 1 2 28460 34971
0 13911 7 2 2 24541 26774
0 13912 7 1 2 33727 36116
0 13913 7 1 2 13910 13912
0 13914 7 1 2 35768 13913
0 13915 5 1 1 13914
0 13916 7 4 2 33412 31956
0 13917 7 1 2 25946 36118
0 13918 7 1 2 35772 13917
0 13919 7 1 2 35766 13918
0 13920 5 1 1 13919
0 13921 7 1 2 13915 13920
0 13922 7 1 2 13909 13921
0 13923 7 1 2 13729 13922
0 13924 7 1 2 12795 13923
0 13925 7 1 2 12352 13924
0 13926 5 1 1 13925
0 13927 7 1 2 22710 13926
0 13928 5 1 1 13927
0 13929 7 2 2 30664 35024
0 13930 7 1 2 26972 36077
0 13931 5 1 1 13930
0 13932 7 6 2 23314 30615
0 13933 7 1 2 29651 36124
0 13934 5 1 1 13933
0 13935 7 1 2 13931 13934
0 13936 5 1 1 13935
0 13937 7 1 2 24967 13936
0 13938 5 1 1 13937
0 13939 7 1 2 22672 10248
0 13940 5 1 1 13939
0 13941 7 1 2 31478 13940
0 13942 5 1 1 13941
0 13943 7 1 2 1924 13942
0 13944 5 1 1 13943
0 13945 7 1 2 23849 13944
0 13946 5 1 1 13945
0 13947 7 1 2 30043 35219
0 13948 5 1 1 13947
0 13949 7 1 2 13946 13948
0 13950 5 1 1 13949
0 13951 7 1 2 26736 13950
0 13952 5 1 1 13951
0 13953 7 1 2 13938 13952
0 13954 5 6 1 13953
0 13955 7 1 2 24230 36130
0 13956 5 1 1 13955
0 13957 7 1 2 31236 35220
0 13958 7 1 2 31676 13957
0 13959 5 1 1 13958
0 13960 7 1 2 13956 13959
0 13961 5 1 1 13960
0 13962 7 1 2 32972 13961
0 13963 5 1 1 13962
0 13964 7 1 2 36131 33241
0 13965 5 1 1 13964
0 13966 7 2 2 28055 34771
0 13967 5 2 1 36136
0 13968 7 2 2 24622 36137
0 13969 5 2 1 36140
0 13970 7 3 2 29712 33254
0 13971 7 1 2 31677 36144
0 13972 7 1 2 36141 13971
0 13973 5 1 1 13972
0 13974 7 1 2 13965 13973
0 13975 7 1 2 13963 13974
0 13976 5 1 1 13975
0 13977 7 1 2 36122 13976
0 13978 5 1 1 13977
0 13979 7 1 2 28584 36132
0 13980 5 2 1 13979
0 13981 7 1 2 30793 35221
0 13982 5 2 1 13981
0 13983 7 2 2 23850 31763
0 13984 5 2 1 36151
0 13985 7 2 2 24623 27307
0 13986 5 1 1 36155
0 13987 7 1 2 36153 13986
0 13988 5 1 1 13987
0 13989 7 1 2 31465 13988
0 13990 5 1 1 13989
0 13991 7 1 2 36149 13990
0 13992 5 1 1 13991
0 13993 7 1 2 25270 13992
0 13994 5 1 1 13993
0 13995 7 2 2 23315 27462
0 13996 7 1 2 31658 36157
0 13997 5 1 1 13996
0 13998 7 1 2 25189 13997
0 13999 7 1 2 13994 13998
0 14000 5 1 1 13999
0 14001 7 1 2 27333 34688
0 14002 5 1 1 14001
0 14003 7 1 2 25271 14002
0 14004 5 1 1 14003
0 14005 7 1 2 31307 32116
0 14006 5 1 1 14005
0 14007 7 1 2 14004 14006
0 14008 5 1 1 14007
0 14009 7 1 2 25090 14008
0 14010 5 1 1 14009
0 14011 7 1 2 30224 29652
0 14012 5 1 1 14011
0 14013 7 1 2 23232 14012
0 14014 7 1 2 14010 14013
0 14015 5 1 1 14014
0 14016 7 1 2 29217 14015
0 14017 7 2 2 14000 14016
0 14018 5 1 1 36159
0 14019 7 1 2 36147 14018
0 14020 5 1 1 14019
0 14021 7 1 2 26590 14020
0 14022 5 1 1 14021
0 14023 7 1 2 22081 31562
0 14024 5 1 1 14023
0 14025 7 1 2 26383 32118
0 14026 7 1 2 14024 14025
0 14027 5 1 1 14026
0 14028 7 1 2 31560 14027
0 14029 5 1 1 14028
0 14030 7 1 2 30176 14029
0 14031 5 1 1 14030
0 14032 7 1 2 26886 35571
0 14033 5 1 1 14032
0 14034 7 1 2 14031 14033
0 14035 5 1 1 14034
0 14036 7 1 2 26923 35957
0 14037 7 1 2 14035 14036
0 14038 5 1 1 14037
0 14039 7 1 2 14022 14038
0 14040 5 1 1 14039
0 14041 7 1 2 24712 14040
0 14042 5 1 1 14041
0 14043 7 1 2 26268 30389
0 14044 5 1 1 14043
0 14045 7 1 2 25190 31760
0 14046 5 2 1 14045
0 14047 7 1 2 26314 36161
0 14048 7 1 2 36152 14047
0 14049 5 1 1 14048
0 14050 7 1 2 14044 14049
0 14051 5 1 1 14050
0 14052 7 1 2 26021 35222
0 14053 7 1 2 14051 14052
0 14054 5 1 1 14053
0 14055 7 1 2 28891 34623
0 14056 5 1 1 14055
0 14057 7 1 2 2907 14056
0 14058 5 1 1 14057
0 14059 7 1 2 14058 35712
0 14060 5 1 1 14059
0 14061 7 1 2 26187 27330
0 14062 5 1 1 14061
0 14063 7 1 2 14060 14062
0 14064 5 1 1 14063
0 14065 7 1 2 31466 14064
0 14066 5 1 1 14065
0 14067 7 2 2 29392 30177
0 14068 7 1 2 29850 36163
0 14069 5 1 1 14068
0 14070 7 1 2 14066 14069
0 14071 7 1 2 14054 14070
0 14072 5 1 1 14071
0 14073 7 1 2 29218 14072
0 14074 5 1 1 14073
0 14075 7 1 2 25508 28077
0 14076 7 2 2 31678 14075
0 14077 5 1 1 36165
0 14078 7 3 2 29926 29460
0 14079 7 1 2 26022 36167
0 14080 7 1 2 36166 14079
0 14081 5 1 1 14080
0 14082 7 1 2 14074 14081
0 14083 5 1 1 14082
0 14084 7 1 2 28519 14083
0 14085 5 1 1 14084
0 14086 7 1 2 29936 32185
0 14087 5 1 1 14086
0 14088 7 1 2 3093 14087
0 14089 5 1 1 14088
0 14090 7 1 2 36158 14089
0 14091 5 1 1 14090
0 14092 7 1 2 830 36154
0 14093 5 1 1 14092
0 14094 7 1 2 31467 14093
0 14095 5 1 1 14094
0 14096 7 1 2 36150 14095
0 14097 5 1 1 14096
0 14098 7 1 2 26737 14097
0 14099 5 1 1 14098
0 14100 7 1 2 14091 14099
0 14101 5 1 1 14100
0 14102 7 1 2 29219 14101
0 14103 5 1 1 14102
0 14104 7 1 2 36148 14103
0 14105 5 1 1 14104
0 14106 7 1 2 24231 14105
0 14107 5 1 1 14106
0 14108 7 1 2 21832 4964
0 14109 5 1 1 14108
0 14110 7 1 2 29220 36162
0 14111 7 1 2 14109 14110
0 14112 5 1 1 14111
0 14113 7 1 2 14077 14112
0 14114 5 1 1 14113
0 14115 7 1 2 29927 14114
0 14116 5 1 1 14115
0 14117 7 2 2 26155 30450
0 14118 7 1 2 35551 36170
0 14119 5 1 1 14118
0 14120 7 1 2 14116 14119
0 14121 5 1 1 14120
0 14122 7 1 2 29461 31134
0 14123 7 1 2 14121 14122
0 14124 5 1 1 14123
0 14125 7 1 2 23553 31327
0 14126 7 1 2 28088 14125
0 14127 7 1 2 30502 14126
0 14128 5 1 1 14127
0 14129 7 1 2 14124 14128
0 14130 5 1 1 14129
0 14131 7 1 2 33030 14130
0 14132 5 1 1 14131
0 14133 7 1 2 14107 14132
0 14134 5 1 1 14133
0 14135 7 1 2 32973 14134
0 14136 5 1 1 14135
0 14137 7 1 2 14085 14136
0 14138 7 1 2 14042 14137
0 14139 5 1 1 14138
0 14140 7 1 2 33413 14139
0 14141 5 1 1 14140
0 14142 7 1 2 13978 14141
0 14143 5 1 1 14142
0 14144 7 1 2 24165 14143
0 14145 5 1 1 14144
0 14146 7 1 2 27525 26901
0 14147 5 1 1 14146
0 14148 7 1 2 30232 14147
0 14149 5 1 1 14148
0 14150 7 2 2 33414 31935
0 14151 7 1 2 36145 33082
0 14152 7 1 2 36172 14151
0 14153 7 1 2 14149 14152
0 14154 5 1 1 14153
0 14155 7 1 2 14145 14154
0 14156 5 1 1 14155
0 14157 7 1 2 23668 14156
0 14158 5 1 1 14157
0 14159 7 1 2 23851 31249
0 14160 7 1 2 31237 14159
0 14161 5 1 1 14160
0 14162 7 3 2 28902 34764
0 14163 5 1 1 36174
0 14164 7 3 2 24232 23125
0 14165 7 1 2 36175 36177
0 14166 5 1 1 14165
0 14167 7 1 2 14161 14166
0 14168 5 1 1 14167
0 14169 7 1 2 34932 14168
0 14170 5 1 1 14169
0 14171 7 1 2 22767 31231
0 14172 7 1 2 27937 14171
0 14173 5 2 1 14172
0 14174 7 1 2 24233 36176
0 14175 5 1 1 14174
0 14176 7 1 2 36180 14175
0 14177 5 1 1 14176
0 14178 7 2 2 25509 14177
0 14179 7 1 2 36182 36090
0 14180 5 1 1 14179
0 14181 7 1 2 14170 14180
0 14182 5 1 1 14181
0 14183 7 1 2 27308 14182
0 14184 5 1 1 14183
0 14185 7 1 2 24234 28401
0 14186 7 1 2 30236 14185
0 14187 5 1 1 14186
0 14188 7 1 2 14187 36181
0 14189 5 1 1 14188
0 14190 7 1 2 34933 14189
0 14191 5 1 1 14190
0 14192 7 2 2 23852 33369
0 14193 7 2 2 26085 36184
0 14194 7 1 2 36183 36186
0 14195 5 1 1 14194
0 14196 7 1 2 14191 14195
0 14197 5 1 1 14196
0 14198 7 1 2 30044 14197
0 14199 5 1 1 14198
0 14200 7 2 2 26287 34731
0 14201 7 1 2 28536 36188
0 14202 7 1 2 33679 14201
0 14203 5 1 1 14202
0 14204 7 1 2 14199 14203
0 14205 7 1 2 14184 14204
0 14206 5 1 1 14205
0 14207 7 1 2 31508 35273
0 14208 7 1 2 14206 14207
0 14209 5 1 1 14208
0 14210 7 1 2 14158 14209
0 14211 5 1 1 14210
0 14212 7 1 2 25412 14211
0 14213 5 1 1 14212
0 14214 7 1 2 28014 36160
0 14215 5 1 1 14214
0 14216 7 1 2 23554 27906
0 14217 5 1 1 14216
0 14218 7 1 2 1354 14217
0 14219 5 1 1 14218
0 14220 7 1 2 36133 14219
0 14221 5 1 1 14220
0 14222 7 1 2 14215 14221
0 14223 5 1 1 14222
0 14224 7 1 2 33320 14223
0 14225 5 1 1 14224
0 14226 7 1 2 28723 36134
0 14227 5 1 1 14226
0 14228 7 2 2 30304 34732
0 14229 7 1 2 26086 35748
0 14230 7 1 2 31756 14229
0 14231 7 1 2 36190 14230
0 14232 5 1 1 14231
0 14233 7 1 2 14227 14232
0 14234 5 1 1 14233
0 14235 7 1 2 33370 14234
0 14236 5 1 1 14235
0 14237 7 1 2 14225 14236
0 14238 5 1 1 14237
0 14239 7 1 2 31178 14238
0 14240 5 1 1 14239
0 14241 7 1 2 27907 30045
0 14242 5 1 1 14241
0 14243 7 1 2 27309 27884
0 14244 5 1 1 14243
0 14245 7 1 2 14242 14244
0 14246 5 1 1 14245
0 14247 7 1 2 24624 14246
0 14248 5 1 1 14247
0 14249 7 1 2 29236 30503
0 14250 5 1 1 14249
0 14251 7 1 2 14248 14250
0 14252 5 1 1 14251
0 14253 7 1 2 25510 14252
0 14254 5 1 1 14253
0 14255 7 1 2 25608 36156
0 14256 7 1 2 29164 14255
0 14257 5 1 1 14256
0 14258 7 1 2 14254 14257
0 14259 5 1 1 14258
0 14260 7 1 2 24108 14259
0 14261 5 1 1 14260
0 14262 7 1 2 28048 29899
0 14263 7 1 2 28659 14262
0 14264 5 1 1 14263
0 14265 7 1 2 14261 14264
0 14266 5 1 1 14265
0 14267 7 1 2 23853 14266
0 14268 5 1 1 14267
0 14269 7 1 2 28724 30046
0 14270 5 1 1 14269
0 14271 7 2 2 27908 29410
0 14272 5 1 1 36192
0 14273 7 1 2 27310 36193
0 14274 5 1 1 14273
0 14275 7 1 2 14270 14274
0 14276 5 1 1 14275
0 14277 7 1 2 29928 14276
0 14278 5 1 1 14277
0 14279 7 1 2 14268 14278
0 14280 5 1 1 14279
0 14281 7 1 2 33321 14280
0 14282 5 1 1 14281
0 14283 7 1 2 23854 30526
0 14284 5 1 1 14283
0 14285 7 1 2 30543 14284
0 14286 5 1 1 14285
0 14287 7 1 2 30047 14286
0 14288 5 1 1 14287
0 14289 7 2 2 28833 29411
0 14290 5 1 1 36194
0 14291 7 1 2 23555 27639
0 14292 5 1 1 14291
0 14293 7 1 2 14290 14292
0 14294 5 1 1 14293
0 14295 7 1 2 27311 14294
0 14296 5 1 1 14295
0 14297 7 1 2 14288 14296
0 14298 5 1 1 14297
0 14299 7 1 2 29929 33711
0 14300 7 1 2 14298 14299
0 14301 5 1 1 14300
0 14302 7 1 2 14282 14301
0 14303 5 1 1 14302
0 14304 7 1 2 29462 14303
0 14305 5 1 1 14304
0 14306 7 1 2 29412 31434
0 14307 7 1 2 34599 14306
0 14308 7 1 2 29199 35181
0 14309 7 1 2 14307 14308
0 14310 5 1 1 14309
0 14311 7 1 2 14305 14310
0 14312 5 1 1 14311
0 14313 7 3 2 33011 35211
0 14314 7 1 2 23380 36196
0 14315 7 1 2 14312 14314
0 14316 5 1 1 14315
0 14317 7 1 2 14240 14316
0 14318 5 1 1 14317
0 14319 7 1 2 28549 14318
0 14320 5 1 1 14319
0 14321 7 1 2 14213 14320
0 14322 5 1 1 14321
0 14323 7 1 2 26211 14322
0 14324 5 1 1 14323
0 14325 7 1 2 26858 36135
0 14326 5 1 1 14325
0 14327 7 1 2 27973 36168
0 14328 7 1 2 31679 14327
0 14329 5 1 1 14328
0 14330 7 1 2 14326 14329
0 14331 5 1 1 14330
0 14332 7 1 2 29221 14331
0 14333 5 1 1 14332
0 14334 7 2 2 24109 28585
0 14335 5 1 1 36199
0 14336 7 1 2 26870 36200
0 14337 7 1 2 34774 14336
0 14338 5 1 1 14337
0 14339 7 1 2 14333 14338
0 14340 5 1 1 14339
0 14341 7 1 2 22768 14340
0 14342 5 1 1 14341
0 14343 7 1 2 28176 30633
0 14344 7 1 2 35223 14343
0 14345 7 1 2 36189 14344
0 14346 5 1 1 14345
0 14347 7 1 2 14342 14346
0 14348 5 1 1 14347
0 14349 7 1 2 22223 14348
0 14350 5 1 1 14349
0 14351 7 1 2 24625 33162
0 14352 7 3 2 35822 14351
0 14353 5 1 1 36201
0 14354 7 1 2 22873 36202
0 14355 5 1 1 14354
0 14356 7 2 2 25413 30634
0 14357 7 1 2 22769 26288
0 14358 5 1 1 14357
0 14359 7 1 2 14163 14358
0 14360 5 3 1 14359
0 14361 7 1 2 36204 36206
0 14362 5 1 1 14361
0 14363 7 1 2 14355 14362
0 14364 5 1 1 14363
0 14365 7 1 2 34775 34564
0 14366 7 1 2 14364 14365
0 14367 5 1 1 14366
0 14368 7 1 2 14350 14367
0 14369 5 1 1 14368
0 14370 7 1 2 22333 14369
0 14371 5 1 1 14370
0 14372 7 2 2 26514 32974
0 14373 5 1 1 36209
0 14374 7 1 2 24713 25191
0 14375 7 1 2 25806 14374
0 14376 5 1 1 14375
0 14377 7 2 2 14373 14376
0 14378 5 1 1 36211
0 14379 7 1 2 22224 36212
0 14380 5 1 1 14379
0 14381 7 2 2 26738 32975
0 14382 5 1 1 36213
0 14383 7 1 2 24235 36142
0 14384 7 1 2 14382 14383
0 14385 5 1 1 14384
0 14386 7 1 2 25414 14385
0 14387 7 1 2 14380 14386
0 14388 5 1 1 14387
0 14389 7 3 2 26775 26859
0 14390 5 1 1 36215
0 14391 7 1 2 26739 36216
0 14392 5 1 1 14391
0 14393 7 1 2 14388 14392
0 14394 5 2 1 14393
0 14395 7 1 2 30665 34733
0 14396 7 2 2 36218 14395
0 14397 7 1 2 32421 36220
0 14398 5 1 1 14397
0 14399 7 1 2 14371 14398
0 14400 5 1 1 14399
0 14401 7 1 2 33322 14400
0 14402 5 1 1 14401
0 14403 7 1 2 35224 33685
0 14404 7 1 2 36221 14403
0 14405 5 1 1 14404
0 14406 7 1 2 14402 14405
0 14407 5 1 1 14406
0 14408 7 1 2 24166 27563
0 14409 7 1 2 14407 14408
0 14410 5 1 1 14409
0 14411 7 1 2 14324 14410
0 14412 5 1 1 14411
0 14413 7 1 2 24654 14412
0 14414 5 1 1 14413
0 14415 7 3 2 27944 36125
0 14416 5 1 1 36222
0 14417 7 3 2 29573 36223
0 14418 5 1 1 36225
0 14419 7 1 2 22151 30701
0 14420 5 1 1 14419
0 14421 7 1 2 23126 30729
0 14422 5 1 1 14421
0 14423 7 1 2 14420 14422
0 14424 5 4 1 14423
0 14425 7 1 2 22564 36228
0 14426 5 1 1 14425
0 14427 7 1 2 31108 14426
0 14428 5 1 1 14427
0 14429 7 1 2 24236 14428
0 14430 5 1 1 14429
0 14431 7 1 2 30748 31534
0 14432 5 2 1 14431
0 14433 7 1 2 22673 30749
0 14434 5 1 1 14433
0 14435 7 2 2 36232 14434
0 14436 7 2 2 27965 27939
0 14437 7 1 2 36234 36236
0 14438 5 1 1 14437
0 14439 7 1 2 14430 14438
0 14440 5 1 1 14439
0 14441 7 1 2 21941 14440
0 14442 5 1 1 14441
0 14443 7 1 2 13652 35829
0 14444 5 2 1 14443
0 14445 7 2 2 29095 36238
0 14446 5 1 1 36240
0 14447 7 1 2 30616 33031
0 14448 5 1 1 14447
0 14449 7 1 2 14446 14448
0 14450 5 1 1 14449
0 14451 7 1 2 26538 14450
0 14452 5 1 1 14451
0 14453 7 1 2 14442 14452
0 14454 5 1 1 14453
0 14455 7 1 2 27463 14454
0 14456 5 1 1 14455
0 14457 7 1 2 22565 31051
0 14458 5 1 1 14457
0 14459 7 1 2 3084 14458
0 14460 5 6 1 14459
0 14461 7 2 2 33032 36242
0 14462 5 1 1 36248
0 14463 7 1 2 14462 35914
0 14464 5 1 1 14463
0 14465 7 1 2 26539 14464
0 14466 5 1 1 14465
0 14467 7 1 2 14456 14466
0 14468 5 1 1 14467
0 14469 7 1 2 24968 14468
0 14470 5 1 1 14469
0 14471 7 1 2 14418 14470
0 14472 5 1 1 14471
0 14473 7 1 2 26408 14472
0 14474 5 1 1 14473
0 14475 7 2 2 25609 35916
0 14476 7 2 2 24167 24866
0 14477 7 2 2 29686 36252
0 14478 7 1 2 36250 36254
0 14479 5 1 1 14478
0 14480 7 1 2 14474 14479
0 14481 5 1 1 14480
0 14482 7 1 2 22407 14481
0 14483 5 1 1 14482
0 14484 7 1 2 22935 26540
0 14485 7 2 2 31908 14484
0 14486 7 1 2 36251 36256
0 14487 5 1 1 14486
0 14488 7 1 2 14483 14487
0 14489 5 1 1 14488
0 14490 7 1 2 33602 14489
0 14491 5 1 1 14490
0 14492 7 1 2 29641 35852
0 14493 7 1 2 27226 14492
0 14494 7 1 2 33084 14493
0 14495 7 1 2 33593 14494
0 14496 5 1 1 14495
0 14497 7 1 2 14491 14496
0 14498 5 1 1 14497
0 14499 7 1 2 34296 14498
0 14500 5 1 1 14499
0 14501 7 1 2 27945 32792
0 14502 5 1 1 14501
0 14503 7 1 2 24237 36229
0 14504 5 1 1 14503
0 14505 7 3 2 24655 23127
0 14506 7 3 2 26269 36258
0 14507 7 1 2 33033 36261
0 14508 5 1 1 14507
0 14509 7 1 2 14504 14508
0 14510 5 1 1 14509
0 14511 7 2 2 22566 14510
0 14512 5 1 1 36264
0 14513 7 1 2 14502 14512
0 14514 5 1 1 14513
0 14515 7 1 2 21942 14514
0 14516 5 1 1 14515
0 14517 7 1 2 30599 31063
0 14518 5 1 1 14517
0 14519 7 1 2 26996 36109
0 14520 7 1 2 14518 14519
0 14521 5 1 1 14520
0 14522 7 1 2 14516 14521
0 14523 5 1 1 14522
0 14524 7 1 2 27464 14523
0 14525 5 1 1 14524
0 14526 7 1 2 26541 36249
0 14527 5 1 1 14526
0 14528 7 1 2 14525 14527
0 14529 5 1 1 14528
0 14530 7 1 2 25343 14529
0 14531 5 1 1 14530
0 14532 7 1 2 26712 36110
0 14533 7 1 2 35754 14532
0 14534 5 1 1 14533
0 14535 7 1 2 14531 14534
0 14536 5 1 1 14535
0 14537 7 1 2 24969 14536
0 14538 5 1 1 14537
0 14539 7 1 2 25344 36226
0 14540 5 1 1 14539
0 14541 7 1 2 14538 14540
0 14542 5 1 1 14541
0 14543 7 1 2 22770 14542
0 14544 5 1 1 14543
0 14545 7 1 2 22225 29642
0 14546 7 1 2 29430 30745
0 14547 7 1 2 14545 14546
0 14548 7 2 2 24656 24714
0 14549 7 2 2 22674 36266
0 14550 7 1 2 30237 36268
0 14551 7 1 2 14547 14550
0 14552 5 1 1 14551
0 14553 7 1 2 14544 14552
0 14554 5 1 1 14553
0 14555 7 1 2 23463 14554
0 14556 5 1 1 14555
0 14557 7 1 2 27465 28177
0 14558 7 1 2 26595 14557
0 14559 7 1 2 35703 14558
0 14560 5 1 1 14559
0 14561 7 1 2 14556 14560
0 14562 5 1 1 14561
0 14563 7 1 2 33594 14562
0 14564 5 1 1 14563
0 14565 7 3 2 24168 34431
0 14566 7 1 2 28508 36270
0 14567 5 1 1 14566
0 14568 7 1 2 1107 33772
0 14569 5 1 1 14568
0 14570 7 1 2 34435 7964
0 14571 5 2 1 14570
0 14572 7 1 2 22567 36273
0 14573 7 1 2 14569 14572
0 14574 5 1 1 14573
0 14575 7 1 2 14567 14574
0 14576 5 1 1 14575
0 14577 7 1 2 34272 14576
0 14578 5 1 1 14577
0 14579 7 1 2 30821 33012
0 14580 7 1 2 35983 14579
0 14581 7 1 2 36235 14580
0 14582 5 1 1 14581
0 14583 7 1 2 14578 14582
0 14584 5 1 1 14583
0 14585 7 1 2 21943 14584
0 14586 5 1 1 14585
0 14587 7 1 2 24238 35793
0 14588 5 1 1 14587
0 14589 7 1 2 35789 14588
0 14590 5 2 1 14589
0 14591 7 2 2 29096 36275
0 14592 5 1 1 36277
0 14593 7 2 2 30617 34829
0 14594 5 1 1 36279
0 14595 7 1 2 14592 14594
0 14596 5 1 1 14595
0 14597 7 1 2 36271 14596
0 14598 5 1 1 14597
0 14599 7 1 2 14586 14598
0 14600 5 1 1 14599
0 14601 7 1 2 27466 14600
0 14602 5 1 1 14601
0 14603 7 2 2 25818 33942
0 14604 7 1 2 36014 36281
0 14605 5 2 1 14604
0 14606 7 1 2 36243 34830
0 14607 5 1 1 14606
0 14608 7 1 2 36283 14607
0 14609 5 1 1 14608
0 14610 7 1 2 36272 14609
0 14611 5 1 1 14610
0 14612 7 1 2 14602 14611
0 14613 5 1 1 14612
0 14614 7 1 2 24970 14613
0 14615 5 1 1 14614
0 14616 7 1 2 34444 32141
0 14617 5 1 1 14616
0 14618 7 1 2 30618 34432
0 14619 5 1 1 14618
0 14620 7 1 2 14617 14619
0 14621 5 1 1 14620
0 14622 7 1 2 29574 14621
0 14623 5 1 1 14622
0 14624 7 1 2 24761 29512
0 14625 7 1 2 34793 14624
0 14626 7 1 2 30659 14625
0 14627 5 1 1 14626
0 14628 7 1 2 14623 14627
0 14629 5 1 1 14628
0 14630 7 1 2 35861 14629
0 14631 5 1 1 14630
0 14632 7 1 2 14615 14631
0 14633 5 1 1 14632
0 14634 7 1 2 24657 14633
0 14635 5 1 1 14634
0 14636 7 7 2 23316 29439
0 14637 7 1 2 33769 35874
0 14638 7 1 2 36274 14637
0 14639 7 1 2 36285 14638
0 14640 5 1 1 14639
0 14641 7 1 2 14635 14640
0 14642 5 1 1 14641
0 14643 7 1 2 22936 14642
0 14644 5 1 1 14643
0 14645 7 1 2 30350 34831
0 14646 5 1 1 14645
0 14647 7 1 2 36284 14646
0 14648 5 1 1 14647
0 14649 7 2 2 30305 14648
0 14650 7 1 2 33323 36255
0 14651 7 1 2 36292 14650
0 14652 5 1 1 14651
0 14653 7 1 2 14644 14652
0 14654 5 1 1 14653
0 14655 7 1 2 22408 14654
0 14656 5 1 1 14655
0 14657 7 1 2 33324 36257
0 14658 7 1 2 36293 14657
0 14659 5 1 1 14658
0 14660 7 1 2 14656 14659
0 14661 5 1 1 14660
0 14662 7 1 2 32976 14661
0 14663 5 1 1 14662
0 14664 7 1 2 14564 14663
0 14665 7 1 2 14500 14664
0 14666 5 1 1 14665
0 14667 7 1 2 28834 14666
0 14668 5 1 1 14667
0 14669 7 2 2 22771 26384
0 14670 7 1 2 31220 36294
0 14671 5 1 1 14670
0 14672 7 1 2 14671 36094
0 14673 5 1 1 14672
0 14674 7 1 2 22675 14673
0 14675 5 1 1 14674
0 14676 7 1 2 27269 28178
0 14677 7 1 2 30697 14676
0 14678 5 1 1 14677
0 14679 7 1 2 14675 14678
0 14680 5 1 1 14679
0 14681 7 1 2 23381 14680
0 14682 5 1 1 14681
0 14683 7 1 2 26860 27966
0 14684 7 1 2 36295 14683
0 14685 5 1 1 14684
0 14686 7 1 2 14682 14685
0 14687 5 1 1 14686
0 14688 7 1 2 34416 14687
0 14689 5 1 1 14688
0 14690 7 1 2 28162 34297
0 14691 7 1 2 35899 14690
0 14692 5 1 1 14691
0 14693 7 1 2 14689 14692
0 14694 5 1 1 14693
0 14695 7 1 2 22226 14694
0 14696 5 1 1 14695
0 14697 7 1 2 30339 31047
0 14698 7 1 2 33216 34369
0 14699 7 1 2 14697 14698
0 14700 5 1 1 14699
0 14701 7 1 2 14696 14700
0 14702 5 1 1 14701
0 14703 7 1 2 29513 14702
0 14704 5 1 1 14703
0 14705 7 2 2 23464 33665
0 14706 7 3 2 22812 25345
0 14707 7 1 2 30722 36298
0 14708 7 1 2 35393 14707
0 14709 7 1 2 36296 14708
0 14710 5 1 1 14709
0 14711 7 1 2 14704 14710
0 14712 5 1 1 14711
0 14713 7 1 2 26542 14712
0 14714 5 1 1 14713
0 14715 7 1 2 36230 34806
0 14716 5 1 1 14715
0 14717 7 2 2 24287 29991
0 14718 7 1 2 24762 25091
0 14719 7 1 2 35692 14718
0 14720 7 1 2 36301 14719
0 14721 5 1 1 14720
0 14722 7 1 2 14716 14721
0 14723 5 1 1 14722
0 14724 7 1 2 14723 33204
0 14725 5 1 1 14724
0 14726 7 1 2 31791 34351
0 14727 5 1 1 14726
0 14728 7 4 2 25272 26311
0 14729 7 1 2 31214 33325
0 14730 7 1 2 36303 14729
0 14731 5 1 1 14730
0 14732 7 1 2 14727 14731
0 14733 5 1 1 14732
0 14734 7 1 2 22227 14733
0 14735 5 1 1 14734
0 14736 7 1 2 24239 36085
0 14737 7 1 2 35246 14736
0 14738 5 1 1 14737
0 14739 7 1 2 14735 14738
0 14740 5 1 1 14739
0 14741 7 1 2 30746 14740
0 14742 5 1 1 14741
0 14743 7 1 2 22813 30708
0 14744 7 1 2 30807 14743
0 14745 7 1 2 35394 14744
0 14746 5 1 1 14745
0 14747 7 1 2 14742 14746
0 14748 5 1 1 14747
0 14749 7 1 2 27080 14748
0 14750 5 1 1 14749
0 14751 7 1 2 14725 14750
0 14752 5 1 1 14751
0 14753 7 1 2 23465 14752
0 14754 5 1 1 14753
0 14755 7 1 2 24240 30358
0 14756 5 1 1 14755
0 14757 7 1 2 28524 14756
0 14758 5 1 1 14757
0 14759 7 1 2 59 756
0 14760 5 1 1 14759
0 14761 7 1 2 25092 25415
0 14762 7 1 2 26543 14761
0 14763 7 1 2 34370 14762
0 14764 7 1 2 14760 14763
0 14765 7 1 2 14758 14764
0 14766 5 1 1 14765
0 14767 7 1 2 14754 14766
0 14768 5 1 1 14767
0 14769 7 1 2 29575 14768
0 14770 5 1 1 14769
0 14771 7 1 2 14714 14770
0 14772 5 1 1 14771
0 14773 7 1 2 27467 14772
0 14774 5 1 1 14773
0 14775 7 1 2 29842 30619
0 14776 5 1 1 14775
0 14777 7 1 2 4140 14776
0 14778 5 1 1 14777
0 14779 7 1 2 26023 14778
0 14780 5 1 1 14779
0 14781 7 1 2 25826 29970
0 14782 5 1 1 14781
0 14783 7 1 2 14780 14782
0 14784 5 1 1 14783
0 14785 7 1 2 21944 14784
0 14786 5 1 1 14785
0 14787 7 1 2 25346 30570
0 14788 7 1 2 36126 14787
0 14789 5 1 1 14788
0 14790 7 1 2 14786 14789
0 14791 5 1 1 14790
0 14792 7 1 2 26544 36070
0 14793 7 1 2 14791 14792
0 14794 5 1 1 14793
0 14795 7 1 2 14774 14794
0 14796 5 1 1 14795
0 14797 7 1 2 28124 14796
0 14798 5 1 1 14797
0 14799 7 1 2 21945 36265
0 14800 5 1 1 14799
0 14801 7 1 2 14416 14800
0 14802 5 1 1 14801
0 14803 7 1 2 33637 14802
0 14804 5 1 1 14803
0 14805 7 1 2 30233 30693
0 14806 5 1 1 14805
0 14807 7 1 2 22152 14806
0 14808 5 1 1 14807
0 14809 7 1 2 23018 30730
0 14810 5 1 1 14809
0 14811 7 1 2 14808 14810
0 14812 5 1 1 14811
0 14813 7 1 2 34417 14812
0 14814 5 1 1 14813
0 14815 7 2 2 28878 33371
0 14816 7 1 2 26545 35693
0 14817 7 1 2 36307 14816
0 14818 5 1 1 14817
0 14819 7 1 2 14814 14818
0 14820 5 2 1 14819
0 14821 7 1 2 24241 36309
0 14822 5 1 1 14821
0 14823 7 1 2 24169 33635
0 14824 5 1 1 14823
0 14825 7 1 2 24626 34447
0 14826 5 1 1 14825
0 14827 7 1 2 14824 14826
0 14828 5 2 1 14827
0 14829 7 1 2 36237 36311
0 14830 5 1 1 14829
0 14831 7 1 2 14822 14830
0 14832 5 1 1 14831
0 14833 7 1 2 29937 14832
0 14834 5 1 1 14833
0 14835 7 1 2 14804 14834
0 14836 5 1 1 14835
0 14837 7 1 2 27468 14836
0 14838 5 1 1 14837
0 14839 7 1 2 36227 34352
0 14840 5 1 1 14839
0 14841 7 1 2 29514 36224
0 14842 5 1 1 14841
0 14843 7 4 2 21946 26546
0 14844 7 1 2 36241 36313
0 14845 5 1 1 14844
0 14846 7 1 2 14842 14845
0 14847 5 1 1 14846
0 14848 7 1 2 33638 14847
0 14849 5 1 1 14848
0 14850 7 1 2 14840 14849
0 14851 7 1 2 14838 14850
0 14852 5 1 1 14851
0 14853 7 1 2 34298 14852
0 14854 5 1 1 14853
0 14855 7 9 2 26547 34854
0 14856 5 1 1 36317
0 14857 7 2 2 36127 36318
0 14858 5 1 1 36326
0 14859 7 1 2 31631 36231
0 14860 5 1 1 14859
0 14861 7 1 2 36262 35850
0 14862 5 1 1 14861
0 14863 7 1 2 14860 14862
0 14864 5 1 1 14863
0 14865 7 1 2 29576 14864
0 14866 5 1 1 14865
0 14867 7 1 2 14858 14866
0 14868 5 1 1 14867
0 14869 7 1 2 27469 14868
0 14870 5 1 1 14869
0 14871 7 1 2 36278 36314
0 14872 5 1 1 14871
0 14873 7 1 2 14870 14872
0 14874 5 1 1 14873
0 14875 7 1 2 33639 14874
0 14876 5 1 1 14875
0 14877 7 1 2 36327 33640
0 14878 5 1 1 14877
0 14879 7 1 2 31632 36310
0 14880 5 1 1 14879
0 14881 7 6 2 24242 24658
0 14882 7 1 2 35794 36328
0 14883 7 1 2 36312 14882
0 14884 5 1 1 14883
0 14885 7 1 2 14880 14884
0 14886 5 1 1 14885
0 14887 7 1 2 29861 14886
0 14888 5 1 1 14887
0 14889 7 1 2 14878 14888
0 14890 5 1 1 14889
0 14891 7 1 2 29515 14890
0 14892 5 1 1 14891
0 14893 7 1 2 22568 34353
0 14894 7 1 2 36315 14893
0 14895 7 1 2 36280 14894
0 14896 5 1 1 14895
0 14897 7 1 2 14892 14896
0 14898 7 1 2 14876 14897
0 14899 5 1 1 14898
0 14900 7 1 2 32977 14899
0 14901 5 1 1 14900
0 14902 7 2 2 26029 35129
0 14903 7 1 2 23556 35946
0 14904 7 1 2 34765 14903
0 14905 7 1 2 26719 14904
0 14906 7 1 2 36334 14905
0 14907 5 1 1 14906
0 14908 7 1 2 14901 14907
0 14909 7 1 2 14854 14908
0 14910 5 1 1 14909
0 14911 7 1 2 28110 14910
0 14912 5 1 1 14911
0 14913 7 1 2 14798 14912
0 14914 7 1 2 14668 14913
0 14915 5 1 1 14914
0 14916 7 1 2 22082 14915
0 14917 5 1 1 14916
0 14918 7 1 2 27273 35154
0 14919 5 1 1 14918
0 14920 7 1 2 26982 35143
0 14921 5 1 1 14920
0 14922 7 1 2 14919 14921
0 14923 5 1 1 14922
0 14924 7 1 2 31135 14923
0 14925 5 1 1 14924
0 14926 7 1 2 25192 30552
0 14927 5 1 1 14926
0 14928 7 1 2 31577 14927
0 14929 5 1 1 14928
0 14930 7 1 2 24110 14929
0 14931 5 1 1 14930
0 14932 7 2 2 25093 26156
0 14933 5 1 1 36336
0 14934 7 1 2 12284 14933
0 14935 5 1 1 14934
0 14936 7 1 2 23855 25821
0 14937 7 1 2 14935 14936
0 14938 5 1 1 14937
0 14939 7 1 2 14931 14938
0 14940 5 1 1 14939
0 14941 7 1 2 35155 14940
0 14942 5 1 1 14941
0 14943 7 1 2 22676 34729
0 14944 5 1 1 14943
0 14945 7 1 2 35749 35144
0 14946 7 1 2 14944 14945
0 14947 5 1 1 14946
0 14948 7 1 2 14942 14947
0 14949 7 1 2 14925 14948
0 14950 5 1 1 14949
0 14951 7 1 2 25273 14950
0 14952 5 1 1 14951
0 14953 7 1 2 33205 36018
0 14954 7 1 2 34734 14953
0 14955 5 1 1 14954
0 14956 7 1 2 14952 14955
0 14957 5 1 1 14956
0 14958 7 1 2 23557 14957
0 14959 5 1 1 14958
0 14960 7 1 2 36178 32240
0 14961 7 1 2 36203 14960
0 14962 5 1 1 14961
0 14963 7 1 2 14959 14962
0 14964 5 1 1 14963
0 14965 7 1 2 25864 14964
0 14966 5 1 1 14965
0 14967 7 1 2 23128 36033
0 14968 7 2 2 36219 14967
0 14969 7 1 2 24111 28835
0 14970 7 1 2 36338 14969
0 14971 5 1 1 14970
0 14972 7 1 2 14966 14971
0 14973 5 1 1 14972
0 14974 7 1 2 33326 14973
0 14975 5 1 1 14974
0 14976 7 1 2 24112 33516
0 14977 7 1 2 36339 14976
0 14978 5 1 1 14977
0 14979 7 1 2 14975 14978
0 14980 5 1 1 14979
0 14981 7 1 2 23669 14980
0 14982 5 1 1 14981
0 14983 7 1 2 26871 35535
0 14984 5 1 1 14983
0 14985 7 1 2 35984 34023
0 14986 7 1 2 33790 14985
0 14987 5 1 1 14986
0 14988 7 1 2 14984 14987
0 14989 5 1 1 14988
0 14990 7 1 2 28836 14989
0 14991 5 1 1 14990
0 14992 7 1 2 23317 28268
0 14993 7 1 2 28914 33372
0 14994 7 1 2 35212 34516
0 14995 7 1 2 14993 14994
0 14996 7 1 2 14992 14995
0 14997 5 1 1 14996
0 14998 7 1 2 34539 35516
0 14999 7 1 2 26872 14998
0 15000 5 1 1 14999
0 15001 7 1 2 14997 15000
0 15002 7 1 2 14991 15001
0 15003 5 1 1 15002
0 15004 7 1 2 29726 15003
0 15005 5 1 1 15004
0 15006 7 1 2 26776 26451
0 15007 7 1 2 28562 15006
0 15008 5 1 1 15007
0 15009 7 1 2 26944 29851
0 15010 7 1 2 36197 15009
0 15011 5 1 1 15010
0 15012 7 1 2 15008 15011
0 15013 5 1 1 15012
0 15014 7 1 2 23466 15013
0 15015 5 1 1 15014
0 15016 7 2 2 30499 31250
0 15017 5 1 1 36340
0 15018 7 1 2 23019 26936
0 15019 5 1 1 15018
0 15020 7 1 2 15017 15019
0 15021 5 1 1 15020
0 15022 7 1 2 22228 15021
0 15023 5 1 1 15022
0 15024 7 1 2 26879 36207
0 15025 5 1 1 15024
0 15026 7 1 2 15023 15025
0 15027 5 1 1 15026
0 15028 7 1 2 26799 15027
0 15029 5 1 1 15028
0 15030 7 1 2 15015 15029
0 15031 5 1 1 15030
0 15032 7 1 2 33737 15031
0 15033 5 1 1 15032
0 15034 7 1 2 32911 32479
0 15035 7 1 2 33529 15034
0 15036 5 1 1 15035
0 15037 7 2 2 34178 35478
0 15038 7 1 2 23020 29974
0 15039 7 1 2 36342 15038
0 15040 5 1 1 15039
0 15041 7 1 2 15036 15040
0 15042 5 1 1 15041
0 15043 7 1 2 26515 15042
0 15044 5 1 1 15043
0 15045 7 1 2 28363 32978
0 15046 7 1 2 35694 35231
0 15047 7 1 2 15045 15046
0 15048 5 1 1 15047
0 15049 7 1 2 15044 15048
0 15050 5 1 1 15049
0 15051 7 1 2 24243 15050
0 15052 5 1 1 15051
0 15053 7 1 2 25416 14378
0 15054 5 1 1 15053
0 15055 7 2 2 26740 34281
0 15056 5 1 1 36344
0 15057 7 1 2 15054 15056
0 15058 5 1 1 15057
0 15059 7 2 2 24342 24763
0 15060 7 1 2 36346 33454
0 15061 7 1 2 32402 15060
0 15062 7 1 2 15058 15061
0 15063 5 1 1 15062
0 15064 7 1 2 15052 15063
0 15065 7 1 2 15033 15064
0 15066 5 1 1 15065
0 15067 7 1 2 27147 15066
0 15068 5 1 1 15067
0 15069 7 1 2 15005 15068
0 15070 5 1 1 15069
0 15071 7 1 2 31442 35627
0 15072 7 1 2 15070 15071
0 15073 5 1 1 15072
0 15074 7 1 2 14982 15073
0 15075 5 1 1 15074
0 15076 7 1 2 26212 15075
0 15077 5 1 1 15076
0 15078 7 1 2 36341 33568
0 15079 5 1 1 15078
0 15080 7 1 2 26937 33694
0 15081 5 1 1 15080
0 15082 7 1 2 15079 15081
0 15083 5 1 1 15082
0 15084 7 1 2 25417 15083
0 15085 5 1 1 15084
0 15086 7 1 2 36345 33569
0 15087 5 1 1 15086
0 15088 7 1 2 15085 15087
0 15089 5 1 1 15088
0 15090 7 1 2 23021 15089
0 15091 5 1 1 15090
0 15092 7 2 2 23558 26873
0 15093 7 1 2 36119 36348
0 15094 5 1 1 15093
0 15095 7 1 2 15091 15094
0 15096 5 1 1 15095
0 15097 7 1 2 27148 15096
0 15098 5 1 1 15097
0 15099 7 1 2 34615 33660
0 15100 7 1 2 36349 15099
0 15101 5 1 1 15100
0 15102 7 1 2 15098 15101
0 15103 5 1 1 15102
0 15104 7 1 2 22229 15103
0 15105 5 1 1 15104
0 15106 7 1 2 36173 32773
0 15107 5 1 1 15106
0 15108 7 1 2 25418 36208
0 15109 7 1 2 33695 15108
0 15110 5 1 1 15109
0 15111 7 1 2 15107 15110
0 15112 5 1 1 15111
0 15113 7 1 2 27149 26880
0 15114 7 1 2 15112 15113
0 15115 5 1 1 15114
0 15116 7 1 2 15105 15115
0 15117 5 1 1 15116
0 15118 7 1 2 27564 31443
0 15119 7 1 2 15117 15118
0 15120 5 1 1 15119
0 15121 7 1 2 15077 15120
0 15122 5 1 1 15121
0 15123 7 1 2 24659 15122
0 15124 5 1 1 15123
0 15125 7 2 2 26438 29316
0 15126 7 1 2 36164 36350
0 15127 7 1 2 36115 35557
0 15128 7 1 2 15126 15127
0 15129 7 1 2 35156 15128
0 15130 5 1 1 15129
0 15131 7 1 2 15124 15130
0 15132 5 1 1 15131
0 15133 7 1 2 24170 15132
0 15134 5 1 1 15133
0 15135 7 1 2 26881 27008
0 15136 7 1 2 36299 33404
0 15137 7 1 2 15135 15136
0 15138 7 1 2 25193 28259
0 15139 7 1 2 36269 15138
0 15140 7 1 2 36351 32786
0 15141 7 1 2 15139 15140
0 15142 7 1 2 15137 15141
0 15143 5 1 1 15142
0 15144 7 1 2 15134 15143
0 15145 5 1 1 15144
0 15146 7 1 2 29602 15145
0 15147 5 1 1 15146
0 15148 7 1 2 27150 35159
0 15149 5 1 1 15148
0 15150 7 1 2 28610 30738
0 15151 5 1 1 15150
0 15152 7 1 2 30544 15151
0 15153 5 1 1 15152
0 15154 7 1 2 28430 33327
0 15155 7 1 2 15153 15154
0 15156 5 1 1 15155
0 15157 7 1 2 15149 15156
0 15158 5 1 1 15157
0 15159 7 1 2 35157 15158
0 15160 5 1 1 15159
0 15161 7 1 2 29229 11490
0 15162 5 2 1 15161
0 15163 7 1 2 21833 32393
0 15164 5 1 1 15163
0 15165 7 2 2 36352 15164
0 15166 5 1 1 36354
0 15167 7 1 2 22334 36355
0 15168 5 1 1 15167
0 15169 7 1 2 25511 32815
0 15170 5 1 1 15169
0 15171 7 1 2 15168 15170
0 15172 5 1 1 15171
0 15173 7 1 2 33328 15172
0 15174 5 1 1 15173
0 15175 7 1 2 27151 33689
0 15176 5 1 1 15175
0 15177 7 1 2 15174 15176
0 15178 5 1 1 15177
0 15179 7 1 2 34855 34254
0 15180 7 1 2 15178 15179
0 15181 5 1 1 15180
0 15182 7 1 2 15160 15181
0 15183 5 1 1 15182
0 15184 7 1 2 23670 15183
0 15185 5 1 1 15184
0 15186 7 1 2 26924 31863
0 15187 7 1 2 32799 15186
0 15188 7 1 2 33749 15187
0 15189 5 1 1 15188
0 15190 7 1 2 15185 15189
0 15191 5 1 1 15190
0 15192 7 1 2 26973 15191
0 15193 5 1 1 15192
0 15194 7 3 2 25419 33217
0 15195 5 1 1 36356
0 15196 7 1 2 35152 15195
0 15197 5 4 1 15196
0 15198 7 1 2 29200 35183
0 15199 7 1 2 36359 15198
0 15200 5 1 1 15199
0 15201 7 1 2 15193 15200
0 15202 5 1 1 15201
0 15203 7 1 2 22937 15202
0 15204 5 1 1 15203
0 15205 7 2 2 24482 22814
0 15206 7 1 2 31172 36363
0 15207 7 1 2 32045 15206
0 15208 7 2 2 23856 22268
0 15209 7 2 2 36365 31961
0 15210 7 1 2 24867 27235
0 15211 7 1 2 30593 15210
0 15212 7 1 2 36367 15211
0 15213 7 1 2 15207 15212
0 15214 5 1 1 15213
0 15215 7 1 2 15204 15214
0 15216 5 1 1 15215
0 15217 7 1 2 22409 15216
0 15218 5 1 1 15217
0 15219 7 1 2 27236 33616
0 15220 7 1 2 35690 15219
0 15221 7 2 2 22772 29399
0 15222 7 1 2 26492 26462
0 15223 7 1 2 36368 15222
0 15224 7 1 2 36369 15223
0 15225 7 1 2 15220 15224
0 15226 5 1 1 15225
0 15227 7 1 2 15218 15226
0 15228 5 1 1 15227
0 15229 7 1 2 26991 35225
0 15230 7 1 2 15228 15229
0 15231 5 1 1 15230
0 15232 7 1 2 15147 15231
0 15233 7 1 2 14917 15232
0 15234 7 1 2 14414 15233
0 15235 5 1 1 15234
0 15236 7 1 2 23766 15235
0 15237 5 1 1 15236
0 15238 7 2 2 25712 26227
0 15239 7 1 2 24244 33166
0 15240 5 1 1 15239
0 15241 7 1 2 30863 33198
0 15242 5 1 1 15241
0 15243 7 1 2 15240 15242
0 15244 5 1 1 15243
0 15245 7 1 2 31654 15244
0 15246 5 1 1 15245
0 15247 7 1 2 26577 28647
0 15248 7 1 2 31885 15247
0 15249 5 1 1 15248
0 15250 7 1 2 15246 15249
0 15251 5 1 1 15250
0 15252 7 1 2 21947 15251
0 15253 5 1 1 15252
0 15254 7 4 2 22773 25512
0 15255 7 5 2 24971 25420
0 15256 7 2 2 36373 36377
0 15257 7 1 2 26591 29407
0 15258 7 1 2 36382 15257
0 15259 5 1 1 15258
0 15260 7 1 2 15253 15259
0 15261 5 1 1 15260
0 15262 7 1 2 26662 15261
0 15263 5 1 1 15262
0 15264 7 2 2 30031 33218
0 15265 5 1 1 36384
0 15266 7 1 2 22230 33167
0 15267 5 1 1 15266
0 15268 7 1 2 15265 15267
0 15269 5 1 1 15268
0 15270 7 1 2 31655 36316
0 15271 7 1 2 15269 15270
0 15272 5 1 1 15271
0 15273 7 1 2 15263 15272
0 15274 5 1 1 15273
0 15275 7 1 2 22486 15274
0 15276 5 1 1 15275
0 15277 7 1 2 26777 31649
0 15278 7 2 2 30831 15277
0 15279 7 1 2 29516 36386
0 15280 5 1 1 15279
0 15281 7 1 2 15276 15280
0 15282 5 1 1 15281
0 15283 7 1 2 21834 15282
0 15284 5 1 1 15283
0 15285 7 1 2 30446 32840
0 15286 5 1 1 15285
0 15287 7 1 2 36387 15286
0 15288 5 1 1 15287
0 15289 7 1 2 15284 15288
0 15290 5 1 1 15289
0 15291 7 1 2 23318 15290
0 15292 5 1 1 15291
0 15293 7 3 2 22711 26950
0 15294 5 1 1 36388
0 15295 7 1 2 759 15294
0 15296 5 27 1 15295
0 15297 7 1 2 36391 33168
0 15298 5 1 1 15297
0 15299 7 10 2 22712 35863
0 15300 7 3 2 32955 36418
0 15301 7 1 2 30864 36428
0 15302 5 1 1 15301
0 15303 7 2 2 15298 15302
0 15304 5 1 1 36431
0 15305 7 1 2 26548 36385
0 15306 5 1 1 15305
0 15307 7 1 2 36432 15306
0 15308 5 2 1 15307
0 15309 7 1 2 25274 27152
0 15310 7 1 2 28988 30891
0 15311 7 2 2 15309 15310
0 15312 7 1 2 36433 36435
0 15313 5 1 1 15312
0 15314 7 1 2 15292 15313
0 15315 5 1 1 15314
0 15316 7 1 2 26120 15315
0 15317 5 1 1 15316
0 15318 7 2 2 29839 35760
0 15319 7 3 2 28450 36437
0 15320 5 2 1 36439
0 15321 7 1 2 33244 36440
0 15322 5 1 1 15321
0 15323 7 1 2 29118 31524
0 15324 5 1 1 15323
0 15325 7 1 2 22487 15324
0 15326 5 1 1 15325
0 15327 7 1 2 33063 15326
0 15328 5 2 1 15327
0 15329 7 6 2 23319 36444
0 15330 5 1 1 36446
0 15331 7 2 2 25347 36447
0 15332 7 1 2 25758 36452
0 15333 5 1 1 15332
0 15334 7 1 2 15322 15333
0 15335 5 1 1 15334
0 15336 7 1 2 26549 15335
0 15337 5 1 1 15336
0 15338 7 2 2 28451 33238
0 15339 7 1 2 25807 28989
0 15340 7 1 2 36389 15339
0 15341 7 1 2 36454 15340
0 15342 5 1 1 15341
0 15343 7 1 2 15337 15342
0 15344 5 1 1 15343
0 15345 7 1 2 32480 34953
0 15346 7 1 2 15344 15345
0 15347 5 1 1 15346
0 15348 7 1 2 15317 15347
0 15349 5 1 1 15348
0 15350 7 1 2 36371 15349
0 15351 5 1 1 15350
0 15352 7 1 2 34767 33838
0 15353 5 1 1 15352
0 15354 7 2 2 35110 34710
0 15355 7 1 2 30977 36456
0 15356 5 1 1 15355
0 15357 7 1 2 15353 15356
0 15358 5 1 1 15357
0 15359 7 1 2 36392 15358
0 15360 5 1 1 15359
0 15361 7 1 2 23320 33135
0 15362 5 1 1 15361
0 15363 7 1 2 28461 36438
0 15364 5 1 1 15363
0 15365 7 1 2 15362 15364
0 15366 5 4 1 15365
0 15367 7 1 2 32956 36458
0 15368 5 1 1 15367
0 15369 7 1 2 30036 30054
0 15370 5 1 1 15369
0 15371 7 1 2 21948 15370
0 15372 5 1 1 15371
0 15373 7 1 2 3266 15372
0 15374 5 1 1 15373
0 15375 7 1 2 22774 27931
0 15376 7 1 2 15374 15375
0 15377 5 1 1 15376
0 15378 7 1 2 15368 15377
0 15379 5 2 1 15378
0 15380 7 1 2 36319 36462
0 15381 5 1 1 15380
0 15382 7 1 2 15360 15381
0 15383 5 1 1 15382
0 15384 7 1 2 34062 15383
0 15385 5 1 1 15384
0 15386 7 2 2 34161 36448
0 15387 7 3 2 26663 34896
0 15388 5 1 1 36466
0 15389 7 1 2 36467 35669
0 15390 7 1 2 36464 15389
0 15391 5 1 1 15390
0 15392 7 1 2 15385 15391
0 15393 5 1 1 15392
0 15394 7 1 2 24400 15393
0 15395 5 1 1 15394
0 15396 7 2 2 28232 35864
0 15397 7 1 2 25886 33373
0 15398 7 2 2 36469 15397
0 15399 7 1 2 36471 36465
0 15400 5 1 1 15399
0 15401 7 1 2 15395 15400
0 15402 5 1 1 15401
0 15403 7 1 2 23671 15402
0 15404 5 1 1 15403
0 15405 7 7 2 34299 36393
0 15406 5 1 1 36473
0 15407 7 1 2 27009 34837
0 15408 5 1 1 15407
0 15409 7 2 2 25275 29145
0 15410 7 1 2 23857 32695
0 15411 7 1 2 36480 15410
0 15412 5 1 1 15411
0 15413 7 1 2 15408 15412
0 15414 5 1 1 15413
0 15415 7 1 2 23022 15414
0 15416 5 1 1 15415
0 15417 7 1 2 26409 36445
0 15418 5 1 1 15417
0 15419 7 1 2 34839 15418
0 15420 5 1 1 15419
0 15421 7 1 2 23321 15420
0 15422 5 1 1 15421
0 15423 7 1 2 15416 15422
0 15424 5 1 1 15423
0 15425 7 1 2 24401 15424
0 15426 5 1 1 15425
0 15427 7 1 2 36442 15330
0 15428 5 2 1 15427
0 15429 7 2 2 23672 36482
0 15430 7 1 2 25887 36484
0 15431 5 1 1 15430
0 15432 7 1 2 15426 15431
0 15433 5 1 1 15432
0 15434 7 1 2 34143 15433
0 15435 5 1 1 15434
0 15436 7 1 2 35473 36449
0 15437 5 1 1 15436
0 15438 7 1 2 15435 15437
0 15439 5 1 1 15438
0 15440 7 1 2 36474 15439
0 15441 5 1 1 15440
0 15442 7 5 2 26664 31633
0 15443 5 4 1 36486
0 15444 7 1 2 14856 36491
0 15445 5 4 1 15444
0 15446 7 1 2 26636 36459
0 15447 5 1 1 15446
0 15448 7 1 2 32469 34648
0 15449 7 1 2 34711 15448
0 15450 5 1 1 15449
0 15451 7 1 2 15447 15450
0 15452 5 1 1 15451
0 15453 7 1 2 24402 15452
0 15454 5 1 1 15453
0 15455 7 1 2 32688 36441
0 15456 5 1 1 15455
0 15457 7 1 2 15454 15456
0 15458 5 1 1 15457
0 15459 7 1 2 36495 15458
0 15460 5 1 1 15459
0 15461 7 1 2 36320 32621
0 15462 7 1 2 36450 15461
0 15463 5 1 1 15462
0 15464 7 1 2 15460 15463
0 15465 5 1 1 15464
0 15466 7 1 2 34144 15465
0 15467 5 1 1 15466
0 15468 7 2 2 22153 34906
0 15469 7 3 2 22713 22815
0 15470 7 1 2 24403 36501
0 15471 7 2 2 36499 15470
0 15472 7 1 2 25513 32075
0 15473 7 1 2 36504 15472
0 15474 7 1 2 36485 15473
0 15475 5 1 1 15474
0 15476 7 1 2 15467 15475
0 15477 5 1 1 15476
0 15478 7 1 2 32979 15477
0 15479 5 1 1 15478
0 15480 7 1 2 15441 15479
0 15481 7 1 2 15404 15480
0 15482 7 1 2 15351 15481
0 15483 5 1 1 15482
0 15484 7 1 2 28837 15483
0 15485 5 1 1 15484
0 15486 7 1 2 26550 28537
0 15487 5 1 1 15486
0 15488 7 1 2 1013 15487
0 15489 5 8 1 15488
0 15490 7 1 2 36460 34134
0 15491 5 1 1 15490
0 15492 7 1 2 25713 29097
0 15493 7 1 2 33070 15492
0 15494 7 1 2 30911 15493
0 15495 5 1 1 15494
0 15496 7 1 2 15491 15495
0 15497 5 1 1 15496
0 15498 7 1 2 36506 15497
0 15499 5 1 1 15498
0 15500 7 5 2 22714 22775
0 15501 5 1 1 36514
0 15502 7 7 2 35865 36515
0 15503 7 2 2 29431 30705
0 15504 5 1 1 36526
0 15505 7 1 2 33856 36527
0 15506 5 1 1 15505
0 15507 7 1 2 30944 33857
0 15508 5 1 1 15507
0 15509 7 1 2 23987 29628
0 15510 5 1 1 15509
0 15511 7 1 2 29531 15510
0 15512 5 1 1 15511
0 15513 7 1 2 36020 15512
0 15514 5 1 1 15513
0 15515 7 1 2 15508 15514
0 15516 5 1 1 15515
0 15517 7 1 2 22569 15516
0 15518 5 1 1 15517
0 15519 7 1 2 15506 15518
0 15520 5 1 1 15519
0 15521 7 1 2 24288 15520
0 15522 5 1 1 15521
0 15523 7 1 2 29701 34722
0 15524 7 1 2 31656 34584
0 15525 7 1 2 15523 15524
0 15526 5 1 1 15525
0 15527 7 1 2 15522 15526
0 15528 5 1 1 15527
0 15529 7 1 2 23322 15528
0 15530 5 1 1 15529
0 15531 7 3 2 28300 33374
0 15532 5 1 1 36528
0 15533 7 1 2 23559 35501
0 15534 5 1 1 15533
0 15535 7 1 2 15532 15534
0 15536 5 1 1 15535
0 15537 7 1 2 36436 15536
0 15538 5 1 1 15537
0 15539 7 1 2 15530 15538
0 15540 5 1 1 15539
0 15541 7 1 2 36519 15540
0 15542 5 1 1 15541
0 15543 7 1 2 15499 15542
0 15544 5 1 1 15543
0 15545 7 1 2 23382 15544
0 15546 5 1 1 15545
0 15547 7 2 2 26665 28538
0 15548 5 2 1 36531
0 15549 7 1 2 761 36533
0 15550 5 5 1 15549
0 15551 7 1 2 35502 36535
0 15552 5 1 1 15551
0 15553 7 1 2 36321 36008
0 15554 5 1 1 15553
0 15555 7 1 2 15552 15554
0 15556 5 1 1 15555
0 15557 7 1 2 26925 36461
0 15558 7 1 2 15556 15557
0 15559 5 1 1 15558
0 15560 7 1 2 15546 15559
0 15561 5 1 1 15560
0 15562 7 1 2 33078 15561
0 15563 5 1 1 15562
0 15564 7 2 2 22269 22776
0 15565 7 3 2 26926 36540
0 15566 5 1 1 36542
0 15567 7 2 2 32912 34122
0 15568 5 1 1 36545
0 15569 7 1 2 15566 15568
0 15570 5 3 1 15569
0 15571 7 1 2 36547 36451
0 15572 5 1 1 15571
0 15573 7 1 2 26452 34723
0 15574 7 1 2 36457 15573
0 15575 5 1 1 15574
0 15576 7 1 2 15572 15575
0 15577 5 1 1 15576
0 15578 7 1 2 34585 15577
0 15579 5 1 1 15578
0 15580 7 2 2 31262 35460
0 15581 5 1 1 36550
0 15582 7 1 2 36551 36481
0 15583 5 1 1 15582
0 15584 7 1 2 33972 33804
0 15585 7 1 2 35926 15584
0 15586 5 1 1 15585
0 15587 7 1 2 15583 15586
0 15588 5 1 1 15587
0 15589 7 1 2 36546 15588
0 15590 5 1 1 15589
0 15591 7 1 2 15579 15590
0 15592 5 1 1 15591
0 15593 7 1 2 36394 15592
0 15594 5 1 1 15593
0 15595 7 25 2 24660 35853
0 15596 7 2 2 33973 34123
0 15597 7 1 2 36552 36577
0 15598 7 1 2 36463 15597
0 15599 5 1 1 15598
0 15600 7 2 2 26666 33455
0 15601 5 1 1 36579
0 15602 7 1 2 26551 34377
0 15603 5 1 1 15602
0 15604 7 1 2 15601 15603
0 15605 5 6 1 15604
0 15606 7 2 2 33858 36581
0 15607 5 1 1 36587
0 15608 7 2 2 36553 34124
0 15609 5 1 1 36589
0 15610 7 1 2 34109 36590
0 15611 5 1 1 15610
0 15612 7 3 2 15607 15611
0 15613 7 2 2 23560 36419
0 15614 7 2 2 36594 35497
0 15615 5 1 1 36596
0 15616 7 1 2 22816 36443
0 15617 5 1 1 15616
0 15618 7 1 2 36597 15617
0 15619 5 1 1 15618
0 15620 7 1 2 36591 15619
0 15621 5 1 1 15620
0 15622 7 1 2 32980 15621
0 15623 5 1 1 15622
0 15624 7 1 2 22270 32913
0 15625 5 1 1 15624
0 15626 7 1 2 24289 31173
0 15627 5 2 1 15626
0 15628 7 1 2 15625 36598
0 15629 5 3 1 15628
0 15630 7 2 2 33859 36600
0 15631 5 1 1 36603
0 15632 7 1 2 36395 36604
0 15633 5 1 1 15632
0 15634 7 1 2 15623 15633
0 15635 5 1 1 15634
0 15636 7 1 2 36483 15635
0 15637 5 1 1 15636
0 15638 7 9 2 22271 36420
0 15639 7 1 2 33617 31889
0 15640 7 3 2 36605 15639
0 15641 7 1 2 36614 36453
0 15642 5 1 1 15641
0 15643 7 1 2 15637 15642
0 15644 7 1 2 15599 15643
0 15645 7 1 2 15594 15644
0 15646 5 1 1 15645
0 15647 7 1 2 33040 15646
0 15648 5 1 1 15647
0 15649 7 1 2 15563 15648
0 15650 7 1 2 15485 15649
0 15651 5 1 1 15650
0 15652 7 1 2 22083 15651
0 15653 5 1 1 15652
0 15654 7 2 2 30073 32731
0 15655 7 2 2 26667 31896
0 15656 7 1 2 36617 36619
0 15657 5 1 1 15656
0 15658 7 2 2 26552 28269
0 15659 7 2 2 36621 31985
0 15660 5 1 1 36623
0 15661 7 1 2 27526 36624
0 15662 5 1 1 15661
0 15663 7 1 2 15657 15662
0 15664 5 2 1 15663
0 15665 7 1 2 33375 36625
0 15666 5 1 1 15665
0 15667 7 3 2 27527 36322
0 15668 5 1 1 36627
0 15669 7 1 2 36628 35251
0 15670 5 1 1 15669
0 15671 7 1 2 15666 15670
0 15672 5 1 1 15671
0 15673 7 1 2 24715 15672
0 15674 5 1 1 15673
0 15675 7 2 2 26599 36396
0 15676 5 1 1 36630
0 15677 7 1 2 35009 36631
0 15678 5 1 1 15677
0 15679 7 1 2 15674 15678
0 15680 5 1 1 15679
0 15681 7 1 2 24868 15680
0 15682 5 1 1 15681
0 15683 7 1 2 24716 36629
0 15684 5 1 1 15683
0 15685 7 1 2 15676 15684
0 15686 5 1 1 15685
0 15687 7 3 2 23673 15686
0 15688 7 1 2 34195 36632
0 15689 5 1 1 15688
0 15690 7 1 2 15682 15689
0 15691 5 1 1 15690
0 15692 7 1 2 24404 15691
0 15693 5 1 1 15692
0 15694 7 1 2 34213 36633
0 15695 5 1 1 15694
0 15696 7 1 2 15693 15695
0 15697 5 1 1 15696
0 15698 7 1 2 25348 15697
0 15699 5 1 1 15698
0 15700 7 3 2 24405 36421
0 15701 7 1 2 25772 28915
0 15702 7 1 2 36343 15701
0 15703 7 1 2 35628 15702
0 15704 7 1 2 36635 15703
0 15705 5 1 1 15704
0 15706 7 1 2 15699 15705
0 15707 5 1 1 15706
0 15708 7 1 2 21949 15707
0 15709 5 1 1 15708
0 15710 7 3 2 26953 36516
0 15711 7 1 2 29800 36638
0 15712 5 2 1 15711
0 15713 7 1 2 29801 31638
0 15714 5 2 1 15713
0 15715 7 1 2 30912 35086
0 15716 5 1 1 15715
0 15717 7 1 2 36643 15716
0 15718 5 1 1 15717
0 15719 7 1 2 26553 15718
0 15720 5 1 1 15719
0 15721 7 1 2 36641 15720
0 15722 5 1 1 15721
0 15723 7 1 2 34222 15722
0 15724 5 1 1 15723
0 15725 7 5 2 22715 24764
0 15726 7 2 2 27066 36645
0 15727 7 2 2 34964 36650
0 15728 7 2 2 27575 35866
0 15729 7 1 2 35039 34017
0 15730 7 1 2 36654 15729
0 15731 7 1 2 36652 15730
0 15732 5 1 1 15731
0 15733 7 1 2 15724 15732
0 15734 5 1 1 15733
0 15735 7 1 2 25349 15734
0 15736 5 1 1 15735
0 15737 7 1 2 15709 15736
0 15738 5 1 1 15737
0 15739 7 1 2 25514 15738
0 15740 5 1 1 15739
0 15741 7 1 2 28367 31729
0 15742 5 1 1 15741
0 15743 7 1 2 23988 31983
0 15744 5 1 1 15743
0 15745 7 1 2 15742 15744
0 15746 5 1 1 15745
0 15747 7 1 2 21835 15746
0 15748 5 1 1 15747
0 15749 7 1 2 25759 36618
0 15750 5 1 1 15749
0 15751 7 1 2 27528 31979
0 15752 5 1 1 15751
0 15753 7 1 2 15750 15752
0 15754 5 1 1 15753
0 15755 7 1 2 21950 15754
0 15756 5 1 1 15755
0 15757 7 1 2 23989 31730
0 15758 7 1 2 31989 15757
0 15759 5 1 1 15758
0 15760 7 1 2 15756 15759
0 15761 7 1 2 15748 15760
0 15762 5 1 1 15761
0 15763 7 1 2 26554 15762
0 15764 5 1 1 15763
0 15765 7 1 2 36532 31986
0 15766 7 1 2 30928 15765
0 15767 5 1 1 15766
0 15768 7 1 2 15764 15767
0 15769 5 1 1 15768
0 15770 7 1 2 24343 15769
0 15771 5 1 1 15770
0 15772 7 1 2 28619 28930
0 15773 7 1 2 36536 15772
0 15774 7 1 2 30929 15773
0 15775 5 1 1 15774
0 15776 7 1 2 15771 15775
0 15777 5 1 1 15776
0 15778 7 1 2 25515 15777
0 15779 5 1 1 15778
0 15780 7 1 2 26087 32607
0 15781 5 1 1 15780
0 15782 7 1 2 7509 15781
0 15783 5 1 1 15782
0 15784 7 1 2 31604 36397
0 15785 7 1 2 15783 15784
0 15786 5 1 1 15785
0 15787 7 1 2 15779 15786
0 15788 5 1 1 15787
0 15789 7 1 2 25350 15788
0 15790 5 1 1 15789
0 15791 7 2 2 24717 36398
0 15792 7 1 2 32451 36656
0 15793 5 1 1 15792
0 15794 7 2 2 22777 36554
0 15795 7 1 2 29034 36658
0 15796 5 1 1 15795
0 15797 7 1 2 15793 15796
0 15798 5 1 1 15797
0 15799 7 1 2 30848 15798
0 15800 5 1 1 15799
0 15801 7 1 2 29165 30913
0 15802 7 1 2 36657 15801
0 15803 5 1 1 15802
0 15804 7 1 2 15800 15803
0 15805 5 1 1 15804
0 15806 7 1 2 25610 15805
0 15807 5 1 1 15806
0 15808 7 4 2 23674 36399
0 15809 7 1 2 26876 33817
0 15810 7 1 2 36660 15809
0 15811 5 1 1 15810
0 15812 7 1 2 15807 15811
0 15813 5 1 1 15812
0 15814 7 1 2 28916 15813
0 15815 5 1 1 15814
0 15816 7 1 2 26121 15815
0 15817 7 1 2 15790 15816
0 15818 5 1 1 15817
0 15819 7 3 2 36400 32926
0 15820 5 1 1 36664
0 15821 7 1 2 24819 36665
0 15822 5 1 1 15821
0 15823 7 7 2 25760 26555
0 15824 7 2 2 26927 36667
0 15825 7 1 2 32046 36674
0 15826 5 1 1 15825
0 15827 7 1 2 15822 15826
0 15828 5 1 1 15827
0 15829 7 1 2 24344 15828
0 15830 5 1 1 15829
0 15831 7 1 2 26556 34159
0 15832 5 1 1 15831
0 15833 7 1 2 15830 15832
0 15834 5 1 1 15833
0 15835 7 1 2 32643 15834
0 15836 5 1 1 15835
0 15837 7 1 2 26136 15836
0 15838 5 1 1 15837
0 15839 7 1 2 36372 15838
0 15840 7 1 2 15818 15839
0 15841 5 1 1 15840
0 15842 7 1 2 36555 35509
0 15843 5 1 1 15842
0 15844 7 1 2 33376 36487
0 15845 5 1 1 15844
0 15846 7 1 2 15843 15845
0 15847 5 1 1 15846
0 15848 7 2 2 32443 15847
0 15849 7 1 2 30930 36676
0 15850 5 1 1 15849
0 15851 7 1 2 24820 35503
0 15852 5 1 1 15851
0 15853 7 1 2 33377 32047
0 15854 5 1 1 15853
0 15855 7 1 2 15852 15854
0 15856 5 1 1 15855
0 15857 7 1 2 36595 15856
0 15858 5 1 1 15857
0 15859 7 1 2 34724 35518
0 15860 5 1 1 15859
0 15861 7 1 2 29222 35507
0 15862 5 1 1 15861
0 15863 7 1 2 15860 15862
0 15864 5 1 1 15863
0 15865 7 1 2 36556 15864
0 15866 5 1 1 15865
0 15867 7 1 2 15858 15866
0 15868 5 2 1 15867
0 15869 7 1 2 30931 36678
0 15870 5 1 1 15869
0 15871 7 7 2 24290 36557
0 15872 7 2 2 28586 33974
0 15873 7 2 2 36680 36687
0 15874 7 1 2 36689 34472
0 15875 5 1 1 15874
0 15876 7 1 2 15870 15875
0 15877 5 1 1 15876
0 15878 7 1 2 24345 15877
0 15879 5 1 1 15878
0 15880 7 1 2 15850 15879
0 15881 5 1 1 15880
0 15882 7 1 2 25611 15881
0 15883 5 1 1 15882
0 15884 7 2 2 25516 32048
0 15885 7 1 2 34540 36691
0 15886 7 1 2 36606 15885
0 15887 5 2 1 15886
0 15888 7 3 2 28301 35525
0 15889 5 1 1 36695
0 15890 7 1 2 36696 36607
0 15891 5 2 1 15890
0 15892 7 1 2 26800 36646
0 15893 7 1 2 36500 15892
0 15894 5 1 1 15893
0 15895 7 1 2 36592 15894
0 15896 5 2 1 15895
0 15897 7 1 2 22874 36700
0 15898 5 1 1 15897
0 15899 7 1 2 36698 15898
0 15900 5 1 1 15899
0 15901 7 1 2 22335 15900
0 15902 5 1 1 15901
0 15903 7 1 2 36693 15902
0 15904 5 1 1 15903
0 15905 7 1 2 32644 15904
0 15906 5 1 1 15905
0 15907 7 1 2 15883 15906
0 15908 5 1 1 15907
0 15909 7 1 2 24406 15908
0 15910 5 1 1 15909
0 15911 7 1 2 25893 15910
0 15912 5 1 1 15911
0 15913 7 1 2 24821 36701
0 15914 5 1 1 15913
0 15915 7 2 2 26801 33511
0 15916 5 1 1 36702
0 15917 7 1 2 36703 36681
0 15918 5 1 1 15917
0 15919 7 1 2 15914 15918
0 15920 5 1 1 15919
0 15921 7 1 2 24346 15920
0 15922 5 1 1 15921
0 15923 7 1 2 36558 34098
0 15924 5 1 1 15923
0 15925 7 1 2 15922 15924
0 15926 5 2 1 15925
0 15927 7 1 2 36704 32645
0 15928 5 1 1 15927
0 15929 7 1 2 26137 15928
0 15930 5 1 1 15929
0 15931 7 1 2 32981 15930
0 15932 7 1 2 15912 15931
0 15933 5 1 1 15932
0 15934 7 1 2 33661 32646
0 15935 5 1 1 15934
0 15936 7 1 2 33738 32608
0 15937 5 1 1 15936
0 15938 7 1 2 15935 15937
0 15939 5 1 1 15938
0 15940 7 1 2 23561 15939
0 15941 5 1 1 15940
0 15942 7 1 2 34475 15941
0 15943 5 1 1 15942
0 15944 7 1 2 26122 15943
0 15945 5 1 1 15944
0 15946 7 1 2 33739 35404
0 15947 5 1 1 15946
0 15948 7 1 2 15945 15947
0 15949 5 1 1 15948
0 15950 7 1 2 26228 36475
0 15951 7 1 2 15949 15950
0 15952 5 1 1 15951
0 15953 7 2 2 23675 35811
0 15954 7 2 2 36706 36429
0 15955 7 1 2 32481 33805
0 15956 7 1 2 36708 15955
0 15957 5 1 1 15956
0 15958 7 1 2 15952 15957
0 15959 7 1 2 15933 15958
0 15960 7 1 2 15841 15959
0 15961 7 1 2 15740 15960
0 15962 5 1 1 15961
0 15963 7 1 2 23323 35981
0 15964 5 1 1 15963
0 15965 7 1 2 35924 15964
0 15966 5 1 1 15965
0 15967 7 1 2 15962 15966
0 15968 5 1 1 15967
0 15969 7 1 2 36286 36548
0 15970 5 1 1 15969
0 15971 7 2 2 23562 34708
0 15972 7 1 2 25276 31174
0 15973 7 1 2 36710 15972
0 15974 7 1 2 34871 15973
0 15975 5 1 1 15974
0 15976 7 1 2 15970 15975
0 15977 5 1 1 15976
0 15978 7 1 2 25094 15977
0 15979 5 1 1 15978
0 15980 7 1 2 29463 32732
0 15981 5 1 1 15980
0 15982 7 1 2 24113 28611
0 15983 5 1 1 15982
0 15984 7 1 2 15981 15983
0 15985 5 1 1 15984
0 15986 7 1 2 36543 35761
0 15987 7 1 2 15985 15986
0 15988 5 1 1 15987
0 15989 7 1 2 15979 15988
0 15990 5 1 1 15989
0 15991 7 1 2 31826 15990
0 15992 5 1 1 15991
0 15993 7 1 2 28990 31028
0 15994 5 1 1 15993
0 15995 7 1 2 25095 34889
0 15996 5 1 1 15995
0 15997 7 1 2 15994 15996
0 15998 5 1 1 15997
0 15999 7 1 2 23990 15998
0 16000 5 1 1 15999
0 16001 7 1 2 16000 6337
0 16002 5 1 1 16001
0 16003 7 1 2 23858 16002
0 16004 5 1 1 16003
0 16005 7 1 2 31535 31505
0 16006 7 1 2 32277 16005
0 16007 7 1 2 34976 16006
0 16008 5 1 1 16007
0 16009 7 1 2 16004 16008
0 16010 5 5 1 16009
0 16011 7 2 2 25947 36712
0 16012 7 2 2 25808 35368
0 16013 7 1 2 29166 36719
0 16014 7 1 2 36717 16013
0 16015 5 1 1 16014
0 16016 7 1 2 15992 16015
0 16017 5 1 1 16016
0 16018 7 1 2 23676 16017
0 16019 5 1 1 16018
0 16020 7 2 2 32914 34027
0 16021 5 1 1 36721
0 16022 7 4 2 25351 36541
0 16023 7 1 2 26088 36723
0 16024 5 1 1 16023
0 16025 7 1 2 16021 16024
0 16026 5 1 1 16025
0 16027 7 2 2 36337 34236
0 16028 7 2 2 35104 36727
0 16029 5 1 1 36729
0 16030 7 1 2 34389 36730
0 16031 7 1 2 16026 16030
0 16032 5 1 1 16031
0 16033 7 1 2 16019 16032
0 16034 5 1 1 16033
0 16035 7 1 2 34586 16034
0 16036 5 1 1 16035
0 16037 7 1 2 23677 36718
0 16038 5 1 1 16037
0 16039 7 1 2 16029 16038
0 16040 5 2 1 16039
0 16041 7 1 2 35520 36731
0 16042 5 1 1 16041
0 16043 7 2 2 23678 36713
0 16044 7 2 2 33994 34499
0 16045 7 1 2 36733 36735
0 16046 5 1 1 16045
0 16047 7 1 2 16042 16046
0 16048 5 1 1 16047
0 16049 7 1 2 23563 16048
0 16050 5 1 1 16049
0 16051 7 1 2 28648 34008
0 16052 7 1 2 31827 16051
0 16053 7 1 2 36714 16052
0 16054 5 1 1 16053
0 16055 7 1 2 16050 16054
0 16056 5 1 1 16055
0 16057 7 1 2 25277 16056
0 16058 5 1 1 16057
0 16059 7 3 2 25096 36287
0 16060 7 1 2 33860 33041
0 16061 7 1 2 36737 16060
0 16062 5 1 1 16061
0 16063 7 1 2 16058 16062
0 16064 5 1 1 16063
0 16065 7 1 2 36601 16064
0 16066 5 1 1 16065
0 16067 7 1 2 16036 16066
0 16068 5 1 1 16067
0 16069 7 1 2 36401 16068
0 16070 5 1 1 16069
0 16071 7 1 2 28991 33809
0 16072 7 1 2 35275 16071
0 16073 5 1 1 16072
0 16074 7 2 2 26123 35652
0 16075 7 1 2 27153 29876
0 16076 7 1 2 36374 16075
0 16077 7 1 2 36740 16076
0 16078 5 1 1 16077
0 16079 7 1 2 16073 16078
0 16080 5 1 1 16079
0 16081 7 1 2 25714 16080
0 16082 5 1 1 16081
0 16083 7 2 2 33329 35959
0 16084 7 1 2 28302 34168
0 16085 7 1 2 36742 16084
0 16086 7 1 2 34875 16085
0 16087 5 1 1 16086
0 16088 7 1 2 16082 16087
0 16089 5 1 1 16088
0 16090 7 1 2 24114 16089
0 16091 5 1 1 16090
0 16092 7 1 2 25352 30963
0 16093 7 1 2 35111 16092
0 16094 7 1 2 35686 16093
0 16095 7 1 2 35350 16094
0 16096 5 1 1 16095
0 16097 7 1 2 16091 16096
0 16098 5 1 1 16097
0 16099 7 1 2 25278 16098
0 16100 5 1 1 16099
0 16101 7 1 2 25948 34145
0 16102 5 1 1 16101
0 16103 7 1 2 7461 16102
0 16104 5 1 1 16103
0 16105 7 1 2 34300 16104
0 16106 7 1 2 36738 16105
0 16107 5 1 1 16106
0 16108 7 1 2 16100 16107
0 16109 5 1 1 16108
0 16110 7 1 2 36402 16109
0 16111 5 1 1 16110
0 16112 7 1 2 32158 36675
0 16113 5 2 1 16112
0 16114 7 3 2 22716 24869
0 16115 7 5 2 35867 36746
0 16116 7 1 2 36749 34225
0 16117 5 1 1 16116
0 16118 7 1 2 36744 16117
0 16119 5 1 1 16118
0 16120 7 1 2 36288 16119
0 16121 5 1 1 16120
0 16122 7 2 2 26453 30245
0 16123 7 2 2 35105 36754
0 16124 7 1 2 24718 26157
0 16125 7 1 2 36750 16124
0 16126 7 1 2 36756 16125
0 16127 5 1 1 16126
0 16128 7 1 2 16121 16127
0 16129 5 1 1 16128
0 16130 7 1 2 25715 16129
0 16131 5 1 1 16130
0 16132 7 2 2 22154 33456
0 16133 7 2 2 23564 36758
0 16134 7 2 2 28233 34047
0 16135 7 1 2 26861 36762
0 16136 7 1 2 36760 16135
0 16137 5 1 1 16136
0 16138 7 2 2 23383 30246
0 16139 7 1 2 36764 34783
0 16140 7 1 2 36659 16139
0 16141 5 1 1 16140
0 16142 7 1 2 16137 16141
0 16143 5 1 1 16142
0 16144 7 1 2 36289 16143
0 16145 5 1 1 16144
0 16146 7 1 2 26617 31543
0 16147 7 1 2 29322 16146
0 16148 7 1 2 36755 16147
0 16149 7 1 2 35134 16148
0 16150 5 1 1 16149
0 16151 7 1 2 16145 16150
0 16152 7 1 2 16131 16151
0 16153 5 1 1 16152
0 16154 7 1 2 25097 16153
0 16155 5 1 1 16154
0 16156 7 1 2 30479 33457
0 16157 7 1 2 36647 16156
0 16158 5 1 1 16157
0 16159 7 1 2 29340 36329
0 16160 7 1 2 25716 16159
0 16161 5 1 1 16160
0 16162 7 1 2 16158 16161
0 16163 5 1 1 16162
0 16164 7 5 2 23129 23565
0 16165 7 1 2 25279 28917
0 16166 7 1 2 36766 16165
0 16167 7 2 2 32637 16166
0 16168 7 1 2 22938 35112
0 16169 7 1 2 36771 16168
0 16170 7 1 2 16163 16169
0 16171 5 1 1 16170
0 16172 7 1 2 16155 16171
0 16173 5 1 1 16172
0 16174 7 1 2 24407 16173
0 16175 5 1 1 16174
0 16176 7 1 2 25809 33806
0 16177 7 1 2 35115 16176
0 16178 5 1 1 16177
0 16179 7 1 2 24719 26024
0 16180 7 1 2 30951 16179
0 16181 7 1 2 29817 16180
0 16182 5 1 1 16181
0 16183 7 1 2 16178 16182
0 16184 5 1 1 16183
0 16185 7 1 2 25717 36559
0 16186 5 1 1 16185
0 16187 7 1 2 15388 16186
0 16188 5 4 1 16187
0 16189 7 1 2 25888 32482
0 16190 7 1 2 36773 16189
0 16191 7 1 2 16184 16190
0 16192 5 1 1 16191
0 16193 7 1 2 16175 16192
0 16194 7 1 2 16111 16193
0 16195 5 1 1 16194
0 16196 7 1 2 28838 16195
0 16197 5 1 1 16196
0 16198 7 1 2 35483 36720
0 16199 7 1 2 36403 16198
0 16200 7 1 2 36715 16199
0 16201 5 1 1 16200
0 16202 7 1 2 25353 36615
0 16203 5 1 1 16202
0 16204 7 1 2 35479 36765
0 16205 7 1 2 36682 16204
0 16206 5 1 1 16205
0 16207 7 1 2 16203 16206
0 16208 5 1 1 16207
0 16209 7 1 2 36290 16208
0 16210 5 1 1 16209
0 16211 7 1 2 26158 33378
0 16212 7 1 2 36668 16211
0 16213 7 1 2 36757 16212
0 16214 5 1 1 16213
0 16215 7 1 2 16210 16214
0 16216 5 1 1 16215
0 16217 7 1 2 25098 16216
0 16218 5 1 1 16217
0 16219 7 2 2 30480 36502
0 16220 7 1 2 24542 35395
0 16221 7 1 2 36777 16220
0 16222 7 1 2 36772 16221
0 16223 5 1 1 16222
0 16224 7 1 2 16218 16223
0 16225 7 1 2 16201 16224
0 16226 5 1 1 16225
0 16227 7 1 2 31828 16226
0 16228 5 1 1 16227
0 16229 7 1 2 16197 16228
0 16230 5 1 1 16229
0 16231 7 1 2 23679 16230
0 16232 5 1 1 16231
0 16233 7 1 2 33503 36560
0 16234 5 1 1 16233
0 16235 7 5 2 22717 34907
0 16236 7 3 2 28751 36779
0 16237 5 1 1 36784
0 16238 7 1 2 16234 16237
0 16239 5 1 1 16238
0 16240 7 1 2 26802 35493
0 16241 5 1 1 16240
0 16242 7 1 2 27684 35484
0 16243 5 1 1 16242
0 16244 7 1 2 16241 16243
0 16245 5 2 1 16244
0 16246 7 1 2 24408 36787
0 16247 5 1 1 16246
0 16248 7 1 2 24870 26803
0 16249 7 1 2 35359 16248
0 16250 5 1 1 16249
0 16251 7 1 2 16247 16250
0 16252 5 1 1 16251
0 16253 7 1 2 16239 16252
0 16254 5 1 1 16253
0 16255 7 1 2 31829 36588
0 16256 5 1 1 16255
0 16257 7 1 2 15916 15889
0 16258 5 1 1 16257
0 16259 7 2 2 25949 36561
0 16260 7 1 2 34179 36789
0 16261 5 1 1 16260
0 16262 7 1 2 36751 35802
0 16263 5 1 1 16262
0 16264 7 1 2 16261 16263
0 16265 5 1 1 16264
0 16266 7 1 2 16258 16265
0 16267 5 1 1 16266
0 16268 7 1 2 16256 16267
0 16269 7 1 2 16254 16268
0 16270 5 2 1 16269
0 16271 7 3 2 23680 36791
0 16272 5 1 1 36793
0 16273 7 1 2 36794 36739
0 16274 5 1 1 16273
0 16275 7 1 2 24822 36785
0 16276 5 1 1 16275
0 16277 7 1 2 36562 34028
0 16278 5 1 1 16277
0 16279 7 1 2 16276 16278
0 16280 5 2 1 16279
0 16281 7 1 2 34587 36796
0 16282 5 1 1 16281
0 16283 7 1 2 36582 35521
0 16284 5 1 1 16283
0 16285 7 1 2 16282 16284
0 16286 5 3 1 16285
0 16287 7 1 2 36798 36732
0 16288 5 1 1 16287
0 16289 7 2 2 27692 36608
0 16290 5 1 1 36801
0 16291 7 2 2 34588 36802
0 16292 5 1 1 36803
0 16293 7 1 2 36583 36736
0 16294 5 1 1 16293
0 16295 7 1 2 16292 16294
0 16296 5 1 1 16295
0 16297 7 1 2 36734 16296
0 16298 5 1 1 16297
0 16299 7 1 2 16288 16298
0 16300 5 1 1 16299
0 16301 7 1 2 23566 16300
0 16302 5 1 1 16301
0 16303 7 1 2 31830 36774
0 16304 5 1 1 16303
0 16305 7 1 2 24871 28839
0 16306 7 1 2 36505 16305
0 16307 5 1 1 16306
0 16308 7 1 2 16304 16307
0 16309 5 2 1 16308
0 16310 7 1 2 28312 36805
0 16311 7 1 2 36716 16310
0 16312 5 1 1 16311
0 16313 7 1 2 16302 16312
0 16314 5 1 1 16313
0 16315 7 1 2 25280 16314
0 16316 5 1 1 16315
0 16317 7 1 2 16274 16316
0 16318 5 1 1 16317
0 16319 7 1 2 32982 16318
0 16320 5 1 1 16319
0 16321 7 1 2 25681 16320
0 16322 7 1 2 16232 16321
0 16323 7 1 2 16070 16322
0 16324 7 1 2 15968 16323
0 16325 7 1 2 15653 16324
0 16326 5 1 1 16325
0 16327 7 1 2 29727 32391
0 16328 5 1 1 16327
0 16329 7 1 2 29603 2565
0 16330 7 1 2 30635 16329
0 16331 5 1 1 16330
0 16332 7 1 2 16328 16331
0 16333 5 1 1 16332
0 16334 7 1 2 26410 16333
0 16335 5 1 1 16334
0 16336 7 5 2 26637 28587
0 16337 7 1 2 36807 32842
0 16338 5 1 1 16337
0 16339 7 1 2 16335 16338
0 16340 5 1 1 16339
0 16341 7 1 2 23859 16340
0 16342 5 1 1 16341
0 16343 7 1 2 26411 30636
0 16344 5 1 1 16343
0 16345 7 1 2 27312 36808
0 16346 5 1 1 16345
0 16347 7 1 2 16344 16346
0 16348 5 1 1 16347
0 16349 7 1 2 31468 16348
0 16350 5 1 1 16349
0 16351 7 1 2 24972 32394
0 16352 5 1 1 16351
0 16353 7 2 2 36353 16352
0 16354 7 1 2 26412 36812
0 16355 5 1 1 16354
0 16356 7 1 2 24115 36809
0 16357 5 1 1 16356
0 16358 7 1 2 16355 16357
0 16359 5 1 1 16358
0 16360 7 1 2 29604 16359
0 16361 5 1 1 16360
0 16362 7 1 2 16350 16361
0 16363 7 1 2 16342 16362
0 16364 5 1 1 16363
0 16365 7 1 2 24171 16364
0 16366 5 1 1 16365
0 16367 7 1 2 24172 36810
0 16368 5 1 1 16367
0 16369 7 2 2 26238 33479
0 16370 7 1 2 24483 36814
0 16371 7 1 2 35185 16370
0 16372 5 1 1 16371
0 16373 7 1 2 16368 16372
0 16374 5 1 1 16373
0 16375 7 1 2 29317 16374
0 16376 5 1 1 16375
0 16377 7 1 2 16366 16376
0 16378 5 1 1 16377
0 16379 7 1 2 22336 16378
0 16380 5 1 1 16379
0 16381 7 1 2 26638 12561
0 16382 5 1 1 16381
0 16383 7 1 2 1977 31454
0 16384 5 1 1 16383
0 16385 7 1 2 26413 16384
0 16386 5 1 1 16385
0 16387 7 1 2 16382 16386
0 16388 5 1 1 16387
0 16389 7 1 2 24173 30734
0 16390 7 1 2 16388 16389
0 16391 5 1 1 16390
0 16392 7 1 2 16380 16391
0 16393 5 1 1 16392
0 16394 7 1 2 23130 16393
0 16395 5 1 1 16394
0 16396 7 1 2 28097 31469
0 16397 5 1 1 16396
0 16398 7 1 2 26639 31184
0 16399 5 1 1 16398
0 16400 7 1 2 16397 16399
0 16401 5 1 1 16400
0 16402 7 1 2 23023 16401
0 16403 5 1 1 16402
0 16404 7 1 2 24872 30767
0 16405 5 1 1 16404
0 16406 7 1 2 26469 31185
0 16407 7 1 2 16405 16406
0 16408 5 1 1 16407
0 16409 7 1 2 16403 16408
0 16410 5 1 1 16409
0 16411 7 1 2 30713 16410
0 16412 5 1 1 16411
0 16413 7 1 2 16395 16412
0 16414 5 1 1 16413
0 16415 7 1 2 22410 16414
0 16416 5 1 1 16415
0 16417 7 1 2 28992 32676
0 16418 5 1 1 16417
0 16419 7 1 2 33159 16418
0 16420 5 1 1 16419
0 16421 7 1 2 25612 25877
0 16422 7 1 2 30714 16421
0 16423 7 1 2 16420 16422
0 16424 5 1 1 16423
0 16425 7 1 2 16416 16424
0 16426 5 1 1 16425
0 16427 7 1 2 22817 36360
0 16428 5 1 1 16427
0 16429 7 1 2 26778 35675
0 16430 5 1 1 16429
0 16431 7 1 2 16428 16430
0 16432 5 1 1 16431
0 16433 7 1 2 22272 16432
0 16434 5 1 1 16433
0 16435 7 1 2 25354 35329
0 16436 7 1 2 35317 16435
0 16437 5 1 1 16436
0 16438 7 1 2 16434 16437
0 16439 5 1 1 16438
0 16440 7 1 2 16426 16439
0 16441 5 1 1 16440
0 16442 7 1 2 29464 33277
0 16443 5 1 1 16442
0 16444 7 1 2 28125 34735
0 16445 5 1 1 16444
0 16446 7 1 2 131 16445
0 16447 5 1 1 16446
0 16448 7 1 2 26933 16447
0 16449 5 1 1 16448
0 16450 7 2 2 23467 33245
0 16451 7 1 2 14272 5226
0 16452 5 1 1 16451
0 16453 7 1 2 22939 16452
0 16454 5 1 1 16453
0 16455 7 2 2 23131 30306
0 16456 7 1 2 32081 36818
0 16457 5 1 1 16456
0 16458 7 1 2 16454 16457
0 16459 5 1 1 16458
0 16460 7 1 2 22411 16459
0 16461 5 1 1 16460
0 16462 7 5 2 28260 27676
0 16463 7 1 2 36820 36819
0 16464 5 1 1 16463
0 16465 7 1 2 16461 16464
0 16466 5 1 1 16465
0 16467 7 1 2 27529 16466
0 16468 5 1 1 16467
0 16469 7 1 2 32362 34532
0 16470 5 1 1 16469
0 16471 7 2 2 26213 29167
0 16472 7 1 2 23132 36825
0 16473 5 1 1 16472
0 16474 7 1 2 16470 16473
0 16475 5 1 1 16474
0 16476 7 1 2 25613 16475
0 16477 5 1 1 16476
0 16478 7 2 2 29179 28649
0 16479 7 1 2 22337 28378
0 16480 7 1 2 36827 16479
0 16481 5 1 1 16480
0 16482 7 1 2 16477 16481
0 16483 7 1 2 16468 16482
0 16484 5 1 1 16483
0 16485 7 1 2 36816 16484
0 16486 5 1 1 16485
0 16487 7 1 2 16449 16486
0 16488 5 1 1 16487
0 16489 7 1 2 31470 16488
0 16490 5 1 1 16489
0 16491 7 1 2 16443 16490
0 16492 5 1 1 16491
0 16493 7 1 2 25718 16492
0 16494 5 1 1 16493
0 16495 7 1 2 22084 31761
0 16496 5 5 1 16495
0 16497 7 1 2 24116 30390
0 16498 5 1 1 16497
0 16499 7 1 2 21836 16498
0 16500 5 1 1 16499
0 16501 7 2 2 36829 16500
0 16502 7 1 2 28126 36834
0 16503 5 1 1 16502
0 16504 7 1 2 749 16503
0 16505 5 1 1 16504
0 16506 7 1 2 26934 16505
0 16507 5 1 1 16506
0 16508 7 1 2 29168 32274
0 16509 5 1 1 16508
0 16510 7 1 2 24117 29035
0 16511 5 1 1 16510
0 16512 7 1 2 16509 16511
0 16513 5 1 1 16512
0 16514 7 1 2 22940 16513
0 16515 5 1 1 16514
0 16516 7 1 2 35175 35354
0 16517 5 1 1 16516
0 16518 7 1 2 16515 16517
0 16519 5 1 1 16518
0 16520 7 1 2 25614 16519
0 16521 5 1 1 16520
0 16522 7 2 2 23860 26414
0 16523 7 1 2 25865 29413
0 16524 7 1 2 36836 16523
0 16525 5 1 1 16524
0 16526 7 1 2 16521 16525
0 16527 5 1 1 16526
0 16528 7 1 2 22412 16527
0 16529 5 1 1 16528
0 16530 7 1 2 32206 36821
0 16531 5 1 1 16530
0 16532 7 1 2 16529 16531
0 16533 5 1 1 16532
0 16534 7 1 2 27313 16533
0 16535 5 1 1 16534
0 16536 7 1 2 23861 33785
0 16537 5 1 1 16536
0 16538 7 1 2 23567 33394
0 16539 5 1 1 16538
0 16540 7 1 2 16537 16539
0 16541 5 1 1 16540
0 16542 7 1 2 25615 16541
0 16543 5 1 1 16542
0 16544 7 1 2 16543 7112
0 16545 5 1 1 16544
0 16546 7 1 2 22413 16545
0 16547 5 1 1 16546
0 16548 7 2 2 23862 30307
0 16549 7 1 2 36838 36822
0 16550 5 1 1 16549
0 16551 7 1 2 16547 16550
0 16552 5 1 1 16551
0 16553 7 1 2 36830 16552
0 16554 5 1 1 16553
0 16555 7 1 2 29414 33274
0 16556 5 1 1 16555
0 16557 7 1 2 16554 16556
0 16558 7 1 2 16535 16557
0 16559 5 1 1 16558
0 16560 7 1 2 36817 16559
0 16561 5 1 1 16560
0 16562 7 1 2 16507 16561
0 16563 5 1 1 16562
0 16564 7 1 2 25719 16563
0 16565 5 1 1 16564
0 16566 7 3 2 36361 33927
0 16567 5 1 1 36840
0 16568 7 1 2 23863 32770
0 16569 5 1 1 16568
0 16570 7 1 2 6860 16569
0 16571 5 1 1 16570
0 16572 7 1 2 27314 16571
0 16573 5 1 1 16572
0 16574 7 2 2 28127 31444
0 16575 5 1 1 36843
0 16576 7 1 2 28113 6838
0 16577 5 1 1 16576
0 16578 7 1 2 36831 16577
0 16579 5 1 1 16578
0 16580 7 1 2 16575 16579
0 16581 7 1 2 16573 16580
0 16582 5 1 1 16581
0 16583 7 1 2 36841 16582
0 16584 5 1 1 16583
0 16585 7 1 2 33712 36826
0 16586 5 1 1 16585
0 16587 7 1 2 28128 34418
0 16588 5 1 1 16587
0 16589 7 1 2 16586 16588
0 16590 5 2 1 16589
0 16591 7 1 2 23864 36362
0 16592 5 1 1 16591
0 16593 7 1 2 14390 16592
0 16594 5 1 1 16593
0 16595 7 1 2 36832 16594
0 16596 5 1 1 16595
0 16597 7 1 2 24118 34822
0 16598 7 1 2 33246 16597
0 16599 5 1 1 16598
0 16600 7 1 2 34282 32275
0 16601 5 1 1 16600
0 16602 7 1 2 24119 34277
0 16603 5 1 1 16602
0 16604 7 1 2 16601 16603
0 16605 5 1 1 16604
0 16606 7 1 2 22231 16605
0 16607 5 1 1 16606
0 16608 7 1 2 24120 36357
0 16609 5 1 1 16608
0 16610 7 1 2 16607 16609
0 16611 5 1 1 16610
0 16612 7 1 2 27315 16611
0 16613 5 1 1 16612
0 16614 7 1 2 16599 16613
0 16615 7 1 2 16596 16614
0 16616 5 1 1 16615
0 16617 7 1 2 36845 16616
0 16618 5 1 1 16617
0 16619 7 1 2 28280 28030
0 16620 7 1 2 28937 34419
0 16621 7 2 2 16619 16620
0 16622 5 1 1 36847
0 16623 7 1 2 27154 36848
0 16624 5 1 1 16623
0 16625 7 1 2 16618 16624
0 16626 7 1 2 16584 16625
0 16627 7 1 2 16565 16626
0 16628 5 1 1 16627
0 16629 7 1 2 29605 16628
0 16630 5 1 1 16629
0 16631 7 1 2 22273 33845
0 16632 7 1 2 33247 16631
0 16633 5 1 1 16632
0 16634 7 1 2 16567 16633
0 16635 5 1 1 16634
0 16636 7 1 2 25990 16635
0 16637 5 1 1 16636
0 16638 7 1 2 26804 28840
0 16639 7 1 2 34462 16638
0 16640 7 1 2 33248 16639
0 16641 5 1 1 16640
0 16642 7 1 2 16637 16641
0 16643 5 1 1 16642
0 16644 7 1 2 36081 16643
0 16645 5 1 1 16644
0 16646 7 1 2 23133 27565
0 16647 5 1 1 16646
0 16648 7 1 2 129 16647
0 16649 5 1 1 16648
0 16650 7 1 2 25866 16649
0 16651 5 1 1 16650
0 16652 7 1 2 25978 28744
0 16653 5 1 1 16652
0 16654 7 1 2 16651 16653
0 16655 5 1 1 16654
0 16656 7 1 2 27530 16655
0 16657 5 1 1 16656
0 16658 7 1 2 28129 32363
0 16659 5 1 1 16658
0 16660 7 1 2 5864 16659
0 16661 7 1 2 16657 16660
0 16662 5 1 1 16661
0 16663 7 1 2 36842 16662
0 16664 5 1 1 16663
0 16665 7 1 2 28179 36001
0 16666 5 1 1 16665
0 16667 7 1 2 12847 16666
0 16668 5 1 1 16667
0 16669 7 1 2 22232 16668
0 16670 5 1 1 16669
0 16671 7 1 2 23134 36358
0 16672 5 1 1 16671
0 16673 7 1 2 16670 16672
0 16674 5 1 1 16673
0 16675 7 1 2 27531 16674
0 16676 5 1 1 16675
0 16677 7 1 2 23135 36217
0 16678 5 1 1 16677
0 16679 7 1 2 25421 32364
0 16680 7 1 2 33249 16679
0 16681 5 1 1 16680
0 16682 7 1 2 16678 16681
0 16683 7 1 2 16676 16682
0 16684 5 1 1 16683
0 16685 7 1 2 36846 16684
0 16686 5 1 1 16685
0 16687 7 1 2 16622 16686
0 16688 7 1 2 16664 16687
0 16689 5 1 1 16688
0 16690 7 1 2 31471 16689
0 16691 5 1 1 16690
0 16692 7 1 2 16645 16691
0 16693 7 1 2 16630 16692
0 16694 7 1 2 16494 16693
0 16695 5 1 1 16694
0 16696 7 1 2 24174 16695
0 16697 5 1 1 16696
0 16698 7 1 2 16441 16697
0 16699 5 1 1 16698
0 16700 7 1 2 24661 16699
0 16701 5 1 1 16700
0 16702 7 2 2 28695 33791
0 16703 7 1 2 27532 36849
0 16704 5 1 1 16703
0 16705 7 2 2 31175 32787
0 16706 7 1 2 22875 36851
0 16707 5 1 1 16706
0 16708 7 1 2 16704 16707
0 16709 5 1 1 16708
0 16710 7 1 2 24245 16709
0 16711 5 1 1 16710
0 16712 7 1 2 22233 27873
0 16713 7 1 2 28180 26928
0 16714 7 1 2 16712 16713
0 16715 5 1 1 16714
0 16716 7 1 2 16711 16715
0 16717 5 1 1 16716
0 16718 7 1 2 22338 16717
0 16719 5 1 1 16718
0 16720 7 2 2 25761 28918
0 16721 7 2 2 29722 36853
0 16722 7 1 2 1771 15166
0 16723 5 1 1 16722
0 16724 7 1 2 36855 16723
0 16725 5 1 1 16724
0 16726 7 1 2 16719 16725
0 16727 5 1 1 16726
0 16728 7 1 2 23024 16727
0 16729 5 1 1 16728
0 16730 7 1 2 25616 11738
0 16731 7 1 2 32445 16730
0 16732 5 1 1 16731
0 16733 7 1 2 28700 16732
0 16734 5 1 1 16733
0 16735 7 1 2 36179 33163
0 16736 7 1 2 16734 16735
0 16737 5 1 1 16736
0 16738 7 1 2 16729 16737
0 16739 5 1 1 16738
0 16740 7 1 2 22941 16739
0 16741 5 1 1 16740
0 16742 7 2 2 30507 31942
0 16743 7 2 2 28919 36191
0 16744 7 1 2 36857 36859
0 16745 5 1 1 16744
0 16746 7 1 2 16741 16745
0 16747 5 1 1 16746
0 16748 7 1 2 22414 16747
0 16749 5 1 1 16748
0 16750 7 2 2 28356 31968
0 16751 7 1 2 36861 36860
0 16752 5 1 1 16751
0 16753 7 1 2 16749 16752
0 16754 5 1 1 16753
0 16755 7 1 2 31472 16754
0 16756 5 1 1 16755
0 16757 7 1 2 30553 36850
0 16758 5 1 1 16757
0 16759 7 2 2 23025 32392
0 16760 7 1 2 36863 36852
0 16761 5 1 1 16760
0 16762 7 1 2 16758 16761
0 16763 5 1 1 16762
0 16764 7 1 2 24246 16763
0 16765 5 1 1 16764
0 16766 7 1 2 33199 32788
0 16767 7 1 2 36864 16766
0 16768 5 1 1 16767
0 16769 7 1 2 16765 16768
0 16770 5 1 1 16769
0 16771 7 1 2 22339 16770
0 16772 5 1 1 16771
0 16773 7 1 2 23136 36813
0 16774 5 1 1 16773
0 16775 7 1 2 14335 16774
0 16776 5 1 1 16775
0 16777 7 1 2 16776 36856
0 16778 5 1 1 16777
0 16779 7 1 2 16772 16778
0 16780 5 1 1 16779
0 16781 7 1 2 23865 16780
0 16782 5 1 1 16781
0 16783 7 1 2 28725 36833
0 16784 5 1 1 16783
0 16785 7 1 2 30391 34057
0 16786 7 1 2 32410 16785
0 16787 5 1 1 16786
0 16788 7 1 2 16784 16787
0 16789 5 1 1 16788
0 16790 7 1 2 36854 16789
0 16791 5 1 1 16790
0 16792 7 1 2 16782 16791
0 16793 5 1 1 16792
0 16794 7 1 2 22942 16793
0 16795 5 1 1 16794
0 16796 7 1 2 27032 26835
0 16797 7 2 2 36835 16796
0 16798 7 1 2 36858 36865
0 16799 5 1 1 16798
0 16800 7 1 2 16795 16799
0 16801 5 1 1 16800
0 16802 7 1 2 22415 16801
0 16803 5 1 1 16802
0 16804 7 1 2 36866 36862
0 16805 5 1 1 16804
0 16806 7 1 2 16803 16805
0 16807 5 1 1 16806
0 16808 7 1 2 29606 16807
0 16809 5 1 1 16808
0 16810 7 1 2 36146 33792
0 16811 7 1 2 35068 16810
0 16812 5 1 1 16811
0 16813 7 1 2 16809 16812
0 16814 7 1 2 16756 16813
0 16815 5 1 1 16814
0 16816 7 1 2 25720 16815
0 16817 5 1 1 16816
0 16818 7 2 2 25762 26578
0 16819 5 1 1 36867
0 16820 7 5 2 22274 35578
0 16821 7 1 2 27920 36869
0 16822 5 1 1 16821
0 16823 7 2 2 25617 33426
0 16824 7 1 2 27384 36874
0 16825 5 1 1 16824
0 16826 7 1 2 16822 16825
0 16827 5 1 1 16826
0 16828 7 1 2 36767 16827
0 16829 5 1 1 16828
0 16830 7 2 2 26159 26428
0 16831 5 1 1 36876
0 16832 7 1 2 33603 36877
0 16833 5 1 1 16832
0 16834 7 3 2 25618 34747
0 16835 7 1 2 36878 32227
0 16836 5 1 1 16835
0 16837 7 1 2 16833 16836
0 16838 5 1 1 16837
0 16839 7 1 2 28841 16838
0 16840 5 1 1 16839
0 16841 7 2 2 25619 32228
0 16842 7 1 2 34749 36881
0 16843 5 1 1 16842
0 16844 7 2 2 28261 33504
0 16845 7 3 2 24484 24765
0 16846 7 1 2 28650 36885
0 16847 7 1 2 32655 16846
0 16848 7 1 2 36883 16847
0 16849 5 1 1 16848
0 16850 7 1 2 16843 16849
0 16851 7 1 2 16840 16850
0 16852 5 2 1 16851
0 16853 7 1 2 29465 36888
0 16854 5 1 1 16853
0 16855 7 1 2 28431 27566
0 16856 5 1 1 16855
0 16857 7 1 2 163 16856
0 16858 5 1 1 16857
0 16859 7 1 2 23137 16858
0 16860 5 1 1 16859
0 16861 7 1 2 23866 26244
0 16862 5 1 1 16861
0 16863 7 1 2 16860 16862
0 16864 5 2 1 16863
0 16865 7 1 2 33530 36890
0 16866 5 1 1 16865
0 16867 7 1 2 27385 28745
0 16868 7 1 2 33542 16867
0 16869 5 1 1 16868
0 16870 7 1 2 16866 16869
0 16871 5 1 1 16870
0 16872 7 1 2 25517 16871
0 16873 5 1 1 16872
0 16874 7 1 2 16854 16873
0 16875 7 1 2 16829 16874
0 16876 5 1 1 16875
0 16877 7 1 2 31473 16876
0 16878 5 1 1 16877
0 16879 7 1 2 23867 36879
0 16880 5 1 1 16879
0 16881 7 1 2 36870 35294
0 16882 5 1 1 16881
0 16883 7 1 2 16880 16882
0 16884 5 1 1 16883
0 16885 7 1 2 28842 16884
0 16886 5 1 1 16885
0 16887 7 1 2 34371 33266
0 16888 5 1 1 16887
0 16889 7 1 2 16888 33613
0 16890 7 1 2 16886 16889
0 16891 5 1 1 16890
0 16892 7 1 2 24121 16891
0 16893 5 1 1 16892
0 16894 7 1 2 35047 16893
0 16895 5 1 1 16894
0 16896 7 1 2 16895 33261
0 16897 5 1 1 16896
0 16898 7 1 2 24122 36880
0 16899 5 1 1 16898
0 16900 7 1 2 23868 36871
0 16901 7 1 2 36828 16900
0 16902 5 1 1 16901
0 16903 7 1 2 16899 16902
0 16904 5 1 1 16903
0 16905 7 1 2 28843 16904
0 16906 5 1 1 16905
0 16907 7 1 2 34372 33275
0 16908 5 1 1 16907
0 16909 7 1 2 23869 34354
0 16910 5 1 1 16909
0 16911 7 1 2 34425 16910
0 16912 5 1 1 16911
0 16913 7 1 2 32771 16912
0 16914 5 1 1 16913
0 16915 7 1 2 16908 16914
0 16916 7 1 2 16906 16915
0 16917 5 1 1 16916
0 16918 7 1 2 27316 16917
0 16919 5 1 1 16918
0 16920 7 1 2 23138 36889
0 16921 5 1 1 16920
0 16922 7 1 2 16919 16921
0 16923 5 1 1 16922
0 16924 7 1 2 29607 16923
0 16925 5 1 1 16924
0 16926 7 1 2 16897 16925
0 16927 7 1 2 16878 16926
0 16928 5 1 1 16927
0 16929 7 1 2 36868 16928
0 16930 5 1 1 16929
0 16931 7 3 2 25422 25721
0 16932 7 1 2 24123 36892
0 16933 5 1 1 16932
0 16934 7 1 2 30892 33824
0 16935 5 1 1 16934
0 16936 7 1 2 16933 16935
0 16937 5 1 1 16936
0 16938 7 1 2 23568 16937
0 16939 5 1 1 16938
0 16940 7 1 2 24124 36529
0 16941 5 1 1 16940
0 16942 7 1 2 16939 16941
0 16943 5 1 1 16942
0 16944 7 1 2 25991 16943
0 16945 5 1 1 16944
0 16946 7 3 2 23569 31972
0 16947 7 1 2 36895 34984
0 16948 5 1 1 16947
0 16949 7 1 2 16945 16948
0 16950 5 1 1 16949
0 16951 7 1 2 25620 16950
0 16952 5 1 1 16951
0 16953 7 1 2 33605 35347
0 16954 7 1 2 28335 16953
0 16955 5 1 1 16954
0 16956 7 1 2 16952 16955
0 16957 5 1 1 16956
0 16958 7 1 2 29119 16957
0 16959 5 1 1 16958
0 16960 7 1 2 23991 36893
0 16961 5 1 1 16960
0 16962 7 1 2 23026 33825
0 16963 5 1 1 16962
0 16964 7 1 2 16961 16963
0 16965 5 1 1 16964
0 16966 7 1 2 23570 16965
0 16967 5 1 1 16966
0 16968 7 1 2 34355 34018
0 16969 5 1 1 16968
0 16970 7 1 2 16967 16969
0 16971 5 1 1 16970
0 16972 7 1 2 25992 16971
0 16973 5 1 1 16972
0 16974 7 2 2 36896 34463
0 16975 5 1 1 36898
0 16976 7 1 2 23027 36899
0 16977 5 1 1 16976
0 16978 7 1 2 16973 16977
0 16979 5 1 1 16978
0 16980 7 1 2 25621 16979
0 16981 5 1 1 16980
0 16982 7 1 2 35291 35343
0 16983 5 1 1 16982
0 16984 7 1 2 16981 16983
0 16985 5 1 1 16984
0 16986 7 1 2 33053 16985
0 16987 5 1 1 16986
0 16988 7 1 2 16959 16987
0 16989 5 1 1 16988
0 16990 7 1 2 27533 16989
0 16991 5 1 1 16990
0 16992 7 2 2 26429 33551
0 16993 5 2 1 36900
0 16994 7 1 2 30527 36891
0 16995 5 1 1 16994
0 16996 7 1 2 36902 16995
0 16997 5 1 1 16996
0 16998 7 1 2 31474 16997
0 16999 5 1 1 16998
0 17000 7 1 2 9708 9475
0 17001 5 1 1 17000
0 17002 7 1 2 30528 17001
0 17003 5 1 1 17002
0 17004 7 1 2 17003 36903
0 17005 5 1 1 17004
0 17006 7 1 2 27317 17005
0 17007 5 1 1 17006
0 17008 7 1 2 25950 36882
0 17009 5 1 1 17008
0 17010 7 1 2 16831 17009
0 17011 5 2 1 17010
0 17012 7 1 2 36195 36904
0 17013 5 1 1 17012
0 17014 7 1 2 17007 17013
0 17015 5 1 1 17014
0 17016 7 1 2 29608 17015
0 17017 5 1 1 17016
0 17018 7 1 2 29466 36905
0 17019 5 1 1 17018
0 17020 7 1 2 24125 33262
0 17021 7 1 2 35052 17020
0 17022 5 1 1 17021
0 17023 7 1 2 17019 17022
0 17024 5 1 1 17023
0 17025 7 1 2 30529 17024
0 17026 5 1 1 17025
0 17027 7 1 2 23870 33263
0 17028 7 1 2 36901 17027
0 17029 5 1 1 17028
0 17030 7 1 2 17026 17029
0 17031 7 1 2 17017 17030
0 17032 7 1 2 16999 17031
0 17033 5 1 1 17032
0 17034 7 1 2 35504 17033
0 17035 5 1 1 17034
0 17036 7 1 2 22085 28893
0 17037 5 1 1 17036
0 17038 7 1 2 31263 34356
0 17039 5 1 1 17038
0 17040 7 1 2 1087 6895
0 17041 5 1 1 17040
0 17042 7 1 2 23571 6899
0 17043 7 1 2 7584 17042
0 17044 7 1 2 17041 17043
0 17045 5 1 1 17044
0 17046 7 1 2 17039 17045
0 17047 5 1 1 17046
0 17048 7 1 2 25993 17047
0 17049 5 1 1 17048
0 17050 7 1 2 16975 17049
0 17051 5 1 1 17050
0 17052 7 1 2 25622 17051
0 17053 5 1 1 17052
0 17054 7 1 2 23468 33611
0 17055 5 1 1 17054
0 17056 7 1 2 17053 17055
0 17057 5 1 1 17056
0 17058 7 1 2 17037 17057
0 17059 5 1 1 17058
0 17060 7 1 2 33866 36844
0 17061 5 1 1 17060
0 17062 7 1 2 17059 17061
0 17063 5 1 1 17062
0 17064 7 1 2 29609 17063
0 17065 5 1 1 17064
0 17066 7 2 2 25994 33867
0 17067 7 1 2 36082 36906
0 17068 5 1 1 17067
0 17069 7 1 2 32365 36907
0 17070 5 1 1 17069
0 17071 7 1 2 23139 32483
0 17072 7 1 2 33427 17071
0 17073 5 1 1 17072
0 17074 7 1 2 17070 17073
0 17075 5 1 1 17074
0 17076 7 1 2 25623 17075
0 17077 5 1 1 17076
0 17078 7 1 2 28313 29180
0 17079 7 1 2 35292 17078
0 17080 5 1 1 17079
0 17081 7 1 2 17077 17080
0 17082 5 1 1 17081
0 17083 7 1 2 31475 17082
0 17084 5 1 1 17083
0 17085 7 1 2 17068 17084
0 17086 7 1 2 17065 17085
0 17087 7 1 2 17035 17086
0 17088 7 1 2 16991 17087
0 17089 5 1 1 17088
0 17090 7 1 2 33206 17089
0 17091 5 1 1 17090
0 17092 7 1 2 16930 17091
0 17093 7 1 2 16817 17092
0 17094 5 1 1 17093
0 17095 7 1 2 26668 17094
0 17096 5 1 1 17095
0 17097 7 1 2 25281 17096
0 17098 7 1 2 16701 17097
0 17099 5 1 1 17098
0 17100 7 1 2 26470 31500
0 17101 5 1 1 17100
0 17102 7 1 2 22488 33086
0 17103 5 1 1 17102
0 17104 7 1 2 24873 32999
0 17105 5 1 1 17104
0 17106 7 1 2 17103 17105
0 17107 5 1 1 17106
0 17108 7 1 2 21837 17107
0 17109 5 1 1 17108
0 17110 7 4 2 22086 24874
0 17111 7 1 2 36908 35033
0 17112 5 1 1 17111
0 17113 7 1 2 17109 17112
0 17114 5 1 1 17113
0 17115 7 1 2 24973 17114
0 17116 5 1 1 17115
0 17117 7 1 2 17101 17116
0 17118 5 1 1 17117
0 17119 7 1 2 22416 17118
0 17120 5 1 1 17119
0 17121 7 2 2 25624 32234
0 17122 7 2 2 22943 32598
0 17123 7 1 2 36912 36914
0 17124 5 1 1 17123
0 17125 7 1 2 17120 17124
0 17126 5 1 1 17125
0 17127 7 2 2 25518 17126
0 17128 7 1 2 36724 36916
0 17129 5 1 1 17128
0 17130 7 5 2 25099 23572
0 17131 7 4 2 22087 24291
0 17132 7 2 2 32915 36923
0 17133 7 1 2 36918 36927
0 17134 7 1 2 35999 17133
0 17135 5 1 1 17134
0 17136 7 1 2 17129 17135
0 17137 5 1 1 17136
0 17138 7 1 2 28844 17137
0 17139 5 1 1 17138
0 17140 7 1 2 35069 36928
0 17141 5 1 1 17140
0 17142 7 2 2 29382 33405
0 17143 7 1 2 35005 32790
0 17144 7 1 2 36929 17143
0 17145 5 1 1 17144
0 17146 7 1 2 17141 17145
0 17147 5 1 1 17146
0 17148 7 1 2 27187 17147
0 17149 5 1 1 17148
0 17150 7 2 2 28651 35931
0 17151 7 1 2 27918 32189
0 17152 7 1 2 34794 17151
0 17153 7 1 2 36931 17152
0 17154 5 1 1 17153
0 17155 7 1 2 17149 17154
0 17156 5 1 1 17155
0 17157 7 1 2 24974 17156
0 17158 5 1 1 17157
0 17159 7 1 2 28130 36549
0 17160 5 1 1 17159
0 17161 7 1 2 36884 36932
0 17162 5 1 1 17161
0 17163 7 1 2 17160 17162
0 17164 5 1 1 17163
0 17165 7 1 2 31501 17164
0 17166 5 1 1 17165
0 17167 7 1 2 17158 17166
0 17168 7 1 2 17139 17167
0 17169 5 1 1 17168
0 17170 7 1 2 29517 17169
0 17171 5 1 1 17170
0 17172 7 1 2 26432 10734
0 17173 5 3 1 17172
0 17174 7 1 2 23384 31936
0 17175 7 2 2 33505 17174
0 17176 5 1 1 36936
0 17177 7 1 2 28845 36725
0 17178 5 1 1 17177
0 17179 7 1 2 17176 17178
0 17180 5 3 1 17179
0 17181 7 1 2 36933 36938
0 17182 5 1 1 17181
0 17183 7 2 2 22944 23385
0 17184 7 2 2 27067 36941
0 17185 7 1 2 35043 36943
0 17186 5 1 1 17185
0 17187 7 1 2 17182 17186
0 17188 5 1 1 17187
0 17189 7 1 2 26178 17188
0 17190 5 1 1 17189
0 17191 7 1 2 21838 26415
0 17192 5 1 1 17191
0 17193 7 1 2 27289 26640
0 17194 5 1 1 17193
0 17195 7 1 2 17192 17194
0 17196 5 1 1 17195
0 17197 7 1 2 22417 17196
0 17198 5 1 1 17197
0 17199 7 2 2 22945 26478
0 17200 7 1 2 32135 36945
0 17201 5 1 1 17200
0 17202 7 1 2 17198 17201
0 17203 5 3 1 17202
0 17204 7 1 2 36947 36939
0 17205 5 1 1 17204
0 17206 7 2 2 26500 34180
0 17207 7 1 2 24975 35034
0 17208 7 1 2 35932 17207
0 17209 7 1 2 36950 17208
0 17210 5 1 1 17209
0 17211 7 1 2 17205 17210
0 17212 7 1 2 17190 17211
0 17213 5 1 1 17212
0 17214 7 1 2 25519 17213
0 17215 5 1 1 17214
0 17216 7 2 2 28262 36930
0 17217 7 1 2 35937 36952
0 17218 5 1 1 17217
0 17219 7 1 2 17215 17218
0 17220 5 1 1 17219
0 17221 7 1 2 35064 17220
0 17222 5 1 1 17221
0 17223 7 1 2 25951 36940
0 17224 5 1 1 17223
0 17225 7 1 2 34201 36944
0 17226 5 1 1 17225
0 17227 7 1 2 17224 17226
0 17228 5 1 1 17227
0 17229 7 1 2 35029 17228
0 17230 5 1 1 17229
0 17231 7 1 2 17222 17230
0 17232 7 1 2 17171 17231
0 17233 5 1 1 17232
0 17234 7 1 2 36404 17233
0 17235 5 1 1 17234
0 17236 7 1 2 36609 36917
0 17237 5 1 1 17236
0 17238 7 1 2 28678 30747
0 17239 7 1 2 36330 34479
0 17240 7 1 2 35057 17239
0 17241 7 1 2 17238 17240
0 17242 5 1 1 17241
0 17243 7 1 2 17237 17242
0 17244 5 1 1 17243
0 17245 7 1 2 28846 17244
0 17246 5 1 1 17245
0 17247 7 1 2 25100 29257
0 17248 7 1 2 34908 17247
0 17249 7 1 2 29273 17248
0 17250 5 1 1 17249
0 17251 7 1 2 36563 36924
0 17252 7 1 2 35070 17251
0 17253 5 1 1 17252
0 17254 7 1 2 17250 17253
0 17255 5 1 1 17254
0 17256 7 1 2 27188 17255
0 17257 5 1 1 17256
0 17258 7 1 2 22946 35854
0 17259 7 1 2 29687 17258
0 17260 7 2 2 28759 30666
0 17261 7 2 2 24292 28950
0 17262 7 1 2 36954 36956
0 17263 7 1 2 17259 17262
0 17264 5 1 1 17263
0 17265 7 1 2 17257 17264
0 17266 5 1 1 17265
0 17267 7 1 2 24976 17266
0 17268 5 1 1 17267
0 17269 7 1 2 23573 36610
0 17270 5 1 1 17269
0 17271 7 1 2 15609 17270
0 17272 5 1 1 17271
0 17273 7 1 2 28131 17272
0 17274 5 1 1 17273
0 17275 7 3 2 22876 36564
0 17276 7 1 2 35295 36957
0 17277 7 1 2 36958 17276
0 17278 5 1 1 17277
0 17279 7 1 2 17274 17278
0 17280 5 1 1 17279
0 17281 7 1 2 31502 17280
0 17282 5 1 1 17281
0 17283 7 1 2 17268 17282
0 17284 7 1 2 17246 17283
0 17285 5 1 1 17284
0 17286 7 1 2 29518 17285
0 17287 5 1 1 17286
0 17288 7 1 2 28847 36611
0 17289 5 1 1 17288
0 17290 7 1 2 25867 36683
0 17291 5 1 1 17290
0 17292 7 1 2 17289 17291
0 17293 5 4 1 17292
0 17294 7 1 2 25952 36961
0 17295 5 1 1 17294
0 17296 7 3 2 22418 36565
0 17297 7 1 2 36951 36965
0 17298 5 1 1 17297
0 17299 7 1 2 17295 17298
0 17300 5 2 1 17299
0 17301 7 1 2 36968 35030
0 17302 5 1 1 17301
0 17303 7 1 2 36962 36934
0 17304 5 1 1 17303
0 17305 7 3 2 31117 35604
0 17306 7 1 2 25625 26501
0 17307 7 1 2 31538 17306
0 17308 7 1 2 36970 17307
0 17309 5 1 1 17308
0 17310 7 1 2 17304 17309
0 17311 5 1 1 17310
0 17312 7 1 2 26179 17311
0 17313 5 1 1 17312
0 17314 7 1 2 36963 36948
0 17315 5 1 1 17314
0 17316 7 1 2 30650 34202
0 17317 7 1 2 36566 36946
0 17318 7 1 2 17316 17317
0 17319 5 1 1 17318
0 17320 7 1 2 17315 17319
0 17321 7 1 2 17313 17320
0 17322 5 1 1 17321
0 17323 7 1 2 25520 17322
0 17324 5 1 1 17323
0 17325 7 1 2 28953 35558
0 17326 7 1 2 36780 17325
0 17327 5 1 1 17326
0 17328 7 1 2 17324 17327
0 17329 5 1 1 17328
0 17330 7 1 2 35065 17329
0 17331 5 1 1 17330
0 17332 7 1 2 17302 17331
0 17333 7 1 2 17287 17332
0 17334 5 1 1 17333
0 17335 7 1 2 32983 17334
0 17336 5 1 1 17335
0 17337 7 1 2 22419 29900
0 17338 7 1 2 36517 17337
0 17339 7 1 2 35773 17338
0 17340 7 1 2 36953 17339
0 17341 5 1 1 17340
0 17342 7 1 2 17336 17341
0 17343 7 1 2 17235 17342
0 17344 5 1 1 17343
0 17345 7 1 2 34589 17344
0 17346 5 1 1 17345
0 17347 7 1 2 27885 33849
0 17348 5 1 1 17347
0 17349 7 1 2 8258 17348
0 17350 5 1 1 17349
0 17351 7 1 2 22489 17350
0 17352 5 1 1 17351
0 17353 7 1 2 22818 33268
0 17354 5 1 1 17353
0 17355 7 1 2 17352 17354
0 17356 5 1 1 17355
0 17357 7 1 2 21839 17356
0 17358 5 1 1 17357
0 17359 7 1 2 33618 35491
0 17360 7 1 2 35973 17359
0 17361 5 1 1 17360
0 17362 7 1 2 17358 17361
0 17363 5 1 1 17362
0 17364 7 1 2 26385 17363
0 17365 5 1 1 17364
0 17366 7 1 2 32484 35977
0 17367 5 1 1 17366
0 17368 7 1 2 24823 33861
0 17369 7 1 2 32235 17368
0 17370 5 1 1 17369
0 17371 7 1 2 17367 17370
0 17372 5 1 1 17371
0 17373 7 1 2 25626 17372
0 17374 5 1 1 17373
0 17375 7 1 2 35330 36955
0 17376 5 1 1 17375
0 17377 7 1 2 24347 17376
0 17378 7 1 2 17374 17377
0 17379 5 1 1 17378
0 17380 7 1 2 28696 34009
0 17381 5 1 1 17380
0 17382 7 1 2 30865 35526
0 17383 5 1 1 17382
0 17384 7 1 2 17381 17383
0 17385 5 1 1 17384
0 17386 7 1 2 25101 17385
0 17387 5 1 1 17386
0 17388 7 1 2 22340 17387
0 17389 5 1 1 17388
0 17390 7 1 2 22088 17389
0 17391 7 1 2 17379 17390
0 17392 5 1 1 17391
0 17393 7 1 2 17365 17392
0 17394 5 1 1 17393
0 17395 7 1 2 22947 17394
0 17396 5 1 1 17395
0 17397 7 2 2 35337 36913
0 17398 7 1 2 36909 36973
0 17399 5 1 1 17398
0 17400 7 1 2 17396 17399
0 17401 5 1 1 17400
0 17402 7 1 2 22420 17401
0 17403 5 1 1 17402
0 17404 7 1 2 36974 36915
0 17405 5 1 1 17404
0 17406 7 1 2 17403 17405
0 17407 5 1 1 17406
0 17408 7 1 2 29519 17407
0 17409 5 1 1 17408
0 17410 7 1 2 31358 35341
0 17411 5 1 1 17410
0 17412 7 1 2 21840 35563
0 17413 5 1 1 17412
0 17414 7 3 2 36378 33834
0 17415 7 1 2 26089 36975
0 17416 5 1 1 17415
0 17417 7 1 2 17413 17416
0 17418 5 1 1 17417
0 17419 7 1 2 22948 17418
0 17420 5 1 1 17419
0 17421 7 1 2 32082 36976
0 17422 5 1 1 17421
0 17423 7 1 2 17420 17422
0 17424 5 1 1 17423
0 17425 7 1 2 22421 17424
0 17426 5 1 1 17425
0 17427 7 1 2 36823 36977
0 17428 5 1 1 17427
0 17429 7 1 2 31973 34048
0 17430 5 1 1 17429
0 17431 7 1 2 21841 35331
0 17432 7 1 2 32093 17431
0 17433 5 1 1 17432
0 17434 7 1 2 17430 17433
0 17435 5 1 1 17434
0 17436 7 1 2 22422 17435
0 17437 5 1 1 17436
0 17438 7 1 2 21842 28340
0 17439 7 1 2 34500 17438
0 17440 5 1 1 17439
0 17441 7 1 2 17437 17440
0 17442 5 1 1 17441
0 17443 7 1 2 26180 17442
0 17444 5 1 1 17443
0 17445 7 1 2 17428 17444
0 17446 7 1 2 17426 17445
0 17447 5 1 1 17446
0 17448 7 1 2 25627 17447
0 17449 5 1 1 17448
0 17450 7 1 2 23574 35581
0 17451 7 1 2 17449 17450
0 17452 5 1 1 17451
0 17453 7 1 2 35588 36935
0 17454 5 1 1 17453
0 17455 7 1 2 27033 34490
0 17456 7 1 2 35287 17455
0 17457 5 1 1 17456
0 17458 7 1 2 17454 17457
0 17459 5 1 1 17458
0 17460 7 1 2 26181 17459
0 17461 5 1 1 17460
0 17462 7 1 2 35589 36949
0 17463 5 1 1 17462
0 17464 7 1 2 27290 34010
0 17465 7 1 2 35060 17464
0 17466 5 1 1 17465
0 17467 7 1 2 25521 17466
0 17468 7 1 2 17463 17467
0 17469 7 1 2 17461 17468
0 17470 5 1 1 17469
0 17471 7 1 2 35066 17470
0 17472 7 1 2 17452 17471
0 17473 5 1 1 17472
0 17474 7 1 2 17411 17473
0 17475 7 1 2 17409 17474
0 17476 5 2 1 17475
0 17477 7 1 2 36584 36978
0 17478 5 1 1 17477
0 17479 7 1 2 26239 26439
0 17480 7 1 2 28897 34649
0 17481 7 1 2 17479 17480
0 17482 7 1 2 36097 17481
0 17483 7 1 2 35307 17482
0 17484 5 1 1 17483
0 17485 7 1 2 27222 31198
0 17486 5 1 1 17485
0 17487 7 1 2 35098 17486
0 17488 5 1 1 17487
0 17489 7 1 2 34110 17488
0 17490 5 1 1 17489
0 17491 7 1 2 31199 33975
0 17492 7 1 2 3008 17491
0 17493 5 1 1 17492
0 17494 7 1 2 17490 17493
0 17495 5 1 1 17494
0 17496 7 1 2 25102 17495
0 17497 5 1 1 17496
0 17498 7 1 2 25423 34796
0 17499 7 1 2 31665 17498
0 17500 5 1 1 17499
0 17501 7 1 2 17497 17500
0 17502 5 2 1 17501
0 17503 7 1 2 36612 32094
0 17504 5 1 1 17503
0 17505 7 1 2 36684 33395
0 17506 5 1 1 17505
0 17507 7 1 2 17504 17506
0 17508 5 1 1 17507
0 17509 7 1 2 22423 17508
0 17510 5 1 1 17509
0 17511 7 1 2 36613 36824
0 17512 5 1 1 17511
0 17513 7 1 2 17510 17512
0 17514 5 1 1 17513
0 17515 7 1 2 25628 17514
0 17516 7 1 2 36980 17515
0 17517 5 1 1 17516
0 17518 7 1 2 17484 17517
0 17519 5 1 1 17518
0 17520 7 1 2 23575 17519
0 17521 5 1 1 17520
0 17522 7 1 2 17478 17521
0 17523 5 1 1 17522
0 17524 7 1 2 32984 17523
0 17525 5 1 1 17524
0 17526 7 1 2 36405 36979
0 17527 5 1 1 17526
0 17528 7 2 2 26805 36503
0 17529 7 1 2 28452 31299
0 17530 7 1 2 31098 17529
0 17531 7 1 2 36982 17530
0 17532 7 1 2 28111 17531
0 17533 5 1 1 17532
0 17534 7 1 2 17527 17533
0 17535 5 1 1 17534
0 17536 7 1 2 36602 17535
0 17537 5 1 1 17536
0 17538 7 1 2 32095 36726
0 17539 5 1 1 17538
0 17540 7 1 2 22949 36722
0 17541 5 1 1 17540
0 17542 7 1 2 17539 17541
0 17543 5 1 1 17542
0 17544 7 1 2 22424 17543
0 17545 5 1 1 17544
0 17546 7 1 2 22950 36370
0 17547 7 1 2 35803 17546
0 17548 5 1 1 17547
0 17549 7 1 2 17545 17548
0 17550 5 1 1 17549
0 17551 7 1 2 28679 36406
0 17552 7 1 2 36981 17551
0 17553 7 1 2 17550 17552
0 17554 5 1 1 17553
0 17555 7 1 2 23324 17554
0 17556 7 1 2 17537 17555
0 17557 7 1 2 17525 17556
0 17558 7 1 2 17346 17557
0 17559 5 1 1 17558
0 17560 7 1 2 17099 17559
0 17561 5 1 1 17560
0 17562 7 1 2 23767 17561
0 17563 5 1 1 17562
0 17564 7 1 2 30146 17563
0 17565 7 1 2 16326 17564
0 17566 5 1 1 17565
0 17567 7 1 2 31232 35950
0 17568 5 1 1 17567
0 17569 7 3 2 25194 30410
0 17570 7 1 2 28539 36984
0 17571 5 1 1 17570
0 17572 7 1 2 17568 17571
0 17573 5 1 1 17572
0 17574 7 1 2 26806 17573
0 17575 5 1 1 17574
0 17576 7 1 2 23469 35213
0 17577 7 2 2 34024 17576
0 17578 7 1 2 36034 36987
0 17579 5 1 1 17578
0 17580 7 1 2 17575 17579
0 17581 5 1 1 17580
0 17582 7 1 2 17581 35140
0 17583 5 1 1 17582
0 17584 7 2 2 25195 26600
0 17585 7 1 2 30784 36989
0 17586 5 2 1 17585
0 17587 7 1 2 36095 36991
0 17588 5 2 1 17587
0 17589 7 2 2 22234 36993
0 17590 5 1 1 36995
0 17591 7 1 2 4178 36023
0 17592 5 3 1 17591
0 17593 7 1 2 34856 36997
0 17594 5 1 1 17593
0 17595 7 1 2 17590 17594
0 17596 5 1 1 17595
0 17597 7 1 2 36919 35831
0 17598 7 1 2 17596 17597
0 17599 5 1 1 17598
0 17600 7 1 2 17583 17599
0 17601 5 2 1 17600
0 17602 7 1 2 33728 37000
0 17603 5 1 1 17602
0 17604 7 3 2 25424 28540
0 17605 7 1 2 31034 36043
0 17606 5 1 1 17605
0 17607 7 1 2 26312 17606
0 17608 5 1 1 17607
0 17609 7 1 2 4245 17608
0 17610 5 1 1 17609
0 17611 7 1 2 23325 17610
0 17612 5 1 1 17611
0 17613 7 1 2 24627 35729
0 17614 5 1 1 17613
0 17615 7 1 2 31106 34700
0 17616 5 1 1 17615
0 17617 7 1 2 17614 17616
0 17618 5 1 1 17617
0 17619 7 1 2 23233 17618
0 17620 5 1 1 17619
0 17621 7 1 2 24628 35954
0 17622 5 1 1 17621
0 17623 7 1 2 17620 17622
0 17624 5 1 1 17623
0 17625 7 1 2 22089 25282
0 17626 7 1 2 17624 17625
0 17627 5 1 1 17626
0 17628 7 1 2 17612 17627
0 17629 5 1 1 17628
0 17630 7 1 2 37002 17629
0 17631 5 1 1 17630
0 17632 7 1 2 36282 31882
0 17633 7 1 2 31844 17632
0 17634 5 1 1 17633
0 17635 7 1 2 17631 17634
0 17636 5 1 1 17635
0 17637 7 1 2 25522 17636
0 17638 5 1 1 17637
0 17639 7 1 2 24629 35725
0 17640 5 1 1 17639
0 17641 7 1 2 22677 32270
0 17642 5 1 1 17641
0 17643 7 1 2 23871 30987
0 17644 7 1 2 17642 17643
0 17645 5 1 1 17644
0 17646 7 1 2 17640 17645
0 17647 5 1 1 17646
0 17648 7 1 2 28993 17647
0 17649 5 1 1 17648
0 17650 7 1 2 28089 35653
0 17651 5 1 1 17650
0 17652 7 1 2 17649 17651
0 17653 5 1 1 17652
0 17654 7 1 2 25283 17653
0 17655 5 1 1 17654
0 17656 7 1 2 30225 35714
0 17657 5 1 1 17656
0 17658 7 1 2 17655 17657
0 17659 5 1 1 17658
0 17660 7 3 2 25523 37003
0 17661 7 1 2 35750 37005
0 17662 7 1 2 17659 17661
0 17663 5 1 1 17662
0 17664 7 1 2 17638 17663
0 17665 5 2 1 17664
0 17666 7 1 2 26090 37008
0 17667 5 1 1 17666
0 17668 7 1 2 31536 12889
0 17669 5 1 1 17668
0 17670 7 1 2 28541 30785
0 17671 7 1 2 17669 17670
0 17672 5 1 1 17671
0 17673 7 1 2 24543 33231
0 17674 7 1 2 34317 17673
0 17675 7 1 2 27354 17674
0 17676 5 1 1 17675
0 17677 7 1 2 17672 17676
0 17678 5 1 1 17677
0 17679 7 2 2 30247 17678
0 17680 7 1 2 26091 37010
0 17681 5 1 1 17680
0 17682 7 3 2 23326 32485
0 17683 7 2 2 30059 37012
0 17684 7 1 2 25763 32418
0 17685 7 1 2 37015 17684
0 17686 5 1 1 17685
0 17687 7 1 2 17681 17686
0 17688 5 1 1 17687
0 17689 7 1 2 23992 17688
0 17690 5 1 1 17689
0 17691 7 1 2 27155 30681
0 17692 5 1 1 17691
0 17693 7 1 2 30795 31418
0 17694 7 1 2 5061 17693
0 17695 5 1 1 17694
0 17696 7 1 2 17692 17695
0 17697 5 1 1 17696
0 17698 7 1 2 22570 17697
0 17699 5 1 1 17698
0 17700 7 1 2 30682 35948
0 17701 5 1 1 17700
0 17702 7 1 2 29393 30156
0 17703 5 1 1 17702
0 17704 7 1 2 1526 17703
0 17705 5 1 1 17704
0 17706 7 1 2 27470 17705
0 17707 5 1 1 17706
0 17708 7 1 2 17701 17707
0 17709 7 1 2 17699 17708
0 17710 5 1 1 17709
0 17711 7 2 2 25284 28542
0 17712 7 1 2 30248 37017
0 17713 7 2 2 17710 17712
0 17714 7 1 2 26092 37019
0 17715 5 1 1 17714
0 17716 7 1 2 24720 26882
0 17717 7 1 2 31082 17716
0 17718 7 2 2 30709 33282
0 17719 7 1 2 32419 37021
0 17720 7 1 2 17717 17719
0 17721 5 1 1 17720
0 17722 7 1 2 17715 17721
0 17723 7 1 2 17690 17722
0 17724 5 1 1 17723
0 17725 7 1 2 31328 17724
0 17726 5 1 1 17725
0 17727 7 1 2 17667 17726
0 17728 5 1 1 17727
0 17729 7 1 2 33379 17728
0 17730 5 1 1 17729
0 17731 7 1 2 17603 17730
0 17732 5 1 1 17731
0 17733 7 1 2 23386 17732
0 17734 5 1 1 17733
0 17735 7 1 2 23993 30414
0 17736 5 1 1 17735
0 17737 7 1 2 32793 35832
0 17738 5 1 1 17737
0 17739 7 1 2 17736 17738
0 17740 5 1 1 17739
0 17741 7 1 2 35078 17740
0 17742 5 1 1 17741
0 17743 7 1 2 35658 36016
0 17744 5 1 1 17743
0 17745 7 1 2 24630 29901
0 17746 7 1 2 35795 17745
0 17747 7 1 2 29678 17746
0 17748 5 1 1 17747
0 17749 7 1 2 17744 17748
0 17750 5 1 1 17749
0 17751 7 1 2 28543 17750
0 17752 5 1 1 17751
0 17753 7 1 2 24544 26160
0 17754 7 1 2 28181 33178
0 17755 7 1 2 17753 17754
0 17756 7 1 2 31113 35106
0 17757 7 1 2 17755 17756
0 17758 5 1 1 17757
0 17759 7 1 2 17752 17758
0 17760 7 1 2 17742 17759
0 17761 5 1 1 17760
0 17762 7 1 2 33928 17761
0 17763 5 1 1 17762
0 17764 7 1 2 36998 35122
0 17765 5 1 1 17764
0 17766 7 2 2 23140 26741
0 17767 7 1 2 22778 37023
0 17768 7 1 2 29679 17767
0 17769 5 1 1 17768
0 17770 7 1 2 17765 17769
0 17771 5 1 1 17770
0 17772 7 1 2 24977 17771
0 17773 5 1 1 17772
0 17774 7 1 2 31548 33232
0 17775 7 1 2 29848 17774
0 17776 5 1 1 17775
0 17777 7 1 2 17773 17776
0 17778 5 1 1 17777
0 17779 7 1 2 23470 17778
0 17780 5 1 1 17779
0 17781 7 1 2 23141 36093
0 17782 7 1 2 36169 17781
0 17783 7 1 2 27355 17782
0 17784 5 1 1 17783
0 17785 7 1 2 22235 17784
0 17786 7 1 2 17780 17785
0 17787 5 1 1 17786
0 17788 7 1 2 36994 35123
0 17789 5 1 1 17788
0 17790 7 1 2 28182 37024
0 17791 7 1 2 29680 17790
0 17792 5 1 1 17791
0 17793 7 1 2 17789 17792
0 17794 5 1 1 17793
0 17795 7 1 2 24978 17794
0 17796 5 1 1 17795
0 17797 7 1 2 22779 30500
0 17798 5 1 1 17797
0 17799 7 1 2 36024 17798
0 17800 5 2 1 17799
0 17801 7 1 2 27860 37025
0 17802 5 1 1 17801
0 17803 7 1 2 28090 31792
0 17804 5 1 1 17803
0 17805 7 1 2 17802 17804
0 17806 5 1 1 17805
0 17807 7 1 2 17806 35227
0 17808 5 1 1 17807
0 17809 7 1 2 24247 17808
0 17810 7 1 2 17796 17809
0 17811 5 1 1 17810
0 17812 7 1 2 34420 17811
0 17813 7 1 2 17787 17812
0 17814 5 1 1 17813
0 17815 7 1 2 17763 17814
0 17816 5 1 1 17815
0 17817 7 2 2 25355 17816
0 17818 7 1 2 26093 37027
0 17819 5 1 1 17818
0 17820 7 1 2 17734 17819
0 17821 5 1 1 17820
0 17822 7 1 2 23681 17821
0 17823 5 1 1 17822
0 17824 7 2 2 24766 26270
0 17825 7 1 2 34912 34513
0 17826 7 1 2 37029 17825
0 17827 7 3 2 27068 27991
0 17828 7 1 2 29902 37031
0 17829 7 1 2 30814 17828
0 17830 7 1 2 17826 17829
0 17831 5 1 1 17830
0 17832 7 1 2 17823 17831
0 17833 5 1 1 17832
0 17834 7 1 2 25953 17833
0 17835 5 1 1 17834
0 17836 7 1 2 35805 37001
0 17837 5 1 1 17836
0 17838 7 1 2 27693 37009
0 17839 5 1 1 17838
0 17840 7 1 2 27694 37011
0 17841 5 1 1 17840
0 17842 7 1 2 28274 27979
0 17843 7 1 2 26508 17842
0 17844 7 1 2 37016 17843
0 17845 5 1 1 17844
0 17846 7 1 2 17841 17845
0 17847 5 1 1 17846
0 17848 7 1 2 23994 17847
0 17849 5 1 1 17848
0 17850 7 1 2 27695 37020
0 17851 5 1 1 17850
0 17852 7 1 2 28027 27069
0 17853 7 1 2 28396 17852
0 17854 7 1 2 37022 35667
0 17855 7 1 2 17853 17854
0 17856 5 1 1 17855
0 17857 7 1 2 17851 17856
0 17858 7 1 2 17849 17857
0 17859 5 1 1 17858
0 17860 7 1 2 31329 17859
0 17861 5 1 1 17860
0 17862 7 1 2 17839 17861
0 17863 5 1 1 17862
0 17864 7 1 2 33380 17863
0 17865 5 1 1 17864
0 17866 7 1 2 17837 17865
0 17867 5 1 1 17866
0 17868 7 1 2 23387 17867
0 17869 5 1 1 17868
0 17870 7 1 2 27696 37028
0 17871 5 1 1 17870
0 17872 7 1 2 17869 17871
0 17873 5 1 1 17872
0 17874 7 1 2 23682 17873
0 17875 5 1 1 17874
0 17876 7 1 2 27249 34881
0 17877 5 1 1 17876
0 17878 7 1 2 24631 35735
0 17879 5 1 1 17878
0 17880 7 1 2 22678 35723
0 17881 5 1 1 17880
0 17882 7 1 2 23234 17881
0 17883 7 1 2 17879 17882
0 17884 5 1 1 17883
0 17885 7 1 2 17877 17884
0 17886 5 1 1 17885
0 17887 7 1 2 25285 17886
0 17888 5 1 1 17887
0 17889 7 1 2 22679 35716
0 17890 5 1 1 17889
0 17891 7 1 2 17888 17890
0 17892 5 1 1 17891
0 17893 7 4 2 25524 33995
0 17894 7 1 2 28544 37034
0 17895 7 1 2 17892 17894
0 17896 5 1 1 17895
0 17897 7 1 2 27967 33255
0 17898 7 1 2 31787 17897
0 17899 7 3 2 23872 32486
0 17900 7 2 2 24632 24721
0 17901 7 2 2 24485 37041
0 17902 7 1 2 37038 37043
0 17903 7 1 2 17898 17902
0 17904 5 1 1 17903
0 17905 7 1 2 17896 17904
0 17906 5 1 1 17905
0 17907 7 1 2 35777 17906
0 17908 5 1 1 17907
0 17909 7 1 2 22680 12119
0 17910 5 1 1 17909
0 17911 7 1 2 30858 17910
0 17912 5 1 1 17911
0 17913 7 1 2 23142 17912
0 17914 5 1 1 17913
0 17915 7 1 2 23995 28432
0 17916 7 1 2 33752 17915
0 17917 5 1 1 17916
0 17918 7 1 2 17914 17917
0 17919 5 1 1 17918
0 17920 7 1 2 34063 17919
0 17921 5 1 1 17920
0 17922 7 2 2 29062 34453
0 17923 7 1 2 33586 37045
0 17924 7 1 2 27361 17923
0 17925 5 1 1 17924
0 17926 7 1 2 17921 17925
0 17927 5 1 1 17926
0 17928 7 1 2 23683 17927
0 17929 5 1 1 17928
0 17930 7 1 2 24875 29728
0 17931 7 2 2 32429 17930
0 17932 7 1 2 34154 37046
0 17933 7 1 2 37047 17932
0 17934 5 1 1 17933
0 17935 7 1 2 17929 17934
0 17936 5 1 1 17935
0 17937 7 1 2 37018 17936
0 17938 5 1 1 17937
0 17939 7 2 2 33381 37048
0 17940 5 1 1 37049
0 17941 7 1 2 23684 30999
0 17942 7 1 2 34081 17941
0 17943 5 1 1 17942
0 17944 7 1 2 17940 17943
0 17945 5 1 1 17944
0 17946 7 1 2 31780 34758
0 17947 7 1 2 17945 17946
0 17948 5 1 1 17947
0 17949 7 1 2 17938 17948
0 17950 5 1 1 17949
0 17951 7 1 2 25425 17950
0 17952 5 1 1 17951
0 17953 7 1 2 26420 292
0 17954 5 1 1 17953
0 17955 7 1 2 34421 17954
0 17956 5 1 1 17955
0 17957 7 1 2 26484 33929
0 17958 5 1 1 17957
0 17959 7 1 2 17956 17958
0 17960 5 1 1 17959
0 17961 7 1 2 23873 17960
0 17962 5 1 1 17961
0 17963 7 1 2 27318 33628
0 17964 5 1 1 17963
0 17965 7 1 2 24486 34988
0 17966 5 1 1 17965
0 17967 7 1 2 17964 17966
0 17968 5 1 1 17967
0 17969 7 1 2 26416 17968
0 17970 5 1 1 17969
0 17971 7 1 2 17962 17970
0 17972 5 1 1 17971
0 17973 7 1 2 30964 17972
0 17974 5 1 1 17973
0 17975 7 1 2 30956 36364
0 17976 7 1 2 36366 17975
0 17977 7 1 2 36815 17976
0 17978 5 1 1 17977
0 17979 7 1 2 17974 17978
0 17980 5 1 1 17979
0 17981 7 1 2 36988 17980
0 17982 5 1 1 17981
0 17983 7 1 2 17952 17982
0 17984 5 1 1 17983
0 17985 7 1 2 24545 17984
0 17986 5 1 1 17985
0 17987 7 1 2 17908 17986
0 17988 5 1 1 17987
0 17989 7 1 2 24126 17988
0 17990 5 1 1 17989
0 17991 7 1 2 36291 34082
0 17992 5 1 1 17991
0 17993 7 1 2 25286 34064
0 17994 7 1 2 30991 17993
0 17995 5 1 1 17994
0 17996 7 1 2 17992 17995
0 17997 5 1 1 17996
0 17998 7 1 2 23235 28545
0 17999 7 1 2 17997 17998
0 18000 5 1 1 17999
0 18001 7 1 2 30374 33382
0 18002 7 1 2 35670 34390
0 18003 7 1 2 18001 18002
0 18004 7 1 2 24248 24979
0 18005 7 1 2 25196 18004
0 18006 7 1 2 29435 18005
0 18007 7 1 2 18003 18006
0 18008 5 1 1 18007
0 18009 7 1 2 18000 18008
0 18010 5 1 1 18009
0 18011 7 1 2 25426 18010
0 18012 5 1 1 18011
0 18013 7 1 2 30085 35091
0 18014 7 1 2 35819 18013
0 18015 5 1 1 18014
0 18016 7 1 2 18012 18015
0 18017 5 1 1 18016
0 18018 7 1 2 25103 18017
0 18019 5 1 1 18018
0 18020 7 1 2 30995 35302
0 18021 5 1 1 18020
0 18022 7 1 2 31003 18021
0 18023 5 1 1 18022
0 18024 7 1 2 23236 18023
0 18025 5 1 1 18024
0 18026 7 1 2 31007 18025
0 18027 5 1 1 18026
0 18028 7 1 2 25287 18027
0 18029 5 1 1 18028
0 18030 7 1 2 24980 30194
0 18031 5 1 1 18030
0 18032 7 1 2 18029 18031
0 18033 5 1 1 18032
0 18034 7 1 2 37006 35739
0 18035 7 1 2 18033 18034
0 18036 5 1 1 18035
0 18037 7 1 2 18019 18036
0 18038 5 1 1 18037
0 18039 7 1 2 22090 18038
0 18040 5 1 1 18039
0 18041 7 2 2 27541 33330
0 18042 7 1 2 26699 37051
0 18043 7 1 2 37007 18042
0 18044 7 1 2 31036 18043
0 18045 5 1 1 18044
0 18046 7 1 2 18040 18045
0 18047 5 1 1 18046
0 18048 7 1 2 23685 18047
0 18049 5 1 1 18048
0 18050 7 1 2 23388 18049
0 18051 7 1 2 17990 18050
0 18052 5 1 1 18051
0 18053 7 1 2 35079 34083
0 18054 5 1 1 18053
0 18055 7 1 2 35087 34073
0 18056 5 1 1 18055
0 18057 7 1 2 18054 18056
0 18058 5 1 1 18057
0 18059 7 1 2 27362 18058
0 18060 5 1 1 18059
0 18061 7 2 2 24722 27156
0 18062 7 1 2 26945 34857
0 18063 7 1 2 37053 18062
0 18064 7 1 2 37052 18063
0 18065 5 1 1 18064
0 18066 7 1 2 18060 18065
0 18067 5 1 1 18066
0 18068 7 1 2 26742 18067
0 18069 5 1 1 18068
0 18070 7 1 2 26182 34077
0 18071 5 1 1 18070
0 18072 7 1 2 27335 34084
0 18073 7 1 2 18071 18072
0 18074 5 1 1 18073
0 18075 7 1 2 29729 36886
0 18076 7 1 2 34480 18075
0 18077 5 1 1 18076
0 18078 7 1 2 18074 18077
0 18079 5 1 1 18078
0 18080 7 1 2 26516 37004
0 18081 7 1 2 18079 18080
0 18082 5 1 1 18081
0 18083 7 1 2 18069 18082
0 18084 5 1 1 18083
0 18085 7 1 2 23686 18084
0 18086 5 1 1 18085
0 18087 7 1 2 34858 37026
0 18088 5 1 1 18087
0 18089 7 1 2 22681 36992
0 18090 5 1 1 18089
0 18091 7 1 2 36996 18090
0 18092 5 1 1 18091
0 18093 7 1 2 18088 18092
0 18094 5 1 1 18093
0 18095 7 1 2 37050 18094
0 18096 5 1 1 18095
0 18097 7 1 2 18086 18096
0 18098 5 1 1 18097
0 18099 7 1 2 35141 18098
0 18100 5 1 1 18099
0 18101 7 1 2 22236 36999
0 18102 5 1 1 18101
0 18103 7 1 2 28520 36304
0 18104 5 1 1 18103
0 18105 7 1 2 18102 18104
0 18106 5 1 1 18105
0 18107 7 1 2 23471 34085
0 18108 7 1 2 18106 18107
0 18109 5 1 1 18108
0 18110 7 1 2 33587 34569
0 18111 7 1 2 36198 18110
0 18112 5 1 1 18111
0 18113 7 1 2 18109 18112
0 18114 5 1 1 18113
0 18115 7 1 2 35834 18114
0 18116 5 1 1 18115
0 18117 7 1 2 25356 18116
0 18118 7 1 2 18100 18117
0 18119 5 1 1 18118
0 18120 7 1 2 24409 18119
0 18121 7 1 2 18052 18120
0 18122 5 1 1 18121
0 18123 7 1 2 24633 22780
0 18124 7 1 2 30473 18123
0 18125 5 1 1 18124
0 18126 7 1 2 32985 36985
0 18127 5 1 1 18126
0 18128 7 1 2 18125 18127
0 18129 5 1 1 18128
0 18130 7 1 2 24293 33976
0 18131 7 1 2 18129 18130
0 18132 5 1 1 18131
0 18133 7 1 2 22819 27968
0 18134 7 1 2 34600 18133
0 18135 7 1 2 27386 33164
0 18136 7 1 2 18134 18135
0 18137 5 1 1 18136
0 18138 7 1 2 18132 18137
0 18139 5 1 1 18138
0 18140 7 1 2 24249 18139
0 18141 5 1 1 18140
0 18142 7 1 2 34301 36986
0 18143 5 1 1 18142
0 18144 7 2 2 25427 36210
0 18145 5 1 1 37055
0 18146 7 1 2 27356 37056
0 18147 5 1 1 18146
0 18148 7 1 2 18143 18147
0 18149 5 1 1 18148
0 18150 7 1 2 34897 18149
0 18151 5 1 1 18150
0 18152 7 1 2 18141 18151
0 18153 5 1 1 18152
0 18154 7 1 2 23576 18153
0 18155 5 1 1 18154
0 18156 7 1 2 30811 31890
0 18157 7 1 2 35561 18156
0 18158 7 1 2 34617 18157
0 18159 7 1 2 27357 18158
0 18160 5 1 1 18159
0 18161 7 1 2 18155 18160
0 18162 5 1 1 18161
0 18163 7 1 2 23143 18162
0 18164 5 1 1 18163
0 18165 7 2 2 27932 37039
0 18166 7 1 2 36335 37044
0 18167 7 1 2 37057 18166
0 18168 5 1 1 18167
0 18169 7 1 2 18164 18168
0 18170 5 1 1 18169
0 18171 7 1 2 29467 18170
0 18172 5 1 1 18171
0 18173 7 1 2 35130 37042
0 18174 7 1 2 36171 18173
0 18175 7 1 2 37058 18174
0 18176 5 1 1 18175
0 18177 7 1 2 18172 18176
0 18178 5 1 1 18177
0 18179 7 1 2 31186 18178
0 18180 5 1 1 18179
0 18181 7 1 2 32986 36276
0 18182 5 1 1 18181
0 18183 7 1 2 34302 36239
0 18184 5 1 1 18183
0 18185 7 1 2 18182 18184
0 18186 5 2 1 18185
0 18187 7 1 2 31272 33383
0 18188 7 1 2 36920 18187
0 18189 7 1 2 29653 18188
0 18190 7 1 2 37059 18189
0 18191 5 1 1 18190
0 18192 7 1 2 18180 18191
0 18193 5 1 1 18192
0 18194 7 1 2 34093 18193
0 18195 5 1 1 18194
0 18196 7 1 2 18122 18195
0 18197 5 1 1 18196
0 18198 7 1 2 28848 18197
0 18199 5 1 1 18198
0 18200 7 1 2 22682 36214
0 18201 5 2 1 18200
0 18202 7 1 2 36143 37061
0 18203 5 1 1 18202
0 18204 7 1 2 26807 18203
0 18205 5 1 1 18204
0 18206 7 1 2 14353 18205
0 18207 5 1 1 18206
0 18208 7 1 2 33729 18207
0 18209 5 1 1 18208
0 18210 7 1 2 37013 37030
0 18211 7 1 2 36937 18210
0 18212 5 1 1 18211
0 18213 7 1 2 18209 18212
0 18214 5 1 1 18213
0 18215 7 1 2 24250 18214
0 18216 5 1 1 18215
0 18217 7 1 2 34303 36305
0 18218 5 2 1 18217
0 18219 7 1 2 37063 18145
0 18220 5 1 1 18219
0 18221 7 1 2 31917 36107
0 18222 7 1 2 18220 18221
0 18223 5 1 1 18222
0 18224 7 1 2 18216 18223
0 18225 5 1 1 18224
0 18226 7 4 2 26641 32554
0 18227 7 1 2 31758 37065
0 18228 7 1 2 34913 18227
0 18229 7 1 2 18225 18228
0 18230 5 1 1 18229
0 18231 7 1 2 18199 18230
0 18232 7 1 2 17875 18231
0 18233 7 1 2 17835 18232
0 18234 5 1 1 18233
0 18235 7 1 2 25682 26557
0 18236 7 1 2 18234 18235
0 18237 5 1 1 18236
0 18238 7 3 2 23327 31348
0 18239 7 4 2 28189 27084
0 18240 7 1 2 34223 37072
0 18241 5 1 1 18240
0 18242 7 1 2 27090 27034
0 18243 7 1 2 35868 34181
0 18244 7 1 2 18242 18243
0 18245 7 2 2 35481 18244
0 18246 5 1 1 37076
0 18247 7 1 2 26124 37077
0 18248 5 1 1 18247
0 18249 7 1 2 18241 18248
0 18250 5 2 1 18249
0 18251 7 1 2 27189 37078
0 18252 5 1 1 18251
0 18253 7 3 2 26642 26862
0 18254 7 1 2 21843 35869
0 18255 7 1 2 37080 18254
0 18256 7 1 2 36653 18255
0 18257 5 1 1 18256
0 18258 7 1 2 18252 18257
0 18259 5 1 1 18258
0 18260 7 1 2 37069 18259
0 18261 5 1 1 18260
0 18262 7 3 2 24348 26493
0 18263 7 2 2 36651 37083
0 18264 7 1 2 28453 30481
0 18265 7 1 2 37081 18264
0 18266 7 1 2 34228 18265
0 18267 7 1 2 37086 18266
0 18268 5 1 1 18267
0 18269 7 1 2 18261 18268
0 18270 5 1 1 18269
0 18271 7 1 2 24981 18270
0 18272 5 1 1 18271
0 18273 7 1 2 27886 28521
0 18274 5 2 1 18273
0 18275 7 1 2 22490 28513
0 18276 7 1 2 35305 18275
0 18277 5 1 1 18276
0 18278 7 1 2 37088 18277
0 18279 5 1 1 18278
0 18280 7 1 2 23874 18279
0 18281 5 2 1 18280
0 18282 7 1 2 24723 31781
0 18283 7 1 2 31794 18282
0 18284 5 1 1 18283
0 18285 7 1 2 37089 18284
0 18286 5 1 1 18285
0 18287 7 1 2 24487 18286
0 18288 5 1 1 18287
0 18289 7 1 2 37090 18288
0 18290 5 1 1 18289
0 18291 7 1 2 33384 18290
0 18292 5 1 1 18291
0 18293 7 2 2 23687 27534
0 18294 7 1 2 28522 37092
0 18295 7 1 2 33519 18294
0 18296 5 1 1 18295
0 18297 7 1 2 18292 18296
0 18298 5 1 1 18297
0 18299 7 1 2 26669 18298
0 18300 5 1 1 18299
0 18301 7 1 2 27952 37093
0 18302 7 1 2 33531 18301
0 18303 5 1 1 18302
0 18304 7 1 2 18300 18303
0 18305 5 1 1 18304
0 18306 7 1 2 23472 18305
0 18307 5 1 1 18306
0 18308 7 1 2 29355 28931
0 18309 7 1 2 36669 18308
0 18310 7 1 2 33532 18309
0 18311 5 1 1 18310
0 18312 7 1 2 18307 18311
0 18313 5 1 1 18312
0 18314 7 1 2 23028 18313
0 18315 5 1 1 18314
0 18316 7 1 2 23996 33533
0 18317 7 1 2 36634 18316
0 18318 5 1 1 18317
0 18319 7 1 2 18315 18318
0 18320 5 1 1 18319
0 18321 7 1 2 24876 18320
0 18322 5 1 1 18321
0 18323 7 1 2 23029 35088
0 18324 5 1 1 18323
0 18325 7 1 2 9826 18324
0 18326 5 1 1 18325
0 18327 7 1 2 23997 18326
0 18328 5 1 1 18327
0 18329 7 1 2 28183 33256
0 18330 5 1 1 18329
0 18331 7 1 2 23030 35080
0 18332 5 1 1 18331
0 18333 7 1 2 18330 18332
0 18334 5 1 1 18333
0 18335 7 1 2 27535 18334
0 18336 5 1 1 18335
0 18337 7 1 2 18328 18336
0 18338 5 1 1 18337
0 18339 7 1 2 26558 18338
0 18340 5 1 1 18339
0 18341 7 2 2 28402 36567
0 18342 7 1 2 25428 26161
0 18343 7 1 2 37094 18342
0 18344 5 1 1 18343
0 18345 7 1 2 32511 36639
0 18346 5 1 1 18345
0 18347 7 1 2 18344 18346
0 18348 7 1 2 18340 18347
0 18349 5 1 1 18348
0 18350 7 2 2 23688 18349
0 18351 7 1 2 34196 37096
0 18352 5 1 1 18351
0 18353 7 1 2 18322 18352
0 18354 5 1 1 18353
0 18355 7 1 2 24410 18354
0 18356 5 1 1 18355
0 18357 7 1 2 34214 37097
0 18358 5 1 1 18357
0 18359 7 1 2 18356 18358
0 18360 5 1 1 18359
0 18361 7 2 2 25357 31319
0 18362 7 1 2 18360 37098
0 18363 5 1 1 18362
0 18364 7 1 2 18272 18363
0 18365 5 1 1 18364
0 18366 7 1 2 25525 18365
0 18367 5 1 1 18366
0 18368 7 2 2 28849 28932
0 18369 7 1 2 36430 37100
0 18370 5 1 1 18369
0 18371 7 2 2 27035 36568
0 18372 7 1 2 26094 31251
0 18373 7 1 2 37102 18372
0 18374 5 1 1 18373
0 18375 7 1 2 18370 18374
0 18376 5 2 1 18375
0 18377 7 1 2 27190 37104
0 18378 5 1 1 18377
0 18379 7 2 2 36569 34231
0 18380 7 1 2 27070 28082
0 18381 7 1 2 37106 18380
0 18382 5 1 1 18381
0 18383 7 1 2 18378 18382
0 18384 5 1 1 18383
0 18385 7 1 2 37070 18384
0 18386 5 1 1 18385
0 18387 7 1 2 28454 31320
0 18388 7 1 2 37032 18387
0 18389 7 1 2 37107 18388
0 18390 5 1 1 18389
0 18391 7 1 2 18386 18390
0 18392 5 1 1 18391
0 18393 7 1 2 24982 18392
0 18394 5 1 1 18393
0 18395 7 3 2 28898 35870
0 18396 7 2 2 27874 37108
0 18397 5 1 1 37111
0 18398 7 1 2 24824 26039
0 18399 7 1 2 37103 18398
0 18400 5 1 1 18399
0 18401 7 1 2 18397 18400
0 18402 5 1 1 18401
0 18403 7 1 2 23875 18402
0 18404 5 1 1 18403
0 18405 7 1 2 27319 37112
0 18406 5 1 1 18405
0 18407 7 1 2 23031 28404
0 18408 7 1 2 29333 28550
0 18409 7 1 2 35040 18408
0 18410 7 1 2 18407 18409
0 18411 5 1 1 18410
0 18412 7 1 2 18406 18411
0 18413 7 1 2 18404 18412
0 18414 5 1 1 18413
0 18415 7 1 2 24349 18414
0 18416 5 1 1 18415
0 18417 7 1 2 28620 37109
0 18418 7 1 2 30870 18417
0 18419 5 1 1 18418
0 18420 7 1 2 18416 18419
0 18421 5 1 1 18420
0 18422 7 1 2 23998 18421
0 18423 5 1 1 18422
0 18424 7 1 2 29745 36422
0 18425 7 1 2 37101 18424
0 18426 5 1 1 18425
0 18427 7 1 2 18423 18426
0 18428 5 1 1 18427
0 18429 7 1 2 24724 37099
0 18430 7 1 2 18428 18429
0 18431 5 1 1 18430
0 18432 7 1 2 18394 18431
0 18433 5 1 1 18432
0 18434 7 1 2 25526 18433
0 18435 5 1 1 18434
0 18436 7 3 2 32512 32470
0 18437 7 4 2 24127 37113
0 18438 7 1 2 25868 37116
0 18439 5 1 1 18438
0 18440 7 1 2 26095 30723
0 18441 7 1 2 33001 18440
0 18442 5 1 1 18441
0 18443 7 1 2 18439 18442
0 18444 5 1 1 18443
0 18445 7 1 2 32927 18444
0 18446 5 1 1 18445
0 18447 7 2 2 28850 33169
0 18448 7 1 2 29629 37071
0 18449 5 1 1 18448
0 18450 7 1 2 28225 31321
0 18451 5 1 1 18450
0 18452 7 1 2 18449 18451
0 18453 5 4 1 18452
0 18454 7 1 2 37120 37122
0 18455 5 1 1 18454
0 18456 7 1 2 25629 26454
0 18457 7 1 2 31605 18456
0 18458 7 1 2 34059 18457
0 18459 7 1 2 28226 18458
0 18460 5 1 1 18459
0 18461 7 1 2 18455 18460
0 18462 7 1 2 18446 18461
0 18463 5 1 1 18462
0 18464 7 1 2 36407 18463
0 18465 5 1 1 18464
0 18466 7 1 2 18435 18465
0 18467 5 1 1 18466
0 18468 7 1 2 24877 18467
0 18469 5 1 1 18468
0 18470 7 1 2 36408 37114
0 18471 7 2 2 34244 18470
0 18472 7 1 2 35215 37126
0 18473 5 1 1 18472
0 18474 7 1 2 18469 18473
0 18475 5 1 1 18474
0 18476 7 1 2 24411 18475
0 18477 5 1 1 18476
0 18478 7 2 2 24878 34972
0 18479 7 1 2 37127 37128
0 18480 5 1 1 18479
0 18481 7 1 2 18477 18480
0 18482 5 1 1 18481
0 18483 7 1 2 25722 18482
0 18484 5 1 1 18483
0 18485 7 1 2 37123 36679
0 18486 5 1 1 18485
0 18487 7 2 2 21951 29540
0 18488 5 1 1 37130
0 18489 7 1 2 30724 37131
0 18490 5 1 1 18489
0 18491 7 1 2 31322 34977
0 18492 5 1 1 18491
0 18493 7 1 2 18490 18492
0 18494 5 1 1 18493
0 18495 7 1 2 21844 18494
0 18496 5 1 1 18495
0 18497 7 1 2 31323 32902
0 18498 5 1 1 18497
0 18499 7 1 2 18496 18498
0 18500 5 2 1 18499
0 18501 7 1 2 36690 37132
0 18502 5 1 1 18501
0 18503 7 1 2 18486 18502
0 18504 5 1 1 18503
0 18505 7 1 2 24350 18504
0 18506 5 1 1 18505
0 18507 7 1 2 37124 36677
0 18508 5 1 1 18507
0 18509 7 1 2 18506 18508
0 18510 5 1 1 18509
0 18511 7 1 2 25630 18510
0 18512 5 1 1 18511
0 18513 7 1 2 15615 36593
0 18514 5 1 1 18513
0 18515 7 1 2 22877 18514
0 18516 5 1 1 18515
0 18517 7 1 2 36699 18516
0 18518 5 1 1 18517
0 18519 7 1 2 22341 18518
0 18520 5 1 1 18519
0 18521 7 1 2 18520 36694
0 18522 5 1 1 18521
0 18523 7 1 2 37117 18522
0 18524 5 1 1 18523
0 18525 7 1 2 18512 18524
0 18526 5 1 1 18525
0 18527 7 1 2 24879 18526
0 18528 5 1 1 18527
0 18529 7 1 2 36570 34148
0 18530 5 1 1 18529
0 18531 7 1 2 31918 31897
0 18532 7 1 2 29365 18531
0 18533 5 1 1 18532
0 18534 7 1 2 18530 18533
0 18535 5 1 1 18534
0 18536 7 1 2 25723 18535
0 18537 5 1 1 18536
0 18538 7 1 2 34934 36496
0 18539 5 1 1 18538
0 18540 7 1 2 28303 35232
0 18541 7 1 2 36423 18540
0 18542 5 1 1 18541
0 18543 7 1 2 18539 18542
0 18544 7 1 2 18537 18543
0 18545 5 1 1 18544
0 18546 7 2 2 37115 18545
0 18547 7 1 2 35216 37134
0 18548 5 1 1 18547
0 18549 7 1 2 18528 18548
0 18550 5 1 1 18549
0 18551 7 1 2 24412 18550
0 18552 5 1 1 18551
0 18553 7 1 2 37129 37135
0 18554 5 1 1 18553
0 18555 7 1 2 18552 18554
0 18556 5 1 1 18555
0 18557 7 1 2 32987 18556
0 18558 5 1 1 18557
0 18559 7 1 2 35800 37118
0 18560 5 1 1 18559
0 18561 7 1 2 33750 37125
0 18562 5 1 1 18561
0 18563 7 1 2 33662 37119
0 18564 5 1 1 18563
0 18565 7 1 2 18562 18564
0 18566 5 1 1 18565
0 18567 7 1 2 26125 18566
0 18568 5 1 1 18567
0 18569 7 1 2 18560 18568
0 18570 5 1 1 18569
0 18571 7 1 2 23577 18570
0 18572 5 1 1 18571
0 18573 7 1 2 26126 34469
0 18574 7 1 2 37133 18573
0 18575 5 1 1 18574
0 18576 7 1 2 18572 18575
0 18577 5 1 1 18576
0 18578 7 1 2 36476 18577
0 18579 5 1 1 18578
0 18580 7 1 2 18558 18579
0 18581 7 1 2 18484 18580
0 18582 7 1 2 18367 18581
0 18583 5 1 1 18582
0 18584 7 1 2 30147 18583
0 18585 5 1 1 18584
0 18586 7 3 2 35960 36752
0 18587 7 3 2 25724 28851
0 18588 7 4 2 27250 28933
0 18589 7 1 2 37139 37142
0 18590 5 1 1 18589
0 18591 7 2 2 23237 30074
0 18592 7 2 2 34155 37146
0 18593 5 1 1 37148
0 18594 7 1 2 34182 37149
0 18595 5 1 1 18594
0 18596 7 1 2 18590 18595
0 18597 5 1 1 18596
0 18598 7 1 2 37136 18597
0 18599 5 1 1 18598
0 18600 7 1 2 37143 34197
0 18601 5 1 1 18600
0 18602 7 1 2 33652 37144
0 18603 5 1 1 18602
0 18604 7 1 2 18593 18603
0 18605 5 1 1 18604
0 18606 7 1 2 24351 18605
0 18607 5 1 1 18606
0 18608 7 1 2 35236 35187
0 18609 7 1 2 35974 18608
0 18610 5 1 1 18609
0 18611 7 1 2 22275 18610
0 18612 7 1 2 18607 18611
0 18613 5 1 1 18612
0 18614 7 1 2 24352 34385
0 18615 7 1 2 37147 18614
0 18616 5 1 1 18615
0 18617 7 1 2 22878 33554
0 18618 7 1 2 37145 18617
0 18619 5 1 1 18618
0 18620 7 1 2 24294 18619
0 18621 7 1 2 18616 18620
0 18622 5 1 1 18621
0 18623 7 1 2 24880 18622
0 18624 7 1 2 18613 18623
0 18625 5 1 1 18624
0 18626 7 1 2 18601 18625
0 18627 5 1 1 18626
0 18628 7 1 2 24413 18627
0 18629 5 1 1 18628
0 18630 7 1 2 28934 34183
0 18631 7 1 2 29279 18630
0 18632 7 1 2 34751 18631
0 18633 5 1 1 18632
0 18634 7 1 2 18629 18633
0 18635 5 1 1 18634
0 18636 7 1 2 36507 18635
0 18637 5 1 1 18636
0 18638 7 1 2 18599 18637
0 18639 5 1 1 18638
0 18640 7 1 2 26836 31324
0 18641 7 2 2 18639 18640
0 18642 5 1 1 37150
0 18643 7 1 2 29356 37151
0 18644 5 1 1 18643
0 18645 7 3 2 33629 32891
0 18646 7 1 2 30190 37152
0 18647 5 1 1 18646
0 18648 7 2 2 26700 37035
0 18649 7 3 2 34386 37155
0 18650 5 1 1 37157
0 18651 7 1 2 23876 24414
0 18652 7 1 2 37158 18651
0 18653 5 1 1 18652
0 18654 7 1 2 23578 35352
0 18655 7 1 2 30191 18654
0 18656 5 1 1 18655
0 18657 7 1 2 18653 18656
0 18658 5 1 1 18657
0 18659 7 1 2 24295 18658
0 18660 5 1 1 18659
0 18661 7 1 2 25693 28004
0 18662 7 1 2 37156 18661
0 18663 5 1 1 18662
0 18664 7 1 2 18660 18663
0 18665 5 1 1 18664
0 18666 7 1 2 28852 18665
0 18667 5 1 1 18666
0 18668 7 1 2 18647 18667
0 18669 5 1 1 18668
0 18670 7 1 2 18669 36520
0 18671 5 1 1 18670
0 18672 7 2 2 30249 31831
0 18673 7 1 2 36185 37160
0 18674 5 1 1 18673
0 18675 7 1 2 33908 36897
0 18676 5 1 1 18675
0 18677 7 1 2 18674 18676
0 18678 5 1 1 18677
0 18679 7 1 2 26887 18678
0 18680 5 1 1 18679
0 18681 7 1 2 28853 33901
0 18682 7 1 2 37159 18681
0 18683 5 2 1 18682
0 18684 7 5 2 30182 32487
0 18685 7 2 2 33909 37164
0 18686 7 1 2 28854 37169
0 18687 5 1 1 18686
0 18688 7 2 2 37162 18687
0 18689 5 1 1 37171
0 18690 7 1 2 23877 18689
0 18691 5 1 1 18690
0 18692 7 1 2 18680 18691
0 18693 5 1 1 18692
0 18694 7 1 2 36508 18693
0 18695 5 1 1 18694
0 18696 7 1 2 18671 18695
0 18697 5 1 1 18696
0 18698 7 1 2 32287 18697
0 18699 5 1 1 18698
0 18700 7 1 2 29357 37079
0 18701 5 1 1 18700
0 18702 7 1 2 31782 35041
0 18703 7 1 2 37033 18702
0 18704 5 1 1 18703
0 18705 7 1 2 37091 18704
0 18706 5 1 1 18705
0 18707 7 1 2 33385 18706
0 18708 5 1 1 18707
0 18709 7 2 2 23878 22781
0 18710 7 1 2 35131 37173
0 18711 7 1 2 28869 18710
0 18712 5 1 1 18711
0 18713 7 1 2 18708 18712
0 18714 5 1 1 18713
0 18715 7 1 2 26670 18714
0 18716 5 1 1 18715
0 18717 7 1 2 23879 27953
0 18718 7 1 2 35010 18717
0 18719 5 1 1 18718
0 18720 7 1 2 18716 18719
0 18721 5 1 1 18720
0 18722 7 1 2 24881 18721
0 18723 5 1 1 18722
0 18724 7 1 2 22782 22951
0 18725 7 1 2 36187 18724
0 18726 7 1 2 36661 18725
0 18727 5 1 1 18726
0 18728 7 1 2 18723 18727
0 18729 5 1 1 18728
0 18730 7 1 2 24415 18729
0 18731 5 1 1 18730
0 18732 7 1 2 34215 37174
0 18733 7 1 2 36662 18732
0 18734 5 1 1 18733
0 18735 7 1 2 18731 18734
0 18736 5 1 1 18735
0 18737 7 1 2 26863 18736
0 18738 5 1 1 18737
0 18739 7 1 2 18701 18738
0 18740 5 1 1 18739
0 18741 7 1 2 25527 18740
0 18742 5 1 1 18741
0 18743 7 3 2 23579 36799
0 18744 5 1 1 37175
0 18745 7 1 2 24488 37176
0 18746 5 1 1 18745
0 18747 7 2 2 29334 30250
0 18748 7 2 2 33989 37178
0 18749 7 3 2 24251 29313
0 18750 7 1 2 34184 37182
0 18751 7 1 2 37180 18750
0 18752 5 1 1 18751
0 18753 7 1 2 18746 18752
0 18754 5 1 1 18753
0 18755 7 1 2 34237 18754
0 18756 5 1 1 18755
0 18757 7 1 2 16272 18756
0 18758 5 1 1 18757
0 18759 7 1 2 23880 18758
0 18760 5 1 1 18759
0 18761 7 1 2 37179 36887
0 18762 7 1 2 36971 18761
0 18763 5 1 1 18762
0 18764 7 1 2 18744 18763
0 18765 5 1 1 18764
0 18766 7 2 2 23999 27323
0 18767 5 1 1 37185
0 18768 7 1 2 18765 37186
0 18769 5 1 1 18768
0 18770 7 1 2 18760 18769
0 18771 5 1 1 18770
0 18772 7 1 2 32988 18771
0 18773 5 1 1 18772
0 18774 7 1 2 29358 34935
0 18775 5 1 1 18774
0 18776 7 1 2 26096 34455
0 18777 7 1 2 35553 18776
0 18778 5 1 1 18777
0 18779 7 1 2 18775 18778
0 18780 5 1 1 18779
0 18781 7 1 2 25631 18780
0 18782 5 1 1 18781
0 18783 7 1 2 23881 35248
0 18784 5 1 1 18783
0 18785 7 1 2 18782 18784
0 18786 5 1 1 18785
0 18787 7 1 2 24882 18786
0 18788 5 1 1 18787
0 18789 7 1 2 34936 36837
0 18790 5 1 1 18789
0 18791 7 1 2 18788 18790
0 18792 5 1 1 18791
0 18793 7 1 2 24416 18792
0 18794 5 1 1 18793
0 18795 7 1 2 23882 32689
0 18796 7 1 2 34937 18795
0 18797 5 1 1 18796
0 18798 7 1 2 18794 18797
0 18799 5 1 1 18798
0 18800 7 1 2 36477 18799
0 18801 5 1 1 18800
0 18802 7 1 2 36709 37040
0 18803 5 1 1 18802
0 18804 7 1 2 26417 34162
0 18805 7 1 2 37095 18804
0 18806 5 1 1 18805
0 18807 7 1 2 24883 29359
0 18808 7 1 2 15304 18807
0 18809 5 1 1 18808
0 18810 7 1 2 18806 18809
0 18811 5 1 1 18810
0 18812 7 1 2 24417 18811
0 18813 5 1 1 18812
0 18814 7 2 2 25764 31539
0 18815 7 1 2 23689 32488
0 18816 7 2 2 23883 24175
0 18817 7 1 2 37189 34169
0 18818 7 1 2 18815 18817
0 18819 7 1 2 37187 18818
0 18820 5 1 1 18819
0 18821 7 1 2 18813 18820
0 18822 5 1 1 18821
0 18823 7 1 2 28855 18822
0 18824 5 1 1 18823
0 18825 7 1 2 23884 32698
0 18826 5 1 1 18825
0 18827 7 1 2 18767 18826
0 18828 5 1 1 18827
0 18829 7 1 2 26097 18828
0 18830 5 1 1 18829
0 18831 7 1 2 655 18830
0 18832 5 1 1 18831
0 18833 7 1 2 36666 18832
0 18834 5 1 1 18833
0 18835 7 1 2 24000 33190
0 18836 5 1 1 18835
0 18837 7 1 2 6393 18836
0 18838 5 1 1 18837
0 18839 7 1 2 23885 18838
0 18840 5 1 1 18839
0 18841 7 1 2 31257 8856
0 18842 5 2 1 18841
0 18843 7 1 2 23886 31258
0 18844 5 1 1 18843
0 18845 7 1 2 24001 18844
0 18846 7 1 2 37191 18845
0 18847 5 1 1 18846
0 18848 7 1 2 18840 18847
0 18849 5 1 1 18848
0 18850 7 1 2 27036 35855
0 18851 7 1 2 33020 18850
0 18852 7 2 2 29337 18851
0 18853 7 1 2 18849 37193
0 18854 5 1 1 18853
0 18855 7 1 2 18834 18854
0 18856 7 1 2 18824 18855
0 18857 5 1 1 18856
0 18858 7 1 2 25725 18857
0 18859 5 1 1 18858
0 18860 7 1 2 18803 18859
0 18861 7 1 2 18801 18860
0 18862 7 1 2 18773 18861
0 18863 7 1 2 18742 18862
0 18864 5 1 1 18863
0 18865 7 1 2 32341 18864
0 18866 5 1 1 18865
0 18867 7 1 2 18699 18866
0 18868 5 1 1 18867
0 18869 7 1 2 22091 18868
0 18870 5 1 1 18869
0 18871 7 1 2 18644 18870
0 18872 5 1 1 18871
0 18873 7 1 2 23032 18872
0 18874 5 1 1 18873
0 18875 7 1 2 32242 36792
0 18876 5 1 1 18875
0 18877 7 1 2 28856 36775
0 18878 5 1 1 18877
0 18879 7 1 2 36786 35527
0 18880 5 1 1 18879
0 18881 7 1 2 18878 18880
0 18882 5 1 1 18881
0 18883 7 1 2 25954 18882
0 18884 5 1 1 18883
0 18885 7 1 2 35806 36424
0 18886 5 1 1 18885
0 18887 7 1 2 18884 18886
0 18888 5 2 1 18887
0 18889 7 1 2 27368 32489
0 18890 7 1 2 37195 18889
0 18891 5 1 1 18890
0 18892 7 1 2 18876 18891
0 18893 5 1 1 18892
0 18894 7 1 2 23690 18893
0 18895 5 1 1 18894
0 18896 7 1 2 33386 37084
0 18897 7 3 2 24662 36379
0 18898 7 2 2 31375 37190
0 18899 7 1 2 37200 36811
0 18900 7 1 2 37197 18899
0 18901 7 1 2 18896 18900
0 18902 5 1 1 18901
0 18903 7 1 2 18895 18902
0 18904 5 1 1 18903
0 18905 7 1 2 32989 18904
0 18906 5 1 1 18905
0 18907 7 1 2 32243 36375
0 18908 7 1 2 36409 18907
0 18909 7 1 2 34218 18908
0 18910 5 1 1 18909
0 18911 7 1 2 26671 31215
0 18912 7 1 2 33108 18911
0 18913 7 1 2 35812 18912
0 18914 5 1 1 18913
0 18915 7 1 2 18910 18914
0 18916 5 1 1 18915
0 18917 7 1 2 23691 18916
0 18918 5 1 1 18917
0 18919 7 1 2 36925 36839
0 18920 7 1 2 36655 18919
0 18921 7 1 2 37087 18920
0 18922 5 1 1 18921
0 18923 7 1 2 18918 18922
0 18924 5 1 1 18923
0 18925 7 1 2 26864 18924
0 18926 5 1 1 18925
0 18927 7 1 2 32244 32928
0 18928 7 1 2 31832 18927
0 18929 5 1 1 18928
0 18930 7 2 2 32490 32036
0 18931 7 1 2 31055 32916
0 18932 7 1 2 37202 18931
0 18933 5 1 1 18932
0 18934 7 1 2 18929 18933
0 18935 5 1 1 18934
0 18936 7 1 2 36410 18935
0 18937 5 1 1 18936
0 18938 7 1 2 36670 34916
0 18939 7 1 2 37203 18938
0 18940 5 1 1 18939
0 18941 7 1 2 18937 18940
0 18942 5 1 1 18941
0 18943 7 1 2 23692 18942
0 18944 5 1 1 18943
0 18945 7 1 2 25773 26877
0 18946 7 1 2 31544 18945
0 18947 7 1 2 25791 34232
0 18948 7 1 2 37201 18947
0 18949 7 1 2 18946 18948
0 18950 5 1 1 18949
0 18951 7 1 2 18944 18950
0 18952 5 1 1 18951
0 18953 7 1 2 25726 18952
0 18954 5 1 1 18953
0 18955 7 1 2 29258 32245
0 18956 7 1 2 35813 18955
0 18957 5 1 1 18956
0 18958 7 1 2 30308 31273
0 18959 7 1 2 35054 18958
0 18960 7 1 2 34208 37085
0 18961 7 1 2 18959 18960
0 18962 5 1 1 18961
0 18963 7 1 2 18957 18962
0 18964 5 1 1 18963
0 18965 7 1 2 36478 18964
0 18966 5 1 1 18965
0 18967 7 1 2 18954 18966
0 18968 7 1 2 18926 18967
0 18969 7 1 2 18906 18968
0 18970 5 1 1 18969
0 18971 7 1 2 32342 18970
0 18972 5 1 1 18971
0 18973 7 1 2 34797 34481
0 18974 7 1 2 37165 18973
0 18975 5 1 1 18974
0 18976 7 1 2 25727 30881
0 18977 7 1 2 37036 18976
0 18978 7 1 2 32246 18977
0 18979 5 1 1 18978
0 18980 7 1 2 18975 18979
0 18981 5 1 1 18980
0 18982 7 1 2 24418 18981
0 18983 5 1 1 18982
0 18984 7 2 2 30178 35361
0 18985 7 1 2 34752 36926
0 18986 7 1 2 37204 18985
0 18987 5 1 1 18986
0 18988 7 1 2 18983 18987
0 18989 5 1 1 18988
0 18990 7 1 2 28857 18989
0 18991 5 1 1 18990
0 18992 7 1 2 37166 35262
0 18993 7 1 2 31833 18992
0 18994 5 1 1 18993
0 18995 7 1 2 18991 18994
0 18996 5 1 1 18995
0 18997 7 1 2 36521 18996
0 18998 5 1 1 18997
0 18999 7 1 2 26888 36578
0 19000 7 1 2 31834 18999
0 19001 5 2 1 19000
0 19002 7 1 2 37163 37206
0 19003 5 1 1 19002
0 19004 7 1 2 32247 19003
0 19005 5 1 1 19004
0 19006 7 1 2 22092 28858
0 19007 7 1 2 37170 19006
0 19008 5 1 1 19007
0 19009 7 1 2 19005 19008
0 19010 5 1 1 19009
0 19011 7 1 2 36509 19010
0 19012 5 1 1 19011
0 19013 7 1 2 18998 19012
0 19014 5 1 1 19013
0 19015 7 1 2 32288 19014
0 19016 5 1 1 19015
0 19017 7 1 2 24002 19016
0 19018 7 1 2 18972 19017
0 19019 5 1 1 19018
0 19020 7 1 2 28938 36671
0 19021 7 2 2 34198 19020
0 19022 5 1 1 37208
0 19023 7 1 2 37073 35011
0 19024 5 1 1 19023
0 19025 7 1 2 25728 37105
0 19026 5 1 1 19025
0 19027 7 1 2 18246 19026
0 19028 7 1 2 19024 19027
0 19029 5 1 1 19028
0 19030 7 1 2 24884 19029
0 19031 5 1 1 19030
0 19032 7 1 2 19022 19031
0 19033 5 1 1 19032
0 19034 7 1 2 24419 19033
0 19035 5 1 1 19034
0 19036 7 1 2 31092 34209
0 19037 7 2 2 28935 31540
0 19038 7 1 2 35372 37210
0 19039 7 1 2 19036 19038
0 19040 5 1 1 19039
0 19041 7 1 2 19035 19040
0 19042 5 1 1 19041
0 19043 7 1 2 27191 19042
0 19044 5 1 1 19043
0 19045 7 1 2 27471 37082
0 19046 7 1 2 32203 19045
0 19047 7 1 2 36776 19046
0 19048 5 1 1 19047
0 19049 7 1 2 19044 19048
0 19050 5 1 1 19049
0 19051 7 1 2 35050 19050
0 19052 5 1 1 19051
0 19053 7 1 2 26929 30282
0 19054 7 2 2 37196 19053
0 19055 7 1 2 37054 37212
0 19056 5 1 1 19055
0 19057 7 1 2 19052 19056
0 19058 5 1 1 19057
0 19059 7 1 2 24983 19058
0 19060 5 1 1 19059
0 19061 7 1 2 34590 36544
0 19062 5 1 1 19061
0 19063 7 1 2 32917 34128
0 19064 5 1 1 19063
0 19065 7 1 2 19062 19064
0 19066 7 1 2 15631 19065
0 19067 5 1 1 19066
0 19068 7 1 2 22879 19067
0 19069 5 1 1 19068
0 19070 7 2 2 28304 31176
0 19071 7 1 2 35531 37214
0 19072 5 1 1 19071
0 19073 7 1 2 19069 19072
0 19074 5 1 1 19073
0 19075 7 1 2 22342 19074
0 19076 5 1 1 19075
0 19077 7 1 2 28710 33331
0 19078 7 1 2 37215 19077
0 19079 5 1 1 19078
0 19080 7 1 2 19076 19079
0 19081 5 1 1 19080
0 19082 7 1 2 32733 19081
0 19083 5 1 1 19082
0 19084 7 1 2 27192 31305
0 19085 7 1 2 36383 19084
0 19086 7 1 2 37140 19085
0 19087 5 1 1 19086
0 19088 7 1 2 19083 19087
0 19089 5 1 1 19088
0 19090 7 1 2 23693 19089
0 19091 5 1 1 19090
0 19092 7 1 2 25729 34245
0 19093 5 1 1 19092
0 19094 7 1 2 34304 34938
0 19095 5 1 1 19094
0 19096 7 1 2 19093 19095
0 19097 5 1 1 19096
0 19098 7 1 2 27193 19097
0 19099 5 1 1 19098
0 19100 7 1 2 34305 35897
0 19101 5 1 1 19100
0 19102 7 1 2 19099 19101
0 19103 5 1 1 19102
0 19104 7 1 2 24128 26479
0 19105 7 1 2 19103 19104
0 19106 5 1 1 19105
0 19107 7 1 2 19091 19106
0 19108 5 1 1 19107
0 19109 7 1 2 26127 19108
0 19110 5 1 1 19109
0 19111 7 1 2 34306 33740
0 19112 5 1 1 19111
0 19113 7 1 2 33814 33782
0 19114 5 1 1 19113
0 19115 7 1 2 19112 19114
0 19116 5 1 1 19115
0 19117 7 1 2 23580 19116
0 19118 5 1 1 19117
0 19119 7 1 2 25696 36599
0 19120 5 1 1 19119
0 19121 7 1 2 25730 6263
0 19122 5 1 1 19121
0 19123 7 1 2 34249 19122
0 19124 7 1 2 19120 19123
0 19125 5 1 1 19124
0 19126 7 1 2 19118 19125
0 19127 5 1 1 19126
0 19128 7 1 2 32734 34954
0 19129 7 1 2 19127 19128
0 19130 5 1 1 19129
0 19131 7 1 2 19110 19130
0 19132 5 1 1 19131
0 19133 7 1 2 26229 36411
0 19134 7 1 2 19132 19133
0 19135 5 1 1 19134
0 19136 7 1 2 36795 32735
0 19137 5 1 1 19136
0 19138 7 1 2 37181 36972
0 19139 5 1 1 19138
0 19140 7 1 2 27194 37177
0 19141 5 1 1 19140
0 19142 7 1 2 19139 19141
0 19143 5 1 1 19142
0 19144 7 1 2 24984 37066
0 19145 7 1 2 19143 19144
0 19146 5 1 1 19145
0 19147 7 1 2 19137 19146
0 19148 5 1 1 19147
0 19149 7 1 2 32990 19148
0 19150 5 1 1 19149
0 19151 7 1 2 35554 33239
0 19152 7 1 2 37213 19151
0 19153 5 1 1 19152
0 19154 7 1 2 19150 19153
0 19155 7 1 2 19135 19154
0 19156 7 1 2 19060 19155
0 19157 5 1 1 19156
0 19158 7 1 2 32343 19157
0 19159 5 1 1 19158
0 19160 7 1 2 30229 33911
0 19161 5 1 1 19160
0 19162 7 2 2 27237 29930
0 19163 7 2 2 25288 30251
0 19164 7 1 2 37218 35687
0 19165 7 1 2 37216 19164
0 19166 5 1 1 19165
0 19167 7 1 2 19161 19166
0 19168 5 1 1 19167
0 19169 7 1 2 28859 19168
0 19170 5 1 1 19169
0 19171 7 1 2 25289 33387
0 19172 7 1 2 37217 19171
0 19173 7 1 2 37161 19172
0 19174 5 1 1 19173
0 19175 7 1 2 19170 19174
0 19176 5 1 1 19175
0 19177 7 1 2 27195 19176
0 19178 5 1 1 19177
0 19179 7 1 2 37172 37207
0 19180 5 1 1 19179
0 19181 7 1 2 32736 19180
0 19182 5 1 1 19181
0 19183 7 1 2 27536 28860
0 19184 7 1 2 30884 19183
0 19185 7 1 2 33912 19184
0 19186 5 1 1 19185
0 19187 7 1 2 19182 19186
0 19188 7 1 2 19178 19187
0 19189 5 1 1 19188
0 19190 7 1 2 36510 19189
0 19191 5 1 1 19190
0 19192 7 1 2 37167 34049
0 19193 5 1 1 19192
0 19194 7 1 2 18650 19193
0 19195 5 1 1 19194
0 19196 7 1 2 24296 19195
0 19197 5 1 1 19196
0 19198 7 1 2 25694 26701
0 19199 7 1 2 27542 30252
0 19200 7 1 2 19198 19199
0 19201 5 1 1 19200
0 19202 7 1 2 19197 19201
0 19203 5 1 1 19202
0 19204 7 1 2 24420 19203
0 19205 5 1 1 19204
0 19206 7 1 2 37205 34754
0 19207 5 1 1 19206
0 19208 7 1 2 19205 19207
0 19209 5 1 1 19208
0 19210 7 1 2 32737 19209
0 19211 5 1 1 19210
0 19212 7 1 2 26702 32491
0 19213 7 1 2 36308 19212
0 19214 7 1 2 35782 19213
0 19215 5 1 1 19214
0 19216 7 1 2 19211 19215
0 19217 5 1 1 19216
0 19218 7 1 2 28861 19217
0 19219 5 1 1 19218
0 19220 7 1 2 23887 30423
0 19221 5 1 1 19220
0 19222 7 1 2 26703 28009
0 19223 5 1 1 19222
0 19224 7 1 2 19221 19223
0 19225 5 1 1 19224
0 19226 7 1 2 24985 19225
0 19227 5 1 1 19226
0 19228 7 1 2 30674 35555
0 19229 5 1 1 19228
0 19230 7 1 2 19227 19229
0 19231 5 1 1 19230
0 19232 7 1 2 37153 19231
0 19233 5 1 1 19232
0 19234 7 1 2 30471 33471
0 19235 7 1 2 36894 19234
0 19236 5 1 1 19235
0 19237 7 4 2 27270 37014
0 19238 7 1 2 24297 22683
0 19239 7 1 2 34050 19238
0 19240 7 1 2 37220 19239
0 19241 5 1 1 19240
0 19242 7 1 2 19236 19241
0 19243 5 1 1 19242
0 19244 7 1 2 24421 19243
0 19245 5 1 1 19244
0 19246 7 1 2 27543 33606
0 19247 7 1 2 37221 19246
0 19248 5 1 1 19247
0 19249 7 1 2 19245 19248
0 19250 5 1 1 19249
0 19251 7 1 2 28862 19250
0 19252 5 1 1 19251
0 19253 7 1 2 30230 37154
0 19254 5 1 1 19253
0 19255 7 1 2 19252 19254
0 19256 5 1 1 19255
0 19257 7 1 2 27196 19256
0 19258 5 1 1 19257
0 19259 7 1 2 19233 19258
0 19260 7 1 2 19219 19259
0 19261 5 1 1 19260
0 19262 7 1 2 36522 19261
0 19263 5 1 1 19262
0 19264 7 1 2 19191 19263
0 19265 5 1 1 19264
0 19266 7 1 2 32289 19265
0 19267 5 1 1 19266
0 19268 7 1 2 21952 19267
0 19269 7 1 2 19159 19268
0 19270 5 1 1 19269
0 19271 7 1 2 19019 19270
0 19272 5 1 1 19271
0 19273 7 1 2 25528 37209
0 19274 5 1 1 19273
0 19275 7 1 2 25731 36434
0 19276 5 1 1 19275
0 19277 7 1 2 32991 36497
0 19278 5 1 1 19277
0 19279 7 1 2 15406 19278
0 19280 5 2 1 19279
0 19281 7 1 2 34445 37224
0 19282 5 1 1 19281
0 19283 7 1 2 34433 37074
0 19284 5 1 1 19283
0 19285 7 1 2 19282 19284
0 19286 7 1 2 19276 19285
0 19287 5 1 1 19286
0 19288 7 1 2 28863 19287
0 19289 5 1 1 19288
0 19290 7 1 2 26808 32992
0 19291 7 1 2 36425 19290
0 19292 5 1 1 19291
0 19293 7 1 2 26601 26837
0 19294 7 1 2 36571 19293
0 19295 5 1 1 19294
0 19296 7 1 2 15820 19295
0 19297 7 1 2 19292 19296
0 19298 5 1 1 19297
0 19299 7 1 2 25732 19298
0 19300 5 1 1 19299
0 19301 7 1 2 31252 33850
0 19302 7 1 2 36580 19301
0 19303 5 1 1 19302
0 19304 7 1 2 34422 37225
0 19305 5 1 1 19304
0 19306 7 1 2 19303 19305
0 19307 7 1 2 19300 19306
0 19308 5 1 1 19307
0 19309 7 1 2 27909 19308
0 19310 5 1 1 19309
0 19311 7 2 2 22343 24663
0 19312 7 1 2 29400 37226
0 19313 7 1 2 34961 19312
0 19314 7 2 2 24176 34510
0 19315 7 1 2 30866 37228
0 19316 7 1 2 19313 19315
0 19317 5 1 1 19316
0 19318 7 1 2 19310 19317
0 19319 7 1 2 19289 19318
0 19320 5 1 1 19319
0 19321 7 1 2 24885 19320
0 19322 5 1 1 19321
0 19323 7 1 2 19274 19322
0 19324 5 1 1 19323
0 19325 7 1 2 24422 19324
0 19326 5 1 1 19325
0 19327 7 1 2 27650 36267
0 19328 7 1 2 31554 19327
0 19329 7 1 2 34210 37229
0 19330 7 1 2 19328 19329
0 19331 5 1 1 19330
0 19332 7 1 2 19326 19331
0 19333 5 1 1 19332
0 19334 7 1 2 22093 32344
0 19335 7 1 2 19333 19334
0 19336 5 1 1 19335
0 19337 7 1 2 18642 19336
0 19338 5 1 1 19337
0 19339 7 1 2 24003 19338
0 19340 5 1 1 19339
0 19341 7 1 2 36511 34219
0 19342 5 1 1 19341
0 19343 7 1 2 37137 37141
0 19344 5 1 1 19343
0 19345 7 1 2 19342 19344
0 19346 5 1 1 19345
0 19347 7 1 2 30672 31620
0 19348 7 1 2 30822 19347
0 19349 7 1 2 32530 19348
0 19350 7 1 2 19346 19349
0 19351 5 1 1 19350
0 19352 7 1 2 19340 19351
0 19353 5 1 1 19352
0 19354 7 1 2 27537 19353
0 19355 5 1 1 19354
0 19356 7 1 2 25683 19355
0 19357 7 1 2 19272 19356
0 19358 7 1 2 18874 19357
0 19359 7 1 2 18585 19358
0 19360 5 1 1 19359
0 19361 7 1 2 36426 35583
0 19362 5 1 1 19361
0 19363 7 1 2 35585 36966
0 19364 5 1 1 19363
0 19365 7 1 2 19362 19364
0 19366 5 1 1 19365
0 19367 7 1 2 25733 19366
0 19368 5 1 1 19367
0 19369 7 1 2 37183 37198
0 19370 5 1 1 19369
0 19371 7 1 2 36492 19370
0 19372 5 1 1 19371
0 19373 7 1 2 27197 19372
0 19374 5 1 1 19373
0 19375 7 1 2 15668 36493
0 19376 5 1 1 19375
0 19377 7 1 2 21953 19376
0 19378 5 1 1 19377
0 19379 7 1 2 28364 35856
0 19380 7 1 2 29688 19379
0 19381 5 2 1 19380
0 19382 7 1 2 19378 37230
0 19383 7 1 2 19374 19382
0 19384 5 1 1 19383
0 19385 7 1 2 33428 19384
0 19386 5 1 1 19385
0 19387 7 1 2 19368 19386
0 19388 5 1 1 19387
0 19389 7 1 2 25632 19388
0 19390 5 1 1 19389
0 19391 7 1 2 22880 28954
0 19392 7 1 2 36781 33962
0 19393 7 1 2 19391 19392
0 19394 5 1 1 19393
0 19395 7 1 2 23581 19394
0 19396 7 1 2 19390 19395
0 19397 5 1 1 19396
0 19398 7 1 2 35593 36964
0 19399 5 1 1 19398
0 19400 7 1 2 32609 36969
0 19401 5 1 1 19400
0 19402 7 1 2 19399 19401
0 19403 5 1 1 19402
0 19404 7 1 2 34591 19403
0 19405 5 1 1 19404
0 19406 7 1 2 35594 35590
0 19407 5 1 1 19406
0 19408 7 1 2 25955 35591
0 19409 5 1 1 19408
0 19410 7 1 2 11700 19409
0 19411 5 1 1 19410
0 19412 7 1 2 32610 19411
0 19413 5 1 1 19412
0 19414 7 1 2 19407 19413
0 19415 5 1 1 19414
0 19416 7 1 2 36585 19415
0 19417 5 1 1 19416
0 19418 7 1 2 25529 19417
0 19419 7 1 2 19405 19418
0 19420 5 1 1 19419
0 19421 7 1 2 32993 19420
0 19422 7 1 2 19397 19421
0 19423 5 1 1 19422
0 19424 7 1 2 34605 35595
0 19425 5 1 1 19424
0 19426 7 1 2 32611 34607
0 19427 5 1 1 19426
0 19428 7 1 2 19425 19427
0 19429 5 1 1 19428
0 19430 7 1 2 25530 19429
0 19431 5 1 1 19430
0 19432 7 1 2 35933 35586
0 19433 5 1 1 19432
0 19434 7 1 2 30932 34609
0 19435 5 1 1 19434
0 19436 7 1 2 19433 19435
0 19437 5 1 1 19436
0 19438 7 1 2 28680 19437
0 19439 5 1 1 19438
0 19440 7 1 2 19431 19439
0 19441 5 1 1 19440
0 19442 7 1 2 36412 19441
0 19443 5 1 1 19442
0 19444 7 1 2 26214 27095
0 19445 7 1 2 31932 19444
0 19446 5 1 1 19445
0 19447 7 1 2 19443 19446
0 19448 5 1 1 19447
0 19449 7 1 2 25734 19448
0 19450 5 1 1 19449
0 19451 7 1 2 32612 34641
0 19452 5 1 1 19451
0 19453 7 1 2 33534 35596
0 19454 5 1 1 19453
0 19455 7 1 2 19452 19454
0 19456 5 1 1 19455
0 19457 7 1 2 25531 19456
0 19458 5 1 1 19457
0 19459 7 1 2 19458 34996
0 19460 5 1 1 19459
0 19461 7 1 2 36479 19460
0 19462 5 1 1 19461
0 19463 7 1 2 28244 35857
0 19464 7 1 2 36942 19463
0 19465 7 1 2 37211 33717
0 19466 7 1 2 19464 19465
0 19467 5 1 1 19466
0 19468 7 1 2 30213 34286
0 19469 5 1 1 19468
0 19470 7 1 2 27198 34307
0 19471 7 1 2 19469 19470
0 19472 5 1 1 19471
0 19473 7 1 2 27472 34287
0 19474 5 1 1 19473
0 19475 7 1 2 21954 34308
0 19476 7 1 2 19474 19475
0 19477 5 1 1 19476
0 19478 7 1 2 23389 28365
0 19479 7 1 2 35094 19478
0 19480 5 1 1 19479
0 19481 7 1 2 19477 19480
0 19482 7 1 2 19472 19481
0 19483 5 1 1 19482
0 19484 7 1 2 36413 19483
0 19485 7 1 2 36875 19484
0 19486 5 1 1 19485
0 19487 7 1 2 19467 19486
0 19488 5 1 1 19487
0 19489 7 1 2 23582 19488
0 19490 5 1 1 19489
0 19491 7 1 2 19462 19490
0 19492 7 1 2 19450 19491
0 19493 7 1 2 19423 19492
0 19494 5 1 1 19493
0 19495 7 1 2 32345 19494
0 19496 5 1 1 19495
0 19497 7 1 2 25735 36537
0 19498 5 1 1 19497
0 19499 7 1 2 36572 36009
0 19500 5 1 1 19499
0 19501 7 1 2 19498 19500
0 19502 5 1 1 19501
0 19503 7 2 2 28438 28961
0 19504 7 1 2 26704 37232
0 19505 7 1 2 33269 19504
0 19506 7 1 2 19502 19505
0 19507 5 1 1 19506
0 19508 7 1 2 23768 19507
0 19509 7 1 2 19496 19508
0 19510 5 1 1 19509
0 19511 7 1 2 32590 19510
0 19512 7 1 2 19360 19511
0 19513 5 1 1 19512
0 19514 7 1 2 25532 35808
0 19515 5 1 1 19514
0 19516 7 1 2 23583 33544
0 19517 5 1 1 19516
0 19518 7 1 2 29270 29373
0 19519 7 1 2 36026 19518
0 19520 7 1 2 19517 19519
0 19521 7 1 2 19515 19520
0 19522 5 1 1 19521
0 19523 7 1 2 30812 30965
0 19524 7 1 2 36087 19523
0 19525 7 1 2 25780 19524
0 19526 7 1 2 35965 19525
0 19527 5 1 1 19526
0 19528 7 1 2 19522 19527
0 19529 5 1 1 19528
0 19530 7 1 2 30757 19529
0 19531 5 1 1 19530
0 19532 7 2 2 27786 31405
0 19533 7 1 2 29520 32496
0 19534 7 1 2 37234 19533
0 19535 7 1 2 33741 19534
0 19536 5 1 1 19535
0 19537 7 1 2 19531 19536
0 19538 5 1 1 19537
0 19539 7 1 2 22783 19538
0 19540 5 1 1 19539
0 19541 7 1 2 28056 31308
0 19542 7 1 2 34939 19541
0 19543 5 1 1 19542
0 19544 7 1 2 34191 32178
0 19545 5 1 1 19544
0 19546 7 1 2 9334 19545
0 19547 5 1 1 19546
0 19548 7 1 2 26188 30438
0 19549 7 1 2 19547 19548
0 19550 5 1 1 19549
0 19551 7 1 2 19543 19550
0 19552 5 1 1 19551
0 19553 7 1 2 33122 31891
0 19554 7 1 2 19552 19553
0 19555 5 1 1 19554
0 19556 7 1 2 19540 19555
0 19557 5 1 1 19556
0 19558 7 1 2 22684 19557
0 19559 5 1 1 19558
0 19560 7 1 2 29063 29521
0 19561 5 1 1 19560
0 19562 7 1 2 30344 19561
0 19563 5 1 1 19562
0 19564 7 1 2 34940 19563
0 19565 5 1 1 19564
0 19566 7 2 2 24353 34813
0 19567 7 1 2 28588 36058
0 19568 7 1 2 30582 19567
0 19569 7 1 2 37236 19568
0 19570 5 1 1 19569
0 19571 7 1 2 19565 19570
0 19572 5 1 1 19571
0 19573 7 1 2 26831 32994
0 19574 7 1 2 33123 19573
0 19575 7 1 2 19572 19574
0 19576 5 1 1 19575
0 19577 7 1 2 19559 19576
0 19578 5 1 1 19577
0 19579 7 1 2 22237 19578
0 19580 5 1 1 19579
0 19581 7 2 2 36128 34283
0 19582 5 1 1 37238
0 19583 7 1 2 31259 7838
0 19584 5 1 1 19583
0 19585 7 1 2 36306 19584
0 19586 5 1 1 19585
0 19587 7 1 2 36138 19586
0 19588 5 1 1 19587
0 19589 7 1 2 23473 19588
0 19590 5 1 1 19589
0 19591 7 2 2 24725 27974
0 19592 5 1 1 37240
0 19593 7 1 2 24986 37241
0 19594 5 1 1 19593
0 19595 7 1 2 19590 19594
0 19596 5 1 1 19595
0 19597 7 1 2 29098 19596
0 19598 5 1 1 19597
0 19599 7 1 2 19582 19598
0 19600 5 2 1 19599
0 19601 7 1 2 34941 37242
0 19602 5 1 1 19601
0 19603 7 1 2 36139 37062
0 19604 5 1 1 19603
0 19605 7 1 2 23474 19604
0 19606 5 1 1 19605
0 19607 7 1 2 19592 19606
0 19608 5 1 1 19607
0 19609 7 1 2 35233 33498
0 19610 7 1 2 19608 19609
0 19611 5 1 1 19610
0 19612 7 1 2 19602 19611
0 19613 5 1 1 19612
0 19614 7 1 2 21955 19613
0 19615 5 1 1 19614
0 19616 7 2 2 22571 37239
0 19617 5 1 1 37244
0 19618 7 1 2 34942 37245
0 19619 5 1 1 19618
0 19620 7 1 2 19615 19619
0 19621 5 1 1 19620
0 19622 7 1 2 27787 31376
0 19623 7 1 2 19621 19622
0 19624 5 1 1 19623
0 19625 7 1 2 19580 19624
0 19626 5 1 1 19625
0 19627 7 1 2 26672 19626
0 19628 5 1 1 19627
0 19629 7 1 2 21956 37243
0 19630 5 1 1 19629
0 19631 7 1 2 19617 19630
0 19632 5 1 1 19631
0 19633 7 1 2 22238 19632
0 19634 5 1 1 19633
0 19635 7 1 2 32995 35796
0 19636 5 1 1 19635
0 19637 7 1 2 19636 37064
0 19638 5 1 1 19637
0 19639 7 1 2 30583 31622
0 19640 7 1 2 19638 19639
0 19641 5 1 1 19640
0 19642 7 1 2 19634 19641
0 19643 5 1 1 19642
0 19644 7 1 2 34943 19643
0 19645 5 1 1 19644
0 19646 7 1 2 30584 35893
0 19647 7 1 2 37237 19646
0 19648 7 1 2 37060 19647
0 19649 5 1 1 19648
0 19650 7 1 2 19645 19649
0 19651 5 1 1 19650
0 19652 7 1 2 26559 33124
0 19653 7 1 2 19651 19652
0 19654 5 1 1 19653
0 19655 7 1 2 25633 19654
0 19656 7 1 2 19628 19655
0 19657 5 1 1 19656
0 19658 7 1 2 30985 33777
0 19659 5 1 1 19658
0 19660 7 1 2 22685 32659
0 19661 5 1 1 19660
0 19662 7 1 2 19659 19661
0 19663 5 2 1 19662
0 19664 7 1 2 24129 37246
0 19665 5 1 1 19664
0 19666 7 1 2 32520 32660
0 19667 5 1 1 19666
0 19668 7 1 2 19665 19667
0 19669 5 2 1 19668
0 19670 7 1 2 30758 37248
0 19671 5 1 1 19670
0 19672 7 1 2 30699 32537
0 19673 5 1 1 19672
0 19674 7 1 2 19671 19673
0 19675 5 1 1 19674
0 19676 7 1 2 27739 19675
0 19677 5 1 1 19676
0 19678 7 1 2 36244 37235
0 19679 5 1 1 19678
0 19680 7 1 2 19677 19679
0 19681 5 1 1 19680
0 19682 7 1 2 26579 19681
0 19683 5 1 1 19682
0 19684 7 1 2 28439 34917
0 19685 7 1 2 32159 19684
0 19686 7 1 2 30439 31556
0 19687 7 1 2 19685 19686
0 19688 5 1 1 19687
0 19689 7 1 2 19683 19688
0 19690 5 1 1 19689
0 19691 7 1 2 36512 19690
0 19692 5 1 1 19691
0 19693 7 1 2 26025 36245
0 19694 5 1 1 19693
0 19695 7 1 2 30327 19694
0 19696 5 2 1 19695
0 19697 7 1 2 23475 36538
0 19698 5 1 1 19697
0 19699 7 2 2 25429 36672
0 19700 5 1 1 37252
0 19701 7 1 2 19698 19700
0 19702 5 2 1 19701
0 19703 7 1 2 37250 37254
0 19704 5 1 1 19703
0 19705 7 1 2 23476 26673
0 19706 7 1 2 36003 19705
0 19707 7 1 2 36246 19706
0 19708 5 1 1 19707
0 19709 7 1 2 19704 19708
0 19710 5 1 1 19709
0 19711 7 1 2 33125 19710
0 19712 5 1 1 19711
0 19713 7 1 2 19692 19712
0 19714 5 1 1 19713
0 19715 7 1 2 25533 19714
0 19716 5 1 1 19715
0 19717 7 1 2 22572 22718
0 19718 7 1 2 28440 19717
0 19719 7 1 2 31349 35871
0 19720 7 2 2 19718 19719
0 19721 7 1 2 28564 30323
0 19722 7 1 2 33815 19721
0 19723 7 1 2 37256 19722
0 19724 5 1 1 19723
0 19725 7 1 2 19716 19724
0 19726 5 1 1 19725
0 19727 7 1 2 22881 19726
0 19728 5 1 1 19727
0 19729 7 2 2 26456 30253
0 19730 7 1 2 36523 35413
0 19731 7 1 2 31361 19730
0 19732 7 1 2 37258 19731
0 19733 5 1 1 19732
0 19734 7 1 2 19728 19733
0 19735 5 1 1 19734
0 19736 7 1 2 35025 19735
0 19737 5 1 1 19736
0 19738 7 2 2 25358 32887
0 19739 7 1 2 26215 29394
0 19740 7 1 2 36673 19739
0 19741 7 1 2 37260 19740
0 19742 5 1 1 19741
0 19743 7 1 2 28770 36747
0 19744 7 1 2 32599 19743
0 19745 7 1 2 36117 35969
0 19746 7 1 2 19744 19745
0 19747 5 1 1 19746
0 19748 7 1 2 19742 19747
0 19749 5 1 1 19748
0 19750 7 1 2 24634 19749
0 19751 5 1 1 19750
0 19752 7 1 2 9931 16819
0 19753 5 1 1 19752
0 19754 7 1 2 22155 31541
0 19755 7 1 2 28733 19754
0 19756 7 1 2 31359 19755
0 19757 7 1 2 19753 19756
0 19758 5 1 1 19757
0 19759 7 1 2 19751 19758
0 19760 5 1 1 19759
0 19761 7 1 2 23238 19760
0 19762 5 1 1 19761
0 19763 7 1 2 29938 36539
0 19764 5 1 1 19763
0 19765 7 1 2 27940 33233
0 19766 5 1 1 19765
0 19767 7 1 2 36534 19766
0 19768 5 1 1 19767
0 19769 7 1 2 29577 19768
0 19770 5 1 1 19769
0 19771 7 1 2 19764 19770
0 19772 5 1 1 19771
0 19773 7 1 2 23390 19772
0 19774 5 1 1 19773
0 19775 7 2 2 25359 29578
0 19776 7 1 2 28514 36259
0 19777 5 1 1 19776
0 19778 7 1 2 26682 6789
0 19779 5 1 1 19778
0 19780 7 1 2 24252 15501
0 19781 7 1 2 19779 19780
0 19782 5 1 1 19781
0 19783 7 1 2 19777 19782
0 19784 5 1 1 19783
0 19785 7 1 2 37262 19784
0 19786 5 1 1 19785
0 19787 7 1 2 19774 19786
0 19788 5 1 1 19787
0 19789 7 1 2 23477 19788
0 19790 5 1 1 19789
0 19791 7 1 2 29130 36331
0 19792 7 1 2 34278 36233
0 19793 7 1 2 19791 19792
0 19794 5 1 1 19793
0 19795 7 1 2 19790 19794
0 19796 5 1 1 19795
0 19797 7 1 2 22686 32254
0 19798 7 1 2 31516 19797
0 19799 7 1 2 19796 19798
0 19800 5 1 1 19799
0 19801 7 1 2 19762 19800
0 19802 5 1 1 19801
0 19803 7 1 2 22882 19802
0 19804 5 1 1 19803
0 19805 7 1 2 29374 35237
0 19806 7 1 2 31901 35006
0 19807 7 1 2 19805 19806
0 19808 7 1 2 37257 19807
0 19809 5 1 1 19808
0 19810 7 1 2 19804 19809
0 19811 5 1 1 19810
0 19812 7 1 2 23584 19811
0 19813 5 1 1 19812
0 19814 7 1 2 24825 28628
0 19815 7 1 2 29771 19814
0 19816 7 2 2 27040 29306
0 19817 7 1 2 37264 35256
0 19818 7 1 2 19815 19817
0 19819 5 1 1 19818
0 19820 7 1 2 35907 35612
0 19821 5 1 1 19820
0 19822 7 1 2 21957 19821
0 19823 5 1 1 19822
0 19824 7 2 2 22573 35903
0 19825 5 1 1 37266
0 19826 7 1 2 19823 19825
0 19827 5 1 1 19826
0 19828 7 2 2 23478 25819
0 19829 7 1 2 23769 37233
0 19830 7 1 2 37268 19829
0 19831 7 1 2 19827 19830
0 19832 5 1 1 19831
0 19833 7 1 2 19819 19832
0 19834 5 1 1 19833
0 19835 7 1 2 22094 19834
0 19836 5 1 1 19835
0 19837 7 1 2 26580 28070
0 19838 7 1 2 32555 19837
0 19839 7 1 2 32179 19838
0 19840 7 1 2 37247 19839
0 19841 5 1 1 19840
0 19842 7 1 2 19836 19841
0 19843 5 1 1 19842
0 19844 7 1 2 36513 19843
0 19845 5 1 1 19844
0 19846 7 1 2 27826 28589
0 19847 7 1 2 31667 19846
0 19848 7 1 2 31778 19847
0 19849 7 1 2 37255 19848
0 19850 5 1 1 19849
0 19851 7 1 2 25290 19850
0 19852 7 1 2 19845 19851
0 19853 7 1 2 19813 19852
0 19854 5 1 1 19853
0 19855 7 1 2 28348 27788
0 19856 7 2 2 27113 19855
0 19857 7 1 2 25104 37270
0 19858 5 1 1 19857
0 19859 7 1 2 37138 35971
0 19860 5 1 1 19859
0 19861 7 1 2 19858 19860
0 19862 5 1 1 19861
0 19863 7 1 2 27238 19862
0 19864 5 1 1 19863
0 19865 7 1 2 28920 30774
0 19866 7 1 2 36518 19865
0 19867 7 1 2 28476 34575
0 19868 7 1 2 19866 19867
0 19869 5 1 1 19868
0 19870 7 1 2 19864 19869
0 19871 5 1 1 19870
0 19872 7 1 2 29522 19871
0 19873 5 1 1 19872
0 19874 7 1 2 22156 31039
0 19875 5 1 1 19874
0 19876 7 1 2 26271 27081
0 19877 5 1 1 19876
0 19878 7 1 2 19875 19877
0 19879 5 1 1 19878
0 19880 7 1 2 29579 19879
0 19881 5 1 1 19880
0 19882 7 1 2 3157 19881
0 19883 5 1 1 19882
0 19884 7 1 2 23144 19883
0 19885 5 1 1 19884
0 19886 7 1 2 28057 29992
0 19887 5 1 1 19886
0 19888 7 1 2 19885 19887
0 19889 5 1 1 19888
0 19890 7 1 2 28349 31517
0 19891 7 1 2 19889 19890
0 19892 5 1 1 19891
0 19893 7 1 2 19873 19892
0 19894 5 1 1 19893
0 19895 7 1 2 22095 19894
0 19896 5 1 1 19895
0 19897 7 1 2 37261 35671
0 19898 7 1 2 32152 19897
0 19899 7 1 2 36967 19898
0 19900 5 1 1 19899
0 19901 7 1 2 27239 27847
0 19902 5 1 1 19901
0 19903 7 1 2 27740 30380
0 19904 5 1 1 19903
0 19905 7 1 2 19902 19904
0 19906 5 1 1 19905
0 19907 7 1 2 35081 19906
0 19908 5 1 1 19907
0 19909 7 1 2 30394 36380
0 19910 7 1 2 31977 19909
0 19911 5 1 1 19910
0 19912 7 1 2 19908 19911
0 19913 5 1 1 19912
0 19914 7 1 2 22096 27096
0 19915 7 1 2 19913 19914
0 19916 5 1 1 19915
0 19917 7 1 2 19900 19916
0 19918 5 1 1 19917
0 19919 7 1 2 29616 19918
0 19920 5 1 1 19919
0 19921 7 1 2 31040 32100
0 19922 7 1 2 36524 19921
0 19923 7 1 2 36741 19922
0 19924 5 1 1 19923
0 19925 7 1 2 28350 27097
0 19926 5 1 1 19925
0 19927 7 1 2 27946 34284
0 19928 5 1 1 19927
0 19929 7 1 2 19926 19928
0 19930 5 1 1 19929
0 19931 7 1 2 30620 19930
0 19932 5 1 1 19931
0 19933 7 1 2 30111 37075
0 19934 5 1 1 19933
0 19935 7 1 2 19932 19934
0 19936 5 1 1 19935
0 19937 7 1 2 28734 31776
0 19938 7 1 2 19936 19937
0 19939 5 1 1 19938
0 19940 7 1 2 19924 19939
0 19941 5 1 1 19940
0 19942 7 1 2 22574 19941
0 19943 5 1 1 19942
0 19944 7 1 2 19920 19943
0 19945 7 1 2 19896 19944
0 19946 5 1 1 19945
0 19947 7 1 2 29223 19946
0 19948 5 1 1 19947
0 19949 7 1 2 32463 7077
0 19950 5 1 1 19949
0 19951 7 1 2 29523 19950
0 19952 5 1 1 19951
0 19953 7 1 2 31049 35611
0 19954 5 1 1 19953
0 19955 7 1 2 19952 19954
0 19956 5 1 1 19955
0 19957 7 1 2 22097 19956
0 19958 5 1 1 19957
0 19959 7 1 2 30081 31200
0 19960 7 1 2 33666 19959
0 19961 5 1 1 19960
0 19962 7 1 2 19958 19961
0 19963 5 1 1 19962
0 19964 7 1 2 31672 19963
0 19965 5 1 1 19964
0 19966 7 1 2 26581 36263
0 19967 5 1 1 19966
0 19968 7 1 2 22719 23239
0 19969 5 1 1 19968
0 19970 7 1 2 33773 19969
0 19971 5 1 1 19970
0 19972 7 1 2 22157 26865
0 19973 7 1 2 19971 19972
0 19974 5 1 1 19973
0 19975 7 1 2 19967 19974
0 19976 5 1 1 19975
0 19977 7 1 2 31706 35904
0 19978 7 1 2 19976 19977
0 19979 5 1 1 19978
0 19980 7 1 2 19965 19979
0 19981 5 1 1 19980
0 19982 7 1 2 27789 19981
0 19983 5 1 1 19982
0 19984 7 1 2 24546 27041
0 19985 7 1 2 25774 32600
0 19986 7 1 2 19984 19985
0 19987 7 1 2 26586 33770
0 19988 7 1 2 19986 19987
0 19989 5 1 1 19988
0 19990 7 1 2 19983 19989
0 19991 5 1 1 19990
0 19992 7 1 2 28546 19991
0 19993 5 1 1 19992
0 19994 7 1 2 36247 37271
0 19995 5 1 1 19994
0 19996 7 1 2 26951 29158
0 19997 7 1 2 29271 19996
0 19998 7 1 2 24726 27091
0 19999 7 1 2 29176 19998
0 20000 7 1 2 19997 19999
0 20001 5 1 1 20000
0 20002 7 1 2 19995 20001
0 20003 5 1 1 20002
0 20004 7 1 2 34274 20003
0 20005 5 1 1 20004
0 20006 7 1 2 23328 20005
0 20007 7 1 2 19993 20006
0 20008 7 1 2 19948 20007
0 20009 5 1 1 20008
0 20010 7 1 2 33415 20009
0 20011 7 1 2 19854 20010
0 20012 5 1 1 20011
0 20013 7 1 2 28711 31350
0 20014 7 1 2 30408 20013
0 20015 7 1 2 36525 34464
0 20016 7 1 2 20014 20015
0 20017 7 1 2 37259 20016
0 20018 5 1 1 20017
0 20019 7 1 2 23694 20018
0 20020 7 1 2 20012 20019
0 20021 7 1 2 19737 20020
0 20022 5 1 1 20021
0 20023 7 1 2 19657 20022
0 20024 5 1 1 20023
0 20025 7 1 2 37263 35258
0 20026 7 1 2 37269 20025
0 20027 7 1 2 32019 20026
0 20028 5 1 1 20027
0 20029 7 1 2 26582 27612
0 20030 7 1 2 37249 20029
0 20031 5 1 1 20030
0 20032 7 1 2 20028 20031
0 20033 5 1 1 20032
0 20034 7 1 2 33388 20033
0 20035 5 1 1 20034
0 20036 7 2 2 22276 22575
0 20037 7 1 2 31351 36300
0 20038 7 1 2 37272 20037
0 20039 7 1 2 28509 20038
0 20040 7 1 2 31993 20039
0 20041 5 1 1 20040
0 20042 7 1 2 20035 20041
0 20043 5 1 1 20042
0 20044 7 1 2 25291 20043
0 20045 5 1 1 20044
0 20046 7 1 2 36027 35665
0 20047 7 1 2 33535 20046
0 20048 5 1 1 20047
0 20049 7 1 2 20045 20048
0 20050 5 1 1 20049
0 20051 7 1 2 26560 20050
0 20052 5 1 1 20051
0 20053 7 1 2 27037 26674
0 20054 7 1 2 34643 20053
0 20055 7 1 2 31147 20054
0 20056 7 1 2 33536 20055
0 20057 5 1 1 20056
0 20058 7 1 2 20052 20057
0 20059 5 1 1 20058
0 20060 7 1 2 25534 20059
0 20061 5 1 1 20060
0 20062 7 1 2 22098 26561
0 20063 7 2 2 27412 20062
0 20064 7 1 2 29224 31143
0 20065 7 1 2 33416 20064
0 20066 7 1 2 37274 20065
0 20067 7 1 2 30982 20066
0 20068 5 1 1 20067
0 20069 7 1 2 20061 20068
0 20070 5 1 1 20069
0 20071 7 1 2 24987 20070
0 20072 5 1 1 20071
0 20073 7 1 2 23329 29064
0 20074 7 1 2 29195 20073
0 20075 7 1 2 36688 35683
0 20076 7 1 2 20074 20075
0 20077 7 1 2 36302 20076
0 20078 5 1 1 20077
0 20079 7 1 2 26675 33663
0 20080 7 1 2 35763 20079
0 20081 7 1 2 37251 20080
0 20082 5 1 1 20081
0 20083 7 1 2 20078 20082
0 20084 5 1 1 20083
0 20085 7 1 2 22099 20084
0 20086 5 1 1 20085
0 20087 7 1 2 20072 20086
0 20088 5 1 1 20087
0 20089 7 1 2 28547 20088
0 20090 5 1 1 20089
0 20091 7 2 2 29524 31391
0 20092 5 1 1 37276
0 20093 7 1 2 29617 32023
0 20094 5 1 1 20093
0 20095 7 1 2 20092 20094
0 20096 5 1 1 20095
0 20097 7 1 2 23330 20096
0 20098 5 1 1 20097
0 20099 7 1 2 23145 30216
0 20100 5 1 1 20099
0 20101 7 1 2 20098 20100
0 20102 5 1 1 20101
0 20103 7 1 2 22100 20102
0 20104 5 1 1 20103
0 20105 7 1 2 28241 30226
0 20106 7 1 2 35654 20105
0 20107 5 1 1 20106
0 20108 7 1 2 20104 20107
0 20109 5 1 1 20108
0 20110 7 1 2 35396 34541
0 20111 5 1 1 20110
0 20112 7 1 2 28468 33389
0 20113 5 1 1 20112
0 20114 7 1 2 20111 20113
0 20115 5 1 1 20114
0 20116 7 1 2 23585 30019
0 20117 7 1 2 20115 20116
0 20118 7 1 2 20109 20117
0 20119 5 1 1 20118
0 20120 7 2 2 22883 26779
0 20121 7 1 2 37168 37278
0 20122 5 1 1 20121
0 20123 7 1 2 28590 35089
0 20124 7 1 2 26902 20123
0 20125 5 1 1 20124
0 20126 7 1 2 20122 20125
0 20127 5 1 1 20126
0 20128 7 1 2 24547 20127
0 20129 5 1 1 20128
0 20130 7 1 2 29618 37279
0 20131 7 1 2 37222 20130
0 20132 5 1 1 20131
0 20133 7 1 2 20129 20132
0 20134 5 1 1 20133
0 20135 7 1 2 23146 20134
0 20136 5 1 1 20135
0 20137 7 1 2 30753 31639
0 20138 7 1 2 37277 20137
0 20139 5 1 1 20138
0 20140 7 1 2 20136 20139
0 20141 5 1 1 20140
0 20142 7 1 2 22101 20141
0 20143 5 1 1 20142
0 20144 7 2 2 27073 37219
0 20145 7 1 2 24988 29931
0 20146 7 1 2 33778 20145
0 20147 7 1 2 37280 20146
0 20148 5 1 1 20147
0 20149 7 1 2 31691 32190
0 20150 7 1 2 37223 20149
0 20151 5 1 1 20150
0 20152 7 1 2 20148 20151
0 20153 5 1 1 20152
0 20154 7 1 2 24004 20153
0 20155 5 1 1 20154
0 20156 7 1 2 24989 32260
0 20157 7 1 2 32661 20156
0 20158 7 1 2 37281 20157
0 20159 5 1 1 20158
0 20160 7 1 2 20155 20159
0 20161 7 1 2 20143 20160
0 20162 5 1 1 20161
0 20163 7 1 2 34192 20162
0 20164 5 1 1 20163
0 20165 7 1 2 20119 20164
0 20166 5 1 1 20165
0 20167 7 1 2 27598 20166
0 20168 5 1 1 20167
0 20169 7 1 2 28351 33570
0 20170 5 1 1 20169
0 20171 7 1 2 26809 28357
0 20172 7 2 2 33718 20171
0 20173 5 1 1 37282
0 20174 7 1 2 20170 20173
0 20175 5 1 1 20174
0 20176 7 1 2 24990 20175
0 20177 5 1 1 20176
0 20178 7 2 2 28469 33719
0 20179 7 1 2 32492 37284
0 20180 5 1 1 20179
0 20181 7 1 2 20177 20180
0 20182 5 1 1 20181
0 20183 7 1 2 29099 20182
0 20184 5 1 1 20183
0 20185 7 1 2 28766 36071
0 20186 5 1 1 20185
0 20187 7 1 2 20184 20186
0 20188 5 1 1 20187
0 20189 7 1 2 23240 20188
0 20190 5 1 1 20189
0 20191 7 1 2 33653 36768
0 20192 7 1 2 35450 20191
0 20193 7 1 2 36990 20192
0 20194 5 1 1 20193
0 20195 7 1 2 20190 20194
0 20196 5 1 1 20195
0 20197 7 1 2 21958 20196
0 20198 5 1 1 20197
0 20199 7 1 2 36120 35919
0 20200 7 1 2 36297 20199
0 20201 5 1 1 20200
0 20202 7 1 2 20198 20201
0 20203 5 1 1 20202
0 20204 7 1 2 27413 31406
0 20205 7 1 2 20203 20204
0 20206 5 1 1 20205
0 20207 7 1 2 20168 20206
0 20208 5 1 1 20207
0 20209 7 1 2 23391 20208
0 20210 5 1 1 20209
0 20211 7 1 2 26918 35026
0 20212 5 1 1 20211
0 20213 7 1 2 28144 33417
0 20214 5 1 1 20213
0 20215 7 1 2 20212 20214
0 20216 5 1 1 20215
0 20217 7 1 2 30637 20216
0 20218 5 1 1 20217
0 20219 7 1 2 28145 36123
0 20220 5 1 1 20219
0 20221 7 1 2 28621 34423
0 20222 5 1 1 20221
0 20223 7 1 2 28712 33930
0 20224 5 1 1 20223
0 20225 7 1 2 20222 20224
0 20226 5 1 1 20225
0 20227 7 1 2 26919 20226
0 20228 5 1 1 20227
0 20229 7 1 2 20220 20228
0 20230 7 1 2 20218 20229
0 20231 5 1 1 20230
0 20232 7 1 2 26480 20231
0 20233 5 1 1 20232
0 20234 7 1 2 30867 37285
0 20235 5 1 1 20234
0 20236 7 1 2 20233 20235
0 20237 5 1 1 20236
0 20238 7 1 2 26457 31362
0 20239 7 1 2 20237 20238
0 20240 5 1 1 20239
0 20241 7 1 2 20210 20240
0 20242 5 1 1 20241
0 20243 7 1 2 26676 20242
0 20244 5 1 1 20243
0 20245 7 1 2 28352 30667
0 20246 7 2 2 30360 20245
0 20247 7 1 2 30587 37286
0 20248 5 1 1 20247
0 20249 7 1 2 31148 32183
0 20250 5 1 1 20249
0 20251 7 1 2 26930 32375
0 20252 7 1 2 36129 20251
0 20253 5 1 1 20252
0 20254 7 1 2 20250 20253
0 20255 5 1 1 20254
0 20256 7 1 2 35082 20255
0 20257 5 1 1 20256
0 20258 7 1 2 25765 29580
0 20259 7 1 2 36205 20258
0 20260 7 1 2 30361 20259
0 20261 5 1 1 20260
0 20262 7 1 2 20257 20261
0 20263 5 1 1 20262
0 20264 7 1 2 22344 20263
0 20265 5 1 1 20264
0 20266 7 1 2 20248 20265
0 20267 5 1 1 20266
0 20268 7 1 2 33332 20267
0 20269 5 1 1 20268
0 20270 7 1 2 37287 33559
0 20271 5 1 1 20270
0 20272 7 1 2 20269 20271
0 20273 5 1 1 20272
0 20274 7 1 2 37275 20273
0 20275 5 1 1 20274
0 20276 7 1 2 20244 20275
0 20277 7 1 2 20090 20276
0 20278 5 1 1 20277
0 20279 7 1 2 25956 20278
0 20280 5 1 1 20279
0 20281 7 1 2 20024 20280
0 20282 5 1 1 20281
0 20283 7 1 2 27199 20282
0 20284 5 1 1 20283
0 20285 7 1 2 31013 35559
0 20286 5 1 1 20285
0 20287 7 9 2 31484 33054
0 20288 7 1 2 24886 34173
0 20289 7 1 2 37288 20288
0 20290 5 1 1 20289
0 20291 7 1 2 20286 20290
0 20292 5 1 1 20291
0 20293 7 1 2 33977 20292
0 20294 5 1 1 20293
0 20295 7 3 2 23695 29100
0 20296 7 1 2 24005 22952
0 20297 7 1 2 36697 20296
0 20298 7 1 2 37297 20297
0 20299 5 1 1 20298
0 20300 7 1 2 20294 20299
0 20301 5 1 1 20300
0 20302 7 1 2 24354 20301
0 20303 5 1 1 20302
0 20304 7 1 2 37298 35348
0 20305 7 1 2 36788 20304
0 20306 5 1 1 20305
0 20307 7 1 2 20303 20306
0 20308 5 1 1 20307
0 20309 7 1 2 24298 20308
0 20310 5 1 1 20309
0 20311 7 1 2 31014 34130
0 20312 7 1 2 34001 20311
0 20313 5 1 1 20312
0 20314 7 1 2 20310 20313
0 20315 5 1 1 20314
0 20316 7 1 2 36573 20315
0 20317 5 1 1 20316
0 20318 7 1 2 32096 33868
0 20319 5 1 1 20318
0 20320 7 1 2 31974 34065
0 20321 5 1 1 20320
0 20322 7 1 2 20319 20321
0 20323 5 1 1 20322
0 20324 7 1 2 26677 31783
0 20325 7 1 2 37299 20324
0 20326 7 1 2 20323 20325
0 20327 5 1 1 20326
0 20328 7 1 2 20317 20327
0 20329 5 1 1 20328
0 20330 7 1 2 24423 20329
0 20331 5 1 1 20330
0 20332 7 1 2 31015 34094
0 20333 7 1 2 36705 20332
0 20334 5 1 1 20333
0 20335 7 1 2 20331 20334
0 20336 5 1 1 20335
0 20337 7 1 2 32738 20336
0 20338 5 1 1 20337
0 20339 7 1 2 25957 33093
0 20340 5 1 1 20339
0 20341 7 1 2 32614 20340
0 20342 5 1 1 20341
0 20343 7 1 2 37289 20342
0 20344 5 1 1 20343
0 20345 7 1 2 32703 36728
0 20346 5 1 1 20345
0 20347 7 1 2 29120 33118
0 20348 5 1 1 20347
0 20349 7 1 2 24130 20348
0 20350 5 1 1 20349
0 20351 7 1 2 36045 20350
0 20352 5 1 1 20351
0 20353 7 1 2 32622 20352
0 20354 5 1 1 20353
0 20355 7 1 2 37067 32710
0 20356 5 1 1 20355
0 20357 7 1 2 20354 20356
0 20358 5 1 1 20357
0 20359 7 1 2 21959 20358
0 20360 5 1 1 20359
0 20361 7 1 2 20346 20360
0 20362 7 1 2 20344 20361
0 20363 5 1 1 20362
0 20364 7 1 2 36800 20363
0 20365 5 1 1 20364
0 20366 7 1 2 24131 29132
0 20367 5 2 1 20366
0 20368 7 1 2 33141 37300
0 20369 5 1 1 20368
0 20370 7 1 2 21845 20369
0 20371 5 1 1 20370
0 20372 7 2 2 28994 29666
0 20373 5 1 1 37302
0 20374 7 1 2 20373 36060
0 20375 5 1 1 20374
0 20376 7 1 2 22102 20375
0 20377 5 1 1 20376
0 20378 7 2 2 20371 20377
0 20379 5 1 1 37304
0 20380 7 1 2 28995 35708
0 20381 5 1 1 20380
0 20382 7 1 2 37301 20381
0 20383 5 1 1 20382
0 20384 7 1 2 24991 20383
0 20385 5 1 1 20384
0 20386 7 4 2 24132 29101
0 20387 7 1 2 21960 37306
0 20388 5 1 1 20387
0 20389 7 1 2 20385 20388
0 20390 5 4 1 20389
0 20391 7 1 2 27697 37310
0 20392 5 1 1 20391
0 20393 7 1 2 37305 20392
0 20394 5 1 1 20393
0 20395 7 1 2 36586 35332
0 20396 7 1 2 33042 20395
0 20397 7 1 2 20394 20396
0 20398 5 1 1 20397
0 20399 7 1 2 25958 36797
0 20400 5 1 1 20399
0 20401 7 1 2 16290 20400
0 20402 5 1 1 20401
0 20403 7 1 2 23696 33978
0 20404 7 1 2 20379 20403
0 20405 7 1 2 20402 20404
0 20406 5 1 1 20405
0 20407 7 1 2 23697 36804
0 20408 7 1 2 37311 20407
0 20409 5 1 1 20408
0 20410 7 1 2 20406 20409
0 20411 7 1 2 20398 20410
0 20412 7 1 2 20365 20411
0 20413 5 1 1 20412
0 20414 7 1 2 23586 20413
0 20415 5 1 1 20414
0 20416 7 1 2 33448 34259
0 20417 7 1 2 33997 20416
0 20418 7 1 2 36685 37290
0 20419 7 1 2 20417 20418
0 20420 5 1 1 20419
0 20421 7 1 2 36046 32718
0 20422 5 1 1 20421
0 20423 7 1 2 21961 20422
0 20424 5 1 1 20423
0 20425 7 1 2 37291 33807
0 20426 5 1 1 20425
0 20427 7 1 2 1484 36061
0 20428 5 1 1 20427
0 20429 7 1 2 22103 20428
0 20430 5 2 1 20429
0 20431 7 1 2 20426 37314
0 20432 7 1 2 20424 20431
0 20433 5 1 1 20432
0 20434 7 1 2 30283 36806
0 20435 7 1 2 20433 20434
0 20436 5 1 1 20435
0 20437 7 1 2 20420 20436
0 20438 5 1 1 20437
0 20439 7 1 2 25535 20438
0 20440 5 1 1 20439
0 20441 7 1 2 20415 20440
0 20442 7 1 2 20338 20441
0 20443 5 1 1 20442
0 20444 7 1 2 25684 20443
0 20445 5 1 1 20444
0 20446 7 3 2 22239 22720
0 20447 5 1 1 37316
0 20448 7 1 2 30482 33979
0 20449 5 1 1 20448
0 20450 7 2 2 28629 34111
0 20451 5 1 1 37319
0 20452 7 1 2 31850 37320
0 20453 5 1 1 20452
0 20454 7 1 2 20449 20453
0 20455 5 1 1 20454
0 20456 7 1 2 21962 20455
0 20457 5 1 1 20456
0 20458 7 1 2 28201 35458
0 20459 5 1 1 20458
0 20460 7 1 2 24133 34592
0 20461 5 1 1 20460
0 20462 7 1 2 28203 33980
0 20463 5 1 1 20462
0 20464 7 1 2 20463 15581
0 20465 7 1 2 20461 20464
0 20466 7 1 2 20459 20465
0 20467 5 1 1 20466
0 20468 7 1 2 25105 20467
0 20469 5 1 1 20468
0 20470 7 1 2 20451 20469
0 20471 5 1 1 20470
0 20472 7 1 2 22158 20471
0 20473 5 1 1 20472
0 20474 7 1 2 20457 20473
0 20475 5 1 1 20474
0 20476 7 1 2 22277 20475
0 20477 5 1 1 20476
0 20478 7 2 2 25106 32677
0 20479 5 1 1 37321
0 20480 7 1 2 20479 32317
0 20481 5 4 1 20480
0 20482 7 2 2 22159 37323
0 20483 7 1 2 35499 37327
0 20484 5 1 1 20483
0 20485 7 1 2 20477 20484
0 20486 5 1 1 20485
0 20487 7 1 2 23587 20486
0 20488 5 1 1 20487
0 20489 7 1 2 37328 36530
0 20490 5 1 1 20489
0 20491 7 1 2 20488 20490
0 20492 5 1 1 20491
0 20493 7 1 2 37317 20492
0 20494 5 1 1 20493
0 20495 7 1 2 34593 34125
0 20496 5 1 1 20495
0 20497 7 1 2 34132 20496
0 20498 5 1 1 20497
0 20499 7 1 2 36574 20498
0 20500 7 1 2 37324 20499
0 20501 5 1 1 20500
0 20502 7 1 2 25869 20501
0 20503 7 1 2 20494 20502
0 20504 5 1 1 20503
0 20505 7 1 2 33333 36323
0 20506 5 1 1 20505
0 20507 7 1 2 36427 35505
0 20508 5 1 1 20507
0 20509 7 1 2 20506 20508
0 20510 5 1 1 20509
0 20511 7 1 2 25536 20510
0 20512 7 1 2 37325 20511
0 20513 5 1 1 20512
0 20514 7 1 2 25873 20513
0 20515 5 1 1 20514
0 20516 7 1 2 22576 26100
0 20517 7 1 2 20515 20516
0 20518 7 1 2 20504 20517
0 20519 5 1 1 20518
0 20520 7 2 2 30004 30578
0 20521 7 1 2 21963 37329
0 20522 5 1 1 20521
0 20523 7 1 2 22104 29610
0 20524 5 1 1 20523
0 20525 7 1 2 20522 20524
0 20526 5 3 1 20525
0 20527 7 1 2 23147 37331
0 20528 5 1 1 20527
0 20529 7 1 2 21964 34665
0 20530 5 2 1 20529
0 20531 7 1 2 22105 29468
0 20532 5 1 1 20531
0 20533 7 2 2 37334 20532
0 20534 7 1 2 20528 37336
0 20535 5 1 1 20534
0 20536 7 1 2 30739 37110
0 20537 5 1 1 20536
0 20538 7 1 2 36692 36622
0 20539 5 1 1 20538
0 20540 7 1 2 20537 20539
0 20541 5 1 1 20540
0 20542 7 1 2 25736 20541
0 20543 5 1 1 20542
0 20544 7 1 2 33571 36498
0 20545 5 1 1 20544
0 20546 7 1 2 20543 20545
0 20547 5 1 1 20546
0 20548 7 1 2 20535 20547
0 20549 5 1 1 20548
0 20550 7 1 2 36324 34666
0 20551 5 1 1 20550
0 20552 7 2 2 24548 35858
0 20553 7 1 2 37199 37338
0 20554 5 1 1 20553
0 20555 7 1 2 36494 20554
0 20556 5 1 1 20555
0 20557 7 1 2 27200 20556
0 20558 5 1 1 20557
0 20559 7 1 2 24992 36488
0 20560 5 1 1 20559
0 20561 7 1 2 37231 20560
0 20562 7 1 2 20558 20561
0 20563 5 1 1 20562
0 20564 7 1 2 23148 20563
0 20565 5 1 1 20564
0 20566 7 1 2 20551 20565
0 20567 5 1 1 20566
0 20568 7 1 2 21965 20567
0 20569 5 1 1 20568
0 20570 7 1 2 5853 35640
0 20571 5 1 1 20570
0 20572 7 1 2 36489 20571
0 20573 5 1 1 20572
0 20574 7 1 2 29125 36325
0 20575 5 1 1 20574
0 20576 7 1 2 25430 36260
0 20577 7 1 2 37339 20576
0 20578 5 1 1 20577
0 20579 7 1 2 20575 20578
0 20580 5 1 1 20579
0 20581 7 1 2 22106 20580
0 20582 5 1 1 20581
0 20583 7 1 2 20573 20582
0 20584 7 1 2 20569 20583
0 20585 5 1 1 20584
0 20586 7 1 2 20585 34950
0 20587 5 1 1 20586
0 20588 7 1 2 20549 20587
0 20589 7 1 2 20519 20588
0 20590 5 1 1 20589
0 20591 7 1 2 25634 20590
0 20592 5 1 1 20591
0 20593 7 1 2 26230 20592
0 20594 5 1 1 20593
0 20595 7 1 2 27336 29843
0 20596 5 2 1 20595
0 20597 7 1 2 26183 31352
0 20598 5 1 1 20597
0 20599 7 1 2 22577 20598
0 20600 5 1 1 20599
0 20601 7 1 2 37340 20600
0 20602 5 1 1 20601
0 20603 7 1 2 25107 20602
0 20604 5 1 1 20603
0 20605 7 3 2 32539 20604
0 20606 5 3 1 37342
0 20607 7 1 2 32546 37343
0 20608 5 3 1 20607
0 20609 7 1 2 22160 37348
0 20610 5 1 1 20609
0 20611 7 1 2 29440 31741
0 20612 5 2 1 20611
0 20613 7 1 2 20610 37351
0 20614 5 2 1 20613
0 20615 7 2 2 28652 36782
0 20616 7 1 2 37353 37355
0 20617 5 1 1 20616
0 20618 7 1 2 23149 37330
0 20619 5 1 1 20618
0 20620 7 1 2 5814 20619
0 20621 5 1 1 20620
0 20622 7 1 2 21966 20621
0 20623 5 2 1 20622
0 20624 7 1 2 22107 30463
0 20625 5 1 1 20624
0 20626 7 2 2 37357 20625
0 20627 7 1 2 22578 37322
0 20628 5 1 1 20627
0 20629 7 1 2 37359 20628
0 20630 5 5 1 20629
0 20631 7 1 2 28681 36686
0 20632 7 1 2 37361 20631
0 20633 5 1 1 20632
0 20634 7 1 2 20617 20633
0 20635 5 1 1 20634
0 20636 7 1 2 24826 20635
0 20637 5 1 1 20636
0 20638 7 1 2 22161 34685
0 20639 5 1 1 20638
0 20640 7 1 2 35638 20639
0 20641 5 2 1 20640
0 20642 7 1 2 29267 36783
0 20643 7 1 2 37366 20642
0 20644 5 1 1 20643
0 20645 7 1 2 20637 20644
0 20646 5 1 1 20645
0 20647 7 1 2 25431 20646
0 20648 5 1 1 20647
0 20649 7 1 2 22721 33458
0 20650 7 2 2 37354 20649
0 20651 5 1 1 37368
0 20652 7 1 2 28305 27875
0 20653 7 1 2 37369 20652
0 20654 5 1 1 20653
0 20655 7 1 2 20648 20654
0 20656 5 1 1 20655
0 20657 7 1 2 24767 20656
0 20658 5 1 1 20657
0 20659 7 1 2 31558 32195
0 20660 5 1 1 20659
0 20661 7 1 2 29418 33700
0 20662 5 1 1 20661
0 20663 7 1 2 20660 20662
0 20664 5 1 1 20663
0 20665 7 1 2 27473 20664
0 20666 5 1 1 20665
0 20667 7 1 2 23150 29346
0 20668 7 1 2 37267 20667
0 20669 5 1 1 20668
0 20670 7 1 2 20666 20669
0 20671 5 1 1 20670
0 20672 7 1 2 22108 20671
0 20673 5 1 1 20672
0 20674 7 1 2 28591 32552
0 20675 5 1 1 20674
0 20676 7 2 2 27201 36769
0 20677 7 1 2 30082 37370
0 20678 5 1 1 20677
0 20679 7 1 2 29230 35613
0 20680 5 1 1 20679
0 20681 7 1 2 3475 20680
0 20682 5 1 1 20681
0 20683 7 1 2 26946 35311
0 20684 5 1 1 20683
0 20685 7 1 2 29231 20684
0 20686 5 1 1 20685
0 20687 7 1 2 27538 20686
0 20688 5 1 1 20687
0 20689 7 1 2 27157 32180
0 20690 5 1 1 20689
0 20691 7 1 2 20688 20690
0 20692 7 1 2 20682 20691
0 20693 5 1 1 20692
0 20694 7 1 2 25108 20693
0 20695 5 1 1 20694
0 20696 7 1 2 20678 20695
0 20697 7 1 2 20675 20696
0 20698 5 1 1 20697
0 20699 7 1 2 22162 20698
0 20700 5 1 1 20699
0 20701 7 1 2 20673 20700
0 20702 5 1 1 20701
0 20703 7 1 2 22722 31634
0 20704 7 1 2 20702 20703
0 20705 5 1 1 20704
0 20706 7 1 2 34824 34686
0 20707 7 1 2 36959 20706
0 20708 5 1 1 20707
0 20709 7 1 2 20705 20708
0 20710 5 1 1 20709
0 20711 7 1 2 35778 20710
0 20712 5 1 1 20711
0 20713 7 1 2 22345 20712
0 20714 7 1 2 20658 20713
0 20715 5 1 1 20714
0 20716 7 1 2 37341 13446
0 20717 5 1 1 20716
0 20718 7 1 2 25109 20717
0 20719 5 1 1 20718
0 20720 7 1 2 32549 20719
0 20721 5 3 1 20720
0 20722 7 1 2 33981 37372
0 20723 5 1 1 20722
0 20724 7 1 2 34112 37307
0 20725 5 1 1 20724
0 20726 7 1 2 20723 20725
0 20727 5 1 1 20726
0 20728 7 1 2 22163 20727
0 20729 5 1 1 20728
0 20730 7 1 2 29544 33982
0 20731 7 1 2 29707 20730
0 20732 5 1 1 20731
0 20733 7 1 2 20729 20732
0 20734 5 1 1 20733
0 20735 7 1 2 37356 20734
0 20736 5 1 1 20735
0 20737 7 1 2 22579 37326
0 20738 5 1 1 20737
0 20739 7 1 2 37337 20738
0 20740 5 2 1 20739
0 20741 7 1 2 33983 37375
0 20742 5 1 1 20741
0 20743 7 1 2 33984 37332
0 20744 5 1 1 20743
0 20745 7 1 2 34113 32543
0 20746 5 1 1 20745
0 20747 7 1 2 20744 20746
0 20748 5 1 1 20747
0 20749 7 1 2 23151 20748
0 20750 5 1 1 20749
0 20751 7 1 2 34114 37345
0 20752 5 1 1 20751
0 20753 7 1 2 20750 20752
0 20754 7 1 2 20742 20753
0 20755 5 1 1 20754
0 20756 7 1 2 24177 20755
0 20757 5 1 1 20756
0 20758 7 2 2 26386 29681
0 20759 5 2 1 37377
0 20760 7 1 2 34115 37378
0 20761 5 1 1 20760
0 20762 7 1 2 20757 20761
0 20763 5 1 1 20762
0 20764 7 2 2 24664 34511
0 20765 7 1 2 28682 37381
0 20766 7 1 2 20763 20765
0 20767 5 1 1 20766
0 20768 7 1 2 20736 20767
0 20769 5 1 1 20768
0 20770 7 1 2 22884 20769
0 20771 5 1 1 20770
0 20772 7 1 2 28306 36468
0 20773 5 1 1 20772
0 20774 7 1 2 22278 26810
0 20775 5 1 1 20774
0 20776 7 1 2 24299 28307
0 20777 5 1 1 20776
0 20778 7 1 2 20775 20777
0 20779 5 2 1 20778
0 20780 7 1 2 22820 36575
0 20781 7 1 2 37383 20780
0 20782 5 2 1 20781
0 20783 7 1 2 20773 37385
0 20784 5 1 1 20783
0 20785 7 1 2 37308 20784
0 20786 5 1 1 20785
0 20787 7 1 2 22580 32303
0 20788 5 2 1 20787
0 20789 7 1 2 37360 37387
0 20790 5 3 1 20789
0 20791 7 1 2 35872 36648
0 20792 7 1 2 37384 20791
0 20793 5 1 1 20792
0 20794 7 1 2 36759 36983
0 20795 5 1 1 20794
0 20796 7 1 2 37386 20795
0 20797 7 1 2 20793 20796
0 20798 5 1 1 20797
0 20799 7 1 2 37389 20798
0 20800 5 1 1 20799
0 20801 7 1 2 20786 20800
0 20802 5 1 1 20801
0 20803 7 1 2 27997 20802
0 20804 5 1 1 20803
0 20805 7 1 2 24355 20804
0 20806 7 1 2 20771 20805
0 20807 5 1 1 20806
0 20808 7 1 2 20715 20807
0 20809 5 1 1 20808
0 20810 7 1 2 22164 37373
0 20811 5 1 1 20810
0 20812 7 1 2 37352 20811
0 20813 5 1 1 20812
0 20814 7 2 2 22723 20813
0 20815 5 1 1 37392
0 20816 7 1 2 35380 37393
0 20817 5 1 1 20816
0 20818 7 1 2 24178 37349
0 20819 5 1 1 20818
0 20820 7 1 2 37379 20819
0 20821 5 2 1 20820
0 20822 7 1 2 22346 37382
0 20823 7 1 2 37394 20822
0 20824 5 1 1 20823
0 20825 7 1 2 20817 20824
0 20826 5 1 1 20825
0 20827 7 1 2 34116 20826
0 20828 5 1 1 20827
0 20829 7 1 2 34909 36347
0 20830 7 1 2 29366 20829
0 20831 7 1 2 37309 20830
0 20832 5 1 1 20831
0 20833 7 1 2 20828 20832
0 20834 5 1 1 20833
0 20835 7 1 2 28697 20834
0 20836 5 1 1 20835
0 20837 7 1 2 35920 36921
0 20838 7 1 2 36778 20837
0 20839 5 1 1 20838
0 20840 7 1 2 33875 36576
0 20841 7 1 2 37362 20840
0 20842 5 1 1 20841
0 20843 7 1 2 20839 20842
0 20844 5 1 1 20843
0 20845 7 1 2 27910 20844
0 20846 5 1 1 20845
0 20847 7 2 2 36332 37395
0 20848 7 1 2 33876 37396
0 20849 5 1 1 20848
0 20850 7 1 2 22821 36770
0 20851 7 1 2 37318 20850
0 20852 7 1 2 37367 20851
0 20853 5 1 1 20852
0 20854 7 1 2 20849 20853
0 20855 5 1 1 20854
0 20856 7 1 2 27716 20855
0 20857 5 1 1 20856
0 20858 7 1 2 20846 20857
0 20859 5 1 1 20858
0 20860 7 1 2 34573 20859
0 20861 5 1 1 20860
0 20862 7 1 2 22279 37397
0 20863 5 1 1 20862
0 20864 7 1 2 20651 20863
0 20865 5 1 1 20864
0 20866 7 1 2 20865 34597
0 20867 5 1 1 20866
0 20868 7 1 2 26216 20867
0 20869 7 1 2 20861 20868
0 20870 7 1 2 20836 20869
0 20871 7 1 2 20809 20870
0 20872 5 1 1 20871
0 20873 7 1 2 20872 36112
0 20874 7 1 2 20594 20873
0 20875 5 1 1 20874
0 20876 7 1 2 20445 20875
0 20877 5 1 1 20876
0 20878 7 1 2 32996 20877
0 20879 5 1 1 20878
0 20880 7 2 2 27941 34667
0 20881 7 1 2 30028 37398
0 20882 5 1 1 20881
0 20883 7 1 2 29643 30726
0 20884 7 1 2 35101 20883
0 20885 5 1 1 20884
0 20886 7 1 2 20882 20885
0 20887 5 2 1 20886
0 20888 7 1 2 33572 37400
0 20889 5 1 1 20888
0 20890 7 1 2 28963 37273
0 20891 7 1 2 35575 20890
0 20892 7 1 2 31750 37371
0 20893 7 1 2 20891 20892
0 20894 5 1 1 20893
0 20895 7 1 2 20889 20894
0 20896 5 1 1 20895
0 20897 7 1 2 24993 20896
0 20898 5 1 1 20897
0 20899 7 1 2 37399 32872
0 20900 5 1 1 20899
0 20901 7 1 2 22724 36099
0 20902 7 1 2 31660 20901
0 20903 5 1 1 20902
0 20904 7 1 2 20900 20903
0 20905 5 1 1 20904
0 20906 7 1 2 34951 20905
0 20907 5 1 1 20906
0 20908 7 1 2 20898 20907
0 20909 5 1 1 20908
0 20910 7 1 2 20909 32066
0 20911 5 1 1 20910
0 20912 7 1 2 32699 34146
0 20913 5 1 1 20912
0 20914 7 1 2 20913 11260
0 20915 5 1 1 20914
0 20916 7 1 2 28864 20915
0 20917 5 1 1 20916
0 20918 7 1 2 23698 34818
0 20919 5 1 1 20918
0 20920 7 1 2 23588 26494
0 20921 7 1 2 26643 20920
0 20922 7 1 2 33730 20921
0 20923 5 1 1 20922
0 20924 7 1 2 20919 20923
0 20925 7 1 2 20917 20924
0 20926 5 1 1 20925
0 20927 7 1 2 36063 20926
0 20928 5 1 1 20927
0 20929 7 1 2 11507 9330
0 20930 5 1 1 20929
0 20931 7 1 2 21967 20930
0 20932 5 1 1 20931
0 20933 7 1 2 35905 34256
0 20934 5 1 1 20933
0 20935 7 1 2 22491 29733
0 20936 5 1 1 20935
0 20937 7 1 2 30214 20936
0 20938 5 1 1 20937
0 20939 7 1 2 21846 35548
0 20940 7 1 2 20938 20939
0 20941 5 1 1 20940
0 20942 7 1 2 20934 20941
0 20943 7 1 2 20932 20942
0 20944 5 1 1 20943
0 20945 7 1 2 34193 20944
0 20946 5 1 1 20945
0 20947 7 1 2 23888 21968
0 20948 5 2 1 20947
0 20949 7 1 2 30915 37402
0 20950 5 1 1 20949
0 20951 7 1 2 35027 31919
0 20952 7 1 2 20950 20951
0 20953 5 1 1 20952
0 20954 7 1 2 20946 20953
0 20955 5 1 1 20954
0 20956 7 1 2 25635 20955
0 20957 5 1 1 20956
0 20958 7 1 2 33630 35297
0 20959 5 1 1 20958
0 20960 7 1 2 26128 20959
0 20961 7 1 2 20957 20960
0 20962 5 1 1 20961
0 20963 7 1 2 34944 32063
0 20964 5 1 1 20963
0 20965 7 1 2 26138 20964
0 20966 5 1 1 20965
0 20967 7 1 2 26231 28996
0 20968 7 1 2 20966 20967
0 20969 7 1 2 20962 20968
0 20970 5 1 1 20969
0 20971 7 1 2 20928 20970
0 20972 5 1 1 20971
0 20973 7 1 2 22109 20972
0 20974 5 1 1 20973
0 20975 7 1 2 36707 36041
0 20976 5 1 1 20975
0 20977 7 1 2 33742 37068
0 20978 7 1 2 30946 20977
0 20979 5 1 1 20978
0 20980 7 1 2 20976 20979
0 20981 5 1 1 20980
0 20982 7 1 2 22581 20981
0 20983 5 1 1 20982
0 20984 7 1 2 32623 36048
0 20985 5 1 1 20984
0 20986 7 1 2 31399 32136
0 20987 7 1 2 33089 20986
0 20988 5 1 1 20987
0 20989 7 1 2 20985 20988
0 20990 5 1 1 20989
0 20991 7 1 2 33743 20990
0 20992 5 1 1 20991
0 20993 7 1 2 36049 35780
0 20994 5 1 1 20993
0 20995 7 1 2 20992 20994
0 20996 5 1 1 20995
0 20997 7 1 2 21969 20996
0 20998 5 1 1 20997
0 20999 7 1 2 20983 20998
0 21000 5 1 1 20999
0 21001 7 1 2 23589 21000
0 21002 5 1 1 21001
0 21003 7 1 2 30533 33877
0 21004 7 1 2 28905 21003
0 21005 7 1 2 35963 21004
0 21006 7 1 2 34473 21005
0 21007 5 1 1 21006
0 21008 7 1 2 21002 21007
0 21009 7 1 2 20974 21008
0 21010 5 1 1 21009
0 21011 7 1 2 25685 21010
0 21012 5 1 1 21011
0 21013 7 1 2 27911 37376
0 21014 5 1 1 21013
0 21015 7 1 2 27717 37346
0 21016 5 1 1 21015
0 21017 7 1 2 21014 21016
0 21018 5 1 1 21017
0 21019 7 1 2 33390 21018
0 21020 5 1 1 21019
0 21021 7 1 2 37347 35252
0 21022 5 1 1 21021
0 21023 7 1 2 35012 32544
0 21024 5 1 1 21023
0 21025 7 1 2 34466 37333
0 21026 5 1 1 21025
0 21027 7 1 2 21024 21026
0 21028 5 1 1 21027
0 21029 7 1 2 23152 21028
0 21030 5 1 1 21029
0 21031 7 1 2 21022 21030
0 21032 7 1 2 21020 21031
0 21033 5 1 1 21032
0 21034 7 1 2 25537 21033
0 21035 5 1 1 21034
0 21036 7 1 2 27892 10821
0 21037 5 1 1 21036
0 21038 7 1 2 33334 21037
0 21039 5 1 1 21038
0 21040 7 1 2 22582 33715
0 21041 5 1 1 21040
0 21042 7 1 2 21039 21041
0 21043 5 1 1 21042
0 21044 7 1 2 24134 21043
0 21045 5 1 1 21044
0 21046 7 1 2 28015 29967
0 21047 7 1 2 33720 21046
0 21048 5 1 1 21047
0 21049 7 1 2 21045 21048
0 21050 5 1 1 21049
0 21051 7 1 2 36922 21050
0 21052 5 1 1 21051
0 21053 7 1 2 35249 35573
0 21054 5 1 1 21053
0 21055 7 1 2 26217 21054
0 21056 7 1 2 21052 21055
0 21057 7 1 2 21035 21056
0 21058 5 1 1 21057
0 21059 7 1 2 33573 37363
0 21060 5 1 1 21059
0 21061 7 1 2 34725 32191
0 21062 7 1 2 35576 35279
0 21063 7 1 2 21061 21062
0 21064 5 1 1 21063
0 21065 7 1 2 21060 21064
0 21066 5 1 1 21065
0 21067 7 1 2 25636 21066
0 21068 5 1 1 21067
0 21069 7 1 2 26232 21068
0 21070 5 1 1 21069
0 21071 7 1 2 36113 21070
0 21072 7 1 2 21058 21071
0 21073 5 1 1 21072
0 21074 7 1 2 21012 21073
0 21075 5 1 1 21074
0 21076 7 1 2 36414 21075
0 21077 5 1 1 21076
0 21078 7 1 2 20911 21077
0 21079 5 1 1 21078
0 21080 7 1 2 34309 21079
0 21081 5 1 1 21080
0 21082 7 1 2 28227 30579
0 21083 5 1 1 21082
0 21084 7 1 2 23153 21083
0 21085 5 1 1 21084
0 21086 7 1 2 37344 21085
0 21087 5 1 1 21086
0 21088 7 1 2 32919 21087
0 21089 5 1 1 21088
0 21090 7 1 2 31419 33235
0 21091 5 1 1 21090
0 21092 7 1 2 21089 21091
0 21093 5 1 1 21092
0 21094 7 1 2 29380 21093
0 21095 5 1 1 21094
0 21096 7 1 2 30309 29877
0 21097 7 2 2 37364 21096
0 21098 7 1 2 24887 35377
0 21099 7 1 2 37404 21098
0 21100 5 1 1 21099
0 21101 7 1 2 21095 21100
0 21102 5 1 1 21101
0 21103 7 1 2 22425 21102
0 21104 5 1 1 21103
0 21105 7 1 2 26502 35961
0 21106 7 1 2 37405 21105
0 21107 5 1 1 21106
0 21108 7 1 2 21104 21107
0 21109 5 1 1 21108
0 21110 7 1 2 22347 21109
0 21111 5 1 1 21110
0 21112 7 1 2 25959 30310
0 21113 7 1 2 34602 21112
0 21114 7 1 2 37365 21113
0 21115 5 1 1 21114
0 21116 7 1 2 21111 21115
0 21117 5 1 1 21116
0 21118 7 1 2 23770 21117
0 21119 5 1 1 21118
0 21120 7 1 2 37292 32650
0 21121 5 1 1 21120
0 21122 7 1 2 37388 32759
0 21123 7 1 2 37358 21122
0 21124 5 2 1 21123
0 21125 7 1 2 27627 37406
0 21126 5 1 1 21125
0 21127 7 1 2 25110 35364
0 21128 5 1 1 21127
0 21129 7 1 2 36037 21128
0 21130 5 1 1 21129
0 21131 7 1 2 22583 21130
0 21132 5 1 1 21131
0 21133 7 1 2 37315 36051
0 21134 7 1 2 21132 21133
0 21135 5 2 1 21134
0 21136 7 1 2 27613 37408
0 21137 5 1 1 21136
0 21138 7 1 2 21126 21137
0 21139 5 1 1 21138
0 21140 7 1 2 25960 21139
0 21141 5 1 1 21140
0 21142 7 1 2 27912 35543
0 21143 5 1 1 21142
0 21144 7 1 2 27718 37409
0 21145 5 1 1 21144
0 21146 7 1 2 21143 21145
0 21147 5 1 1 21146
0 21148 7 1 2 27741 21147
0 21149 5 1 1 21148
0 21150 7 1 2 27913 37407
0 21151 5 1 1 21150
0 21152 7 1 2 27719 31742
0 21153 5 1 1 21152
0 21154 7 1 2 21151 21153
0 21155 5 1 1 21154
0 21156 7 1 2 27790 21155
0 21157 5 1 1 21156
0 21158 7 1 2 21149 21157
0 21159 7 1 2 21141 21158
0 21160 7 1 2 21121 21159
0 21161 5 1 1 21160
0 21162 7 1 2 32929 21161
0 21163 5 1 1 21162
0 21164 7 1 2 31218 33793
0 21165 7 1 2 32037 21164
0 21166 7 1 2 37312 21165
0 21167 5 1 1 21166
0 21168 7 1 2 21163 21167
0 21169 7 1 2 21119 21168
0 21170 5 1 1 21169
0 21171 7 1 2 36415 21170
0 21172 5 1 1 21171
0 21173 7 1 2 30288 35859
0 21174 7 2 2 34170 21173
0 21175 7 1 2 35312 37410
0 21176 5 1 1 21175
0 21177 7 1 2 28263 26592
0 21178 7 1 2 29713 34343
0 21179 7 1 2 21177 21178
0 21180 5 1 1 21179
0 21181 7 1 2 21176 21180
0 21182 5 1 1 21181
0 21183 7 1 2 30686 31380
0 21184 7 1 2 21182 21183
0 21185 5 1 1 21184
0 21186 7 1 2 24253 29415
0 21187 7 1 2 33704 21186
0 21188 7 1 2 28966 21187
0 21189 7 1 2 35636 21188
0 21190 5 1 1 21189
0 21191 7 1 2 21185 21190
0 21192 5 1 1 21191
0 21193 7 1 2 24994 21192
0 21194 5 1 1 21193
0 21195 7 1 2 29525 31400
0 21196 5 2 1 21195
0 21197 7 1 2 29318 1801
0 21198 5 1 1 21197
0 21199 7 1 2 21847 12145
0 21200 5 2 1 21199
0 21201 7 1 2 30893 37414
0 21202 7 1 2 21198 21201
0 21203 5 1 1 21202
0 21204 7 1 2 37412 21203
0 21205 5 1 1 21204
0 21206 7 1 2 25111 21205
0 21207 5 1 1 21206
0 21208 7 1 2 22110 37303
0 21209 5 1 1 21208
0 21210 7 1 2 21848 31201
0 21211 7 1 2 33055 21210
0 21212 5 2 1 21211
0 21213 7 1 2 21209 37416
0 21214 7 1 2 21207 21213
0 21215 5 1 1 21214
0 21216 7 1 2 29335 37411
0 21217 7 1 2 21215 21216
0 21218 5 1 1 21217
0 21219 7 1 2 21194 21218
0 21220 5 1 1 21219
0 21221 7 1 2 22426 21220
0 21222 5 1 1 21221
0 21223 7 1 2 24995 35719
0 21224 5 1 1 21223
0 21225 7 2 2 32663 21224
0 21226 5 1 1 37418
0 21227 7 1 2 23889 37419
0 21228 5 1 1 21227
0 21229 7 1 2 24006 28418
0 21230 7 1 2 37415 21229
0 21231 7 1 2 21228 21230
0 21232 5 1 1 21231
0 21233 7 1 2 37413 21232
0 21234 5 1 1 21233
0 21235 7 1 2 25112 21234
0 21236 5 1 1 21235
0 21237 7 1 2 29102 33796
0 21238 5 1 1 21237
0 21239 7 1 2 33142 21238
0 21240 5 1 1 21239
0 21241 7 1 2 22492 21240
0 21242 5 1 1 21241
0 21243 7 1 2 22111 31020
0 21244 5 1 1 21243
0 21245 7 2 2 21242 21244
0 21246 7 1 2 37420 37417
0 21247 7 1 2 21236 21246
0 21248 5 1 1 21247
0 21249 7 1 2 25878 31212
0 21250 7 1 2 31920 21249
0 21251 7 1 2 27085 21250
0 21252 7 1 2 21248 21251
0 21253 5 1 1 21252
0 21254 7 1 2 21222 21253
0 21255 5 1 1 21254
0 21256 7 1 2 23479 21255
0 21257 5 1 1 21256
0 21258 7 1 2 30933 37293
0 21259 5 1 1 21258
0 21260 7 1 2 35541 21259
0 21261 5 3 1 21260
0 21262 7 2 2 27042 37422
0 21263 7 1 2 34171 31948
0 21264 7 1 2 36636 21263
0 21265 7 1 2 37425 21264
0 21266 5 1 1 21265
0 21267 7 1 2 21257 21266
0 21268 5 1 1 21267
0 21269 7 1 2 24727 21268
0 21270 5 1 1 21269
0 21271 7 2 2 26618 32218
0 21272 7 1 2 27043 32070
0 21273 7 1 2 37427 21272
0 21274 5 1 1 21273
0 21275 7 1 2 33468 21274
0 21276 5 1 1 21275
0 21277 7 1 2 23890 21276
0 21278 5 1 1 21277
0 21279 7 2 2 22953 33433
0 21280 7 2 2 18488 37429
0 21281 7 1 2 28379 37431
0 21282 5 1 1 21281
0 21283 7 1 2 25113 21282
0 21284 7 1 2 21278 21283
0 21285 5 1 1 21284
0 21286 7 1 2 29630 33464
0 21287 5 1 1 21286
0 21288 7 1 2 28074 36910
0 21289 7 1 2 37265 21288
0 21290 5 1 1 21289
0 21291 7 1 2 23154 21290
0 21292 7 1 2 21287 21291
0 21293 5 1 1 21292
0 21294 7 1 2 22165 21293
0 21295 7 1 2 21285 21294
0 21296 5 1 1 21295
0 21297 7 1 2 29528 29939
0 21298 5 1 1 21297
0 21299 7 1 2 33132 21298
0 21300 5 1 1 21299
0 21301 7 1 2 22112 33465
0 21302 7 1 2 21300 21301
0 21303 5 1 1 21302
0 21304 7 1 2 21296 21303
0 21305 5 1 1 21304
0 21306 7 1 2 26593 21305
0 21307 5 1 1 21306
0 21308 7 1 2 31743 35997
0 21309 7 1 2 29654 21308
0 21310 7 1 2 33466 21309
0 21311 5 1 1 21310
0 21312 7 1 2 21307 21311
0 21313 5 1 1 21312
0 21314 7 1 2 22725 31902
0 21315 7 1 2 21313 21314
0 21316 5 1 1 21315
0 21317 7 1 2 21270 21316
0 21318 5 1 1 21317
0 21319 7 1 2 22348 21318
0 21320 5 1 1 21319
0 21321 7 1 2 30254 36753
0 21322 7 1 2 37192 21321
0 21323 5 1 1 21322
0 21324 7 1 2 36745 21323
0 21325 5 1 1 21324
0 21326 7 1 2 24424 21325
0 21327 5 1 1 21326
0 21328 7 1 2 36253 34163
0 21329 7 1 2 37188 21328
0 21330 5 1 1 21329
0 21331 7 1 2 21327 21330
0 21332 5 1 1 21331
0 21333 7 1 2 36064 21332
0 21334 5 1 1 21333
0 21335 7 2 2 32493 36790
0 21336 5 1 1 37433
0 21337 7 2 2 31715 36748
0 21338 7 1 2 30874 36381
0 21339 7 1 2 37435 21338
0 21340 5 1 1 21339
0 21341 7 1 2 21336 21340
0 21342 5 1 1 21341
0 21343 7 1 2 27202 21342
0 21344 5 1 1 21343
0 21345 7 1 2 29532 37403
0 21346 5 1 1 21345
0 21347 7 1 2 37037 36637
0 21348 7 1 2 21346 21347
0 21349 5 1 1 21348
0 21350 7 1 2 21344 21349
0 21351 5 1 1 21350
0 21352 7 1 2 28997 32957
0 21353 7 1 2 21351 21352
0 21354 5 1 1 21353
0 21355 7 1 2 21334 21354
0 21356 5 1 1 21355
0 21357 7 1 2 22113 21356
0 21358 5 1 1 21357
0 21359 7 1 2 37434 35646
0 21360 5 1 1 21359
0 21361 7 1 2 22584 30947
0 21362 5 1 1 21361
0 21363 7 1 2 21362 15504
0 21364 5 1 1 21363
0 21365 7 1 2 30484 37436
0 21366 7 1 2 21364 21365
0 21367 5 1 1 21366
0 21368 7 1 2 21360 21367
0 21369 5 1 1 21368
0 21370 7 1 2 32958 21369
0 21371 5 1 1 21370
0 21372 7 1 2 21358 21371
0 21373 5 1 1 21372
0 21374 7 1 2 25686 28713
0 21375 7 1 2 21373 21374
0 21376 5 1 1 21375
0 21377 7 1 2 21320 21376
0 21378 5 1 1 21377
0 21379 7 1 2 23699 21378
0 21380 5 1 1 21379
0 21381 7 1 2 27742 37423
0 21382 5 1 1 21381
0 21383 7 1 2 27791 37350
0 21384 5 1 1 21383
0 21385 7 1 2 21382 21384
0 21386 5 1 1 21385
0 21387 7 1 2 36416 21386
0 21388 5 1 1 21387
0 21389 7 1 2 31518 37401
0 21390 5 1 1 21389
0 21391 7 1 2 21388 21390
0 21392 5 1 1 21391
0 21393 7 1 2 37121 21392
0 21394 5 1 1 21393
0 21395 7 1 2 32959 32739
0 21396 5 1 1 21395
0 21397 7 1 2 7844 21396
0 21398 5 1 1 21397
0 21399 7 1 2 21970 21398
0 21400 5 1 1 21399
0 21401 7 1 2 30210 33192
0 21402 5 1 1 21401
0 21403 7 1 2 26040 31253
0 21404 5 1 1 21403
0 21405 7 1 2 21402 21404
0 21406 5 1 1 21405
0 21407 7 1 2 21849 21406
0 21408 5 1 1 21407
0 21409 7 1 2 23392 31883
0 21410 7 1 2 34257 21409
0 21411 5 1 1 21410
0 21412 7 1 2 21408 21411
0 21413 7 1 2 21400 21412
0 21414 5 1 1 21413
0 21415 7 1 2 37294 21414
0 21416 5 1 1 21415
0 21417 7 1 2 31254 35544
0 21418 5 1 1 21417
0 21419 7 1 2 21416 21418
0 21420 5 1 1 21419
0 21421 7 1 2 25687 37194
0 21422 7 1 2 21420 21421
0 21423 5 1 1 21422
0 21424 7 1 2 21394 21423
0 21425 7 1 2 21380 21424
0 21426 7 1 2 21172 21425
0 21427 5 1 1 21426
0 21428 7 1 2 25737 21427
0 21429 5 1 1 21428
0 21430 7 1 2 25766 33831
0 21431 5 1 1 21430
0 21432 7 1 2 36644 21431
0 21433 5 1 1 21432
0 21434 7 1 2 26562 21433
0 21435 5 1 1 21434
0 21436 7 1 2 36642 21435
0 21437 5 1 1 21436
0 21438 7 1 2 33931 21437
0 21439 5 1 1 21438
0 21440 7 1 2 21850 33335
0 21441 7 1 2 32494 21440
0 21442 7 1 2 36470 21441
0 21443 5 1 1 21442
0 21444 7 1 2 21439 21443
0 21445 5 1 1 21444
0 21446 7 1 2 37295 21445
0 21447 5 1 1 21446
0 21448 7 1 2 32318 11057
0 21449 5 1 1 21448
0 21450 7 1 2 22585 36039
0 21451 7 1 2 21449 21450
0 21452 5 1 1 21451
0 21453 7 2 2 36052 21452
0 21454 5 1 1 37437
0 21455 7 1 2 35083 21454
0 21456 5 1 1 21455
0 21457 7 1 2 35096 35539
0 21458 5 1 1 21457
0 21459 7 1 2 31635 30940
0 21460 7 1 2 35113 21459
0 21461 5 1 1 21460
0 21462 7 1 2 28737 34859
0 21463 7 1 2 36455 21462
0 21464 5 1 1 21463
0 21465 7 1 2 21461 21464
0 21466 5 1 1 21465
0 21467 7 1 2 22114 21466
0 21468 5 1 1 21467
0 21469 7 1 2 21458 21468
0 21470 7 1 2 21456 21469
0 21471 5 1 1 21470
0 21472 7 1 2 26563 21471
0 21473 5 1 1 21472
0 21474 7 1 2 29038 31744
0 21475 5 2 1 21474
0 21476 7 1 2 37438 37439
0 21477 5 1 1 21476
0 21478 7 1 2 36640 21477
0 21479 5 1 1 21478
0 21480 7 1 2 21473 21479
0 21481 5 1 1 21480
0 21482 7 1 2 33932 21481
0 21483 5 1 1 21482
0 21484 7 1 2 31017 32750
0 21485 5 1 1 21484
0 21486 7 1 2 21851 21485
0 21487 5 1 1 21486
0 21488 7 1 2 25114 28455
0 21489 7 1 2 21226 21488
0 21490 5 1 1 21489
0 21491 7 1 2 21487 21490
0 21492 7 1 2 37421 21491
0 21493 5 1 1 21492
0 21494 7 1 2 36616 21493
0 21495 5 1 1 21494
0 21496 7 2 2 21483 21495
0 21497 5 1 1 37441
0 21498 7 1 2 21447 37442
0 21499 5 1 1 21498
0 21500 7 1 2 27614 21499
0 21501 5 1 1 21500
0 21502 7 1 2 24179 37374
0 21503 5 1 1 21502
0 21504 7 1 2 37380 21503
0 21505 5 1 1 21504
0 21506 7 1 2 22240 21505
0 21507 5 1 1 21506
0 21508 7 1 2 20815 21507
0 21509 5 1 1 21508
0 21510 7 1 2 35764 20447
0 21511 7 2 2 21509 21510
0 21512 7 1 2 36121 37443
0 21513 5 1 1 21512
0 21514 7 1 2 21501 21513
0 21515 5 1 1 21514
0 21516 7 1 2 25961 21515
0 21517 5 1 1 21516
0 21518 7 2 2 22954 37444
0 21519 7 1 2 35939 37445
0 21520 5 1 1 21519
0 21521 7 1 2 21971 36626
0 21522 5 1 1 21521
0 21523 7 1 2 36620 31981
0 21524 5 1 1 21523
0 21525 7 1 2 15660 21524
0 21526 5 1 1 21525
0 21527 7 1 2 30211 21526
0 21528 5 1 1 21527
0 21529 7 1 2 26041 35975
0 21530 7 1 2 36960 21529
0 21531 5 1 1 21530
0 21532 7 1 2 21528 21531
0 21533 5 1 1 21532
0 21534 7 1 2 21852 21533
0 21535 5 1 1 21534
0 21536 7 1 2 27291 37227
0 21537 7 1 2 37184 21536
0 21538 7 1 2 31987 21537
0 21539 5 1 1 21538
0 21540 7 1 2 21535 21539
0 21541 7 1 2 21522 21540
0 21542 5 1 1 21541
0 21543 7 1 2 24728 21542
0 21544 5 1 1 21543
0 21545 7 1 2 28245 29802
0 21546 7 1 2 32049 21545
0 21547 7 1 2 36663 21546
0 21548 5 1 1 21547
0 21549 7 1 2 21544 21548
0 21550 5 1 1 21549
0 21551 7 1 2 33933 21550
0 21552 5 1 1 21551
0 21553 7 1 2 29261 31799
0 21554 7 1 2 36490 36010
0 21555 7 1 2 21553 21554
0 21556 5 1 1 21555
0 21557 7 1 2 21552 21556
0 21558 5 1 1 21557
0 21559 7 1 2 37296 21558
0 21560 5 1 1 21559
0 21561 7 1 2 27720 21497
0 21562 5 1 1 21561
0 21563 7 1 2 21560 21562
0 21564 5 1 1 21563
0 21565 7 1 2 27743 21564
0 21566 5 1 1 21565
0 21567 7 1 2 21520 21566
0 21568 7 1 2 21517 21567
0 21569 5 1 1 21568
0 21570 7 1 2 25360 21569
0 21571 5 1 1 21570
0 21572 7 1 2 37446 35770
0 21573 5 1 1 21572
0 21574 7 2 2 36376 33954
0 21575 7 1 2 34378 37447
0 21576 5 1 1 21575
0 21577 7 1 2 28515 34074
0 21578 5 1 1 21577
0 21579 7 1 2 21576 21578
0 21580 5 1 1 21579
0 21581 7 1 2 26678 21580
0 21582 5 1 1 21581
0 21583 7 1 2 22280 27947
0 21584 7 1 2 37448 21583
0 21585 5 1 1 21584
0 21586 7 1 2 21582 21585
0 21587 5 1 1 21586
0 21588 7 1 2 24425 21587
0 21589 5 1 1 21588
0 21590 7 1 2 23590 36472
0 21591 5 1 1 21590
0 21592 7 1 2 21589 21591
0 21593 5 1 1 21592
0 21594 7 1 2 33143 37335
0 21595 5 1 1 21594
0 21596 7 1 2 21853 21595
0 21597 5 1 1 21596
0 21598 7 1 2 37440 21597
0 21599 7 1 2 35642 21598
0 21600 5 1 1 21599
0 21601 7 1 2 21593 21600
0 21602 5 1 1 21601
0 21603 7 2 2 36761 36068
0 21604 7 1 2 37449 36763
0 21605 5 1 1 21604
0 21606 7 1 2 22784 34066
0 21607 7 1 2 36417 21606
0 21608 7 1 2 37313 21607
0 21609 5 1 1 21608
0 21610 7 1 2 21605 21609
0 21611 5 1 1 21610
0 21612 7 1 2 24426 21611
0 21613 5 1 1 21612
0 21614 7 1 2 24729 25889
0 21615 7 1 2 36649 21614
0 21616 7 1 2 37450 21615
0 21617 5 1 1 21616
0 21618 7 1 2 21613 21617
0 21619 7 1 2 21602 21618
0 21620 5 1 1 21619
0 21621 7 1 2 23480 21620
0 21622 5 1 1 21621
0 21623 7 1 2 37253 33905
0 21624 7 1 2 37424 21623
0 21625 5 1 1 21624
0 21626 7 1 2 21622 21625
0 21627 5 1 1 21626
0 21628 7 1 2 27599 21627
0 21629 5 1 1 21628
0 21630 7 1 2 21573 21629
0 21631 5 1 1 21630
0 21632 7 1 2 25361 21631
0 21633 5 1 1 21632
0 21634 7 3 2 23771 37390
0 21635 7 1 2 31696 34962
0 21636 7 2 2 37451 21635
0 21637 7 1 2 22427 33459
0 21638 7 1 2 37454 21637
0 21639 5 1 1 21638
0 21640 7 1 2 24254 36911
0 21641 7 1 2 36743 21640
0 21642 7 1 2 35433 21641
0 21643 7 1 2 36065 21642
0 21644 5 1 1 21643
0 21645 7 1 2 21639 21644
0 21646 5 1 1 21645
0 21647 7 1 2 26564 21646
0 21648 5 1 1 21647
0 21649 7 1 2 33584 36390
0 21650 7 1 2 37455 21649
0 21651 5 1 1 21650
0 21652 7 1 2 21648 21651
0 21653 5 1 1 21652
0 21654 7 1 2 26583 21653
0 21655 5 1 1 21654
0 21656 7 1 2 21633 21655
0 21657 5 1 1 21656
0 21658 7 1 2 28865 21657
0 21659 5 1 1 21658
0 21660 7 1 2 23481 31716
0 21661 7 1 2 34206 35315
0 21662 7 1 2 21660 21661
0 21663 7 1 2 37426 21662
0 21664 5 1 1 21663
0 21665 7 1 2 28275 34726
0 21666 7 1 2 34860 33959
0 21667 7 1 2 21665 21666
0 21668 7 1 2 37452 21667
0 21669 5 1 1 21668
0 21670 7 1 2 21664 21669
0 21671 5 1 1 21670
0 21672 7 1 2 26098 21671
0 21673 5 1 1 21672
0 21674 7 1 2 25962 37283
0 21675 7 1 2 37453 21674
0 21676 5 1 1 21675
0 21677 7 1 2 21673 21676
0 21678 5 1 1 21677
0 21679 7 1 2 26679 21678
0 21680 5 1 1 21679
0 21681 7 1 2 35333 35320
0 21682 7 1 2 33434 21681
0 21683 7 1 2 27948 21682
0 21684 7 1 2 25995 21683
0 21685 7 1 2 37391 21684
0 21686 5 1 1 21685
0 21687 7 1 2 21680 21686
0 21688 5 1 1 21687
0 21689 7 1 2 25637 21688
0 21690 5 1 1 21689
0 21691 7 2 2 37430 36872
0 21692 5 1 1 37456
0 21693 7 2 2 27549 34126
0 21694 7 1 2 24768 37428
0 21695 7 1 2 37458 21694
0 21696 5 1 1 21695
0 21697 7 1 2 21692 21696
0 21698 5 1 1 21697
0 21699 7 1 2 23891 21698
0 21700 5 1 1 21699
0 21701 7 1 2 37432 36873
0 21702 5 1 1 21701
0 21703 7 1 2 25115 21702
0 21704 7 1 2 21700 21703
0 21705 5 1 1 21704
0 21706 7 1 2 31694 36088
0 21707 7 1 2 37459 21706
0 21708 5 1 1 21707
0 21709 7 1 2 29631 37457
0 21710 5 1 1 21709
0 21711 7 1 2 23155 21710
0 21712 7 1 2 21708 21711
0 21713 5 1 1 21712
0 21714 7 1 2 24180 21713
0 21715 7 1 2 21705 21714
0 21716 5 1 1 21715
0 21717 7 1 2 35007 35579
0 21718 7 1 2 36711 21717
0 21719 7 1 2 32889 21718
0 21720 5 1 1 21719
0 21721 7 1 2 21716 21720
0 21722 5 1 1 21721
0 21723 7 1 2 25870 21722
0 21724 5 1 1 21723
0 21725 7 1 2 27044 25963
0 21726 7 1 2 29331 34336
0 21727 7 1 2 21725 21726
0 21728 7 1 2 36066 21727
0 21729 5 1 1 21728
0 21730 7 1 2 21724 21729
0 21731 5 1 1 21730
0 21732 7 1 2 23700 36333
0 21733 7 1 2 31903 21732
0 21734 7 1 2 21731 21733
0 21735 5 1 1 21734
0 21736 7 1 2 21690 21735
0 21737 5 1 1 21736
0 21738 7 1 2 23393 21737
0 21739 5 1 1 21738
0 21740 7 1 2 21659 21739
0 21741 7 1 2 21571 21740
0 21742 7 1 2 21429 21741
0 21743 7 1 2 21081 21742
0 21744 7 1 2 20879 21743
0 21745 5 1 1 21744
0 21746 7 1 2 32346 21745
0 21747 5 1 1 21746
0 21748 7 1 2 20284 21747
0 21749 7 1 2 19513 21748
0 21750 7 1 2 18237 21749
0 21751 7 1 2 17566 21750
0 21752 7 1 2 15237 21751
0 21753 7 1 2 13928 21752
0 21754 7 1 2 11905 21753
0 21755 7 1 2 4263 21754
3 49999 5 0 1 21755
