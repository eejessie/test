1 0 0 8 0
2 32 1 0
2 1985 1 0
2 1986 1 0
2 1987 1 0
2 1988 1 0
2 1989 1 0
2 1990 1 0
2 1991 1 0
1 1 0 10 0
2 1992 1 1
2 1993 1 1
2 1994 1 1
2 1995 1 1
2 1996 1 1
2 1997 1 1
2 1998 1 1
2 1999 1 1
2 2000 1 1
2 2001 1 1
1 2 0 10 0
2 2002 1 2
2 2003 1 2
2 2004 1 2
2 2005 1 2
2 2006 1 2
2 2007 1 2
2 2008 1 2
2 2009 1 2
2 2010 1 2
2 2011 1 2
1 3 0 11 0
2 2012 1 3
2 2013 1 3
2 2014 1 3
2 2015 1 3
2 2016 1 3
2 2017 1 3
2 2018 1 3
2 2019 1 3
2 2020 1 3
2 2021 1 3
2 2022 1 3
1 4 0 10 0
2 2023 1 4
2 2024 1 4
2 2025 1 4
2 2026 1 4
2 2027 1 4
2 2028 1 4
2 2029 1 4
2 2030 1 4
2 2031 1 4
2 2032 1 4
1 5 0 11 0
2 2033 1 5
2 2034 1 5
2 2035 1 5
2 2036 1 5
2 2037 1 5
2 2038 1 5
2 2039 1 5
2 2040 1 5
2 2041 1 5
2 2042 1 5
2 2043 1 5
1 6 0 10 0
2 2044 1 6
2 2045 1 6
2 2046 1 6
2 2047 1 6
2 2048 1 6
2 2049 1 6
2 2050 1 6
2 2051 1 6
2 2052 1 6
2 2053 1 6
1 7 0 10 0
2 2054 1 7
2 2055 1 7
2 2056 1 7
2 2057 1 7
2 2058 1 7
2 2059 1 7
2 2060 1 7
2 2061 1 7
2 2062 1 7
2 2063 1 7
1 8 0 10 0
2 2064 1 8
2 2065 1 8
2 2066 1 8
2 2067 1 8
2 2068 1 8
2 2069 1 8
2 2070 1 8
2 2071 1 8
2 2072 1 8
2 2073 1 8
1 9 0 10 0
2 2074 1 9
2 2075 1 9
2 2076 1 9
2 2077 1 9
2 2078 1 9
2 2079 1 9
2 2080 1 9
2 2081 1 9
2 2082 1 9
2 2083 1 9
1 10 0 11 0
2 2084 1 10
2 2085 1 10
2 2086 1 10
2 2087 1 10
2 2088 1 10
2 2089 1 10
2 2090 1 10
2 2091 1 10
2 2092 1 10
2 2093 1 10
2 2094 1 10
1 11 0 10 0
2 2095 1 11
2 2096 1 11
2 2097 1 11
2 2098 1 11
2 2099 1 11
2 2100 1 11
2 2101 1 11
2 2102 1 11
2 2103 1 11
2 2104 1 11
1 12 0 10 0
2 2105 1 12
2 2106 1 12
2 2107 1 12
2 2108 1 12
2 2109 1 12
2 2110 1 12
2 2111 1 12
2 2112 1 12
2 2113 1 12
2 2114 1 12
1 13 0 10 0
2 2115 1 13
2 2116 1 13
2 2117 1 13
2 2118 1 13
2 2119 1 13
2 2120 1 13
2 2121 1 13
2 2122 1 13
2 2123 1 13
2 2124 1 13
1 14 0 10 0
2 2125 1 14
2 2126 1 14
2 2127 1 14
2 2128 1 14
2 2129 1 14
2 2130 1 14
2 2131 1 14
2 2132 1 14
2 2133 1 14
2 2134 1 14
1 15 0 10 0
2 2135 1 15
2 2136 1 15
2 2137 1 15
2 2138 1 15
2 2139 1 15
2 2140 1 15
2 2141 1 15
2 2142 1 15
2 2143 1 15
2 2144 1 15
1 16 0 3 0
2 2145 1 16
2 2146 1 16
2 2147 1 16
1 17 0 3 0
2 2148 1 17
2 2149 1 17
2 2150 1 17
1 18 0 3 0
2 2151 1 18
2 2152 1 18
2 2153 1 18
1 19 0 3 0
2 2154 1 19
2 2155 1 19
2 2156 1 19
1 20 0 3 0
2 2157 1 20
2 2158 1 20
2 2159 1 20
1 21 0 3 0
2 2160 1 21
2 2161 1 21
2 2162 1 21
1 22 0 3 0
2 2163 1 22
2 2164 1 22
2 2165 1 22
1 23 0 3 0
2 2166 1 23
2 2167 1 23
2 2168 1 23
1 24 0 3 0
2 2169 1 24
2 2170 1 24
2 2171 1 24
1 25 0 3 0
2 2172 1 25
2 2173 1 25
2 2174 1 25
1 26 0 3 0
2 2175 1 26
2 2176 1 26
2 2177 1 26
1 27 0 3 0
2 2178 1 27
2 2179 1 27
2 2180 1 27
1 28 0 4 0
2 2181 1 28
2 2182 1 28
2 2183 1 28
2 2184 1 28
1 29 0 3 0
2 2185 1 29
2 2186 1 29
2 2187 1 29
1 30 0 4 0
2 2188 1 30
2 2189 1 30
2 2190 1 30
2 2191 1 30
1 31 0 4 0
2 2192 1 31
2 2193 1 31
2 2194 1 31
2 2195 1 31
2 2196 1 34
2 2197 1 34
2 2198 1 35
2 2199 1 35
2 2200 1 36
2 2201 1 36
2 2202 1 37
2 2203 1 37
2 2204 1 38
2 2205 1 38
2 2206 1 39
2 2207 1 39
2 2208 1 40
2 2209 1 40
2 2210 1 41
2 2211 1 41
2 2212 1 42
2 2213 1 42
2 2214 1 43
2 2215 1 43
2 2216 1 44
2 2217 1 44
2 2218 1 45
2 2219 1 45
2 2220 1 46
2 2221 1 46
2 2222 1 47
2 2223 1 47
2 2224 1 48
2 2225 1 48
2 2226 1 48
2 2227 1 49
2 2228 1 49
2 2229 1 49
2 2230 1 50
2 2231 1 50
2 2232 1 50
2 2233 1 51
2 2234 1 51
2 2235 1 51
2 2236 1 52
2 2237 1 52
2 2238 1 52
2 2239 1 53
2 2240 1 53
2 2241 1 53
2 2242 1 54
2 2243 1 54
2 2244 1 54
2 2245 1 55
2 2246 1 55
2 2247 1 55
2 2248 1 56
2 2249 1 56
2 2250 1 56
2 2251 1 57
2 2252 1 57
2 2253 1 57
2 2254 1 58
2 2255 1 58
2 2256 1 58
2 2257 1 59
2 2258 1 59
2 2259 1 59
2 2260 1 60
2 2261 1 60
2 2262 1 60
2 2263 1 60
2 2264 1 61
2 2265 1 61
2 2266 1 61
2 2267 1 62
2 2268 1 62
2 2269 1 63
2 2270 1 63
2 2271 1 64
2 2272 1 64
2 2273 1 66
2 2274 1 66
2 2275 1 66
2 2276 1 68
2 2277 1 68
2 2278 1 74
2 2279 1 74
2 2280 1 76
2 2281 1 76
2 2282 1 81
2 2283 1 81
2 2284 1 84
2 2285 1 84
2 2286 1 87
2 2287 1 87
2 2288 1 89
2 2289 1 89
2 2290 1 90
2 2291 1 90
2 2292 1 95
2 2293 1 95
2 2294 1 98
2 2295 1 98
2 2296 1 103
2 2297 1 103
2 2298 1 104
2 2299 1 104
2 2300 1 105
2 2301 1 105
2 2302 1 108
2 2303 1 108
2 2304 1 111
2 2305 1 111
2 2306 1 113
2 2307 1 113
2 2308 1 114
2 2309 1 114
2 2310 1 119
2 2311 1 119
2 2312 1 122
2 2313 1 122
2 2314 1 127
2 2315 1 127
2 2316 1 127
2 2317 1 129
2 2318 1 129
2 2319 1 132
2 2320 1 132
2 2321 1 135
2 2322 1 135
2 2323 1 137
2 2324 1 137
2 2325 1 138
2 2326 1 138
2 2327 1 143
2 2328 1 143
2 2329 1 146
2 2330 1 146
2 2331 1 151
2 2332 1 151
2 2333 1 151
2 2334 1 153
2 2335 1 153
2 2336 1 156
2 2337 1 156
2 2338 1 159
2 2339 1 159
2 2340 1 161
2 2341 1 161
2 2342 1 162
2 2343 1 162
2 2344 1 167
2 2345 1 167
2 2346 1 170
2 2347 1 170
2 2348 1 175
2 2349 1 175
2 2350 1 175
2 2351 1 177
2 2352 1 177
2 2353 1 180
2 2354 1 180
2 2355 1 183
2 2356 1 183
2 2357 1 185
2 2358 1 185
2 2359 1 186
2 2360 1 186
2 2361 1 191
2 2362 1 191
2 2363 1 194
2 2364 1 194
2 2365 1 199
2 2366 1 199
2 2367 1 199
2 2368 1 201
2 2369 1 201
2 2370 1 204
2 2371 1 204
2 2372 1 207
2 2373 1 207
2 2374 1 209
2 2375 1 209
2 2376 1 210
2 2377 1 210
2 2378 1 215
2 2379 1 215
2 2380 1 218
2 2381 1 218
2 2382 1 223
2 2383 1 223
2 2384 1 223
2 2385 1 225
2 2386 1 225
2 2387 1 228
2 2388 1 228
2 2389 1 231
2 2390 1 231
2 2391 1 233
2 2392 1 233
2 2393 1 234
2 2394 1 234
2 2395 1 239
2 2396 1 239
2 2397 1 242
2 2398 1 242
2 2399 1 247
2 2400 1 247
2 2401 1 247
2 2402 1 249
2 2403 1 249
2 2404 1 252
2 2405 1 252
2 2406 1 255
2 2407 1 255
2 2408 1 257
2 2409 1 257
2 2410 1 258
2 2411 1 258
2 2412 1 263
2 2413 1 263
2 2414 1 266
2 2415 1 266
2 2416 1 271
2 2417 1 271
2 2418 1 271
2 2419 1 273
2 2420 1 273
2 2421 1 276
2 2422 1 276
2 2423 1 279
2 2424 1 279
2 2425 1 281
2 2426 1 281
2 2427 1 282
2 2428 1 282
2 2429 1 287
2 2430 1 287
2 2431 1 290
2 2432 1 290
2 2433 1 295
2 2434 1 295
2 2435 1 295
2 2436 1 297
2 2437 1 297
2 2438 1 300
2 2439 1 300
2 2440 1 303
2 2441 1 303
2 2442 1 305
2 2443 1 305
2 2444 1 306
2 2445 1 306
2 2446 1 311
2 2447 1 311
2 2448 1 314
2 2449 1 314
2 2450 1 319
2 2451 1 319
2 2452 1 319
2 2453 1 321
2 2454 1 321
2 2455 1 324
2 2456 1 324
2 2457 1 327
2 2458 1 327
2 2459 1 329
2 2460 1 329
2 2461 1 330
2 2462 1 330
2 2463 1 335
2 2464 1 335
2 2465 1 338
2 2466 1 338
2 2467 1 343
2 2468 1 343
2 2469 1 343
2 2470 1 345
2 2471 1 345
2 2472 1 348
2 2473 1 348
2 2474 1 351
2 2475 1 351
2 2476 1 353
2 2477 1 353
2 2478 1 354
2 2479 1 354
2 2480 1 359
2 2481 1 359
2 2482 1 362
2 2483 1 362
2 2484 1 367
2 2485 1 367
2 2486 1 367
2 2487 1 369
2 2488 1 369
2 2489 1 372
2 2490 1 372
2 2491 1 375
2 2492 1 375
2 2493 1 377
2 2494 1 377
2 2495 1 378
2 2496 1 378
2 2497 1 383
2 2498 1 383
2 2499 1 386
2 2500 1 386
2 2501 1 391
2 2502 1 391
2 2503 1 391
2 2504 1 393
2 2505 1 393
2 2506 1 396
2 2507 1 396
2 2508 1 399
2 2509 1 399
2 2510 1 401
2 2511 1 401
2 2512 1 402
2 2513 1 402
2 2514 1 407
2 2515 1 407
2 2516 1 410
2 2517 1 410
2 2518 1 415
2 2519 1 415
2 2520 1 415
2 2521 1 417
2 2522 1 417
2 2523 1 420
2 2524 1 420
2 2525 1 423
2 2526 1 423
2 2527 1 425
2 2528 1 425
2 2529 1 426
2 2530 1 426
2 2531 1 431
2 2532 1 431
2 2533 1 434
2 2534 1 434
2 2535 1 439
2 2536 1 439
2 2537 1 439
2 2538 1 441
2 2539 1 441
2 2540 1 444
2 2541 1 444
2 2542 1 447
2 2543 1 447
2 2544 1 449
2 2545 1 449
2 2546 1 450
2 2547 1 450
2 2548 1 455
2 2549 1 455
2 2550 1 458
2 2551 1 458
2 2552 1 463
2 2553 1 463
2 2554 1 463
2 2555 1 465
2 2556 1 465
2 2557 1 468
2 2558 1 468
2 2559 1 471
2 2560 1 471
2 2561 1 473
2 2562 1 473
2 2563 1 474
2 2564 1 474
2 2565 1 479
2 2566 1 479
2 2567 1 482
2 2568 1 482
2 2569 1 487
2 2570 1 487
2 2571 1 487
2 2572 1 489
2 2573 1 489
2 2574 1 492
2 2575 1 492
2 2576 1 495
2 2577 1 495
2 2578 1 497
2 2579 1 497
2 2580 1 498
2 2581 1 498
2 2582 1 503
2 2583 1 503
2 2584 1 506
2 2585 1 506
2 2586 1 511
2 2587 1 511
2 2588 1 511
2 2589 1 513
2 2590 1 513
2 2591 1 516
2 2592 1 516
2 2593 1 519
2 2594 1 519
2 2595 1 521
2 2596 1 521
2 2597 1 522
2 2598 1 522
2 2599 1 527
2 2600 1 527
2 2601 1 530
2 2602 1 530
2 2603 1 535
2 2604 1 535
2 2605 1 535
2 2606 1 537
2 2607 1 537
2 2608 1 540
2 2609 1 540
2 2610 1 543
2 2611 1 543
2 2612 1 545
2 2613 1 545
2 2614 1 546
2 2615 1 546
2 2616 1 551
2 2617 1 551
2 2618 1 554
2 2619 1 554
2 2620 1 559
2 2621 1 559
2 2622 1 559
2 2623 1 561
2 2624 1 561
2 2625 1 564
2 2626 1 564
2 2627 1 567
2 2628 1 567
2 2629 1 569
2 2630 1 569
2 2631 1 570
2 2632 1 570
2 2633 1 575
2 2634 1 575
2 2635 1 578
2 2636 1 578
2 2637 1 583
2 2638 1 583
2 2639 1 583
2 2640 1 585
2 2641 1 585
2 2642 1 588
2 2643 1 588
2 2644 1 591
2 2645 1 591
2 2646 1 593
2 2647 1 593
2 2648 1 594
2 2649 1 594
2 2650 1 599
2 2651 1 599
2 2652 1 602
2 2653 1 602
2 2654 1 607
2 2655 1 607
2 2656 1 607
2 2657 1 609
2 2658 1 609
2 2659 1 612
2 2660 1 612
2 2661 1 615
2 2662 1 615
2 2663 1 617
2 2664 1 617
2 2665 1 618
2 2666 1 618
2 2667 1 623
2 2668 1 623
2 2669 1 626
2 2670 1 626
2 2671 1 631
2 2672 1 631
2 2673 1 631
2 2674 1 633
2 2675 1 633
2 2676 1 636
2 2677 1 636
2 2678 1 639
2 2679 1 639
2 2680 1 641
2 2681 1 641
2 2682 1 642
2 2683 1 642
2 2684 1 647
2 2685 1 647
2 2686 1 650
2 2687 1 650
2 2688 1 655
2 2689 1 655
2 2690 1 655
2 2691 1 657
2 2692 1 657
2 2693 1 660
2 2694 1 660
2 2695 1 663
2 2696 1 663
2 2697 1 665
2 2698 1 665
2 2699 1 666
2 2700 1 666
2 2701 1 671
2 2702 1 671
2 2703 1 674
2 2704 1 674
2 2705 1 679
2 2706 1 679
2 2707 1 679
2 2708 1 681
2 2709 1 681
2 2710 1 686
2 2711 1 686
2 2712 1 687
2 2713 1 687
2 2714 1 689
2 2715 1 689
2 2716 1 690
2 2717 1 690
2 2718 1 695
2 2719 1 695
2 2720 1 698
2 2721 1 698
2 2722 1 703
2 2723 1 703
2 2724 1 703
2 2725 1 711
2 2726 1 711
2 2727 1 714
2 2728 1 714
2 2729 1 717
2 2730 1 717
2 2731 1 727
2 2732 1 727
2 2733 1 734
2 2734 1 734
2 2735 1 736
2 2736 1 736
2 2737 1 738
2 2738 1 738
2 2739 1 739
2 2740 1 739
2 2741 1 740
2 2742 1 740
2 2743 1 742
2 2744 1 742
2 2745 1 745
2 2746 1 745
2 2747 1 748
2 2748 1 748
2 2749 1 751
2 2750 1 751
2 2751 1 752
2 2752 1 752
2 2753 1 754
2 2754 1 754
2 2755 1 756
2 2756 1 756
2 2757 1 762
2 2758 1 762
2 2759 1 765
2 2760 1 765
2 2761 1 765
2 2762 1 769
2 2763 1 769
2 2764 1 770
2 2765 1 770
2 2766 1 772
2 2767 1 772
2 2768 1 775
2 2769 1 775
2 2770 1 776
2 2771 1 776
2 2772 1 780
2 2773 1 780
2 2774 1 783
2 2775 1 783
2 2776 1 784
2 2777 1 784
2 2778 1 788
2 2779 1 788
2 2780 1 791
2 2781 1 791
2 2782 1 792
2 2783 1 792
2 2784 1 796
2 2785 1 796
2 2786 1 799
2 2787 1 799
2 2788 1 800
2 2789 1 800
2 2790 1 802
2 2791 1 802
2 2792 1 805
2 2793 1 805
2 2794 1 806
2 2795 1 806
2 2796 1 810
2 2797 1 810
2 2798 1 813
2 2799 1 813
2 2800 1 814
2 2801 1 814
2 2802 1 818
2 2803 1 818
2 2804 1 821
2 2805 1 821
2 2806 1 822
2 2807 1 822
2 2808 1 826
2 2809 1 826
2 2810 1 829
2 2811 1 829
2 2812 1 830
2 2813 1 830
2 2814 1 834
2 2815 1 834
2 2816 1 837
2 2817 1 837
2 2818 1 838
2 2819 1 838
2 2820 1 842
2 2821 1 842
2 2822 1 845
2 2823 1 845
2 2824 1 846
2 2825 1 846
2 2826 1 850
2 2827 1 850
2 2828 1 853
2 2829 1 853
2 2830 1 854
2 2831 1 854
2 2832 1 858
2 2833 1 858
2 2834 1 861
2 2835 1 861
2 2836 1 862
2 2837 1 862
2 2838 1 864
2 2839 1 864
2 2840 1 866
2 2841 1 866
2 2842 1 867
2 2843 1 867
2 2844 1 868
2 2845 1 868
2 2846 1 869
2 2847 1 869
2 2848 1 870
2 2849 1 870
2 2850 1 873
2 2851 1 873
2 2852 1 874
2 2853 1 874
2 2854 1 878
2 2855 1 878
2 2856 1 881
2 2857 1 881
2 2858 1 882
2 2859 1 882
2 2860 1 886
2 2861 1 886
2 2862 1 889
2 2863 1 889
2 2864 1 890
2 2865 1 890
2 2866 1 894
2 2867 1 894
2 2868 1 897
2 2869 1 897
2 2870 1 898
2 2871 1 898
2 2872 1 902
2 2873 1 902
2 2874 1 905
2 2875 1 905
2 2876 1 906
2 2877 1 906
2 2878 1 910
2 2879 1 910
2 2880 1 913
2 2881 1 913
2 2882 1 914
2 2883 1 914
2 2884 1 918
2 2885 1 918
2 2886 1 921
2 2887 1 921
2 2888 1 922
2 2889 1 922
2 2890 1 926
2 2891 1 926
2 2892 1 929
2 2893 1 929
2 2894 1 930
2 2895 1 930
2 2896 1 932
2 2897 1 932
2 2898 1 935
2 2899 1 935
2 2900 1 938
2 2901 1 938
2 2902 1 942
2 2903 1 942
2 2904 1 945
2 2905 1 945
2 2906 1 946
2 2907 1 946
2 2908 1 950
2 2909 1 950
2 2910 1 953
2 2911 1 953
2 2912 1 954
2 2913 1 954
2 2914 1 956
2 2915 1 956
2 2916 1 959
2 2917 1 959
2 2918 1 960
2 2919 1 960
2 2920 1 962
2 2921 1 962
2 2922 1 968
2 2923 1 968
2 2924 1 971
2 2925 1 971
2 2926 1 974
2 2927 1 974
2 2928 1 977
2 2929 1 977
2 2930 1 980
2 2931 1 980
2 2932 1 984
2 2933 1 984
2 2934 1 987
2 2935 1 987
2 2936 1 988
2 2937 1 988
2 2938 1 992
2 2939 1 992
2 2940 1 995
2 2941 1 995
2 2942 1 996
2 2943 1 996
2 2944 1 998
2 2945 1 998
2 2946 1 1001
2 2947 1 1001
2 2948 1 1004
2 2949 1 1004
2 2950 1 1008
2 2951 1 1008
2 2952 1 1011
2 2953 1 1011
2 2954 1 1012
2 2955 1 1012
2 2956 1 1016
2 2957 1 1016
2 2958 1 1019
2 2959 1 1019
2 2960 1 1020
2 2961 1 1020
2 2962 1 1024
2 2963 1 1024
2 2964 1 1027
2 2965 1 1027
2 2966 1 1028
2 2967 1 1028
2 2968 1 1032
2 2969 1 1032
2 2970 1 1035
2 2971 1 1035
2 2972 1 1036
2 2973 1 1036
2 2974 1 1040
2 2975 1 1040
2 2976 1 1043
2 2977 1 1043
2 2978 1 1044
2 2979 1 1044
2 2980 1 1046
2 2981 1 1046
2 2982 1 1049
2 2983 1 1049
2 2984 1 1050
2 2985 1 1050
2 2986 1 1054
2 2987 1 1054
2 2988 1 1057
2 2989 1 1057
2 2990 1 1058
2 2991 1 1058
2 2992 1 1060
2 2993 1 1060
2 2994 1 1062
2 2995 1 1062
2 2996 1 1065
2 2997 1 1065
2 2998 1 1066
2 2999 1 1066
2 3000 1 1068
2 3001 1 1068
2 3002 1 1070
2 3003 1 1070
2 3004 1 1072
2 3005 1 1072
2 3006 1 1074
2 3007 1 1074
2 3008 1 1075
2 3009 1 1075
2 3010 1 1076
2 3011 1 1076
2 3012 1 1077
2 3013 1 1077
2 3014 1 1078
2 3015 1 1078
2 3016 1 1079
2 3017 1 1079
2 3018 1 1080
2 3019 1 1080
2 3020 1 1081
2 3021 1 1081
2 3022 1 1083
2 3023 1 1083
2 3024 1 1086
2 3025 1 1086
2 3026 1 1090
2 3027 1 1090
2 3028 1 1093
2 3029 1 1093
2 3030 1 1096
2 3031 1 1096
2 3032 1 1100
2 3033 1 1100
2 3034 1 1103
2 3035 1 1103
2 3036 1 1104
2 3037 1 1104
2 3038 1 1107
2 3039 1 1107
2 3040 1 1108
2 3041 1 1108
2 3042 1 1112
2 3043 1 1112
2 3044 1 1115
2 3045 1 1115
2 3046 1 1116
2 3047 1 1116
2 3048 1 1120
2 3049 1 1120
2 3050 1 1123
2 3051 1 1123
2 3052 1 1124
2 3053 1 1124
2 3054 1 1128
2 3055 1 1128
2 3056 1 1131
2 3057 1 1131
2 3058 1 1134
2 3059 1 1134
2 3060 1 1138
2 3061 1 1138
2 3062 1 1141
2 3063 1 1141
2 3064 1 1144
2 3065 1 1144
2 3066 1 1148
2 3067 1 1148
2 3068 1 1151
2 3069 1 1151
2 3070 1 1152
2 3071 1 1152
2 3072 1 1154
2 3073 1 1154
2 3074 1 1157
2 3075 1 1157
2 3076 1 1158
2 3077 1 1158
2 3078 1 1162
2 3079 1 1162
2 3080 1 1165
2 3081 1 1165
2 3082 1 1166
2 3083 1 1166
2 3084 1 1170
2 3085 1 1170
2 3086 1 1173
2 3087 1 1173
2 3088 1 1174
2 3089 1 1174
2 3090 1 1178
2 3091 1 1178
2 3092 1 1181
2 3093 1 1181
2 3094 1 1182
2 3095 1 1182
2 3096 1 1186
2 3097 1 1186
2 3098 1 1189
2 3099 1 1189
2 3100 1 1190
2 3101 1 1190
2 3102 1 1194
2 3103 1 1194
2 3104 1 1197
2 3105 1 1197
2 3106 1 1198
2 3107 1 1198
2 3108 1 1200
2 3109 1 1200
2 3110 1 1206
2 3111 1 1206
2 3112 1 1209
2 3113 1 1209
2 3114 1 1212
2 3115 1 1212
2 3116 1 1215
2 3117 1 1215
2 3118 1 1218
2 3119 1 1218
2 3120 1 1222
2 3121 1 1222
2 3122 1 1225
2 3123 1 1225
2 3124 1 1226
2 3125 1 1226
2 3126 1 1230
2 3127 1 1230
2 3128 1 1233
2 3129 1 1233
2 3130 1 1234
2 3131 1 1234
2 3132 1 1238
2 3133 1 1238
2 3134 1 1241
2 3135 1 1241
2 3136 1 1242
2 3137 1 1242
2 3138 1 1246
2 3139 1 1246
2 3140 1 1249
2 3141 1 1249
2 3142 1 1250
2 3143 1 1250
2 3144 1 1254
2 3145 1 1254
2 3146 1 1257
2 3147 1 1257
2 3148 1 1258
2 3149 1 1258
2 3150 1 1262
2 3151 1 1262
2 3152 1 1265
2 3153 1 1265
2 3154 1 1266
2 3155 1 1266
2 3156 1 1270
2 3157 1 1270
2 3158 1 1273
2 3159 1 1273
2 3160 1 1274
2 3161 1 1274
2 3162 1 1276
2 3163 1 1276
2 3164 1 1279
2 3165 1 1279
2 3166 1 1282
2 3167 1 1282
2 3168 1 1286
2 3169 1 1286
2 3170 1 1289
2 3171 1 1289
2 3172 1 1290
2 3173 1 1290
2 3174 1 1294
2 3175 1 1294
2 3176 1 1297
2 3177 1 1297
2 3178 1 1298
2 3179 1 1298
2 3180 1 1302
2 3181 1 1302
2 3182 1 1305
2 3183 1 1305
2 3184 1 1306
2 3185 1 1306
2 3186 1 1310
2 3187 1 1310
2 3188 1 1313
2 3189 1 1313
2 3190 1 1314
2 3191 1 1314
2 3192 1 1320
2 3193 1 1320
2 3194 1 1323
2 3195 1 1323
2 3196 1 1324
2 3197 1 1324
2 3198 1 1328
2 3199 1 1328
2 3200 1 1331
2 3201 1 1331
2 3202 1 1332
2 3203 1 1332
2 3204 1 1336
2 3205 1 1336
2 3206 1 1339
2 3207 1 1339
2 3208 1 1340
2 3209 1 1340
2 3210 1 1344
2 3211 1 1344
2 3212 1 1347
2 3213 1 1347
2 3214 1 1348
2 3215 1 1348
2 3216 1 1350
2 3217 1 1350
2 3218 1 1353
2 3219 1 1353
2 3220 1 1356
2 3221 1 1356
2 3222 1 1360
2 3223 1 1360
2 3224 1 1363
2 3225 1 1363
2 3226 1 1364
2 3227 1 1364
2 3228 1 1368
2 3229 1 1368
2 3230 1 1371
2 3231 1 1371
2 3232 1 1374
2 3233 1 1374
2 3234 1 1376
2 3235 1 1376
2 3236 1 1378
2 3237 1 1378
2 3238 1 1380
2 3239 1 1380
2 3240 1 1382
2 3241 1 1382
2 3242 1 1384
2 3243 1 1384
2 3244 1 1386
2 3245 1 1386
2 3246 1 1387
2 3247 1 1387
2 3248 1 1388
2 3249 1 1388
2 3250 1 1388
2 3251 1 1391
2 3252 1 1391
2 3253 1 1394
2 3254 1 1394
2 3255 1 1402
2 3256 1 1402
2 3257 1 1405
2 3258 1 1405
2 3259 1 1406
2 3260 1 1406
2 3261 1 1410
2 3262 1 1410
2 3263 1 1413
2 3264 1 1413
2 3265 1 1416
2 3266 1 1416
2 3267 1 1418
2 3268 1 1418
2 3269 1 1420
2 3270 1 1420
2 3271 1 1422
2 3272 1 1422
2 3273 1 1423
2 3274 1 1423
2 3275 1 1425
2 3276 1 1425
2 3277 1 1426
2 3278 1 1426
2 3279 1 1430
2 3280 1 1430
2 3281 1 1433
2 3282 1 1433
2 3283 1 1434
2 3284 1 1434
2 3285 1 1438
2 3286 1 1438
2 3287 1 1441
2 3288 1 1441
2 3289 1 1442
2 3290 1 1442
2 3291 1 1446
2 3292 1 1446
2 3293 1 1449
2 3294 1 1449
2 3295 1 1450
2 3296 1 1450
2 3297 1 1454
2 3298 1 1454
2 3299 1 1457
2 3300 1 1457
2 3301 1 1458
2 3302 1 1458
2 3303 1 1462
2 3304 1 1462
2 3305 1 1465
2 3306 1 1465
2 3307 1 1466
2 3308 1 1466
2 3309 1 1470
2 3310 1 1470
2 3311 1 1473
2 3312 1 1473
2 3313 1 1474
2 3314 1 1474
2 3315 1 1478
2 3316 1 1478
2 3317 1 1481
2 3318 1 1481
2 3319 1 1482
2 3320 1 1482
2 3321 1 1486
2 3322 1 1486
2 3323 1 1489
2 3324 1 1489
2 3325 1 1490
2 3326 1 1490
2 3327 1 1494
2 3328 1 1494
2 3329 1 1497
2 3330 1 1497
2 3331 1 1498
2 3332 1 1498
2 3333 1 1502
2 3334 1 1502
2 3335 1 1505
2 3336 1 1505
2 3337 1 1506
2 3338 1 1506
2 3339 1 1510
2 3340 1 1510
2 3341 1 1513
2 3342 1 1513
2 3343 1 1514
2 3344 1 1514
2 3345 1 1518
2 3346 1 1518
2 3347 1 1521
2 3348 1 1521
2 3349 1 1522
2 3350 1 1522
2 3351 1 1524
2 3352 1 1524
2 3353 1 1525
2 3354 1 1525
2 3355 1 1525
2 3356 1 1528
2 3357 1 1528
2 3358 1 1530
2 3359 1 1530
2 3360 1 1531
2 3361 1 1531
2 3362 1 1531
2 3363 1 1532
2 3364 1 1532
2 3365 1 1533
2 3366 1 1533
2 3367 1 1534
2 3368 1 1534
2 3369 1 1537
2 3370 1 1537
2 3371 1 1540
2 3372 1 1540
2 3373 1 1540
2 3374 1 1542
2 3375 1 1542
2 3376 1 1542
2 3377 1 1542
2 3378 1 1545
2 3379 1 1545
2 3380 1 1548
2 3381 1 1548
2 3382 1 1548
2 3383 1 1548
2 3384 1 1550
2 3385 1 1550
2 3386 1 1553
2 3387 1 1553
2 3388 1 1556
2 3389 1 1556
2 3390 1 1556
2 3391 1 1557
2 3392 1 1557
2 3393 1 1557
2 3394 1 1558
2 3395 1 1558
2 3396 1 1559
2 3397 1 1559
2 3398 1 1559
2 3399 1 1559
2 3400 1 1562
2 3401 1 1562
2 3402 1 1565
2 3403 1 1565
2 3404 1 1565
2 3405 1 1567
2 3406 1 1567
2 3407 1 1567
2 3408 1 1570
2 3409 1 1570
2 3410 1 1573
2 3411 1 1573
2 3412 1 1573
2 3413 1 1574
2 3414 1 1574
2 3415 1 1575
2 3416 1 1575
2 3417 1 1576
2 3418 1 1576
2 3419 1 1576
2 3420 1 1576
2 3421 1 1579
2 3422 1 1579
2 3423 1 1582
2 3424 1 1582
2 3425 1 1582
2 3426 1 1584
2 3427 1 1584
2 3428 1 1584
2 3429 1 1584
2 3430 1 1587
2 3431 1 1587
2 3432 1 1590
2 3433 1 1590
2 3434 1 1590
2 3435 1 1592
2 3436 1 1592
2 3437 1 1592
2 3438 1 1592
2 3439 1 1595
2 3440 1 1595
2 3441 1 1598
2 3442 1 1598
2 3443 1 1598
2 3444 1 1600
2 3445 1 1600
2 3446 1 1600
2 3447 1 1600
2 3448 1 1603
2 3449 1 1603
2 3450 1 1606
2 3451 1 1606
2 3452 1 1606
2 3453 1 1606
2 3454 1 1608
2 3455 1 1608
2 3456 1 1608
2 3457 1 1608
2 3458 1 1611
2 3459 1 1611
2 3460 1 1614
2 3461 1 1614
2 3462 1 1614
2 3463 1 1614
2 3464 1 1616
2 3465 1 1616
2 3466 1 1616
2 3467 1 1616
2 3468 1 1619
2 3469 1 1619
2 3470 1 1622
2 3471 1 1622
2 3472 1 1622
2 3473 1 1622
2 3474 1 1624
2 3475 1 1624
2 3476 1 1624
2 3477 1 1627
2 3478 1 1627
2 3479 1 1630
2 3480 1 1630
2 3481 1 1630
2 3482 1 1632
2 3483 1 1632
2 3484 1 1632
2 3485 1 1632
2 3486 1 1635
2 3487 1 1635
2 3488 1 1638
2 3489 1 1638
2 3490 1 1640
2 3491 1 1640
2 3492 1 1641
2 3493 1 1641
2 3494 1 1645
2 3495 1 1645
2 3496 1 1648
2 3497 1 1648
2 3498 1 1648
2 3499 1 1651
2 3500 1 1651
2 3501 1 1651
2 3502 1 1655
2 3503 1 1655
2 3504 1 1657
2 3505 1 1657
2 3506 1 1659
2 3507 1 1659
2 3508 1 1660
2 3509 1 1660
2 3510 1 1663
2 3511 1 1663
2 3512 1 1664
2 3513 1 1664
2 3514 1 1667
2 3515 1 1667
2 3516 1 1668
2 3517 1 1668
2 3518 1 1671
2 3519 1 1671
2 3520 1 1672
2 3521 1 1672
2 3522 1 1675
2 3523 1 1675
2 3524 1 1675
2 3525 1 1681
2 3526 1 1681
2 3527 1 1681
2 3528 1 1687
2 3529 1 1687
2 3530 1 1688
2 3531 1 1688
2 3532 1 1691
2 3533 1 1691
2 3534 1 1692
2 3535 1 1692
2 3536 1 1694
2 3537 1 1694
2 3538 1 1694
2 3539 1 1694
2 3540 1 1699
2 3541 1 1699
2 3542 1 1700
2 3543 1 1700
2 3544 1 1703
2 3545 1 1703
2 3546 1 1703
2 3547 1 1704
2 3548 1 1704
2 3549 1 1705
2 3550 1 1705
2 3551 1 1708
2 3552 1 1708
2 3553 1 1709
2 3554 1 1709
2 3555 1 1711
2 3556 1 1711
2 3557 1 1712
2 3558 1 1712
2 3559 1 1715
2 3560 1 1715
2 3561 1 1717
2 3562 1 1717
2 3563 1 1719
2 3564 1 1719
2 3565 1 1720
2 3566 1 1720
2 3567 1 1723
2 3568 1 1723
2 3569 1 1724
2 3570 1 1724
2 3571 1 1727
2 3572 1 1727
2 3573 1 1728
2 3574 1 1728
2 3575 1 1731
2 3576 1 1731
2 3577 1 1732
2 3578 1 1732
2 3579 1 1735
2 3580 1 1735
2 3581 1 1736
2 3582 1 1736
2 3583 1 1739
2 3584 1 1739
2 3585 1 1739
2 3586 1 1740
2 3587 1 1740
2 3588 1 1743
2 3589 1 1743
2 3590 1 1745
2 3591 1 1745
2 3592 1 1746
2 3593 1 1746
2 3594 1 1747
2 3595 1 1747
2 3596 1 1747
2 3597 1 1748
2 3598 1 1748
2 3599 1 1757
2 3600 1 1757
2 3601 1 1759
2 3602 1 1759
2 3603 1 1769
2 3604 1 1769
2 3605 1 1769
2 3606 1 1770
2 3607 1 1770
2 3608 1 1777
2 3609 1 1777
2 3610 1 1777
2 3611 1 1778
2 3612 1 1778
2 3613 1 1783
2 3614 1 1783
2 3615 1 1783
2 3616 1 1784
2 3617 1 1784
2 3618 1 1791
2 3619 1 1791
2 3620 1 1791
2 3621 1 1792
2 3622 1 1792
2 3623 1 1795
2 3624 1 1795
2 3625 1 1795
2 3626 1 1796
2 3627 1 1796
2 3628 1 1801
2 3629 1 1801
2 3630 1 1801
2 3631 1 1802
2 3632 1 1802
2 3633 1 1807
2 3634 1 1807
2 3635 1 1808
2 3636 1 1808
2 3637 1 1811
2 3638 1 1811
2 3639 1 1812
2 3640 1 1812
2 3641 1 1817
2 3642 1 1817
2 3643 1 1818
2 3644 1 1818
2 3645 1 1823
2 3646 1 1823
2 3647 1 1824
2 3648 1 1824
2 3649 1 1860
2 3650 1 1860
2 3651 1 1864
2 3652 1 1864
2 3653 1 1865
2 3654 1 1865
0 33 5 1 1 1992
0 34 5 2 1 2002
0 35 5 2 1 2012
0 36 5 2 1 2023
0 37 5 2 1 2033
0 38 5 2 1 2044
0 39 5 2 1 2054
0 40 5 2 1 2064
0 41 5 2 1 2074
0 42 5 2 1 2084
0 43 5 2 1 2095
0 44 5 2 1 2105
0 45 5 2 1 2115
0 46 5 2 1 2125
0 47 5 2 1 2135
0 48 5 3 1 2145
0 49 5 3 1 2148
0 50 5 3 1 2151
0 51 5 3 1 2154
0 52 5 3 1 2157
0 53 5 3 1 2160
0 54 5 3 1 2163
0 55 5 3 1 2166
0 56 5 3 1 2169
0 57 5 3 1 2172
0 58 5 3 1 2175
0 59 5 3 1 2178
0 60 5 4 1 2181
0 61 5 3 1 2185
0 62 5 2 1 2188
0 63 5 2 1 2192
0 64 7 2 2 2264 2267
0 65 5 1 1 2271
0 66 7 3 2 2193 2272
0 67 5 1 1 2273
0 68 7 2 2 2265 2194
0 69 5 1 1 2276
0 70 7 1 2 65 2277
0 71 5 1 1 70
0 72 7 1 2 2186 2269
0 73 5 1 1 72
0 74 7 2 2 71 73
0 75 5 1 1 2278
0 76 7 2 2 2260 2279
0 77 5 1 1 2280
0 78 7 1 2 2189 69
0 79 7 1 2 77 78
0 80 5 1 1 79
0 81 7 2 2 67 80
0 82 5 1 1 2282
0 83 7 1 2 2261 82
0 84 5 2 1 83
0 85 7 1 2 2182 2283
0 86 5 1 1 85
0 87 7 2 2 2284 86
0 88 5 1 1 2286
0 89 7 2 2 2257 2287
0 90 5 2 1 2288
0 91 7 1 2 75 2285
0 92 5 1 1 91
0 93 7 1 2 2262 2274
0 94 5 1 1 93
0 95 7 2 2 92 94
0 96 5 1 1 2292
0 97 7 1 2 2290 96
0 98 5 2 1 97
0 99 7 1 2 2190 2281
0 100 5 1 1 99
0 101 7 1 2 2183 2275
0 102 5 1 1 101
0 103 7 2 2 100 102
0 104 5 2 1 2296
0 105 7 2 2 2294 2297
0 106 5 1 1 2300
0 107 7 1 2 2258 106
0 108 5 2 1 107
0 109 7 1 2 2179 2301
0 110 5 1 1 109
0 111 7 2 2 2302 110
0 112 5 1 1 2304
0 113 7 2 2 2254 2305
0 114 5 2 1 2306
0 115 7 1 2 88 2303
0 116 5 1 1 115
0 117 7 1 2 2289 2298
0 118 5 1 1 117
0 119 7 2 2 116 118
0 120 5 1 1 2310
0 121 7 1 2 2308 120
0 122 5 2 1 121
0 123 7 1 2 2291 2299
0 124 5 1 1 123
0 125 7 1 2 2293 124
0 126 5 1 1 125
0 127 7 3 2 2295 126
0 128 5 1 1 2314
0 129 7 2 2 2312 128
0 130 5 1 1 2317
0 131 7 1 2 2255 130
0 132 5 2 1 131
0 133 7 1 2 2176 2318
0 134 5 1 1 133
0 135 7 2 2 2319 134
0 136 5 1 1 2321
0 137 7 2 2 2251 2322
0 138 5 2 1 2323
0 139 7 1 2 112 2320
0 140 5 1 1 139
0 141 7 1 2 2307 2315
0 142 5 1 1 141
0 143 7 2 2 140 142
0 144 5 1 1 2327
0 145 7 1 2 2325 144
0 146 5 2 1 145
0 147 7 1 2 2309 2316
0 148 5 1 1 147
0 149 7 1 2 2311 148
0 150 5 1 1 149
0 151 7 3 2 2313 150
0 152 5 1 1 2331
0 153 7 2 2 2329 152
0 154 5 1 1 2334
0 155 7 1 2 2252 154
0 156 5 2 1 155
0 157 7 1 2 2173 2335
0 158 5 1 1 157
0 159 7 2 2 2336 158
0 160 5 1 1 2338
0 161 7 2 2 2248 2339
0 162 5 2 1 2340
0 163 7 1 2 136 2337
0 164 5 1 1 163
0 165 7 1 2 2324 2332
0 166 5 1 1 165
0 167 7 2 2 164 166
0 168 5 1 1 2344
0 169 7 1 2 2342 168
0 170 5 2 1 169
0 171 7 1 2 2326 2333
0 172 5 1 1 171
0 173 7 1 2 2328 172
0 174 5 1 1 173
0 175 7 3 2 2330 174
0 176 5 1 1 2348
0 177 7 2 2 2346 176
0 178 5 1 1 2351
0 179 7 1 2 2249 178
0 180 5 2 1 179
0 181 7 1 2 2170 2352
0 182 5 1 1 181
0 183 7 2 2 2353 182
0 184 5 1 1 2355
0 185 7 2 2 2245 2356
0 186 5 2 1 2357
0 187 7 1 2 160 2354
0 188 5 1 1 187
0 189 7 1 2 2341 2349
0 190 5 1 1 189
0 191 7 2 2 188 190
0 192 5 1 1 2361
0 193 7 1 2 2359 192
0 194 5 2 1 193
0 195 7 1 2 2343 2350
0 196 5 1 1 195
0 197 7 1 2 2345 196
0 198 5 1 1 197
0 199 7 3 2 2347 198
0 200 5 1 1 2365
0 201 7 2 2 2363 200
0 202 5 1 1 2368
0 203 7 1 2 2246 202
0 204 5 2 1 203
0 205 7 1 2 2167 2369
0 206 5 1 1 205
0 207 7 2 2 2370 206
0 208 5 1 1 2372
0 209 7 2 2 2242 2373
0 210 5 2 1 2374
0 211 7 1 2 184 2371
0 212 5 1 1 211
0 213 7 1 2 2358 2366
0 214 5 1 1 213
0 215 7 2 2 212 214
0 216 5 1 1 2378
0 217 7 1 2 2376 216
0 218 5 2 1 217
0 219 7 1 2 2360 2367
0 220 5 1 1 219
0 221 7 1 2 2362 220
0 222 5 1 1 221
0 223 7 3 2 2364 222
0 224 5 1 1 2382
0 225 7 2 2 2380 224
0 226 5 1 1 2385
0 227 7 1 2 2243 226
0 228 5 2 1 227
0 229 7 1 2 2164 2386
0 230 5 1 1 229
0 231 7 2 2 2387 230
0 232 5 1 1 2389
0 233 7 2 2 2239 2390
0 234 5 2 1 2391
0 235 7 1 2 208 2388
0 236 5 1 1 235
0 237 7 1 2 2375 2383
0 238 5 1 1 237
0 239 7 2 2 236 238
0 240 5 1 1 2395
0 241 7 1 2 2393 240
0 242 5 2 1 241
0 243 7 1 2 2377 2384
0 244 5 1 1 243
0 245 7 1 2 2379 244
0 246 5 1 1 245
0 247 7 3 2 2381 246
0 248 5 1 1 2399
0 249 7 2 2 2397 248
0 250 5 1 1 2402
0 251 7 1 2 2240 250
0 252 5 2 1 251
0 253 7 1 2 2161 2403
0 254 5 1 1 253
0 255 7 2 2 2404 254
0 256 5 1 1 2406
0 257 7 2 2 2236 2407
0 258 5 2 1 2408
0 259 7 1 2 232 2405
0 260 5 1 1 259
0 261 7 1 2 2392 2400
0 262 5 1 1 261
0 263 7 2 2 260 262
0 264 5 1 1 2412
0 265 7 1 2 2410 264
0 266 5 2 1 265
0 267 7 1 2 2394 2401
0 268 5 1 1 267
0 269 7 1 2 2396 268
0 270 5 1 1 269
0 271 7 3 2 2398 270
0 272 5 1 1 2416
0 273 7 2 2 2414 272
0 274 5 1 1 2419
0 275 7 1 2 2237 274
0 276 5 2 1 275
0 277 7 1 2 2158 2420
0 278 5 1 1 277
0 279 7 2 2 2421 278
0 280 5 1 1 2423
0 281 7 2 2 2233 2424
0 282 5 2 1 2425
0 283 7 1 2 256 2422
0 284 5 1 1 283
0 285 7 1 2 2409 2417
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 2429
0 289 7 1 2 2427 288
0 290 5 2 1 289
0 291 7 1 2 2411 2418
0 292 5 1 1 291
0 293 7 1 2 2413 292
0 294 5 1 1 293
0 295 7 3 2 2415 294
0 296 5 1 1 2433
0 297 7 2 2 2431 296
0 298 5 1 1 2436
0 299 7 1 2 2234 298
0 300 5 2 1 299
0 301 7 1 2 2155 2437
0 302 5 1 1 301
0 303 7 2 2 2438 302
0 304 5 1 1 2440
0 305 7 2 2 2230 2441
0 306 5 2 1 2442
0 307 7 1 2 280 2439
0 308 5 1 1 307
0 309 7 1 2 2426 2434
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 2446
0 313 7 1 2 2444 312
0 314 5 2 1 313
0 315 7 1 2 2428 2435
0 316 5 1 1 315
0 317 7 1 2 2430 316
0 318 5 1 1 317
0 319 7 3 2 2432 318
0 320 5 1 1 2450
0 321 7 2 2 2448 320
0 322 5 1 1 2453
0 323 7 1 2 2231 322
0 324 5 2 1 323
0 325 7 1 2 2152 2454
0 326 5 1 1 325
0 327 7 2 2 2455 326
0 328 5 1 1 2457
0 329 7 2 2 2227 2458
0 330 5 2 1 2459
0 331 7 1 2 304 2456
0 332 5 1 1 331
0 333 7 1 2 2443 2451
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 2463
0 337 7 1 2 2461 336
0 338 5 2 1 337
0 339 7 1 2 2445 2452
0 340 5 1 1 339
0 341 7 1 2 2447 340
0 342 5 1 1 341
0 343 7 3 2 2449 342
0 344 5 1 1 2467
0 345 7 2 2 2465 344
0 346 5 1 1 2470
0 347 7 1 2 2228 346
0 348 5 2 1 347
0 349 7 1 2 2149 2471
0 350 5 1 1 349
0 351 7 2 2 2472 350
0 352 5 1 1 2474
0 353 7 2 2 2224 2475
0 354 5 2 1 2476
0 355 7 1 2 328 2473
0 356 5 1 1 355
0 357 7 1 2 2460 2468
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 2480
0 361 7 1 2 2478 360
0 362 5 2 1 361
0 363 7 1 2 2462 2469
0 364 5 1 1 363
0 365 7 1 2 2464 364
0 366 5 1 1 365
0 367 7 3 2 2466 366
0 368 5 1 1 2484
0 369 7 2 2 2482 368
0 370 5 1 1 2487
0 371 7 1 2 2225 370
0 372 5 2 1 371
0 373 7 1 2 2146 2488
0 374 5 1 1 373
0 375 7 2 2 2489 374
0 376 5 1 1 2491
0 377 7 2 2 2222 2492
0 378 5 2 1 2493
0 379 7 1 2 352 2490
0 380 5 1 1 379
0 381 7 1 2 2477 2485
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 2497
0 385 7 1 2 2495 384
0 386 5 2 1 385
0 387 7 1 2 2479 2486
0 388 5 1 1 387
0 389 7 1 2 2481 388
0 390 5 1 1 389
0 391 7 3 2 2483 390
0 392 5 1 1 2501
0 393 7 2 2 2499 392
0 394 5 1 1 2504
0 395 7 1 2 2223 394
0 396 5 2 1 395
0 397 7 1 2 2136 2505
0 398 5 1 1 397
0 399 7 2 2 2506 398
0 400 5 1 1 2508
0 401 7 2 2 2220 2509
0 402 5 2 1 2510
0 403 7 1 2 376 2507
0 404 5 1 1 403
0 405 7 1 2 2494 2502
0 406 5 1 1 405
0 407 7 2 2 404 406
0 408 5 1 1 2514
0 409 7 1 2 2512 408
0 410 5 2 1 409
0 411 7 1 2 2496 2503
0 412 5 1 1 411
0 413 7 1 2 2498 412
0 414 5 1 1 413
0 415 7 3 2 2500 414
0 416 5 1 1 2518
0 417 7 2 2 2516 416
0 418 5 1 1 2521
0 419 7 1 2 2221 418
0 420 5 2 1 419
0 421 7 1 2 2126 2522
0 422 5 1 1 421
0 423 7 2 2 2523 422
0 424 5 1 1 2525
0 425 7 2 2 2218 2526
0 426 5 2 1 2527
0 427 7 1 2 400 2524
0 428 5 1 1 427
0 429 7 1 2 2511 2519
0 430 5 1 1 429
0 431 7 2 2 428 430
0 432 5 1 1 2531
0 433 7 1 2 2529 432
0 434 5 2 1 433
0 435 7 1 2 2513 2520
0 436 5 1 1 435
0 437 7 1 2 2515 436
0 438 5 1 1 437
0 439 7 3 2 2517 438
0 440 5 1 1 2535
0 441 7 2 2 2533 440
0 442 5 1 1 2538
0 443 7 1 2 2219 442
0 444 5 2 1 443
0 445 7 1 2 2116 2539
0 446 5 1 1 445
0 447 7 2 2 2540 446
0 448 5 1 1 2542
0 449 7 2 2 2216 2543
0 450 5 2 1 2544
0 451 7 1 2 424 2541
0 452 5 1 1 451
0 453 7 1 2 2528 2536
0 454 5 1 1 453
0 455 7 2 2 452 454
0 456 5 1 1 2548
0 457 7 1 2 2546 456
0 458 5 2 1 457
0 459 7 1 2 2530 2537
0 460 5 1 1 459
0 461 7 1 2 2532 460
0 462 5 1 1 461
0 463 7 3 2 2534 462
0 464 5 1 1 2552
0 465 7 2 2 2550 464
0 466 5 1 1 2555
0 467 7 1 2 2217 466
0 468 5 2 1 467
0 469 7 1 2 2106 2556
0 470 5 1 1 469
0 471 7 2 2 2557 470
0 472 5 1 1 2559
0 473 7 2 2 2214 2560
0 474 5 2 1 2561
0 475 7 1 2 448 2558
0 476 5 1 1 475
0 477 7 1 2 2545 2553
0 478 5 1 1 477
0 479 7 2 2 476 478
0 480 5 1 1 2565
0 481 7 1 2 2563 480
0 482 5 2 1 481
0 483 7 1 2 2547 2554
0 484 5 1 1 483
0 485 7 1 2 2549 484
0 486 5 1 1 485
0 487 7 3 2 2551 486
0 488 5 1 1 2569
0 489 7 2 2 2567 488
0 490 5 1 1 2572
0 491 7 1 2 2215 490
0 492 5 2 1 491
0 493 7 1 2 2096 2573
0 494 5 1 1 493
0 495 7 2 2 2574 494
0 496 5 1 1 2576
0 497 7 2 2 2212 2577
0 498 5 2 1 2578
0 499 7 1 2 472 2575
0 500 5 1 1 499
0 501 7 1 2 2562 2570
0 502 5 1 1 501
0 503 7 2 2 500 502
0 504 5 1 1 2582
0 505 7 1 2 2580 504
0 506 5 2 1 505
0 507 7 1 2 2564 2571
0 508 5 1 1 507
0 509 7 1 2 2566 508
0 510 5 1 1 509
0 511 7 3 2 2568 510
0 512 5 1 1 2586
0 513 7 2 2 2584 512
0 514 5 1 1 2589
0 515 7 1 2 2213 514
0 516 5 2 1 515
0 517 7 1 2 2085 2590
0 518 5 1 1 517
0 519 7 2 2 2591 518
0 520 5 1 1 2593
0 521 7 2 2 2210 2594
0 522 5 2 1 2595
0 523 7 1 2 496 2592
0 524 5 1 1 523
0 525 7 1 2 2579 2587
0 526 5 1 1 525
0 527 7 2 2 524 526
0 528 5 1 1 2599
0 529 7 1 2 2597 528
0 530 5 2 1 529
0 531 7 1 2 2581 2588
0 532 5 1 1 531
0 533 7 1 2 2583 532
0 534 5 1 1 533
0 535 7 3 2 2585 534
0 536 5 1 1 2603
0 537 7 2 2 2601 536
0 538 5 1 1 2606
0 539 7 1 2 2211 538
0 540 5 2 1 539
0 541 7 1 2 2075 2607
0 542 5 1 1 541
0 543 7 2 2 2608 542
0 544 5 1 1 2610
0 545 7 2 2 2208 2611
0 546 5 2 1 2612
0 547 7 1 2 520 2609
0 548 5 1 1 547
0 549 7 1 2 2596 2604
0 550 5 1 1 549
0 551 7 2 2 548 550
0 552 5 1 1 2616
0 553 7 1 2 2614 552
0 554 5 2 1 553
0 555 7 1 2 2598 2605
0 556 5 1 1 555
0 557 7 1 2 2600 556
0 558 5 1 1 557
0 559 7 3 2 2602 558
0 560 5 1 1 2620
0 561 7 2 2 2618 560
0 562 5 1 1 2623
0 563 7 1 2 2209 562
0 564 5 2 1 563
0 565 7 1 2 2065 2624
0 566 5 1 1 565
0 567 7 2 2 2625 566
0 568 5 1 1 2627
0 569 7 2 2 2206 2628
0 570 5 2 1 2629
0 571 7 1 2 544 2626
0 572 5 1 1 571
0 573 7 1 2 2613 2621
0 574 5 1 1 573
0 575 7 2 2 572 574
0 576 5 1 1 2633
0 577 7 1 2 2631 576
0 578 5 2 1 577
0 579 7 1 2 2615 2622
0 580 5 1 1 579
0 581 7 1 2 2617 580
0 582 5 1 1 581
0 583 7 3 2 2619 582
0 584 5 1 1 2637
0 585 7 2 2 2635 584
0 586 5 1 1 2640
0 587 7 1 2 2207 586
0 588 5 2 1 587
0 589 7 1 2 2055 2641
0 590 5 1 1 589
0 591 7 2 2 2642 590
0 592 5 1 1 2644
0 593 7 2 2 2204 2645
0 594 5 2 1 2646
0 595 7 1 2 568 2643
0 596 5 1 1 595
0 597 7 1 2 2630 2638
0 598 5 1 1 597
0 599 7 2 2 596 598
0 600 5 1 1 2650
0 601 7 1 2 2648 600
0 602 5 2 1 601
0 603 7 1 2 2632 2639
0 604 5 1 1 603
0 605 7 1 2 2634 604
0 606 5 1 1 605
0 607 7 3 2 2636 606
0 608 5 1 1 2654
0 609 7 2 2 2652 608
0 610 5 1 1 2657
0 611 7 1 2 2205 610
0 612 5 2 1 611
0 613 7 1 2 2045 2658
0 614 5 1 1 613
0 615 7 2 2 2659 614
0 616 5 1 1 2661
0 617 7 2 2 2202 2662
0 618 5 2 1 2663
0 619 7 1 2 592 2660
0 620 5 1 1 619
0 621 7 1 2 2647 2655
0 622 5 1 1 621
0 623 7 2 2 620 622
0 624 5 1 1 2667
0 625 7 1 2 2665 624
0 626 5 2 1 625
0 627 7 1 2 2649 2656
0 628 5 1 1 627
0 629 7 1 2 2651 628
0 630 5 1 1 629
0 631 7 3 2 2653 630
0 632 5 1 1 2671
0 633 7 2 2 2669 632
0 634 5 1 1 2674
0 635 7 1 2 2203 634
0 636 5 2 1 635
0 637 7 1 2 2034 2675
0 638 5 1 1 637
0 639 7 2 2 2676 638
0 640 5 1 1 2678
0 641 7 2 2 2200 2679
0 642 5 2 1 2680
0 643 7 1 2 616 2677
0 644 5 1 1 643
0 645 7 1 2 2664 2672
0 646 5 1 1 645
0 647 7 2 2 644 646
0 648 5 1 1 2684
0 649 7 1 2 2682 648
0 650 5 2 1 649
0 651 7 1 2 2666 2673
0 652 5 1 1 651
0 653 7 1 2 2668 652
0 654 5 1 1 653
0 655 7 3 2 2670 654
0 656 5 1 1 2688
0 657 7 2 2 2686 656
0 658 5 1 1 2691
0 659 7 1 2 2201 658
0 660 5 2 1 659
0 661 7 1 2 2024 2692
0 662 5 1 1 661
0 663 7 2 2 2693 662
0 664 5 1 1 2695
0 665 7 2 2 2198 2696
0 666 5 2 1 2697
0 667 7 1 2 640 2694
0 668 5 1 1 667
0 669 7 1 2 2681 2689
0 670 5 1 1 669
0 671 7 2 2 668 670
0 672 5 1 1 2701
0 673 7 1 2 2699 672
0 674 5 2 1 673
0 675 7 1 2 2683 2690
0 676 5 1 1 675
0 677 7 1 2 2685 676
0 678 5 1 1 677
0 679 7 3 2 2687 678
0 680 5 1 1 2705
0 681 7 2 2 2703 680
0 682 5 1 1 2708
0 683 7 1 2 2013 2709
0 684 5 1 1 683
0 685 7 1 2 2199 682
0 686 5 2 1 685
0 687 7 2 2 684 2710
0 688 5 1 1 2712
0 689 7 2 2 2196 2713
0 690 5 2 1 2714
0 691 7 1 2 664 2711
0 692 5 1 1 691
0 693 7 1 2 2698 2706
0 694 5 1 1 693
0 695 7 2 2 692 694
0 696 5 1 1 2718
0 697 7 1 2 2716 696
0 698 5 2 1 697
0 699 7 1 2 2700 2707
0 700 5 1 1 699
0 701 7 1 2 2702 700
0 702 5 1 1 701
0 703 7 3 2 2704 702
0 704 5 1 1 2722
0 705 7 1 2 2717 2723
0 706 5 1 1 705
0 707 7 1 2 2719 706
0 708 5 1 1 707
0 709 7 1 2 2720 708
0 710 5 1 1 709
0 711 7 2 2 2721 704
0 712 5 1 1 2725
0 713 7 1 2 2197 712
0 714 5 2 1 713
0 715 7 1 2 2003 2726
0 716 5 1 1 715
0 717 7 2 2 2727 716
0 718 5 1 1 2729
0 719 7 1 2 1993 718
0 720 5 1 1 719
0 721 7 1 2 710 720
0 722 5 1 1 721
0 723 7 1 2 688 2728
0 724 5 1 1 723
0 725 7 1 2 2715 2724
0 726 5 1 1 725
0 727 7 2 2 724 726
0 728 5 1 1 2731
0 729 7 1 2 722 2732
0 730 5 1 1 729
0 731 7 1 2 33 2730
0 732 7 1 2 728 731
0 733 5 1 1 732
0 734 7 2 2 730 733
0 735 5 1 1 2733
0 736 7 2 2 2056 2137
0 737 5 1 1 2735
0 738 7 2 2 2046 2127
0 739 5 2 1 2737
0 740 7 2 2 2057 2117
0 741 5 1 1 2741
0 742 7 2 2 2035 2138
0 743 5 1 1 2743
0 744 7 1 2 2742 2744
0 745 5 2 1 744
0 746 7 1 2 741 743
0 747 5 1 1 746
0 748 7 2 2 747 2745
0 749 5 1 1 2747
0 750 7 1 2 2738 2748
0 751 5 2 1 750
0 752 7 2 2 2746 2749
0 753 5 1 1 2751
0 754 7 2 2 2047 2139
0 755 5 1 1 2753
0 756 7 2 2 2058 2128
0 757 5 1 1 2755
0 758 7 1 2 755 2756
0 759 5 1 1 758
0 760 7 1 2 2754 757
0 761 5 1 1 760
0 762 7 2 2 759 761
0 763 5 1 1 2757
0 764 7 1 2 753 763
0 765 5 3 1 764
0 766 7 1 2 2739 2759
0 767 5 1 1 766
0 768 7 1 2 2736 767
0 769 5 2 1 768
0 770 7 2 2 2025 2140
0 771 5 1 1 2764
0 772 7 2 2 2059 2107
0 773 5 1 1 2766
0 774 7 1 2 2765 2767
0 775 5 2 1 774
0 776 7 2 2 2048 2118
0 777 5 1 1 2770
0 778 7 1 2 771 773
0 779 5 1 1 778
0 780 7 2 2 2768 779
0 781 5 1 1 2772
0 782 7 1 2 2771 2773
0 783 5 2 1 782
0 784 7 2 2 2769 2774
0 785 5 1 1 2776
0 786 7 1 2 2740 749
0 787 5 1 1 786
0 788 7 2 2 2750 787
0 789 5 1 1 2778
0 790 7 1 2 785 2779
0 791 5 2 1 790
0 792 7 2 2 2036 2129
0 793 5 1 1 2782
0 794 7 1 2 777 781
0 795 5 1 1 794
0 796 7 2 2 2775 795
0 797 5 1 1 2784
0 798 7 1 2 2783 2785
0 799 5 2 1 798
0 800 7 2 2 2014 2141
0 801 5 1 1 2788
0 802 7 2 2 2060 2097
0 803 5 1 1 2790
0 804 7 1 2 2789 2791
0 805 5 2 1 804
0 806 7 2 2 2049 2108
0 807 5 1 1 2794
0 808 7 1 2 801 803
0 809 5 1 1 808
0 810 7 2 2 2792 809
0 811 5 1 1 2796
0 812 7 1 2 2795 2797
0 813 5 2 1 812
0 814 7 2 2 2793 2798
0 815 5 1 1 2800
0 816 7 1 2 793 797
0 817 5 1 1 816
0 818 7 2 2 2786 817
0 819 5 1 1 2802
0 820 7 1 2 815 2803
0 821 5 2 1 820
0 822 7 2 2 2787 2804
0 823 5 1 1 2806
0 824 7 1 2 2777 789
0 825 5 1 1 824
0 826 7 2 2 2780 825
0 827 5 1 1 2808
0 828 7 1 2 823 2809
0 829 5 2 1 828
0 830 7 2 2 2781 2810
0 831 5 1 1 2812
0 832 7 1 2 2752 2758
0 833 5 1 1 832
0 834 7 2 2 2760 833
0 835 5 1 1 2814
0 836 7 1 2 831 2815
0 837 5 2 1 836
0 838 7 2 2 2026 2130
0 839 5 1 1 2818
0 840 7 1 2 807 811
0 841 5 1 1 840
0 842 7 2 2 2799 841
0 843 5 1 1 2820
0 844 7 1 2 2819 2821
0 845 5 2 1 844
0 846 7 2 2 2037 2119
0 847 5 1 1 2824
0 848 7 1 2 839 843
0 849 5 1 1 848
0 850 7 2 2 2822 849
0 851 5 1 1 2826
0 852 7 1 2 2825 2827
0 853 5 2 1 852
0 854 7 2 2 2823 2828
0 855 5 1 1 2830
0 856 7 1 2 2801 819
0 857 5 1 1 856
0 858 7 2 2 2805 857
0 859 5 1 1 2832
0 860 7 1 2 855 2833
0 861 5 2 1 860
0 862 7 2 2 2061 2066
0 863 5 1 1 2836
0 864 7 2 2 2050 2076
0 865 5 1 1 2838
0 866 7 2 2 2837 2839
0 867 5 2 1 2840
0 868 7 2 2 2086 2841
0 869 5 2 1 2844
0 870 7 2 2 2004 2142
0 871 5 1 1 2848
0 872 7 1 2 2845 2849
0 873 5 2 1 872
0 874 7 2 2 2062 2087
0 875 5 1 1 2852
0 876 7 1 2 2846 871
0 877 5 1 1 876
0 878 7 2 2 2850 877
0 879 5 1 1 2854
0 880 7 1 2 2853 2855
0 881 5 2 1 880
0 882 7 2 2 2851 2856
0 883 5 1 1 2858
0 884 7 1 2 847 851
0 885 5 1 1 884
0 886 7 2 2 2829 885
0 887 5 1 1 2860
0 888 7 1 2 883 2861
0 889 5 2 1 888
0 890 7 2 2 2038 2109
0 891 5 1 1 2864
0 892 7 1 2 875 879
0 893 5 1 1 892
0 894 7 2 2 2857 893
0 895 5 1 1 2866
0 896 7 1 2 2865 2867
0 897 5 2 1 896
0 898 7 2 2 2051 2098
0 899 5 1 1 2870
0 900 7 1 2 891 895
0 901 5 1 1 900
0 902 7 2 2 2868 901
0 903 5 1 1 2872
0 904 7 1 2 2871 2873
0 905 5 2 1 904
0 906 7 2 2 2869 2874
0 907 5 1 1 2876
0 908 7 1 2 2859 887
0 909 5 1 1 908
0 910 7 2 2 2862 909
0 911 5 1 1 2878
0 912 7 1 2 907 2879
0 913 5 2 1 912
0 914 7 2 2 2863 2880
0 915 5 1 1 2882
0 916 7 1 2 2831 859
0 917 5 1 1 916
0 918 7 2 2 2834 917
0 919 5 1 1 2884
0 920 7 1 2 915 2885
0 921 5 2 1 920
0 922 7 2 2 2835 2886
0 923 5 1 1 2888
0 924 7 1 2 2807 827
0 925 5 1 1 924
0 926 7 2 2 2811 925
0 927 5 1 1 2890
0 928 7 1 2 923 2891
0 929 5 2 1 928
0 930 7 2 2 2015 2131
0 931 5 1 1 2894
0 932 7 2 2 2027 2120
0 933 5 1 1 2896
0 934 7 1 2 2895 2897
0 935 5 2 1 934
0 936 7 1 2 899 903
0 937 5 1 1 936
0 938 7 2 2 2875 937
0 939 5 1 1 2900
0 940 7 1 2 931 933
0 941 5 1 1 940
0 942 7 2 2 2898 941
0 943 5 1 1 2902
0 944 7 1 2 2901 2903
0 945 5 2 1 944
0 946 7 2 2 2899 2904
0 947 5 1 1 2906
0 948 7 1 2 2877 911
0 949 5 1 1 948
0 950 7 2 2 2881 949
0 951 5 1 1 2908
0 952 7 1 2 947 2909
0 953 5 2 1 952
0 954 7 2 2 2039 2099
0 955 5 1 1 2912
0 956 7 2 2 2005 2132
0 957 5 1 1 2914
0 958 7 1 2 2913 2915
0 959 5 2 1 958
0 960 7 2 2 1994 2143
0 961 5 1 1 2918
0 962 7 2 2 2028 2110
0 963 5 1 1 2920
0 964 7 1 2 2052 2088
0 965 5 1 1 964
0 966 7 1 2 2842 965
0 967 5 1 1 966
0 968 7 2 2 2847 967
0 969 5 1 1 2922
0 970 7 1 2 2921 2923
0 971 5 2 1 970
0 972 7 1 2 963 969
0 973 5 1 1 972
0 974 7 2 2 2924 973
0 975 5 1 1 2926
0 976 7 1 2 2919 2927
0 977 5 2 1 976
0 978 7 1 2 961 975
0 979 5 1 1 978
0 980 7 2 2 2928 979
0 981 5 1 1 2930
0 982 7 1 2 955 957
0 983 5 1 1 982
0 984 7 2 2 2916 983
0 985 5 1 1 2932
0 986 7 1 2 2931 2933
0 987 5 2 1 986
0 988 7 2 2 2917 2934
0 989 5 1 1 2936
0 990 7 1 2 939 943
0 991 5 1 1 990
0 992 7 2 2 2905 991
0 993 5 1 1 2938
0 994 7 1 2 989 2939
0 995 5 2 1 994
0 996 7 2 2 2063 2077
0 997 5 1 1 2942
0 998 7 2 2 2016 2121
0 999 5 1 1 2944
0 1000 7 1 2 2943 2945
0 1001 5 2 1 1000
0 1002 7 1 2 981 985
0 1003 5 1 1 1002
0 1004 7 2 2 2935 1003
0 1005 5 1 1 2948
0 1006 7 1 2 997 999
0 1007 5 1 1 1006
0 1008 7 2 2 2946 1007
0 1009 5 1 1 2950
0 1010 7 1 2 2949 2951
0 1011 5 2 1 1010
0 1012 7 2 2 2947 2952
0 1013 5 1 1 2954
0 1014 7 1 2 2937 993
0 1015 5 1 1 1014
0 1016 7 2 2 2940 1015
0 1017 5 1 1 2956
0 1018 7 1 2 1013 2957
0 1019 5 2 1 1018
0 1020 7 2 2 2941 2958
0 1021 5 1 1 2960
0 1022 7 1 2 2907 951
0 1023 5 1 1 1022
0 1024 7 2 2 2910 1023
0 1025 5 1 1 2962
0 1026 7 1 2 1021 2963
0 1027 5 2 1 1026
0 1028 7 2 2 2911 2964
0 1029 5 1 1 2966
0 1030 7 1 2 2883 919
0 1031 5 1 1 1030
0 1032 7 2 2 2887 1031
0 1033 5 1 1 2968
0 1034 7 1 2 1029 2969
0 1035 5 2 1 1034
0 1036 7 2 2 2925 2929
0 1037 5 1 1 2972
0 1038 7 1 2 2955 1017
0 1039 5 1 1 1038
0 1040 7 2 2 2959 1039
0 1041 5 1 1 2974
0 1042 7 1 2 1037 2975
0 1043 5 2 1 1042
0 1044 7 2 2 2040 2089
0 1045 5 1 1 2978
0 1046 7 2 2 2029 2100
0 1047 5 1 1 2980
0 1048 7 1 2 2979 2981
0 1049 5 2 1 1048
0 1050 7 2 2 1995 2133
0 1051 5 1 1 2984
0 1052 7 1 2 1045 1047
0 1053 5 1 1 1052
0 1054 7 2 2 2982 1053
0 1055 5 1 1 2986
0 1056 7 1 2 2985 2987
0 1057 5 2 1 1056
0 1058 7 2 2 2983 2988
0 1059 5 1 1 2990
0 1060 7 2 2 2006 2122
0 1061 5 1 1 2992
0 1062 7 2 2 32 2144
0 1063 5 1 1 2994
0 1064 7 1 2 2993 2995
0 1065 5 2 1 1064
0 1066 7 2 2 2017 2111
0 1067 5 1 1 2998
0 1068 7 2 2 2030 2078
0 1069 5 1 1 3000
0 1070 7 2 2 1985 2101
0 1071 5 1 1 3002
0 1072 7 2 2 2007 2079
0 1073 5 1 1 3004
0 1074 7 2 2 3003 3005
0 1075 5 2 1 3006
0 1076 7 2 2 2018 3007
0 1077 5 2 1 3010
0 1078 7 2 2 3001 3011
0 1079 5 2 1 3014
0 1080 7 2 2 2041 3015
0 1081 5 2 1 3018
0 1082 7 1 2 2999 3019
0 1083 5 2 1 1082
0 1084 7 1 2 1067 3020
0 1085 5 1 1 1084
0 1086 7 2 2 3022 1085
0 1087 5 1 1 3024
0 1088 7 1 2 863 865
0 1089 5 1 1 1088
0 1090 7 2 2 2843 1089
0 1091 5 1 1 3026
0 1092 7 1 2 3025 3027
0 1093 5 2 1 1092
0 1094 7 1 2 1087 1091
0 1095 5 1 1 1094
0 1096 7 2 2 3028 1095
0 1097 5 1 1 3030
0 1098 7 1 2 1061 1063
0 1099 5 1 1 1098
0 1100 7 2 2 2996 1099
0 1101 5 1 1 3032
0 1102 7 1 2 3031 3033
0 1103 5 2 1 1102
0 1104 7 2 2 2997 3034
0 1105 5 1 1 3036
0 1106 7 1 2 1059 1105
0 1107 5 2 1 1106
0 1108 7 2 2 3023 3029
0 1109 5 1 1 3040
0 1110 7 1 2 2991 3037
0 1111 5 1 1 1110
0 1112 7 2 2 3038 1111
0 1113 5 1 1 3042
0 1114 7 1 2 1109 3043
0 1115 5 2 1 1114
0 1116 7 2 2 3039 3044
0 1117 5 1 1 3046
0 1118 7 1 2 2973 1041
0 1119 5 1 1 1118
0 1120 7 2 2 2976 1119
0 1121 5 1 1 3048
0 1122 7 1 2 1117 3049
0 1123 5 2 1 1122
0 1124 7 2 2 2977 3050
0 1125 5 1 1 3052
0 1126 7 1 2 2961 1025
0 1127 5 1 1 1126
0 1128 7 2 2 2965 1127
0 1129 5 1 1 3054
0 1130 7 1 2 1125 3055
0 1131 5 2 1 1130
0 1132 7 1 2 1005 1009
0 1133 5 1 1 1132
0 1134 7 2 2 2953 1133
0 1135 5 1 1 3058
0 1136 7 1 2 3041 1113
0 1137 5 1 1 1136
0 1138 7 2 2 3045 1137
0 1139 5 1 1 3060
0 1140 7 1 2 3059 3061
0 1141 5 2 1 1140
0 1142 7 1 2 1051 1055
0 1143 5 1 1 1142
0 1144 7 2 2 2989 1143
0 1145 5 1 1 3064
0 1146 7 1 2 1097 1101
0 1147 5 1 1 1146
0 1148 7 2 2 3035 1147
0 1149 5 1 1 3066
0 1150 7 1 2 3065 3067
0 1151 5 2 1 1150
0 1152 7 2 2 2019 2102
0 1153 5 1 1 3070
0 1154 7 2 2 2008 2112
0 1155 5 1 1 3072
0 1156 7 1 2 3071 3073
0 1157 5 2 1 1156
0 1158 7 2 2 1996 2123
0 1159 5 1 1 3076
0 1160 7 1 2 1153 1155
0 1161 5 1 1 1160
0 1162 7 2 2 3074 1161
0 1163 5 1 1 3078
0 1164 7 1 2 3077 3079
0 1165 5 2 1 1164
0 1166 7 2 2 3075 3080
0 1167 5 1 1 3082
0 1168 7 1 2 1145 1149
0 1169 5 1 1 1168
0 1170 7 2 2 3068 1169
0 1171 5 1 1 3084
0 1172 7 1 2 1167 3085
0 1173 5 2 1 1172
0 1174 7 2 2 3069 3086
0 1175 5 1 1 3088
0 1176 7 1 2 1135 1139
0 1177 5 1 1 1176
0 1178 7 2 2 3062 1177
0 1179 5 1 1 3090
0 1180 7 1 2 1175 3091
0 1181 5 2 1 1180
0 1182 7 2 2 3063 3092
0 1183 5 1 1 3094
0 1184 7 1 2 3047 1121
0 1185 5 1 1 1184
0 1186 7 2 2 3051 1185
0 1187 5 1 1 3096
0 1188 7 1 2 1183 3097
0 1189 5 2 1 1188
0 1190 7 2 2 1986 2134
0 1191 5 1 1 3100
0 1192 7 1 2 1159 1163
0 1193 5 1 1 1192
0 1194 7 2 2 3081 1193
0 1195 5 1 1 3102
0 1196 7 1 2 3101 3103
0 1197 5 2 1 1196
0 1198 7 2 2 2053 2067
0 1199 5 1 1 3106
0 1200 7 2 2 2031 2090
0 1201 5 1 1 3108
0 1202 7 1 2 2042 2080
0 1203 5 1 1 1202
0 1204 7 1 2 3016 1203
0 1205 5 1 1 1204
0 1206 7 2 2 3021 1205
0 1207 5 1 1 3110
0 1208 7 1 2 3109 3111
0 1209 5 2 1 1208
0 1210 7 1 2 1201 1207
0 1211 5 1 1 1210
0 1212 7 2 2 3112 1211
0 1213 5 1 1 3114
0 1214 7 1 2 3107 3115
0 1215 5 2 1 1214
0 1216 7 1 2 1199 1213
0 1217 5 1 1 1216
0 1218 7 2 2 3116 1217
0 1219 5 1 1 3118
0 1220 7 1 2 1191 1195
0 1221 5 1 1 1220
0 1222 7 2 2 3104 1221
0 1223 5 1 1 3120
0 1224 7 1 2 3119 3121
0 1225 5 2 1 1224
0 1226 7 2 2 3105 3122
0 1227 5 1 1 3124
0 1228 7 1 2 3083 1171
0 1229 5 1 1 1228
0 1230 7 2 2 3087 1229
0 1231 5 1 1 3126
0 1232 7 1 2 1227 3127
0 1233 5 2 1 1232
0 1234 7 2 2 3113 3117
0 1235 5 1 1 3130
0 1236 7 1 2 3125 1231
0 1237 5 1 1 1236
0 1238 7 2 2 3128 1237
0 1239 5 1 1 3132
0 1240 7 1 2 1235 3133
0 1241 5 2 1 1240
0 1242 7 2 2 3129 3134
0 1243 5 1 1 3136
0 1244 7 1 2 3089 1179
0 1245 5 1 1 1244
0 1246 7 2 2 3093 1245
0 1247 5 1 1 3138
0 1248 7 1 2 1243 3139
0 1249 5 2 1 1248
0 1250 7 2 2 2020 2091
0 1251 5 1 1 3142
0 1252 7 1 2 1069 3012
0 1253 5 1 1 1252
0 1254 7 2 2 3017 1253
0 1255 5 1 1 3144
0 1256 7 1 2 3143 3145
0 1257 5 2 1 1256
0 1258 7 2 2 2043 2068
0 1259 5 1 1 3148
0 1260 7 1 2 1251 1255
0 1261 5 1 1 1260
0 1262 7 2 2 3146 1261
0 1263 5 1 1 3150
0 1264 7 1 2 3149 3151
0 1265 5 2 1 1264
0 1266 7 2 2 3147 3152
0 1267 5 1 1 3154
0 1268 7 1 2 1219 1223
0 1269 5 1 1 1268
0 1270 7 2 2 3123 1269
0 1271 5 1 1 3156
0 1272 7 1 2 1267 3157
0 1273 5 2 1 1272
0 1274 7 2 2 2009 2103
0 1275 5 1 1 3160
0 1276 7 2 2 1987 2124
0 1277 5 1 1 3162
0 1278 7 1 2 3161 3163
0 1279 5 2 1 1278
0 1280 7 1 2 1259 1263
0 1281 5 1 1 1280
0 1282 7 2 2 3153 1281
0 1283 5 1 1 3166
0 1284 7 1 2 1275 1277
0 1285 5 1 1 1284
0 1286 7 2 2 3164 1285
0 1287 5 1 1 3168
0 1288 7 1 2 3167 3169
0 1289 5 2 1 1288
0 1290 7 2 2 3165 3170
0 1291 5 1 1 3172
0 1292 7 1 2 3155 1271
0 1293 5 1 1 1292
0 1294 7 2 2 3158 1293
0 1295 5 1 1 3174
0 1296 7 1 2 1291 3175
0 1297 5 2 1 1296
0 1298 7 2 2 3159 3176
0 1299 5 1 1 3178
0 1300 7 1 2 3131 1239
0 1301 5 1 1 1300
0 1302 7 2 2 3135 1301
0 1303 5 1 1 3180
0 1304 7 1 2 1299 3181
0 1305 5 2 1 1304
0 1306 7 2 2 1997 2113
0 1307 5 1 1 3184
0 1308 7 1 2 1283 1287
0 1309 5 1 1 1308
0 1310 7 2 2 3171 1309
0 1311 5 1 1 3186
0 1312 7 1 2 3185 3187
0 1313 5 2 1 1312
0 1314 7 2 2 2010 2092
0 1315 5 1 1 3190
0 1316 7 1 2 2021 2081
0 1317 5 1 1 1316
0 1318 7 1 2 3008 1317
0 1319 5 1 1 1318
0 1320 7 2 2 3013 1319
0 1321 5 1 1 3192
0 1322 7 1 2 3191 3193
0 1323 5 2 1 1322
0 1324 7 2 2 2032 2069
0 1325 5 1 1 3196
0 1326 7 1 2 1315 1321
0 1327 5 1 1 1326
0 1328 7 2 2 3194 1327
0 1329 5 1 1 3198
0 1330 7 1 2 3197 3199
0 1331 5 2 1 1330
0 1332 7 2 2 3195 3200
0 1333 5 1 1 3202
0 1334 7 1 2 1307 1311
0 1335 5 1 1 1334
0 1336 7 2 2 3188 1335
0 1337 5 1 1 3204
0 1338 7 1 2 1333 3205
0 1339 5 2 1 1338
0 1340 7 2 2 3189 3206
0 1341 5 1 1 3208
0 1342 7 1 2 3173 1295
0 1343 5 1 1 1342
0 1344 7 2 2 3177 1343
0 1345 5 1 1 3210
0 1346 7 1 2 1341 3211
0 1347 5 2 1 1346
0 1348 7 2 2 1988 2114
0 1349 5 1 1 3214
0 1350 7 2 2 1998 2104
0 1351 5 1 1 3216
0 1352 7 1 2 3215 3217
0 1353 5 2 1 1352
0 1354 7 1 2 1325 1329
0 1355 5 1 1 1354
0 1356 7 2 2 3201 1355
0 1357 5 1 1 3220
0 1358 7 1 2 1349 1351
0 1359 5 1 1 1358
0 1360 7 2 2 3218 1359
0 1361 5 1 1 3222
0 1362 7 1 2 3221 3223
0 1363 5 2 1 1362
0 1364 7 2 2 3219 3224
0 1365 5 1 1 3226
0 1366 7 1 2 3203 1337
0 1367 5 1 1 1366
0 1368 7 2 2 3207 1367
0 1369 5 1 1 3228
0 1370 7 1 2 1365 3229
0 1371 5 2 1 1370
0 1372 7 1 2 1357 1361
0 1373 5 1 1 1372
0 1374 7 2 2 3225 1373
0 1375 5 1 1 3232
0 1376 7 2 2 1999 2093
0 1377 5 1 1 3234
0 1378 7 2 2 2022 2070
0 1379 5 1 1 3236
0 1380 7 2 2 3235 3237
0 1381 5 1 1 3238
0 1382 7 2 2 2000 2082
0 1383 5 1 1 3240
0 1384 7 2 2 1989 2094
0 1385 5 1 1 3242
0 1386 7 2 2 3241 3243
0 1387 5 2 1 3244
0 1388 7 3 2 1381 3246
0 1389 5 1 1 3248
0 1390 7 1 2 3233 1389
0 1391 5 2 1 1390
0 1392 7 1 2 1071 1073
0 1393 5 1 1 1392
0 1394 7 2 2 3009 1393
0 1395 5 1 1 3253
0 1396 7 1 2 1377 1379
0 1397 5 1 1 1396
0 1398 7 1 2 3249 1397
0 1399 5 1 1 1398
0 1400 7 1 2 3239 3245
0 1401 5 1 1 1400
0 1402 7 2 2 1399 1401
0 1403 5 1 1 3255
0 1404 7 1 2 3254 1403
0 1405 5 2 1 1404
0 1406 7 2 2 2011 2071
0 1407 5 1 1 3259
0 1408 7 1 2 1383 1385
0 1409 5 1 1 1408
0 1410 7 2 2 3247 1409
0 1411 5 1 1 3261
0 1412 7 1 2 3260 3262
0 1413 5 2 1 1412
0 1414 7 1 2 1407 1411
0 1415 5 1 1 1414
0 1416 7 2 2 3263 1415
0 1417 5 1 1 3265
0 1418 7 2 2 1990 2083
0 1419 5 1 1 3267
0 1420 7 2 2 2001 2072
0 1421 5 1 1 3269
0 1422 7 2 2 3268 3270
0 1423 5 2 1 3271
0 1424 7 1 2 3266 3272
0 1425 5 2 1 1424
0 1426 7 2 2 3264 3275
0 1427 5 1 1 3277
0 1428 7 1 2 1395 3256
0 1429 5 1 1 1428
0 1430 7 2 2 3257 1429
0 1431 5 1 1 3279
0 1432 7 1 2 1427 3280
0 1433 5 2 1 1432
0 1434 7 2 2 3258 3281
0 1435 5 1 1 3283
0 1436 7 1 2 1375 3250
0 1437 5 1 1 1436
0 1438 7 2 2 3251 1437
0 1439 5 1 1 3285
0 1440 7 1 2 1435 3286
0 1441 5 2 1 1440
0 1442 7 2 2 3252 3287
0 1443 5 1 1 3289
0 1444 7 1 2 3227 1369
0 1445 5 1 1 1444
0 1446 7 2 2 3230 1445
0 1447 5 1 1 3291
0 1448 7 1 2 1443 3292
0 1449 5 2 1 1448
0 1450 7 2 2 3231 3293
0 1451 5 1 1 3295
0 1452 7 1 2 3209 1345
0 1453 5 1 1 1452
0 1454 7 2 2 3212 1453
0 1455 5 1 1 3297
0 1456 7 1 2 1451 3298
0 1457 5 2 1 1456
0 1458 7 2 2 3213 3299
0 1459 5 1 1 3301
0 1460 7 1 2 3179 1303
0 1461 5 1 1 1460
0 1462 7 2 2 3182 1461
0 1463 5 1 1 3303
0 1464 7 1 2 1459 3304
0 1465 5 2 1 1464
0 1466 7 2 2 3183 3305
0 1467 5 1 1 3307
0 1468 7 1 2 3137 1247
0 1469 5 1 1 1468
0 1470 7 2 2 3140 1469
0 1471 5 1 1 3309
0 1472 7 1 2 1467 3310
0 1473 5 2 1 1472
0 1474 7 2 2 3141 3311
0 1475 5 1 1 3313
0 1476 7 1 2 3095 1187
0 1477 5 1 1 1476
0 1478 7 2 2 3098 1477
0 1479 5 1 1 3315
0 1480 7 1 2 1475 3316
0 1481 5 2 1 1480
0 1482 7 2 2 3099 3317
0 1483 5 1 1 3319
0 1484 7 1 2 3053 1129
0 1485 5 1 1 1484
0 1486 7 2 2 3056 1485
0 1487 5 1 1 3321
0 1488 7 1 2 1483 3322
0 1489 5 2 1 1488
0 1490 7 2 2 3057 3323
0 1491 5 1 1 3325
0 1492 7 1 2 2967 1033
0 1493 5 1 1 1492
0 1494 7 2 2 2970 1493
0 1495 5 1 1 3327
0 1496 7 1 2 1491 3328
0 1497 5 2 1 1496
0 1498 7 2 2 2971 3329
0 1499 5 1 1 3331
0 1500 7 1 2 2889 927
0 1501 5 1 1 1500
0 1502 7 2 2 2892 1501
0 1503 5 1 1 3333
0 1504 7 1 2 1499 3334
0 1505 5 2 1 1504
0 1506 7 2 2 2893 3335
0 1507 5 1 1 3337
0 1508 7 1 2 2813 835
0 1509 5 1 1 1508
0 1510 7 2 2 2816 1509
0 1511 5 1 1 3339
0 1512 7 1 2 1507 3340
0 1513 5 2 1 1512
0 1514 7 2 2 2817 3341
0 1515 5 1 1 3343
0 1516 7 1 2 2761 737
0 1517 5 1 1 1516
0 1518 7 2 2 2762 1517
0 1519 5 1 1 3345
0 1520 7 1 2 1515 3346
0 1521 5 2 1 1520
0 1522 7 2 2 2763 3347
0 1523 5 1 1 3349
0 1524 7 2 2 2270 1523
0 1525 5 3 1 3351
0 1526 7 1 2 3344 1519
0 1527 5 1 1 1526
0 1528 7 2 2 3348 1527
0 1529 5 1 1 3356
0 1530 7 2 2 2191 1529
0 1531 5 3 1 3358
0 1532 7 2 2 2195 3350
0 1533 5 2 1 3363
0 1534 7 2 2 3360 3365
0 1535 7 1 2 3338 1511
0 1536 5 1 1 1535
0 1537 7 2 2 3342 1536
0 1538 5 1 1 3369
0 1539 7 1 2 2187 1538
0 1540 5 3 1 1539
0 1541 7 1 2 2266 3370
0 1542 5 4 1 1541
0 1543 7 1 2 3332 1503
0 1544 5 1 1 1543
0 1545 7 2 2 3336 1544
0 1546 5 1 1 3378
0 1547 7 1 2 2184 1546
0 1548 5 4 1 1547
0 1549 7 1 2 2263 3379
0 1550 5 2 1 1549
0 1551 7 1 2 3326 1495
0 1552 5 1 1 1551
0 1553 7 2 2 3330 1552
0 1554 5 1 1 3386
0 1555 7 1 2 2259 3387
0 1556 5 3 1 1555
0 1557 7 3 2 3384 3388
0 1558 7 2 2 2180 1554
0 1559 5 4 1 3394
0 1560 7 1 2 3320 1487
0 1561 5 1 1 1560
0 1562 7 2 2 3324 1561
0 1563 5 1 1 3400
0 1564 7 1 2 2177 1563
0 1565 5 3 1 1564
0 1566 7 1 2 2256 3401
0 1567 5 3 1 1566
0 1568 7 1 2 3314 1479
0 1569 5 1 1 1568
0 1570 7 2 2 3318 1569
0 1571 5 1 1 3408
0 1572 7 1 2 2253 3409
0 1573 5 3 1 1572
0 1574 7 2 2 3405 3410
0 1575 7 2 2 2174 1571
0 1576 5 4 1 3415
0 1577 7 1 2 3308 1471
0 1578 5 1 1 1577
0 1579 7 2 2 3312 1578
0 1580 5 1 1 3421
0 1581 7 1 2 2171 1580
0 1582 5 3 1 1581
0 1583 7 1 2 2250 3422
0 1584 5 4 1 1583
0 1585 7 1 2 3302 1463
0 1586 5 1 1 1585
0 1587 7 2 2 3306 1586
0 1588 5 1 1 3430
0 1589 7 1 2 2168 1588
0 1590 5 3 1 1589
0 1591 7 1 2 2247 3431
0 1592 5 4 1 1591
0 1593 7 1 2 3296 1455
0 1594 5 1 1 1593
0 1595 7 2 2 3300 1594
0 1596 5 1 1 3439
0 1597 7 1 2 2165 1596
0 1598 5 3 1 1597
0 1599 7 1 2 2244 3440
0 1600 5 4 1 1599
0 1601 7 1 2 3290 1447
0 1602 5 1 1 1601
0 1603 7 2 2 3294 1602
0 1604 5 1 1 3448
0 1605 7 1 2 2162 1604
0 1606 5 4 1 1605
0 1607 7 1 2 2241 3449
0 1608 5 4 1 1607
0 1609 7 1 2 3284 1439
0 1610 5 1 1 1609
0 1611 7 2 2 3288 1610
0 1612 5 1 1 3458
0 1613 7 1 2 2159 1612
0 1614 5 4 1 1613
0 1615 7 1 2 2238 3459
0 1616 5 4 1 1615
0 1617 7 1 2 3278 1431
0 1618 5 1 1 1617
0 1619 7 2 2 3282 1618
0 1620 5 1 1 3468
0 1621 7 1 2 2156 1620
0 1622 5 4 1 1621
0 1623 7 1 2 2235 3469
0 1624 5 3 1 1623
0 1625 7 1 2 1417 3273
0 1626 5 1 1 1625
0 1627 7 2 2 3276 1626
0 1628 5 1 1 3477
0 1629 7 1 2 2232 3478
0 1630 5 3 1 1629
0 1631 7 1 2 2153 1628
0 1632 5 4 1 1631
0 1633 7 1 2 1419 1421
0 1634 5 1 1 1633
0 1635 7 2 2 3274 1634
0 1636 5 1 1 3486
0 1637 7 1 2 2229 3487
0 1638 5 2 1 1637
0 1639 7 1 2 2150 1636
0 1640 5 2 1 1639
0 1641 7 2 2 1991 2073
0 1642 5 1 1 3492
0 1643 7 1 2 2147 1642
0 1644 5 1 1 1643
0 1645 7 2 2 3490 1644
0 1646 5 1 1 3494
0 1647 7 1 2 3488 1646
0 1648 5 3 1 1647
0 1649 7 1 2 3482 3496
0 1650 5 1 1 1649
0 1651 7 3 2 3479 1650
0 1652 5 1 1 3499
0 1653 7 1 2 3474 3500
0 1654 5 1 1 1653
0 1655 7 2 2 3470 1654
0 1656 5 1 1 3502
0 1657 7 2 2 3464 1656
0 1658 5 1 1 3504
0 1659 7 2 2 3460 1658
0 1660 5 2 1 3506
0 1661 7 1 2 3454 3508
0 1662 5 1 1 1661
0 1663 7 2 2 3450 1662
0 1664 5 2 1 3510
0 1665 7 1 2 3444 3512
0 1666 5 1 1 1665
0 1667 7 2 2 3441 1666
0 1668 5 2 1 3514
0 1669 7 1 2 3435 3516
0 1670 5 1 1 1669
0 1671 7 2 2 3432 1670
0 1672 5 2 1 3518
0 1673 7 1 2 3426 3520
0 1674 5 1 1 1673
0 1675 7 3 2 3423 1674
0 1676 5 1 1 3522
0 1677 7 1 2 3417 3523
0 1678 5 1 1 1677
0 1679 7 1 2 3413 1678
0 1680 5 1 1 1679
0 1681 7 3 2 3402 1680
0 1682 5 1 1 3525
0 1683 7 1 2 3396 3526
0 1684 5 1 1 1683
0 1685 7 1 2 3391 1684
0 1686 5 1 1 1685
0 1687 7 2 2 3380 1686
0 1688 5 2 1 3528
0 1689 7 1 2 3374 3530
0 1690 5 1 1 1689
0 1691 7 2 2 3371 1690
0 1692 5 2 1 3532
0 1693 7 1 2 2268 3357
0 1694 5 4 1 1693
0 1695 7 1 2 3534 3536
0 1696 5 1 1 1695
0 1697 7 1 2 3367 1696
0 1698 5 1 1 1697
0 1699 7 2 2 3353 1698
0 1700 5 2 1 3540
0 1701 7 1 2 2226 3493
0 1702 5 1 1 1701
0 1703 7 3 2 3489 1702
0 1704 5 2 1 3544
0 1705 7 2 2 3491 3547
0 1706 7 1 2 3483 3549
0 1707 5 1 1 1706
0 1708 7 2 2 3475 3480
0 1709 7 2 2 1707 3551
0 1710 5 1 1 3553
0 1711 7 2 2 3471 1710
0 1712 5 2 1 3555
0 1713 7 1 2 3465 3557
0 1714 5 1 1 1713
0 1715 7 2 2 3461 1714
0 1716 5 1 1 3559
0 1717 7 2 2 3455 1716
0 1718 5 1 1 3561
0 1719 7 2 2 3451 1718
0 1720 5 2 1 3563
0 1721 7 1 2 3445 3565
0 1722 5 1 1 1721
0 1723 7 2 2 3442 1722
0 1724 5 2 1 3567
0 1725 7 1 2 3436 3569
0 1726 5 1 1 1725
0 1727 7 2 2 3433 1726
0 1728 5 2 1 3571
0 1729 7 1 2 3427 3573
0 1730 5 1 1 1729
0 1731 7 2 2 3424 1730
0 1732 5 2 1 3575
0 1733 7 1 2 3411 3577
0 1734 5 1 1 1733
0 1735 7 2 2 3418 1734
0 1736 5 2 1 3579
0 1737 7 1 2 3406 3581
0 1738 5 1 1 1737
0 1739 7 3 2 3403 1738
0 1740 5 2 1 3583
0 1741 7 1 2 3397 3584
0 1742 5 1 1 1741
0 1743 7 2 2 3392 1742
0 1744 5 1 1 3588
0 1745 7 2 2 3381 1744
0 1746 5 2 1 3590
0 1747 7 3 2 3372 3375
0 1748 5 2 1 3594
0 1749 7 1 2 3591 3597
0 1750 5 1 1 1749
0 1751 7 1 2 3592 3595
0 1752 5 1 1 1751
0 1753 7 1 2 1750 1752
0 1754 5 1 1 1753
0 1755 7 1 2 3364 3537
0 1756 5 1 1 1755
0 1757 7 2 2 3382 3385
0 1758 5 1 1 3599
0 1759 7 2 2 3398 1758
0 1760 5 1 1 3601
0 1761 7 1 2 3389 3586
0 1762 5 1 1 1761
0 1763 7 1 2 3602 1762
0 1764 5 1 1 1763
0 1765 7 1 2 3383 3589
0 1766 5 1 1 1765
0 1767 7 1 2 1764 1766
0 1768 5 1 1 1767
0 1769 7 3 2 3390 3399
0 1770 5 2 1 3603
0 1771 7 1 2 3587 3604
0 1772 5 1 1 1771
0 1773 7 1 2 3585 3606
0 1774 5 1 1 1773
0 1775 7 1 2 1772 1774
0 1776 5 1 1 1775
0 1777 7 3 2 3404 3407
0 1778 5 2 1 3608
0 1779 7 1 2 3582 3611
0 1780 5 1 1 1779
0 1781 7 1 2 3580 3609
0 1782 5 1 1 1781
0 1783 7 3 2 3419 3412
0 1784 5 2 1 3613
0 1785 7 1 2 3578 3614
0 1786 5 1 1 1785
0 1787 7 1 2 3576 3616
0 1788 5 1 1 1787
0 1789 7 1 2 1786 1788
0 1790 5 1 1 1789
0 1791 7 3 2 3425 3428
0 1792 5 2 1 3618
0 1793 7 1 2 3572 3621
0 1794 5 1 1 1793
0 1795 7 3 2 3434 3437
0 1796 5 2 1 3623
0 1797 7 1 2 3568 3624
0 1798 5 1 1 1797
0 1799 7 1 2 3570 3626
0 1800 5 1 1 1799
0 1801 7 3 2 3443 3446
0 1802 5 2 1 3628
0 1803 7 1 2 3564 3629
0 1804 5 1 1 1803
0 1805 7 1 2 3452 3562
0 1806 5 1 1 1805
0 1807 7 2 2 3453 3456
0 1808 5 2 1 3633
0 1809 7 1 2 3560 3635
0 1810 5 1 1 1809
0 1811 7 2 2 3462 3466
0 1812 5 2 1 3637
0 1813 7 1 2 3556 3638
0 1814 5 1 1 1813
0 1815 7 1 2 3472 3554
0 1816 5 1 1 1815
0 1817 7 2 2 3473 3476
0 1818 5 2 1 3641
0 1819 7 1 2 3484 3643
0 1820 5 1 1 1819
0 1821 7 1 2 3545 3495
0 1822 5 1 1 1821
0 1823 7 2 2 3485 3481
0 1824 5 2 1 3645
0 1825 7 1 2 3550 3647
0 1826 5 1 1 1825
0 1827 7 1 2 1822 1826
0 1828 7 1 2 1820 1827
0 1829 7 1 2 1816 1828
0 1830 5 1 1 1829
0 1831 7 1 2 3558 3639
0 1832 5 1 1 1831
0 1833 7 1 2 1830 1832
0 1834 7 1 2 1814 1833
0 1835 5 1 1 1834
0 1836 7 1 2 1810 1835
0 1837 7 1 2 1806 1836
0 1838 5 1 1 1837
0 1839 7 1 2 3566 3631
0 1840 5 1 1 1839
0 1841 7 1 2 1838 1840
0 1842 7 1 2 1804 1841
0 1843 7 1 2 1800 1842
0 1844 7 1 2 1798 1843
0 1845 5 1 1 1844
0 1846 7 1 2 3574 3619
0 1847 5 1 1 1846
0 1848 7 1 2 1845 1847
0 1849 7 1 2 1794 1848
0 1850 5 1 1 1849
0 1851 7 1 2 1790 1850
0 1852 7 1 2 1782 1851
0 1853 7 1 2 1780 1852
0 1854 7 1 2 1776 1853
0 1855 7 1 2 1768 1854
0 1856 7 1 2 1756 1855
0 1857 7 1 2 1754 1856
0 1858 7 1 2 3376 3593
0 1859 5 1 1 1858
0 1860 7 2 2 3373 1859
0 1861 5 1 1 3649
0 1862 7 1 2 3368 3650
0 1863 5 1 1 1862
0 1864 7 2 2 3361 3538
0 1865 5 2 1 3651
0 1866 7 1 2 1861 3653
0 1867 5 1 1 1866
0 1868 7 1 2 1863 1867
0 1869 7 1 2 1857 1868
0 1870 7 1 2 3541 1869
0 1871 5 1 1 1870
0 1872 7 1 2 3362 3354
0 1873 5 1 1 1872
0 1874 7 1 2 3359 3352
0 1875 5 1 1 1874
0 1876 7 1 2 1873 1875
0 1877 5 1 1 1876
0 1878 7 1 2 3531 3598
0 1879 5 1 1 1878
0 1880 7 1 2 3529 3596
0 1881 5 1 1 1880
0 1882 7 1 2 1879 1881
0 1883 5 1 1 1882
0 1884 7 1 2 3395 3600
0 1885 5 1 1 1884
0 1886 7 1 2 1682 3605
0 1887 5 1 1 1886
0 1888 7 1 2 3527 3607
0 1889 5 1 1 1888
0 1890 7 1 2 3416 3610
0 1891 5 1 1 1890
0 1892 7 1 2 3420 3612
0 1893 5 1 1 1892
0 1894 7 1 2 1676 3617
0 1895 5 1 1 1894
0 1896 7 1 2 3524 3615
0 1897 5 1 1 1896
0 1898 7 1 2 1895 1897
0 1899 5 1 1 1898
0 1900 7 1 2 3515 3627
0 1901 5 1 1 1900
0 1902 7 1 2 3517 3625
0 1903 5 1 1 1902
0 1904 7 1 2 3513 3630
0 1905 5 1 1 1904
0 1906 7 1 2 3507 3634
0 1907 5 1 1 1906
0 1908 7 1 2 3463 3505
0 1909 5 1 1 1908
0 1910 7 1 2 3503 3640
0 1911 5 1 1 1910
0 1912 7 1 2 1652 3642
0 1913 5 1 1 1912
0 1914 7 1 2 3501 3644
0 1915 5 1 1 1914
0 1916 7 1 2 3548 3497
0 1917 5 1 1 1916
0 1918 7 1 2 3648 1917
0 1919 5 1 1 1918
0 1920 7 1 2 3498 3646
0 1921 5 1 1 1920
0 1922 7 1 2 1919 1921
0 1923 7 1 2 1915 1922
0 1924 7 1 2 1913 1923
0 1925 5 1 1 1924
0 1926 7 1 2 1911 1925
0 1927 7 1 2 1909 1926
0 1928 5 1 1 1927
0 1929 7 1 2 3509 3636
0 1930 5 1 1 1929
0 1931 7 1 2 1928 1930
0 1932 7 1 2 1907 1931
0 1933 5 1 1 1932
0 1934 7 1 2 3511 3632
0 1935 5 1 1 1934
0 1936 7 1 2 1933 1935
0 1937 7 1 2 1905 1936
0 1938 7 1 2 1903 1937
0 1939 7 1 2 1901 1938
0 1940 5 1 1 1939
0 1941 7 1 2 3519 3622
0 1942 5 1 1 1941
0 1943 7 1 2 3521 3620
0 1944 5 1 1 1943
0 1945 7 1 2 1942 1944
0 1946 5 1 1 1945
0 1947 7 1 2 1940 1946
0 1948 5 1 1 1947
0 1949 7 1 2 1899 1948
0 1950 7 1 2 1893 1949
0 1951 7 1 2 1891 1950
0 1952 7 1 2 1889 1951
0 1953 7 1 2 1887 1952
0 1954 7 1 2 1760 1953
0 1955 7 1 2 1885 1954
0 1956 7 1 2 3366 1955
0 1957 7 1 2 1883 1956
0 1958 7 1 2 1877 1957
0 1959 7 1 2 3533 3654
0 1960 5 1 1 1959
0 1961 7 1 2 3535 3652
0 1962 5 1 1 1961
0 1963 7 1 2 1960 1962
0 1964 7 1 2 1958 1963
0 1965 7 1 2 3542 1964
0 1966 5 1 1 1965
0 1967 7 1 2 1871 1966
0 1968 7 1 2 2734 1967
0 1969 5 1 1 1968
0 1970 7 1 2 3546 3552
0 1971 7 1 2 3467 1970
0 1972 7 1 2 3457 1971
0 1973 7 1 2 3447 1972
0 1974 7 1 2 3438 1973
0 1975 7 1 2 3429 1974
0 1976 7 1 2 3414 1975
0 1977 7 1 2 3393 1976
0 1978 7 1 2 3377 1977
0 1979 7 1 2 3355 1978
0 1980 7 1 2 3539 1979
0 1981 7 1 2 3543 1980
0 1982 5 1 1 1981
0 1983 7 1 2 735 1982
0 1984 5 1 1 1983
3 4099 7 0 2 1969 1984
