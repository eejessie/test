1 0 0 119 0
2 25 1 0
2 26 1 0
2 63719 1 0
2 63720 1 0
2 63721 1 0
2 63722 1 0
2 63723 1 0
2 63724 1 0
2 63725 1 0
2 63726 1 0
2 63727 1 0
2 63728 1 0
2 63729 1 0
2 63730 1 0
2 63731 1 0
2 63732 1 0
2 63733 1 0
2 63734 1 0
2 63735 1 0
2 63736 1 0
2 63737 1 0
2 63738 1 0
2 63739 1 0
2 63740 1 0
2 63741 1 0
2 63742 1 0
2 63743 1 0
2 63744 1 0
2 63745 1 0
2 63746 1 0
2 63747 1 0
2 63748 1 0
2 63749 1 0
2 63750 1 0
2 63751 1 0
2 63752 1 0
2 63753 1 0
2 63754 1 0
2 63755 1 0
2 63756 1 0
2 63757 1 0
2 63758 1 0
2 63759 1 0
2 63760 1 0
2 63761 1 0
2 63762 1 0
2 63763 1 0
2 63764 1 0
2 63765 1 0
2 63766 1 0
2 63767 1 0
2 63768 1 0
2 63769 1 0
2 63770 1 0
2 63771 1 0
2 63772 1 0
2 63773 1 0
2 63774 1 0
2 63775 1 0
2 63776 1 0
2 63777 1 0
2 63778 1 0
2 63779 1 0
2 63780 1 0
2 63781 1 0
2 63782 1 0
2 63783 1 0
2 63784 1 0
2 63785 1 0
2 63786 1 0
2 63787 1 0
2 63788 1 0
2 63789 1 0
2 63790 1 0
2 63791 1 0
2 63792 1 0
2 63793 1 0
2 63794 1 0
2 63795 1 0
2 63796 1 0
2 63797 1 0
2 63798 1 0
2 63799 1 0
2 63800 1 0
2 63801 1 0
2 63802 1 0
2 63803 1 0
2 63804 1 0
2 63805 1 0
2 63806 1 0
2 63807 1 0
2 63808 1 0
2 63809 1 0
2 63810 1 0
2 63811 1 0
2 63812 1 0
2 63813 1 0
2 63814 1 0
2 63815 1 0
2 63816 1 0
2 63817 1 0
2 63818 1 0
2 63819 1 0
2 63820 1 0
2 63821 1 0
2 63822 1 0
2 63823 1 0
2 63824 1 0
2 63825 1 0
2 63826 1 0
2 63827 1 0
2 63828 1 0
2 63829 1 0
2 63830 1 0
2 63831 1 0
2 63832 1 0
2 63833 1 0
2 63834 1 0
2 63835 1 0
1 1 0 114 0
2 63836 1 1
2 63837 1 1
2 63838 1 1
2 63839 1 1
2 63840 1 1
2 63841 1 1
2 63842 1 1
2 63843 1 1
2 63844 1 1
2 63845 1 1
2 63846 1 1
2 63847 1 1
2 63848 1 1
2 63849 1 1
2 63850 1 1
2 63851 1 1
2 63852 1 1
2 63853 1 1
2 63854 1 1
2 63855 1 1
2 63856 1 1
2 63857 1 1
2 63858 1 1
2 63859 1 1
2 63860 1 1
2 63861 1 1
2 63862 1 1
2 63863 1 1
2 63864 1 1
2 63865 1 1
2 63866 1 1
2 63867 1 1
2 63868 1 1
2 63869 1 1
2 63870 1 1
2 63871 1 1
2 63872 1 1
2 63873 1 1
2 63874 1 1
2 63875 1 1
2 63876 1 1
2 63877 1 1
2 63878 1 1
2 63879 1 1
2 63880 1 1
2 63881 1 1
2 63882 1 1
2 63883 1 1
2 63884 1 1
2 63885 1 1
2 63886 1 1
2 63887 1 1
2 63888 1 1
2 63889 1 1
2 63890 1 1
2 63891 1 1
2 63892 1 1
2 63893 1 1
2 63894 1 1
2 63895 1 1
2 63896 1 1
2 63897 1 1
2 63898 1 1
2 63899 1 1
2 63900 1 1
2 63901 1 1
2 63902 1 1
2 63903 1 1
2 63904 1 1
2 63905 1 1
2 63906 1 1
2 63907 1 1
2 63908 1 1
2 63909 1 1
2 63910 1 1
2 63911 1 1
2 63912 1 1
2 63913 1 1
2 63914 1 1
2 63915 1 1
2 63916 1 1
2 63917 1 1
2 63918 1 1
2 63919 1 1
2 63920 1 1
2 63921 1 1
2 63922 1 1
2 63923 1 1
2 63924 1 1
2 63925 1 1
2 63926 1 1
2 63927 1 1
2 63928 1 1
2 63929 1 1
2 63930 1 1
2 63931 1 1
2 63932 1 1
2 63933 1 1
2 63934 1 1
2 63935 1 1
2 63936 1 1
2 63937 1 1
2 63938 1 1
2 63939 1 1
2 63940 1 1
2 63941 1 1
2 63942 1 1
2 63943 1 1
2 63944 1 1
2 63945 1 1
2 63946 1 1
2 63947 1 1
2 63948 1 1
2 63949 1 1
1 2 0 60 0
2 63950 1 2
2 63951 1 2
2 63952 1 2
2 63953 1 2
2 63954 1 2
2 63955 1 2
2 63956 1 2
2 63957 1 2
2 63958 1 2
2 63959 1 2
2 63960 1 2
2 63961 1 2
2 63962 1 2
2 63963 1 2
2 63964 1 2
2 63965 1 2
2 63966 1 2
2 63967 1 2
2 63968 1 2
2 63969 1 2
2 63970 1 2
2 63971 1 2
2 63972 1 2
2 63973 1 2
2 63974 1 2
2 63975 1 2
2 63976 1 2
2 63977 1 2
2 63978 1 2
2 63979 1 2
2 63980 1 2
2 63981 1 2
2 63982 1 2
2 63983 1 2
2 63984 1 2
2 63985 1 2
2 63986 1 2
2 63987 1 2
2 63988 1 2
2 63989 1 2
2 63990 1 2
2 63991 1 2
2 63992 1 2
2 63993 1 2
2 63994 1 2
2 63995 1 2
2 63996 1 2
2 63997 1 2
2 63998 1 2
2 63999 1 2
2 64000 1 2
2 64001 1 2
2 64002 1 2
2 64003 1 2
2 64004 1 2
2 64005 1 2
2 64006 1 2
2 64007 1 2
2 64008 1 2
2 64009 1 2
1 3 0 219 0
2 64010 1 3
2 64011 1 3
2 64012 1 3
2 64013 1 3
2 64014 1 3
2 64015 1 3
2 64016 1 3
2 64017 1 3
2 64018 1 3
2 64019 1 3
2 64020 1 3
2 64021 1 3
2 64022 1 3
2 64023 1 3
2 64024 1 3
2 64025 1 3
2 64026 1 3
2 64027 1 3
2 64028 1 3
2 64029 1 3
2 64030 1 3
2 64031 1 3
2 64032 1 3
2 64033 1 3
2 64034 1 3
2 64035 1 3
2 64036 1 3
2 64037 1 3
2 64038 1 3
2 64039 1 3
2 64040 1 3
2 64041 1 3
2 64042 1 3
2 64043 1 3
2 64044 1 3
2 64045 1 3
2 64046 1 3
2 64047 1 3
2 64048 1 3
2 64049 1 3
2 64050 1 3
2 64051 1 3
2 64052 1 3
2 64053 1 3
2 64054 1 3
2 64055 1 3
2 64056 1 3
2 64057 1 3
2 64058 1 3
2 64059 1 3
2 64060 1 3
2 64061 1 3
2 64062 1 3
2 64063 1 3
2 64064 1 3
2 64065 1 3
2 64066 1 3
2 64067 1 3
2 64068 1 3
2 64069 1 3
2 64070 1 3
2 64071 1 3
2 64072 1 3
2 64073 1 3
2 64074 1 3
2 64075 1 3
2 64076 1 3
2 64077 1 3
2 64078 1 3
2 64079 1 3
2 64080 1 3
2 64081 1 3
2 64082 1 3
2 64083 1 3
2 64084 1 3
2 64085 1 3
2 64086 1 3
2 64087 1 3
2 64088 1 3
2 64089 1 3
2 64090 1 3
2 64091 1 3
2 64092 1 3
2 64093 1 3
2 64094 1 3
2 64095 1 3
2 64096 1 3
2 64097 1 3
2 64098 1 3
2 64099 1 3
2 64100 1 3
2 64101 1 3
2 64102 1 3
2 64103 1 3
2 64104 1 3
2 64105 1 3
2 64106 1 3
2 64107 1 3
2 64108 1 3
2 64109 1 3
2 64110 1 3
2 64111 1 3
2 64112 1 3
2 64113 1 3
2 64114 1 3
2 64115 1 3
2 64116 1 3
2 64117 1 3
2 64118 1 3
2 64119 1 3
2 64120 1 3
2 64121 1 3
2 64122 1 3
2 64123 1 3
2 64124 1 3
2 64125 1 3
2 64126 1 3
2 64127 1 3
2 64128 1 3
2 64129 1 3
2 64130 1 3
2 64131 1 3
2 64132 1 3
2 64133 1 3
2 64134 1 3
2 64135 1 3
2 64136 1 3
2 64137 1 3
2 64138 1 3
2 64139 1 3
2 64140 1 3
2 64141 1 3
2 64142 1 3
2 64143 1 3
2 64144 1 3
2 64145 1 3
2 64146 1 3
2 64147 1 3
2 64148 1 3
2 64149 1 3
2 64150 1 3
2 64151 1 3
2 64152 1 3
2 64153 1 3
2 64154 1 3
2 64155 1 3
2 64156 1 3
2 64157 1 3
2 64158 1 3
2 64159 1 3
2 64160 1 3
2 64161 1 3
2 64162 1 3
2 64163 1 3
2 64164 1 3
2 64165 1 3
2 64166 1 3
2 64167 1 3
2 64168 1 3
2 64169 1 3
2 64170 1 3
2 64171 1 3
2 64172 1 3
2 64173 1 3
2 64174 1 3
2 64175 1 3
2 64176 1 3
2 64177 1 3
2 64178 1 3
2 64179 1 3
2 64180 1 3
2 64181 1 3
2 64182 1 3
2 64183 1 3
2 64184 1 3
2 64185 1 3
2 64186 1 3
2 64187 1 3
2 64188 1 3
2 64189 1 3
2 64190 1 3
2 64191 1 3
2 64192 1 3
2 64193 1 3
2 64194 1 3
2 64195 1 3
2 64196 1 3
2 64197 1 3
2 64198 1 3
2 64199 1 3
2 64200 1 3
2 64201 1 3
2 64202 1 3
2 64203 1 3
2 64204 1 3
2 64205 1 3
2 64206 1 3
2 64207 1 3
2 64208 1 3
2 64209 1 3
2 64210 1 3
2 64211 1 3
2 64212 1 3
2 64213 1 3
2 64214 1 3
2 64215 1 3
2 64216 1 3
2 64217 1 3
2 64218 1 3
2 64219 1 3
2 64220 1 3
2 64221 1 3
2 64222 1 3
2 64223 1 3
2 64224 1 3
2 64225 1 3
2 64226 1 3
2 64227 1 3
2 64228 1 3
1 4 0 307 0
2 64229 1 4
2 64230 1 4
2 64231 1 4
2 64232 1 4
2 64233 1 4
2 64234 1 4
2 64235 1 4
2 64236 1 4
2 64237 1 4
2 64238 1 4
2 64239 1 4
2 64240 1 4
2 64241 1 4
2 64242 1 4
2 64243 1 4
2 64244 1 4
2 64245 1 4
2 64246 1 4
2 64247 1 4
2 64248 1 4
2 64249 1 4
2 64250 1 4
2 64251 1 4
2 64252 1 4
2 64253 1 4
2 64254 1 4
2 64255 1 4
2 64256 1 4
2 64257 1 4
2 64258 1 4
2 64259 1 4
2 64260 1 4
2 64261 1 4
2 64262 1 4
2 64263 1 4
2 64264 1 4
2 64265 1 4
2 64266 1 4
2 64267 1 4
2 64268 1 4
2 64269 1 4
2 64270 1 4
2 64271 1 4
2 64272 1 4
2 64273 1 4
2 64274 1 4
2 64275 1 4
2 64276 1 4
2 64277 1 4
2 64278 1 4
2 64279 1 4
2 64280 1 4
2 64281 1 4
2 64282 1 4
2 64283 1 4
2 64284 1 4
2 64285 1 4
2 64286 1 4
2 64287 1 4
2 64288 1 4
2 64289 1 4
2 64290 1 4
2 64291 1 4
2 64292 1 4
2 64293 1 4
2 64294 1 4
2 64295 1 4
2 64296 1 4
2 64297 1 4
2 64298 1 4
2 64299 1 4
2 64300 1 4
2 64301 1 4
2 64302 1 4
2 64303 1 4
2 64304 1 4
2 64305 1 4
2 64306 1 4
2 64307 1 4
2 64308 1 4
2 64309 1 4
2 64310 1 4
2 64311 1 4
2 64312 1 4
2 64313 1 4
2 64314 1 4
2 64315 1 4
2 64316 1 4
2 64317 1 4
2 64318 1 4
2 64319 1 4
2 64320 1 4
2 64321 1 4
2 64322 1 4
2 64323 1 4
2 64324 1 4
2 64325 1 4
2 64326 1 4
2 64327 1 4
2 64328 1 4
2 64329 1 4
2 64330 1 4
2 64331 1 4
2 64332 1 4
2 64333 1 4
2 64334 1 4
2 64335 1 4
2 64336 1 4
2 64337 1 4
2 64338 1 4
2 64339 1 4
2 64340 1 4
2 64341 1 4
2 64342 1 4
2 64343 1 4
2 64344 1 4
2 64345 1 4
2 64346 1 4
2 64347 1 4
2 64348 1 4
2 64349 1 4
2 64350 1 4
2 64351 1 4
2 64352 1 4
2 64353 1 4
2 64354 1 4
2 64355 1 4
2 64356 1 4
2 64357 1 4
2 64358 1 4
2 64359 1 4
2 64360 1 4
2 64361 1 4
2 64362 1 4
2 64363 1 4
2 64364 1 4
2 64365 1 4
2 64366 1 4
2 64367 1 4
2 64368 1 4
2 64369 1 4
2 64370 1 4
2 64371 1 4
2 64372 1 4
2 64373 1 4
2 64374 1 4
2 64375 1 4
2 64376 1 4
2 64377 1 4
2 64378 1 4
2 64379 1 4
2 64380 1 4
2 64381 1 4
2 64382 1 4
2 64383 1 4
2 64384 1 4
2 64385 1 4
2 64386 1 4
2 64387 1 4
2 64388 1 4
2 64389 1 4
2 64390 1 4
2 64391 1 4
2 64392 1 4
2 64393 1 4
2 64394 1 4
2 64395 1 4
2 64396 1 4
2 64397 1 4
2 64398 1 4
2 64399 1 4
2 64400 1 4
2 64401 1 4
2 64402 1 4
2 64403 1 4
2 64404 1 4
2 64405 1 4
2 64406 1 4
2 64407 1 4
2 64408 1 4
2 64409 1 4
2 64410 1 4
2 64411 1 4
2 64412 1 4
2 64413 1 4
2 64414 1 4
2 64415 1 4
2 64416 1 4
2 64417 1 4
2 64418 1 4
2 64419 1 4
2 64420 1 4
2 64421 1 4
2 64422 1 4
2 64423 1 4
2 64424 1 4
2 64425 1 4
2 64426 1 4
2 64427 1 4
2 64428 1 4
2 64429 1 4
2 64430 1 4
2 64431 1 4
2 64432 1 4
2 64433 1 4
2 64434 1 4
2 64435 1 4
2 64436 1 4
2 64437 1 4
2 64438 1 4
2 64439 1 4
2 64440 1 4
2 64441 1 4
2 64442 1 4
2 64443 1 4
2 64444 1 4
2 64445 1 4
2 64446 1 4
2 64447 1 4
2 64448 1 4
2 64449 1 4
2 64450 1 4
2 64451 1 4
2 64452 1 4
2 64453 1 4
2 64454 1 4
2 64455 1 4
2 64456 1 4
2 64457 1 4
2 64458 1 4
2 64459 1 4
2 64460 1 4
2 64461 1 4
2 64462 1 4
2 64463 1 4
2 64464 1 4
2 64465 1 4
2 64466 1 4
2 64467 1 4
2 64468 1 4
2 64469 1 4
2 64470 1 4
2 64471 1 4
2 64472 1 4
2 64473 1 4
2 64474 1 4
2 64475 1 4
2 64476 1 4
2 64477 1 4
2 64478 1 4
2 64479 1 4
2 64480 1 4
2 64481 1 4
2 64482 1 4
2 64483 1 4
2 64484 1 4
2 64485 1 4
2 64486 1 4
2 64487 1 4
2 64488 1 4
2 64489 1 4
2 64490 1 4
2 64491 1 4
2 64492 1 4
2 64493 1 4
2 64494 1 4
2 64495 1 4
2 64496 1 4
2 64497 1 4
2 64498 1 4
2 64499 1 4
2 64500 1 4
2 64501 1 4
2 64502 1 4
2 64503 1 4
2 64504 1 4
2 64505 1 4
2 64506 1 4
2 64507 1 4
2 64508 1 4
2 64509 1 4
2 64510 1 4
2 64511 1 4
2 64512 1 4
2 64513 1 4
2 64514 1 4
2 64515 1 4
2 64516 1 4
2 64517 1 4
2 64518 1 4
2 64519 1 4
2 64520 1 4
2 64521 1 4
2 64522 1 4
2 64523 1 4
2 64524 1 4
2 64525 1 4
2 64526 1 4
2 64527 1 4
2 64528 1 4
2 64529 1 4
2 64530 1 4
2 64531 1 4
2 64532 1 4
2 64533 1 4
2 64534 1 4
2 64535 1 4
1 5 0 384 0
2 64536 1 5
2 64537 1 5
2 64538 1 5
2 64539 1 5
2 64540 1 5
2 64541 1 5
2 64542 1 5
2 64543 1 5
2 64544 1 5
2 64545 1 5
2 64546 1 5
2 64547 1 5
2 64548 1 5
2 64549 1 5
2 64550 1 5
2 64551 1 5
2 64552 1 5
2 64553 1 5
2 64554 1 5
2 64555 1 5
2 64556 1 5
2 64557 1 5
2 64558 1 5
2 64559 1 5
2 64560 1 5
2 64561 1 5
2 64562 1 5
2 64563 1 5
2 64564 1 5
2 64565 1 5
2 64566 1 5
2 64567 1 5
2 64568 1 5
2 64569 1 5
2 64570 1 5
2 64571 1 5
2 64572 1 5
2 64573 1 5
2 64574 1 5
2 64575 1 5
2 64576 1 5
2 64577 1 5
2 64578 1 5
2 64579 1 5
2 64580 1 5
2 64581 1 5
2 64582 1 5
2 64583 1 5
2 64584 1 5
2 64585 1 5
2 64586 1 5
2 64587 1 5
2 64588 1 5
2 64589 1 5
2 64590 1 5
2 64591 1 5
2 64592 1 5
2 64593 1 5
2 64594 1 5
2 64595 1 5
2 64596 1 5
2 64597 1 5
2 64598 1 5
2 64599 1 5
2 64600 1 5
2 64601 1 5
2 64602 1 5
2 64603 1 5
2 64604 1 5
2 64605 1 5
2 64606 1 5
2 64607 1 5
2 64608 1 5
2 64609 1 5
2 64610 1 5
2 64611 1 5
2 64612 1 5
2 64613 1 5
2 64614 1 5
2 64615 1 5
2 64616 1 5
2 64617 1 5
2 64618 1 5
2 64619 1 5
2 64620 1 5
2 64621 1 5
2 64622 1 5
2 64623 1 5
2 64624 1 5
2 64625 1 5
2 64626 1 5
2 64627 1 5
2 64628 1 5
2 64629 1 5
2 64630 1 5
2 64631 1 5
2 64632 1 5
2 64633 1 5
2 64634 1 5
2 64635 1 5
2 64636 1 5
2 64637 1 5
2 64638 1 5
2 64639 1 5
2 64640 1 5
2 64641 1 5
2 64642 1 5
2 64643 1 5
2 64644 1 5
2 64645 1 5
2 64646 1 5
2 64647 1 5
2 64648 1 5
2 64649 1 5
2 64650 1 5
2 64651 1 5
2 64652 1 5
2 64653 1 5
2 64654 1 5
2 64655 1 5
2 64656 1 5
2 64657 1 5
2 64658 1 5
2 64659 1 5
2 64660 1 5
2 64661 1 5
2 64662 1 5
2 64663 1 5
2 64664 1 5
2 64665 1 5
2 64666 1 5
2 64667 1 5
2 64668 1 5
2 64669 1 5
2 64670 1 5
2 64671 1 5
2 64672 1 5
2 64673 1 5
2 64674 1 5
2 64675 1 5
2 64676 1 5
2 64677 1 5
2 64678 1 5
2 64679 1 5
2 64680 1 5
2 64681 1 5
2 64682 1 5
2 64683 1 5
2 64684 1 5
2 64685 1 5
2 64686 1 5
2 64687 1 5
2 64688 1 5
2 64689 1 5
2 64690 1 5
2 64691 1 5
2 64692 1 5
2 64693 1 5
2 64694 1 5
2 64695 1 5
2 64696 1 5
2 64697 1 5
2 64698 1 5
2 64699 1 5
2 64700 1 5
2 64701 1 5
2 64702 1 5
2 64703 1 5
2 64704 1 5
2 64705 1 5
2 64706 1 5
2 64707 1 5
2 64708 1 5
2 64709 1 5
2 64710 1 5
2 64711 1 5
2 64712 1 5
2 64713 1 5
2 64714 1 5
2 64715 1 5
2 64716 1 5
2 64717 1 5
2 64718 1 5
2 64719 1 5
2 64720 1 5
2 64721 1 5
2 64722 1 5
2 64723 1 5
2 64724 1 5
2 64725 1 5
2 64726 1 5
2 64727 1 5
2 64728 1 5
2 64729 1 5
2 64730 1 5
2 64731 1 5
2 64732 1 5
2 64733 1 5
2 64734 1 5
2 64735 1 5
2 64736 1 5
2 64737 1 5
2 64738 1 5
2 64739 1 5
2 64740 1 5
2 64741 1 5
2 64742 1 5
2 64743 1 5
2 64744 1 5
2 64745 1 5
2 64746 1 5
2 64747 1 5
2 64748 1 5
2 64749 1 5
2 64750 1 5
2 64751 1 5
2 64752 1 5
2 64753 1 5
2 64754 1 5
2 64755 1 5
2 64756 1 5
2 64757 1 5
2 64758 1 5
2 64759 1 5
2 64760 1 5
2 64761 1 5
2 64762 1 5
2 64763 1 5
2 64764 1 5
2 64765 1 5
2 64766 1 5
2 64767 1 5
2 64768 1 5
2 64769 1 5
2 64770 1 5
2 64771 1 5
2 64772 1 5
2 64773 1 5
2 64774 1 5
2 64775 1 5
2 64776 1 5
2 64777 1 5
2 64778 1 5
2 64779 1 5
2 64780 1 5
2 64781 1 5
2 64782 1 5
2 64783 1 5
2 64784 1 5
2 64785 1 5
2 64786 1 5
2 64787 1 5
2 64788 1 5
2 64789 1 5
2 64790 1 5
2 64791 1 5
2 64792 1 5
2 64793 1 5
2 64794 1 5
2 64795 1 5
2 64796 1 5
2 64797 1 5
2 64798 1 5
2 64799 1 5
2 64800 1 5
2 64801 1 5
2 64802 1 5
2 64803 1 5
2 64804 1 5
2 64805 1 5
2 64806 1 5
2 64807 1 5
2 64808 1 5
2 64809 1 5
2 64810 1 5
2 64811 1 5
2 64812 1 5
2 64813 1 5
2 64814 1 5
2 64815 1 5
2 64816 1 5
2 64817 1 5
2 64818 1 5
2 64819 1 5
2 64820 1 5
2 64821 1 5
2 64822 1 5
2 64823 1 5
2 64824 1 5
2 64825 1 5
2 64826 1 5
2 64827 1 5
2 64828 1 5
2 64829 1 5
2 64830 1 5
2 64831 1 5
2 64832 1 5
2 64833 1 5
2 64834 1 5
2 64835 1 5
2 64836 1 5
2 64837 1 5
2 64838 1 5
2 64839 1 5
2 64840 1 5
2 64841 1 5
2 64842 1 5
2 64843 1 5
2 64844 1 5
2 64845 1 5
2 64846 1 5
2 64847 1 5
2 64848 1 5
2 64849 1 5
2 64850 1 5
2 64851 1 5
2 64852 1 5
2 64853 1 5
2 64854 1 5
2 64855 1 5
2 64856 1 5
2 64857 1 5
2 64858 1 5
2 64859 1 5
2 64860 1 5
2 64861 1 5
2 64862 1 5
2 64863 1 5
2 64864 1 5
2 64865 1 5
2 64866 1 5
2 64867 1 5
2 64868 1 5
2 64869 1 5
2 64870 1 5
2 64871 1 5
2 64872 1 5
2 64873 1 5
2 64874 1 5
2 64875 1 5
2 64876 1 5
2 64877 1 5
2 64878 1 5
2 64879 1 5
2 64880 1 5
2 64881 1 5
2 64882 1 5
2 64883 1 5
2 64884 1 5
2 64885 1 5
2 64886 1 5
2 64887 1 5
2 64888 1 5
2 64889 1 5
2 64890 1 5
2 64891 1 5
2 64892 1 5
2 64893 1 5
2 64894 1 5
2 64895 1 5
2 64896 1 5
2 64897 1 5
2 64898 1 5
2 64899 1 5
2 64900 1 5
2 64901 1 5
2 64902 1 5
2 64903 1 5
2 64904 1 5
2 64905 1 5
2 64906 1 5
2 64907 1 5
2 64908 1 5
2 64909 1 5
2 64910 1 5
2 64911 1 5
2 64912 1 5
2 64913 1 5
2 64914 1 5
2 64915 1 5
2 64916 1 5
2 64917 1 5
2 64918 1 5
2 64919 1 5
1 6 0 322 0
2 64920 1 6
2 64921 1 6
2 64922 1 6
2 64923 1 6
2 64924 1 6
2 64925 1 6
2 64926 1 6
2 64927 1 6
2 64928 1 6
2 64929 1 6
2 64930 1 6
2 64931 1 6
2 64932 1 6
2 64933 1 6
2 64934 1 6
2 64935 1 6
2 64936 1 6
2 64937 1 6
2 64938 1 6
2 64939 1 6
2 64940 1 6
2 64941 1 6
2 64942 1 6
2 64943 1 6
2 64944 1 6
2 64945 1 6
2 64946 1 6
2 64947 1 6
2 64948 1 6
2 64949 1 6
2 64950 1 6
2 64951 1 6
2 64952 1 6
2 64953 1 6
2 64954 1 6
2 64955 1 6
2 64956 1 6
2 64957 1 6
2 64958 1 6
2 64959 1 6
2 64960 1 6
2 64961 1 6
2 64962 1 6
2 64963 1 6
2 64964 1 6
2 64965 1 6
2 64966 1 6
2 64967 1 6
2 64968 1 6
2 64969 1 6
2 64970 1 6
2 64971 1 6
2 64972 1 6
2 64973 1 6
2 64974 1 6
2 64975 1 6
2 64976 1 6
2 64977 1 6
2 64978 1 6
2 64979 1 6
2 64980 1 6
2 64981 1 6
2 64982 1 6
2 64983 1 6
2 64984 1 6
2 64985 1 6
2 64986 1 6
2 64987 1 6
2 64988 1 6
2 64989 1 6
2 64990 1 6
2 64991 1 6
2 64992 1 6
2 64993 1 6
2 64994 1 6
2 64995 1 6
2 64996 1 6
2 64997 1 6
2 64998 1 6
2 64999 1 6
2 65000 1 6
2 65001 1 6
2 65002 1 6
2 65003 1 6
2 65004 1 6
2 65005 1 6
2 65006 1 6
2 65007 1 6
2 65008 1 6
2 65009 1 6
2 65010 1 6
2 65011 1 6
2 65012 1 6
2 65013 1 6
2 65014 1 6
2 65015 1 6
2 65016 1 6
2 65017 1 6
2 65018 1 6
2 65019 1 6
2 65020 1 6
2 65021 1 6
2 65022 1 6
2 65023 1 6
2 65024 1 6
2 65025 1 6
2 65026 1 6
2 65027 1 6
2 65028 1 6
2 65029 1 6
2 65030 1 6
2 65031 1 6
2 65032 1 6
2 65033 1 6
2 65034 1 6
2 65035 1 6
2 65036 1 6
2 65037 1 6
2 65038 1 6
2 65039 1 6
2 65040 1 6
2 65041 1 6
2 65042 1 6
2 65043 1 6
2 65044 1 6
2 65045 1 6
2 65046 1 6
2 65047 1 6
2 65048 1 6
2 65049 1 6
2 65050 1 6
2 65051 1 6
2 65052 1 6
2 65053 1 6
2 65054 1 6
2 65055 1 6
2 65056 1 6
2 65057 1 6
2 65058 1 6
2 65059 1 6
2 65060 1 6
2 65061 1 6
2 65062 1 6
2 65063 1 6
2 65064 1 6
2 65065 1 6
2 65066 1 6
2 65067 1 6
2 65068 1 6
2 65069 1 6
2 65070 1 6
2 65071 1 6
2 65072 1 6
2 65073 1 6
2 65074 1 6
2 65075 1 6
2 65076 1 6
2 65077 1 6
2 65078 1 6
2 65079 1 6
2 65080 1 6
2 65081 1 6
2 65082 1 6
2 65083 1 6
2 65084 1 6
2 65085 1 6
2 65086 1 6
2 65087 1 6
2 65088 1 6
2 65089 1 6
2 65090 1 6
2 65091 1 6
2 65092 1 6
2 65093 1 6
2 65094 1 6
2 65095 1 6
2 65096 1 6
2 65097 1 6
2 65098 1 6
2 65099 1 6
2 65100 1 6
2 65101 1 6
2 65102 1 6
2 65103 1 6
2 65104 1 6
2 65105 1 6
2 65106 1 6
2 65107 1 6
2 65108 1 6
2 65109 1 6
2 65110 1 6
2 65111 1 6
2 65112 1 6
2 65113 1 6
2 65114 1 6
2 65115 1 6
2 65116 1 6
2 65117 1 6
2 65118 1 6
2 65119 1 6
2 65120 1 6
2 65121 1 6
2 65122 1 6
2 65123 1 6
2 65124 1 6
2 65125 1 6
2 65126 1 6
2 65127 1 6
2 65128 1 6
2 65129 1 6
2 65130 1 6
2 65131 1 6
2 65132 1 6
2 65133 1 6
2 65134 1 6
2 65135 1 6
2 65136 1 6
2 65137 1 6
2 65138 1 6
2 65139 1 6
2 65140 1 6
2 65141 1 6
2 65142 1 6
2 65143 1 6
2 65144 1 6
2 65145 1 6
2 65146 1 6
2 65147 1 6
2 65148 1 6
2 65149 1 6
2 65150 1 6
2 65151 1 6
2 65152 1 6
2 65153 1 6
2 65154 1 6
2 65155 1 6
2 65156 1 6
2 65157 1 6
2 65158 1 6
2 65159 1 6
2 65160 1 6
2 65161 1 6
2 65162 1 6
2 65163 1 6
2 65164 1 6
2 65165 1 6
2 65166 1 6
2 65167 1 6
2 65168 1 6
2 65169 1 6
2 65170 1 6
2 65171 1 6
2 65172 1 6
2 65173 1 6
2 65174 1 6
2 65175 1 6
2 65176 1 6
2 65177 1 6
2 65178 1 6
2 65179 1 6
2 65180 1 6
2 65181 1 6
2 65182 1 6
2 65183 1 6
2 65184 1 6
2 65185 1 6
2 65186 1 6
2 65187 1 6
2 65188 1 6
2 65189 1 6
2 65190 1 6
2 65191 1 6
2 65192 1 6
2 65193 1 6
2 65194 1 6
2 65195 1 6
2 65196 1 6
2 65197 1 6
2 65198 1 6
2 65199 1 6
2 65200 1 6
2 65201 1 6
2 65202 1 6
2 65203 1 6
2 65204 1 6
2 65205 1 6
2 65206 1 6
2 65207 1 6
2 65208 1 6
2 65209 1 6
2 65210 1 6
2 65211 1 6
2 65212 1 6
2 65213 1 6
2 65214 1 6
2 65215 1 6
2 65216 1 6
2 65217 1 6
2 65218 1 6
2 65219 1 6
2 65220 1 6
2 65221 1 6
2 65222 1 6
2 65223 1 6
2 65224 1 6
2 65225 1 6
2 65226 1 6
2 65227 1 6
2 65228 1 6
2 65229 1 6
2 65230 1 6
2 65231 1 6
2 65232 1 6
2 65233 1 6
2 65234 1 6
2 65235 1 6
2 65236 1 6
2 65237 1 6
2 65238 1 6
2 65239 1 6
2 65240 1 6
2 65241 1 6
1 7 0 306 0
2 65242 1 7
2 65243 1 7
2 65244 1 7
2 65245 1 7
2 65246 1 7
2 65247 1 7
2 65248 1 7
2 65249 1 7
2 65250 1 7
2 65251 1 7
2 65252 1 7
2 65253 1 7
2 65254 1 7
2 65255 1 7
2 65256 1 7
2 65257 1 7
2 65258 1 7
2 65259 1 7
2 65260 1 7
2 65261 1 7
2 65262 1 7
2 65263 1 7
2 65264 1 7
2 65265 1 7
2 65266 1 7
2 65267 1 7
2 65268 1 7
2 65269 1 7
2 65270 1 7
2 65271 1 7
2 65272 1 7
2 65273 1 7
2 65274 1 7
2 65275 1 7
2 65276 1 7
2 65277 1 7
2 65278 1 7
2 65279 1 7
2 65280 1 7
2 65281 1 7
2 65282 1 7
2 65283 1 7
2 65284 1 7
2 65285 1 7
2 65286 1 7
2 65287 1 7
2 65288 1 7
2 65289 1 7
2 65290 1 7
2 65291 1 7
2 65292 1 7
2 65293 1 7
2 65294 1 7
2 65295 1 7
2 65296 1 7
2 65297 1 7
2 65298 1 7
2 65299 1 7
2 65300 1 7
2 65301 1 7
2 65302 1 7
2 65303 1 7
2 65304 1 7
2 65305 1 7
2 65306 1 7
2 65307 1 7
2 65308 1 7
2 65309 1 7
2 65310 1 7
2 65311 1 7
2 65312 1 7
2 65313 1 7
2 65314 1 7
2 65315 1 7
2 65316 1 7
2 65317 1 7
2 65318 1 7
2 65319 1 7
2 65320 1 7
2 65321 1 7
2 65322 1 7
2 65323 1 7
2 65324 1 7
2 65325 1 7
2 65326 1 7
2 65327 1 7
2 65328 1 7
2 65329 1 7
2 65330 1 7
2 65331 1 7
2 65332 1 7
2 65333 1 7
2 65334 1 7
2 65335 1 7
2 65336 1 7
2 65337 1 7
2 65338 1 7
2 65339 1 7
2 65340 1 7
2 65341 1 7
2 65342 1 7
2 65343 1 7
2 65344 1 7
2 65345 1 7
2 65346 1 7
2 65347 1 7
2 65348 1 7
2 65349 1 7
2 65350 1 7
2 65351 1 7
2 65352 1 7
2 65353 1 7
2 65354 1 7
2 65355 1 7
2 65356 1 7
2 65357 1 7
2 65358 1 7
2 65359 1 7
2 65360 1 7
2 65361 1 7
2 65362 1 7
2 65363 1 7
2 65364 1 7
2 65365 1 7
2 65366 1 7
2 65367 1 7
2 65368 1 7
2 65369 1 7
2 65370 1 7
2 65371 1 7
2 65372 1 7
2 65373 1 7
2 65374 1 7
2 65375 1 7
2 65376 1 7
2 65377 1 7
2 65378 1 7
2 65379 1 7
2 65380 1 7
2 65381 1 7
2 65382 1 7
2 65383 1 7
2 65384 1 7
2 65385 1 7
2 65386 1 7
2 65387 1 7
2 65388 1 7
2 65389 1 7
2 65390 1 7
2 65391 1 7
2 65392 1 7
2 65393 1 7
2 65394 1 7
2 65395 1 7
2 65396 1 7
2 65397 1 7
2 65398 1 7
2 65399 1 7
2 65400 1 7
2 65401 1 7
2 65402 1 7
2 65403 1 7
2 65404 1 7
2 65405 1 7
2 65406 1 7
2 65407 1 7
2 65408 1 7
2 65409 1 7
2 65410 1 7
2 65411 1 7
2 65412 1 7
2 65413 1 7
2 65414 1 7
2 65415 1 7
2 65416 1 7
2 65417 1 7
2 65418 1 7
2 65419 1 7
2 65420 1 7
2 65421 1 7
2 65422 1 7
2 65423 1 7
2 65424 1 7
2 65425 1 7
2 65426 1 7
2 65427 1 7
2 65428 1 7
2 65429 1 7
2 65430 1 7
2 65431 1 7
2 65432 1 7
2 65433 1 7
2 65434 1 7
2 65435 1 7
2 65436 1 7
2 65437 1 7
2 65438 1 7
2 65439 1 7
2 65440 1 7
2 65441 1 7
2 65442 1 7
2 65443 1 7
2 65444 1 7
2 65445 1 7
2 65446 1 7
2 65447 1 7
2 65448 1 7
2 65449 1 7
2 65450 1 7
2 65451 1 7
2 65452 1 7
2 65453 1 7
2 65454 1 7
2 65455 1 7
2 65456 1 7
2 65457 1 7
2 65458 1 7
2 65459 1 7
2 65460 1 7
2 65461 1 7
2 65462 1 7
2 65463 1 7
2 65464 1 7
2 65465 1 7
2 65466 1 7
2 65467 1 7
2 65468 1 7
2 65469 1 7
2 65470 1 7
2 65471 1 7
2 65472 1 7
2 65473 1 7
2 65474 1 7
2 65475 1 7
2 65476 1 7
2 65477 1 7
2 65478 1 7
2 65479 1 7
2 65480 1 7
2 65481 1 7
2 65482 1 7
2 65483 1 7
2 65484 1 7
2 65485 1 7
2 65486 1 7
2 65487 1 7
2 65488 1 7
2 65489 1 7
2 65490 1 7
2 65491 1 7
2 65492 1 7
2 65493 1 7
2 65494 1 7
2 65495 1 7
2 65496 1 7
2 65497 1 7
2 65498 1 7
2 65499 1 7
2 65500 1 7
2 65501 1 7
2 65502 1 7
2 65503 1 7
2 65504 1 7
2 65505 1 7
2 65506 1 7
2 65507 1 7
2 65508 1 7
2 65509 1 7
2 65510 1 7
2 65511 1 7
2 65512 1 7
2 65513 1 7
2 65514 1 7
2 65515 1 7
2 65516 1 7
2 65517 1 7
2 65518 1 7
2 65519 1 7
2 65520 1 7
2 65521 1 7
2 65522 1 7
2 65523 1 7
2 65524 1 7
2 65525 1 7
2 65526 1 7
2 65527 1 7
2 65528 1 7
2 65529 1 7
2 65530 1 7
2 65531 1 7
2 65532 1 7
2 65533 1 7
2 65534 1 7
2 65535 1 7
2 65536 1 7
2 65537 1 7
2 65538 1 7
2 65539 1 7
2 65540 1 7
2 65541 1 7
2 65542 1 7
2 65543 1 7
2 65544 1 7
2 65545 1 7
2 65546 1 7
2 65547 1 7
1 8 0 69 0
2 65548 1 8
2 65549 1 8
2 65550 1 8
2 65551 1 8
2 65552 1 8
2 65553 1 8
2 65554 1 8
2 65555 1 8
2 65556 1 8
2 65557 1 8
2 65558 1 8
2 65559 1 8
2 65560 1 8
2 65561 1 8
2 65562 1 8
2 65563 1 8
2 65564 1 8
2 65565 1 8
2 65566 1 8
2 65567 1 8
2 65568 1 8
2 65569 1 8
2 65570 1 8
2 65571 1 8
2 65572 1 8
2 65573 1 8
2 65574 1 8
2 65575 1 8
2 65576 1 8
2 65577 1 8
2 65578 1 8
2 65579 1 8
2 65580 1 8
2 65581 1 8
2 65582 1 8
2 65583 1 8
2 65584 1 8
2 65585 1 8
2 65586 1 8
2 65587 1 8
2 65588 1 8
2 65589 1 8
2 65590 1 8
2 65591 1 8
2 65592 1 8
2 65593 1 8
2 65594 1 8
2 65595 1 8
2 65596 1 8
2 65597 1 8
2 65598 1 8
2 65599 1 8
2 65600 1 8
2 65601 1 8
2 65602 1 8
2 65603 1 8
2 65604 1 8
2 65605 1 8
2 65606 1 8
2 65607 1 8
2 65608 1 8
2 65609 1 8
2 65610 1 8
2 65611 1 8
2 65612 1 8
2 65613 1 8
2 65614 1 8
2 65615 1 8
2 65616 1 8
1 9 0 52 0
2 65617 1 9
2 65618 1 9
2 65619 1 9
2 65620 1 9
2 65621 1 9
2 65622 1 9
2 65623 1 9
2 65624 1 9
2 65625 1 9
2 65626 1 9
2 65627 1 9
2 65628 1 9
2 65629 1 9
2 65630 1 9
2 65631 1 9
2 65632 1 9
2 65633 1 9
2 65634 1 9
2 65635 1 9
2 65636 1 9
2 65637 1 9
2 65638 1 9
2 65639 1 9
2 65640 1 9
2 65641 1 9
2 65642 1 9
2 65643 1 9
2 65644 1 9
2 65645 1 9
2 65646 1 9
2 65647 1 9
2 65648 1 9
2 65649 1 9
2 65650 1 9
2 65651 1 9
2 65652 1 9
2 65653 1 9
2 65654 1 9
2 65655 1 9
2 65656 1 9
2 65657 1 9
2 65658 1 9
2 65659 1 9
2 65660 1 9
2 65661 1 9
2 65662 1 9
2 65663 1 9
2 65664 1 9
2 65665 1 9
2 65666 1 9
2 65667 1 9
2 65668 1 9
1 10 0 39 0
2 65669 1 10
2 65670 1 10
2 65671 1 10
2 65672 1 10
2 65673 1 10
2 65674 1 10
2 65675 1 10
2 65676 1 10
2 65677 1 10
2 65678 1 10
2 65679 1 10
2 65680 1 10
2 65681 1 10
2 65682 1 10
2 65683 1 10
2 65684 1 10
2 65685 1 10
2 65686 1 10
2 65687 1 10
2 65688 1 10
2 65689 1 10
2 65690 1 10
2 65691 1 10
2 65692 1 10
2 65693 1 10
2 65694 1 10
2 65695 1 10
2 65696 1 10
2 65697 1 10
2 65698 1 10
2 65699 1 10
2 65700 1 10
2 65701 1 10
2 65702 1 10
2 65703 1 10
2 65704 1 10
2 65705 1 10
2 65706 1 10
2 65707 1 10
1 11 0 158 0
2 65708 1 11
2 65709 1 11
2 65710 1 11
2 65711 1 11
2 65712 1 11
2 65713 1 11
2 65714 1 11
2 65715 1 11
2 65716 1 11
2 65717 1 11
2 65718 1 11
2 65719 1 11
2 65720 1 11
2 65721 1 11
2 65722 1 11
2 65723 1 11
2 65724 1 11
2 65725 1 11
2 65726 1 11
2 65727 1 11
2 65728 1 11
2 65729 1 11
2 65730 1 11
2 65731 1 11
2 65732 1 11
2 65733 1 11
2 65734 1 11
2 65735 1 11
2 65736 1 11
2 65737 1 11
2 65738 1 11
2 65739 1 11
2 65740 1 11
2 65741 1 11
2 65742 1 11
2 65743 1 11
2 65744 1 11
2 65745 1 11
2 65746 1 11
2 65747 1 11
2 65748 1 11
2 65749 1 11
2 65750 1 11
2 65751 1 11
2 65752 1 11
2 65753 1 11
2 65754 1 11
2 65755 1 11
2 65756 1 11
2 65757 1 11
2 65758 1 11
2 65759 1 11
2 65760 1 11
2 65761 1 11
2 65762 1 11
2 65763 1 11
2 65764 1 11
2 65765 1 11
2 65766 1 11
2 65767 1 11
2 65768 1 11
2 65769 1 11
2 65770 1 11
2 65771 1 11
2 65772 1 11
2 65773 1 11
2 65774 1 11
2 65775 1 11
2 65776 1 11
2 65777 1 11
2 65778 1 11
2 65779 1 11
2 65780 1 11
2 65781 1 11
2 65782 1 11
2 65783 1 11
2 65784 1 11
2 65785 1 11
2 65786 1 11
2 65787 1 11
2 65788 1 11
2 65789 1 11
2 65790 1 11
2 65791 1 11
2 65792 1 11
2 65793 1 11
2 65794 1 11
2 65795 1 11
2 65796 1 11
2 65797 1 11
2 65798 1 11
2 65799 1 11
2 65800 1 11
2 65801 1 11
2 65802 1 11
2 65803 1 11
2 65804 1 11
2 65805 1 11
2 65806 1 11
2 65807 1 11
2 65808 1 11
2 65809 1 11
2 65810 1 11
2 65811 1 11
2 65812 1 11
2 65813 1 11
2 65814 1 11
2 65815 1 11
2 65816 1 11
2 65817 1 11
2 65818 1 11
2 65819 1 11
2 65820 1 11
2 65821 1 11
2 65822 1 11
2 65823 1 11
2 65824 1 11
2 65825 1 11
2 65826 1 11
2 65827 1 11
2 65828 1 11
2 65829 1 11
2 65830 1 11
2 65831 1 11
2 65832 1 11
2 65833 1 11
2 65834 1 11
2 65835 1 11
2 65836 1 11
2 65837 1 11
2 65838 1 11
2 65839 1 11
2 65840 1 11
2 65841 1 11
2 65842 1 11
2 65843 1 11
2 65844 1 11
2 65845 1 11
2 65846 1 11
2 65847 1 11
2 65848 1 11
2 65849 1 11
2 65850 1 11
2 65851 1 11
2 65852 1 11
2 65853 1 11
2 65854 1 11
2 65855 1 11
2 65856 1 11
2 65857 1 11
2 65858 1 11
2 65859 1 11
2 65860 1 11
2 65861 1 11
2 65862 1 11
2 65863 1 11
2 65864 1 11
2 65865 1 11
1 12 0 230 0
2 65866 1 12
2 65867 1 12
2 65868 1 12
2 65869 1 12
2 65870 1 12
2 65871 1 12
2 65872 1 12
2 65873 1 12
2 65874 1 12
2 65875 1 12
2 65876 1 12
2 65877 1 12
2 65878 1 12
2 65879 1 12
2 65880 1 12
2 65881 1 12
2 65882 1 12
2 65883 1 12
2 65884 1 12
2 65885 1 12
2 65886 1 12
2 65887 1 12
2 65888 1 12
2 65889 1 12
2 65890 1 12
2 65891 1 12
2 65892 1 12
2 65893 1 12
2 65894 1 12
2 65895 1 12
2 65896 1 12
2 65897 1 12
2 65898 1 12
2 65899 1 12
2 65900 1 12
2 65901 1 12
2 65902 1 12
2 65903 1 12
2 65904 1 12
2 65905 1 12
2 65906 1 12
2 65907 1 12
2 65908 1 12
2 65909 1 12
2 65910 1 12
2 65911 1 12
2 65912 1 12
2 65913 1 12
2 65914 1 12
2 65915 1 12
2 65916 1 12
2 65917 1 12
2 65918 1 12
2 65919 1 12
2 65920 1 12
2 65921 1 12
2 65922 1 12
2 65923 1 12
2 65924 1 12
2 65925 1 12
2 65926 1 12
2 65927 1 12
2 65928 1 12
2 65929 1 12
2 65930 1 12
2 65931 1 12
2 65932 1 12
2 65933 1 12
2 65934 1 12
2 65935 1 12
2 65936 1 12
2 65937 1 12
2 65938 1 12
2 65939 1 12
2 65940 1 12
2 65941 1 12
2 65942 1 12
2 65943 1 12
2 65944 1 12
2 65945 1 12
2 65946 1 12
2 65947 1 12
2 65948 1 12
2 65949 1 12
2 65950 1 12
2 65951 1 12
2 65952 1 12
2 65953 1 12
2 65954 1 12
2 65955 1 12
2 65956 1 12
2 65957 1 12
2 65958 1 12
2 65959 1 12
2 65960 1 12
2 65961 1 12
2 65962 1 12
2 65963 1 12
2 65964 1 12
2 65965 1 12
2 65966 1 12
2 65967 1 12
2 65968 1 12
2 65969 1 12
2 65970 1 12
2 65971 1 12
2 65972 1 12
2 65973 1 12
2 65974 1 12
2 65975 1 12
2 65976 1 12
2 65977 1 12
2 65978 1 12
2 65979 1 12
2 65980 1 12
2 65981 1 12
2 65982 1 12
2 65983 1 12
2 65984 1 12
2 65985 1 12
2 65986 1 12
2 65987 1 12
2 65988 1 12
2 65989 1 12
2 65990 1 12
2 65991 1 12
2 65992 1 12
2 65993 1 12
2 65994 1 12
2 65995 1 12
2 65996 1 12
2 65997 1 12
2 65998 1 12
2 65999 1 12
2 66000 1 12
2 66001 1 12
2 66002 1 12
2 66003 1 12
2 66004 1 12
2 66005 1 12
2 66006 1 12
2 66007 1 12
2 66008 1 12
2 66009 1 12
2 66010 1 12
2 66011 1 12
2 66012 1 12
2 66013 1 12
2 66014 1 12
2 66015 1 12
2 66016 1 12
2 66017 1 12
2 66018 1 12
2 66019 1 12
2 66020 1 12
2 66021 1 12
2 66022 1 12
2 66023 1 12
2 66024 1 12
2 66025 1 12
2 66026 1 12
2 66027 1 12
2 66028 1 12
2 66029 1 12
2 66030 1 12
2 66031 1 12
2 66032 1 12
2 66033 1 12
2 66034 1 12
2 66035 1 12
2 66036 1 12
2 66037 1 12
2 66038 1 12
2 66039 1 12
2 66040 1 12
2 66041 1 12
2 66042 1 12
2 66043 1 12
2 66044 1 12
2 66045 1 12
2 66046 1 12
2 66047 1 12
2 66048 1 12
2 66049 1 12
2 66050 1 12
2 66051 1 12
2 66052 1 12
2 66053 1 12
2 66054 1 12
2 66055 1 12
2 66056 1 12
2 66057 1 12
2 66058 1 12
2 66059 1 12
2 66060 1 12
2 66061 1 12
2 66062 1 12
2 66063 1 12
2 66064 1 12
2 66065 1 12
2 66066 1 12
2 66067 1 12
2 66068 1 12
2 66069 1 12
2 66070 1 12
2 66071 1 12
2 66072 1 12
2 66073 1 12
2 66074 1 12
2 66075 1 12
2 66076 1 12
2 66077 1 12
2 66078 1 12
2 66079 1 12
2 66080 1 12
2 66081 1 12
2 66082 1 12
2 66083 1 12
2 66084 1 12
2 66085 1 12
2 66086 1 12
2 66087 1 12
2 66088 1 12
2 66089 1 12
2 66090 1 12
2 66091 1 12
2 66092 1 12
2 66093 1 12
2 66094 1 12
2 66095 1 12
1 13 0 319 0
2 66096 1 13
2 66097 1 13
2 66098 1 13
2 66099 1 13
2 66100 1 13
2 66101 1 13
2 66102 1 13
2 66103 1 13
2 66104 1 13
2 66105 1 13
2 66106 1 13
2 66107 1 13
2 66108 1 13
2 66109 1 13
2 66110 1 13
2 66111 1 13
2 66112 1 13
2 66113 1 13
2 66114 1 13
2 66115 1 13
2 66116 1 13
2 66117 1 13
2 66118 1 13
2 66119 1 13
2 66120 1 13
2 66121 1 13
2 66122 1 13
2 66123 1 13
2 66124 1 13
2 66125 1 13
2 66126 1 13
2 66127 1 13
2 66128 1 13
2 66129 1 13
2 66130 1 13
2 66131 1 13
2 66132 1 13
2 66133 1 13
2 66134 1 13
2 66135 1 13
2 66136 1 13
2 66137 1 13
2 66138 1 13
2 66139 1 13
2 66140 1 13
2 66141 1 13
2 66142 1 13
2 66143 1 13
2 66144 1 13
2 66145 1 13
2 66146 1 13
2 66147 1 13
2 66148 1 13
2 66149 1 13
2 66150 1 13
2 66151 1 13
2 66152 1 13
2 66153 1 13
2 66154 1 13
2 66155 1 13
2 66156 1 13
2 66157 1 13
2 66158 1 13
2 66159 1 13
2 66160 1 13
2 66161 1 13
2 66162 1 13
2 66163 1 13
2 66164 1 13
2 66165 1 13
2 66166 1 13
2 66167 1 13
2 66168 1 13
2 66169 1 13
2 66170 1 13
2 66171 1 13
2 66172 1 13
2 66173 1 13
2 66174 1 13
2 66175 1 13
2 66176 1 13
2 66177 1 13
2 66178 1 13
2 66179 1 13
2 66180 1 13
2 66181 1 13
2 66182 1 13
2 66183 1 13
2 66184 1 13
2 66185 1 13
2 66186 1 13
2 66187 1 13
2 66188 1 13
2 66189 1 13
2 66190 1 13
2 66191 1 13
2 66192 1 13
2 66193 1 13
2 66194 1 13
2 66195 1 13
2 66196 1 13
2 66197 1 13
2 66198 1 13
2 66199 1 13
2 66200 1 13
2 66201 1 13
2 66202 1 13
2 66203 1 13
2 66204 1 13
2 66205 1 13
2 66206 1 13
2 66207 1 13
2 66208 1 13
2 66209 1 13
2 66210 1 13
2 66211 1 13
2 66212 1 13
2 66213 1 13
2 66214 1 13
2 66215 1 13
2 66216 1 13
2 66217 1 13
2 66218 1 13
2 66219 1 13
2 66220 1 13
2 66221 1 13
2 66222 1 13
2 66223 1 13
2 66224 1 13
2 66225 1 13
2 66226 1 13
2 66227 1 13
2 66228 1 13
2 66229 1 13
2 66230 1 13
2 66231 1 13
2 66232 1 13
2 66233 1 13
2 66234 1 13
2 66235 1 13
2 66236 1 13
2 66237 1 13
2 66238 1 13
2 66239 1 13
2 66240 1 13
2 66241 1 13
2 66242 1 13
2 66243 1 13
2 66244 1 13
2 66245 1 13
2 66246 1 13
2 66247 1 13
2 66248 1 13
2 66249 1 13
2 66250 1 13
2 66251 1 13
2 66252 1 13
2 66253 1 13
2 66254 1 13
2 66255 1 13
2 66256 1 13
2 66257 1 13
2 66258 1 13
2 66259 1 13
2 66260 1 13
2 66261 1 13
2 66262 1 13
2 66263 1 13
2 66264 1 13
2 66265 1 13
2 66266 1 13
2 66267 1 13
2 66268 1 13
2 66269 1 13
2 66270 1 13
2 66271 1 13
2 66272 1 13
2 66273 1 13
2 66274 1 13
2 66275 1 13
2 66276 1 13
2 66277 1 13
2 66278 1 13
2 66279 1 13
2 66280 1 13
2 66281 1 13
2 66282 1 13
2 66283 1 13
2 66284 1 13
2 66285 1 13
2 66286 1 13
2 66287 1 13
2 66288 1 13
2 66289 1 13
2 66290 1 13
2 66291 1 13
2 66292 1 13
2 66293 1 13
2 66294 1 13
2 66295 1 13
2 66296 1 13
2 66297 1 13
2 66298 1 13
2 66299 1 13
2 66300 1 13
2 66301 1 13
2 66302 1 13
2 66303 1 13
2 66304 1 13
2 66305 1 13
2 66306 1 13
2 66307 1 13
2 66308 1 13
2 66309 1 13
2 66310 1 13
2 66311 1 13
2 66312 1 13
2 66313 1 13
2 66314 1 13
2 66315 1 13
2 66316 1 13
2 66317 1 13
2 66318 1 13
2 66319 1 13
2 66320 1 13
2 66321 1 13
2 66322 1 13
2 66323 1 13
2 66324 1 13
2 66325 1 13
2 66326 1 13
2 66327 1 13
2 66328 1 13
2 66329 1 13
2 66330 1 13
2 66331 1 13
2 66332 1 13
2 66333 1 13
2 66334 1 13
2 66335 1 13
2 66336 1 13
2 66337 1 13
2 66338 1 13
2 66339 1 13
2 66340 1 13
2 66341 1 13
2 66342 1 13
2 66343 1 13
2 66344 1 13
2 66345 1 13
2 66346 1 13
2 66347 1 13
2 66348 1 13
2 66349 1 13
2 66350 1 13
2 66351 1 13
2 66352 1 13
2 66353 1 13
2 66354 1 13
2 66355 1 13
2 66356 1 13
2 66357 1 13
2 66358 1 13
2 66359 1 13
2 66360 1 13
2 66361 1 13
2 66362 1 13
2 66363 1 13
2 66364 1 13
2 66365 1 13
2 66366 1 13
2 66367 1 13
2 66368 1 13
2 66369 1 13
2 66370 1 13
2 66371 1 13
2 66372 1 13
2 66373 1 13
2 66374 1 13
2 66375 1 13
2 66376 1 13
2 66377 1 13
2 66378 1 13
2 66379 1 13
2 66380 1 13
2 66381 1 13
2 66382 1 13
2 66383 1 13
2 66384 1 13
2 66385 1 13
2 66386 1 13
2 66387 1 13
2 66388 1 13
2 66389 1 13
2 66390 1 13
2 66391 1 13
2 66392 1 13
2 66393 1 13
2 66394 1 13
2 66395 1 13
2 66396 1 13
2 66397 1 13
2 66398 1 13
2 66399 1 13
2 66400 1 13
2 66401 1 13
2 66402 1 13
2 66403 1 13
2 66404 1 13
2 66405 1 13
2 66406 1 13
2 66407 1 13
2 66408 1 13
2 66409 1 13
2 66410 1 13
2 66411 1 13
2 66412 1 13
2 66413 1 13
2 66414 1 13
1 14 0 206 0
2 66415 1 14
2 66416 1 14
2 66417 1 14
2 66418 1 14
2 66419 1 14
2 66420 1 14
2 66421 1 14
2 66422 1 14
2 66423 1 14
2 66424 1 14
2 66425 1 14
2 66426 1 14
2 66427 1 14
2 66428 1 14
2 66429 1 14
2 66430 1 14
2 66431 1 14
2 66432 1 14
2 66433 1 14
2 66434 1 14
2 66435 1 14
2 66436 1 14
2 66437 1 14
2 66438 1 14
2 66439 1 14
2 66440 1 14
2 66441 1 14
2 66442 1 14
2 66443 1 14
2 66444 1 14
2 66445 1 14
2 66446 1 14
2 66447 1 14
2 66448 1 14
2 66449 1 14
2 66450 1 14
2 66451 1 14
2 66452 1 14
2 66453 1 14
2 66454 1 14
2 66455 1 14
2 66456 1 14
2 66457 1 14
2 66458 1 14
2 66459 1 14
2 66460 1 14
2 66461 1 14
2 66462 1 14
2 66463 1 14
2 66464 1 14
2 66465 1 14
2 66466 1 14
2 66467 1 14
2 66468 1 14
2 66469 1 14
2 66470 1 14
2 66471 1 14
2 66472 1 14
2 66473 1 14
2 66474 1 14
2 66475 1 14
2 66476 1 14
2 66477 1 14
2 66478 1 14
2 66479 1 14
2 66480 1 14
2 66481 1 14
2 66482 1 14
2 66483 1 14
2 66484 1 14
2 66485 1 14
2 66486 1 14
2 66487 1 14
2 66488 1 14
2 66489 1 14
2 66490 1 14
2 66491 1 14
2 66492 1 14
2 66493 1 14
2 66494 1 14
2 66495 1 14
2 66496 1 14
2 66497 1 14
2 66498 1 14
2 66499 1 14
2 66500 1 14
2 66501 1 14
2 66502 1 14
2 66503 1 14
2 66504 1 14
2 66505 1 14
2 66506 1 14
2 66507 1 14
2 66508 1 14
2 66509 1 14
2 66510 1 14
2 66511 1 14
2 66512 1 14
2 66513 1 14
2 66514 1 14
2 66515 1 14
2 66516 1 14
2 66517 1 14
2 66518 1 14
2 66519 1 14
2 66520 1 14
2 66521 1 14
2 66522 1 14
2 66523 1 14
2 66524 1 14
2 66525 1 14
2 66526 1 14
2 66527 1 14
2 66528 1 14
2 66529 1 14
2 66530 1 14
2 66531 1 14
2 66532 1 14
2 66533 1 14
2 66534 1 14
2 66535 1 14
2 66536 1 14
2 66537 1 14
2 66538 1 14
2 66539 1 14
2 66540 1 14
2 66541 1 14
2 66542 1 14
2 66543 1 14
2 66544 1 14
2 66545 1 14
2 66546 1 14
2 66547 1 14
2 66548 1 14
2 66549 1 14
2 66550 1 14
2 66551 1 14
2 66552 1 14
2 66553 1 14
2 66554 1 14
2 66555 1 14
2 66556 1 14
2 66557 1 14
2 66558 1 14
2 66559 1 14
2 66560 1 14
2 66561 1 14
2 66562 1 14
2 66563 1 14
2 66564 1 14
2 66565 1 14
2 66566 1 14
2 66567 1 14
2 66568 1 14
2 66569 1 14
2 66570 1 14
2 66571 1 14
2 66572 1 14
2 66573 1 14
2 66574 1 14
2 66575 1 14
2 66576 1 14
2 66577 1 14
2 66578 1 14
2 66579 1 14
2 66580 1 14
2 66581 1 14
2 66582 1 14
2 66583 1 14
2 66584 1 14
2 66585 1 14
2 66586 1 14
2 66587 1 14
2 66588 1 14
2 66589 1 14
2 66590 1 14
2 66591 1 14
2 66592 1 14
2 66593 1 14
2 66594 1 14
2 66595 1 14
2 66596 1 14
2 66597 1 14
2 66598 1 14
2 66599 1 14
2 66600 1 14
2 66601 1 14
2 66602 1 14
2 66603 1 14
2 66604 1 14
2 66605 1 14
2 66606 1 14
2 66607 1 14
2 66608 1 14
2 66609 1 14
2 66610 1 14
2 66611 1 14
2 66612 1 14
2 66613 1 14
2 66614 1 14
2 66615 1 14
2 66616 1 14
2 66617 1 14
2 66618 1 14
2 66619 1 14
2 66620 1 14
1 15 0 190 0
2 66621 1 15
2 66622 1 15
2 66623 1 15
2 66624 1 15
2 66625 1 15
2 66626 1 15
2 66627 1 15
2 66628 1 15
2 66629 1 15
2 66630 1 15
2 66631 1 15
2 66632 1 15
2 66633 1 15
2 66634 1 15
2 66635 1 15
2 66636 1 15
2 66637 1 15
2 66638 1 15
2 66639 1 15
2 66640 1 15
2 66641 1 15
2 66642 1 15
2 66643 1 15
2 66644 1 15
2 66645 1 15
2 66646 1 15
2 66647 1 15
2 66648 1 15
2 66649 1 15
2 66650 1 15
2 66651 1 15
2 66652 1 15
2 66653 1 15
2 66654 1 15
2 66655 1 15
2 66656 1 15
2 66657 1 15
2 66658 1 15
2 66659 1 15
2 66660 1 15
2 66661 1 15
2 66662 1 15
2 66663 1 15
2 66664 1 15
2 66665 1 15
2 66666 1 15
2 66667 1 15
2 66668 1 15
2 66669 1 15
2 66670 1 15
2 66671 1 15
2 66672 1 15
2 66673 1 15
2 66674 1 15
2 66675 1 15
2 66676 1 15
2 66677 1 15
2 66678 1 15
2 66679 1 15
2 66680 1 15
2 66681 1 15
2 66682 1 15
2 66683 1 15
2 66684 1 15
2 66685 1 15
2 66686 1 15
2 66687 1 15
2 66688 1 15
2 66689 1 15
2 66690 1 15
2 66691 1 15
2 66692 1 15
2 66693 1 15
2 66694 1 15
2 66695 1 15
2 66696 1 15
2 66697 1 15
2 66698 1 15
2 66699 1 15
2 66700 1 15
2 66701 1 15
2 66702 1 15
2 66703 1 15
2 66704 1 15
2 66705 1 15
2 66706 1 15
2 66707 1 15
2 66708 1 15
2 66709 1 15
2 66710 1 15
2 66711 1 15
2 66712 1 15
2 66713 1 15
2 66714 1 15
2 66715 1 15
2 66716 1 15
2 66717 1 15
2 66718 1 15
2 66719 1 15
2 66720 1 15
2 66721 1 15
2 66722 1 15
2 66723 1 15
2 66724 1 15
2 66725 1 15
2 66726 1 15
2 66727 1 15
2 66728 1 15
2 66729 1 15
2 66730 1 15
2 66731 1 15
2 66732 1 15
2 66733 1 15
2 66734 1 15
2 66735 1 15
2 66736 1 15
2 66737 1 15
2 66738 1 15
2 66739 1 15
2 66740 1 15
2 66741 1 15
2 66742 1 15
2 66743 1 15
2 66744 1 15
2 66745 1 15
2 66746 1 15
2 66747 1 15
2 66748 1 15
2 66749 1 15
2 66750 1 15
2 66751 1 15
2 66752 1 15
2 66753 1 15
2 66754 1 15
2 66755 1 15
2 66756 1 15
2 66757 1 15
2 66758 1 15
2 66759 1 15
2 66760 1 15
2 66761 1 15
2 66762 1 15
2 66763 1 15
2 66764 1 15
2 66765 1 15
2 66766 1 15
2 66767 1 15
2 66768 1 15
2 66769 1 15
2 66770 1 15
2 66771 1 15
2 66772 1 15
2 66773 1 15
2 66774 1 15
2 66775 1 15
2 66776 1 15
2 66777 1 15
2 66778 1 15
2 66779 1 15
2 66780 1 15
2 66781 1 15
2 66782 1 15
2 66783 1 15
2 66784 1 15
2 66785 1 15
2 66786 1 15
2 66787 1 15
2 66788 1 15
2 66789 1 15
2 66790 1 15
2 66791 1 15
2 66792 1 15
2 66793 1 15
2 66794 1 15
2 66795 1 15
2 66796 1 15
2 66797 1 15
2 66798 1 15
2 66799 1 15
2 66800 1 15
2 66801 1 15
2 66802 1 15
2 66803 1 15
2 66804 1 15
2 66805 1 15
2 66806 1 15
2 66807 1 15
2 66808 1 15
2 66809 1 15
2 66810 1 15
1 16 0 98 0
2 66811 1 16
2 66812 1 16
2 66813 1 16
2 66814 1 16
2 66815 1 16
2 66816 1 16
2 66817 1 16
2 66818 1 16
2 66819 1 16
2 66820 1 16
2 66821 1 16
2 66822 1 16
2 66823 1 16
2 66824 1 16
2 66825 1 16
2 66826 1 16
2 66827 1 16
2 66828 1 16
2 66829 1 16
2 66830 1 16
2 66831 1 16
2 66832 1 16
2 66833 1 16
2 66834 1 16
2 66835 1 16
2 66836 1 16
2 66837 1 16
2 66838 1 16
2 66839 1 16
2 66840 1 16
2 66841 1 16
2 66842 1 16
2 66843 1 16
2 66844 1 16
2 66845 1 16
2 66846 1 16
2 66847 1 16
2 66848 1 16
2 66849 1 16
2 66850 1 16
2 66851 1 16
2 66852 1 16
2 66853 1 16
2 66854 1 16
2 66855 1 16
2 66856 1 16
2 66857 1 16
2 66858 1 16
2 66859 1 16
2 66860 1 16
2 66861 1 16
2 66862 1 16
2 66863 1 16
2 66864 1 16
2 66865 1 16
2 66866 1 16
2 66867 1 16
2 66868 1 16
2 66869 1 16
2 66870 1 16
2 66871 1 16
2 66872 1 16
2 66873 1 16
2 66874 1 16
2 66875 1 16
2 66876 1 16
2 66877 1 16
2 66878 1 16
2 66879 1 16
2 66880 1 16
2 66881 1 16
2 66882 1 16
2 66883 1 16
2 66884 1 16
2 66885 1 16
2 66886 1 16
2 66887 1 16
2 66888 1 16
2 66889 1 16
2 66890 1 16
2 66891 1 16
2 66892 1 16
2 66893 1 16
2 66894 1 16
2 66895 1 16
2 66896 1 16
2 66897 1 16
2 66898 1 16
2 66899 1 16
2 66900 1 16
2 66901 1 16
2 66902 1 16
2 66903 1 16
2 66904 1 16
2 66905 1 16
2 66906 1 16
2 66907 1 16
2 66908 1 16
1 17 0 108 0
2 66909 1 17
2 66910 1 17
2 66911 1 17
2 66912 1 17
2 66913 1 17
2 66914 1 17
2 66915 1 17
2 66916 1 17
2 66917 1 17
2 66918 1 17
2 66919 1 17
2 66920 1 17
2 66921 1 17
2 66922 1 17
2 66923 1 17
2 66924 1 17
2 66925 1 17
2 66926 1 17
2 66927 1 17
2 66928 1 17
2 66929 1 17
2 66930 1 17
2 66931 1 17
2 66932 1 17
2 66933 1 17
2 66934 1 17
2 66935 1 17
2 66936 1 17
2 66937 1 17
2 66938 1 17
2 66939 1 17
2 66940 1 17
2 66941 1 17
2 66942 1 17
2 66943 1 17
2 66944 1 17
2 66945 1 17
2 66946 1 17
2 66947 1 17
2 66948 1 17
2 66949 1 17
2 66950 1 17
2 66951 1 17
2 66952 1 17
2 66953 1 17
2 66954 1 17
2 66955 1 17
2 66956 1 17
2 66957 1 17
2 66958 1 17
2 66959 1 17
2 66960 1 17
2 66961 1 17
2 66962 1 17
2 66963 1 17
2 66964 1 17
2 66965 1 17
2 66966 1 17
2 66967 1 17
2 66968 1 17
2 66969 1 17
2 66970 1 17
2 66971 1 17
2 66972 1 17
2 66973 1 17
2 66974 1 17
2 66975 1 17
2 66976 1 17
2 66977 1 17
2 66978 1 17
2 66979 1 17
2 66980 1 17
2 66981 1 17
2 66982 1 17
2 66983 1 17
2 66984 1 17
2 66985 1 17
2 66986 1 17
2 66987 1 17
2 66988 1 17
2 66989 1 17
2 66990 1 17
2 66991 1 17
2 66992 1 17
2 66993 1 17
2 66994 1 17
2 66995 1 17
2 66996 1 17
2 66997 1 17
2 66998 1 17
2 66999 1 17
2 67000 1 17
2 67001 1 17
2 67002 1 17
2 67003 1 17
2 67004 1 17
2 67005 1 17
2 67006 1 17
2 67007 1 17
2 67008 1 17
2 67009 1 17
2 67010 1 17
2 67011 1 17
2 67012 1 17
2 67013 1 17
2 67014 1 17
2 67015 1 17
2 67016 1 17
1 18 0 135 0
2 67017 1 18
2 67018 1 18
2 67019 1 18
2 67020 1 18
2 67021 1 18
2 67022 1 18
2 67023 1 18
2 67024 1 18
2 67025 1 18
2 67026 1 18
2 67027 1 18
2 67028 1 18
2 67029 1 18
2 67030 1 18
2 67031 1 18
2 67032 1 18
2 67033 1 18
2 67034 1 18
2 67035 1 18
2 67036 1 18
2 67037 1 18
2 67038 1 18
2 67039 1 18
2 67040 1 18
2 67041 1 18
2 67042 1 18
2 67043 1 18
2 67044 1 18
2 67045 1 18
2 67046 1 18
2 67047 1 18
2 67048 1 18
2 67049 1 18
2 67050 1 18
2 67051 1 18
2 67052 1 18
2 67053 1 18
2 67054 1 18
2 67055 1 18
2 67056 1 18
2 67057 1 18
2 67058 1 18
2 67059 1 18
2 67060 1 18
2 67061 1 18
2 67062 1 18
2 67063 1 18
2 67064 1 18
2 67065 1 18
2 67066 1 18
2 67067 1 18
2 67068 1 18
2 67069 1 18
2 67070 1 18
2 67071 1 18
2 67072 1 18
2 67073 1 18
2 67074 1 18
2 67075 1 18
2 67076 1 18
2 67077 1 18
2 67078 1 18
2 67079 1 18
2 67080 1 18
2 67081 1 18
2 67082 1 18
2 67083 1 18
2 67084 1 18
2 67085 1 18
2 67086 1 18
2 67087 1 18
2 67088 1 18
2 67089 1 18
2 67090 1 18
2 67091 1 18
2 67092 1 18
2 67093 1 18
2 67094 1 18
2 67095 1 18
2 67096 1 18
2 67097 1 18
2 67098 1 18
2 67099 1 18
2 67100 1 18
2 67101 1 18
2 67102 1 18
2 67103 1 18
2 67104 1 18
2 67105 1 18
2 67106 1 18
2 67107 1 18
2 67108 1 18
2 67109 1 18
2 67110 1 18
2 67111 1 18
2 67112 1 18
2 67113 1 18
2 67114 1 18
2 67115 1 18
2 67116 1 18
2 67117 1 18
2 67118 1 18
2 67119 1 18
2 67120 1 18
2 67121 1 18
2 67122 1 18
2 67123 1 18
2 67124 1 18
2 67125 1 18
2 67126 1 18
2 67127 1 18
2 67128 1 18
2 67129 1 18
2 67130 1 18
2 67131 1 18
2 67132 1 18
2 67133 1 18
2 67134 1 18
2 67135 1 18
2 67136 1 18
2 67137 1 18
2 67138 1 18
2 67139 1 18
2 67140 1 18
2 67141 1 18
2 67142 1 18
2 67143 1 18
2 67144 1 18
2 67145 1 18
2 67146 1 18
2 67147 1 18
2 67148 1 18
2 67149 1 18
2 67150 1 18
2 67151 1 18
1 19 0 99 0
2 67152 1 19
2 67153 1 19
2 67154 1 19
2 67155 1 19
2 67156 1 19
2 67157 1 19
2 67158 1 19
2 67159 1 19
2 67160 1 19
2 67161 1 19
2 67162 1 19
2 67163 1 19
2 67164 1 19
2 67165 1 19
2 67166 1 19
2 67167 1 19
2 67168 1 19
2 67169 1 19
2 67170 1 19
2 67171 1 19
2 67172 1 19
2 67173 1 19
2 67174 1 19
2 67175 1 19
2 67176 1 19
2 67177 1 19
2 67178 1 19
2 67179 1 19
2 67180 1 19
2 67181 1 19
2 67182 1 19
2 67183 1 19
2 67184 1 19
2 67185 1 19
2 67186 1 19
2 67187 1 19
2 67188 1 19
2 67189 1 19
2 67190 1 19
2 67191 1 19
2 67192 1 19
2 67193 1 19
2 67194 1 19
2 67195 1 19
2 67196 1 19
2 67197 1 19
2 67198 1 19
2 67199 1 19
2 67200 1 19
2 67201 1 19
2 67202 1 19
2 67203 1 19
2 67204 1 19
2 67205 1 19
2 67206 1 19
2 67207 1 19
2 67208 1 19
2 67209 1 19
2 67210 1 19
2 67211 1 19
2 67212 1 19
2 67213 1 19
2 67214 1 19
2 67215 1 19
2 67216 1 19
2 67217 1 19
2 67218 1 19
2 67219 1 19
2 67220 1 19
2 67221 1 19
2 67222 1 19
2 67223 1 19
2 67224 1 19
2 67225 1 19
2 67226 1 19
2 67227 1 19
2 67228 1 19
2 67229 1 19
2 67230 1 19
2 67231 1 19
2 67232 1 19
2 67233 1 19
2 67234 1 19
2 67235 1 19
2 67236 1 19
2 67237 1 19
2 67238 1 19
2 67239 1 19
2 67240 1 19
2 67241 1 19
2 67242 1 19
2 67243 1 19
2 67244 1 19
2 67245 1 19
2 67246 1 19
2 67247 1 19
2 67248 1 19
2 67249 1 19
2 67250 1 19
1 20 0 244 0
2 67251 1 20
2 67252 1 20
2 67253 1 20
2 67254 1 20
2 67255 1 20
2 67256 1 20
2 67257 1 20
2 67258 1 20
2 67259 1 20
2 67260 1 20
2 67261 1 20
2 67262 1 20
2 67263 1 20
2 67264 1 20
2 67265 1 20
2 67266 1 20
2 67267 1 20
2 67268 1 20
2 67269 1 20
2 67270 1 20
2 67271 1 20
2 67272 1 20
2 67273 1 20
2 67274 1 20
2 67275 1 20
2 67276 1 20
2 67277 1 20
2 67278 1 20
2 67279 1 20
2 67280 1 20
2 67281 1 20
2 67282 1 20
2 67283 1 20
2 67284 1 20
2 67285 1 20
2 67286 1 20
2 67287 1 20
2 67288 1 20
2 67289 1 20
2 67290 1 20
2 67291 1 20
2 67292 1 20
2 67293 1 20
2 67294 1 20
2 67295 1 20
2 67296 1 20
2 67297 1 20
2 67298 1 20
2 67299 1 20
2 67300 1 20
2 67301 1 20
2 67302 1 20
2 67303 1 20
2 67304 1 20
2 67305 1 20
2 67306 1 20
2 67307 1 20
2 67308 1 20
2 67309 1 20
2 67310 1 20
2 67311 1 20
2 67312 1 20
2 67313 1 20
2 67314 1 20
2 67315 1 20
2 67316 1 20
2 67317 1 20
2 67318 1 20
2 67319 1 20
2 67320 1 20
2 67321 1 20
2 67322 1 20
2 67323 1 20
2 67324 1 20
2 67325 1 20
2 67326 1 20
2 67327 1 20
2 67328 1 20
2 67329 1 20
2 67330 1 20
2 67331 1 20
2 67332 1 20
2 67333 1 20
2 67334 1 20
2 67335 1 20
2 67336 1 20
2 67337 1 20
2 67338 1 20
2 67339 1 20
2 67340 1 20
2 67341 1 20
2 67342 1 20
2 67343 1 20
2 67344 1 20
2 67345 1 20
2 67346 1 20
2 67347 1 20
2 67348 1 20
2 67349 1 20
2 67350 1 20
2 67351 1 20
2 67352 1 20
2 67353 1 20
2 67354 1 20
2 67355 1 20
2 67356 1 20
2 67357 1 20
2 67358 1 20
2 67359 1 20
2 67360 1 20
2 67361 1 20
2 67362 1 20
2 67363 1 20
2 67364 1 20
2 67365 1 20
2 67366 1 20
2 67367 1 20
2 67368 1 20
2 67369 1 20
2 67370 1 20
2 67371 1 20
2 67372 1 20
2 67373 1 20
2 67374 1 20
2 67375 1 20
2 67376 1 20
2 67377 1 20
2 67378 1 20
2 67379 1 20
2 67380 1 20
2 67381 1 20
2 67382 1 20
2 67383 1 20
2 67384 1 20
2 67385 1 20
2 67386 1 20
2 67387 1 20
2 67388 1 20
2 67389 1 20
2 67390 1 20
2 67391 1 20
2 67392 1 20
2 67393 1 20
2 67394 1 20
2 67395 1 20
2 67396 1 20
2 67397 1 20
2 67398 1 20
2 67399 1 20
2 67400 1 20
2 67401 1 20
2 67402 1 20
2 67403 1 20
2 67404 1 20
2 67405 1 20
2 67406 1 20
2 67407 1 20
2 67408 1 20
2 67409 1 20
2 67410 1 20
2 67411 1 20
2 67412 1 20
2 67413 1 20
2 67414 1 20
2 67415 1 20
2 67416 1 20
2 67417 1 20
2 67418 1 20
2 67419 1 20
2 67420 1 20
2 67421 1 20
2 67422 1 20
2 67423 1 20
2 67424 1 20
2 67425 1 20
2 67426 1 20
2 67427 1 20
2 67428 1 20
2 67429 1 20
2 67430 1 20
2 67431 1 20
2 67432 1 20
2 67433 1 20
2 67434 1 20
2 67435 1 20
2 67436 1 20
2 67437 1 20
2 67438 1 20
2 67439 1 20
2 67440 1 20
2 67441 1 20
2 67442 1 20
2 67443 1 20
2 67444 1 20
2 67445 1 20
2 67446 1 20
2 67447 1 20
2 67448 1 20
2 67449 1 20
2 67450 1 20
2 67451 1 20
2 67452 1 20
2 67453 1 20
2 67454 1 20
2 67455 1 20
2 67456 1 20
2 67457 1 20
2 67458 1 20
2 67459 1 20
2 67460 1 20
2 67461 1 20
2 67462 1 20
2 67463 1 20
2 67464 1 20
2 67465 1 20
2 67466 1 20
2 67467 1 20
2 67468 1 20
2 67469 1 20
2 67470 1 20
2 67471 1 20
2 67472 1 20
2 67473 1 20
2 67474 1 20
2 67475 1 20
2 67476 1 20
2 67477 1 20
2 67478 1 20
2 67479 1 20
2 67480 1 20
2 67481 1 20
2 67482 1 20
2 67483 1 20
2 67484 1 20
2 67485 1 20
2 67486 1 20
2 67487 1 20
2 67488 1 20
2 67489 1 20
2 67490 1 20
2 67491 1 20
2 67492 1 20
2 67493 1 20
2 67494 1 20
1 21 0 344 0
2 67495 1 21
2 67496 1 21
2 67497 1 21
2 67498 1 21
2 67499 1 21
2 67500 1 21
2 67501 1 21
2 67502 1 21
2 67503 1 21
2 67504 1 21
2 67505 1 21
2 67506 1 21
2 67507 1 21
2 67508 1 21
2 67509 1 21
2 67510 1 21
2 67511 1 21
2 67512 1 21
2 67513 1 21
2 67514 1 21
2 67515 1 21
2 67516 1 21
2 67517 1 21
2 67518 1 21
2 67519 1 21
2 67520 1 21
2 67521 1 21
2 67522 1 21
2 67523 1 21
2 67524 1 21
2 67525 1 21
2 67526 1 21
2 67527 1 21
2 67528 1 21
2 67529 1 21
2 67530 1 21
2 67531 1 21
2 67532 1 21
2 67533 1 21
2 67534 1 21
2 67535 1 21
2 67536 1 21
2 67537 1 21
2 67538 1 21
2 67539 1 21
2 67540 1 21
2 67541 1 21
2 67542 1 21
2 67543 1 21
2 67544 1 21
2 67545 1 21
2 67546 1 21
2 67547 1 21
2 67548 1 21
2 67549 1 21
2 67550 1 21
2 67551 1 21
2 67552 1 21
2 67553 1 21
2 67554 1 21
2 67555 1 21
2 67556 1 21
2 67557 1 21
2 67558 1 21
2 67559 1 21
2 67560 1 21
2 67561 1 21
2 67562 1 21
2 67563 1 21
2 67564 1 21
2 67565 1 21
2 67566 1 21
2 67567 1 21
2 67568 1 21
2 67569 1 21
2 67570 1 21
2 67571 1 21
2 67572 1 21
2 67573 1 21
2 67574 1 21
2 67575 1 21
2 67576 1 21
2 67577 1 21
2 67578 1 21
2 67579 1 21
2 67580 1 21
2 67581 1 21
2 67582 1 21
2 67583 1 21
2 67584 1 21
2 67585 1 21
2 67586 1 21
2 67587 1 21
2 67588 1 21
2 67589 1 21
2 67590 1 21
2 67591 1 21
2 67592 1 21
2 67593 1 21
2 67594 1 21
2 67595 1 21
2 67596 1 21
2 67597 1 21
2 67598 1 21
2 67599 1 21
2 67600 1 21
2 67601 1 21
2 67602 1 21
2 67603 1 21
2 67604 1 21
2 67605 1 21
2 67606 1 21
2 67607 1 21
2 67608 1 21
2 67609 1 21
2 67610 1 21
2 67611 1 21
2 67612 1 21
2 67613 1 21
2 67614 1 21
2 67615 1 21
2 67616 1 21
2 67617 1 21
2 67618 1 21
2 67619 1 21
2 67620 1 21
2 67621 1 21
2 67622 1 21
2 67623 1 21
2 67624 1 21
2 67625 1 21
2 67626 1 21
2 67627 1 21
2 67628 1 21
2 67629 1 21
2 67630 1 21
2 67631 1 21
2 67632 1 21
2 67633 1 21
2 67634 1 21
2 67635 1 21
2 67636 1 21
2 67637 1 21
2 67638 1 21
2 67639 1 21
2 67640 1 21
2 67641 1 21
2 67642 1 21
2 67643 1 21
2 67644 1 21
2 67645 1 21
2 67646 1 21
2 67647 1 21
2 67648 1 21
2 67649 1 21
2 67650 1 21
2 67651 1 21
2 67652 1 21
2 67653 1 21
2 67654 1 21
2 67655 1 21
2 67656 1 21
2 67657 1 21
2 67658 1 21
2 67659 1 21
2 67660 1 21
2 67661 1 21
2 67662 1 21
2 67663 1 21
2 67664 1 21
2 67665 1 21
2 67666 1 21
2 67667 1 21
2 67668 1 21
2 67669 1 21
2 67670 1 21
2 67671 1 21
2 67672 1 21
2 67673 1 21
2 67674 1 21
2 67675 1 21
2 67676 1 21
2 67677 1 21
2 67678 1 21
2 67679 1 21
2 67680 1 21
2 67681 1 21
2 67682 1 21
2 67683 1 21
2 67684 1 21
2 67685 1 21
2 67686 1 21
2 67687 1 21
2 67688 1 21
2 67689 1 21
2 67690 1 21
2 67691 1 21
2 67692 1 21
2 67693 1 21
2 67694 1 21
2 67695 1 21
2 67696 1 21
2 67697 1 21
2 67698 1 21
2 67699 1 21
2 67700 1 21
2 67701 1 21
2 67702 1 21
2 67703 1 21
2 67704 1 21
2 67705 1 21
2 67706 1 21
2 67707 1 21
2 67708 1 21
2 67709 1 21
2 67710 1 21
2 67711 1 21
2 67712 1 21
2 67713 1 21
2 67714 1 21
2 67715 1 21
2 67716 1 21
2 67717 1 21
2 67718 1 21
2 67719 1 21
2 67720 1 21
2 67721 1 21
2 67722 1 21
2 67723 1 21
2 67724 1 21
2 67725 1 21
2 67726 1 21
2 67727 1 21
2 67728 1 21
2 67729 1 21
2 67730 1 21
2 67731 1 21
2 67732 1 21
2 67733 1 21
2 67734 1 21
2 67735 1 21
2 67736 1 21
2 67737 1 21
2 67738 1 21
2 67739 1 21
2 67740 1 21
2 67741 1 21
2 67742 1 21
2 67743 1 21
2 67744 1 21
2 67745 1 21
2 67746 1 21
2 67747 1 21
2 67748 1 21
2 67749 1 21
2 67750 1 21
2 67751 1 21
2 67752 1 21
2 67753 1 21
2 67754 1 21
2 67755 1 21
2 67756 1 21
2 67757 1 21
2 67758 1 21
2 67759 1 21
2 67760 1 21
2 67761 1 21
2 67762 1 21
2 67763 1 21
2 67764 1 21
2 67765 1 21
2 67766 1 21
2 67767 1 21
2 67768 1 21
2 67769 1 21
2 67770 1 21
2 67771 1 21
2 67772 1 21
2 67773 1 21
2 67774 1 21
2 67775 1 21
2 67776 1 21
2 67777 1 21
2 67778 1 21
2 67779 1 21
2 67780 1 21
2 67781 1 21
2 67782 1 21
2 67783 1 21
2 67784 1 21
2 67785 1 21
2 67786 1 21
2 67787 1 21
2 67788 1 21
2 67789 1 21
2 67790 1 21
2 67791 1 21
2 67792 1 21
2 67793 1 21
2 67794 1 21
2 67795 1 21
2 67796 1 21
2 67797 1 21
2 67798 1 21
2 67799 1 21
2 67800 1 21
2 67801 1 21
2 67802 1 21
2 67803 1 21
2 67804 1 21
2 67805 1 21
2 67806 1 21
2 67807 1 21
2 67808 1 21
2 67809 1 21
2 67810 1 21
2 67811 1 21
2 67812 1 21
2 67813 1 21
2 67814 1 21
2 67815 1 21
2 67816 1 21
2 67817 1 21
2 67818 1 21
2 67819 1 21
2 67820 1 21
2 67821 1 21
2 67822 1 21
2 67823 1 21
2 67824 1 21
2 67825 1 21
2 67826 1 21
2 67827 1 21
2 67828 1 21
2 67829 1 21
2 67830 1 21
2 67831 1 21
2 67832 1 21
2 67833 1 21
2 67834 1 21
2 67835 1 21
2 67836 1 21
2 67837 1 21
2 67838 1 21
1 22 0 392 0
2 67839 1 22
2 67840 1 22
2 67841 1 22
2 67842 1 22
2 67843 1 22
2 67844 1 22
2 67845 1 22
2 67846 1 22
2 67847 1 22
2 67848 1 22
2 67849 1 22
2 67850 1 22
2 67851 1 22
2 67852 1 22
2 67853 1 22
2 67854 1 22
2 67855 1 22
2 67856 1 22
2 67857 1 22
2 67858 1 22
2 67859 1 22
2 67860 1 22
2 67861 1 22
2 67862 1 22
2 67863 1 22
2 67864 1 22
2 67865 1 22
2 67866 1 22
2 67867 1 22
2 67868 1 22
2 67869 1 22
2 67870 1 22
2 67871 1 22
2 67872 1 22
2 67873 1 22
2 67874 1 22
2 67875 1 22
2 67876 1 22
2 67877 1 22
2 67878 1 22
2 67879 1 22
2 67880 1 22
2 67881 1 22
2 67882 1 22
2 67883 1 22
2 67884 1 22
2 67885 1 22
2 67886 1 22
2 67887 1 22
2 67888 1 22
2 67889 1 22
2 67890 1 22
2 67891 1 22
2 67892 1 22
2 67893 1 22
2 67894 1 22
2 67895 1 22
2 67896 1 22
2 67897 1 22
2 67898 1 22
2 67899 1 22
2 67900 1 22
2 67901 1 22
2 67902 1 22
2 67903 1 22
2 67904 1 22
2 67905 1 22
2 67906 1 22
2 67907 1 22
2 67908 1 22
2 67909 1 22
2 67910 1 22
2 67911 1 22
2 67912 1 22
2 67913 1 22
2 67914 1 22
2 67915 1 22
2 67916 1 22
2 67917 1 22
2 67918 1 22
2 67919 1 22
2 67920 1 22
2 67921 1 22
2 67922 1 22
2 67923 1 22
2 67924 1 22
2 67925 1 22
2 67926 1 22
2 67927 1 22
2 67928 1 22
2 67929 1 22
2 67930 1 22
2 67931 1 22
2 67932 1 22
2 67933 1 22
2 67934 1 22
2 67935 1 22
2 67936 1 22
2 67937 1 22
2 67938 1 22
2 67939 1 22
2 67940 1 22
2 67941 1 22
2 67942 1 22
2 67943 1 22
2 67944 1 22
2 67945 1 22
2 67946 1 22
2 67947 1 22
2 67948 1 22
2 67949 1 22
2 67950 1 22
2 67951 1 22
2 67952 1 22
2 67953 1 22
2 67954 1 22
2 67955 1 22
2 67956 1 22
2 67957 1 22
2 67958 1 22
2 67959 1 22
2 67960 1 22
2 67961 1 22
2 67962 1 22
2 67963 1 22
2 67964 1 22
2 67965 1 22
2 67966 1 22
2 67967 1 22
2 67968 1 22
2 67969 1 22
2 67970 1 22
2 67971 1 22
2 67972 1 22
2 67973 1 22
2 67974 1 22
2 67975 1 22
2 67976 1 22
2 67977 1 22
2 67978 1 22
2 67979 1 22
2 67980 1 22
2 67981 1 22
2 67982 1 22
2 67983 1 22
2 67984 1 22
2 67985 1 22
2 67986 1 22
2 67987 1 22
2 67988 1 22
2 67989 1 22
2 67990 1 22
2 67991 1 22
2 67992 1 22
2 67993 1 22
2 67994 1 22
2 67995 1 22
2 67996 1 22
2 67997 1 22
2 67998 1 22
2 67999 1 22
2 68000 1 22
2 68001 1 22
2 68002 1 22
2 68003 1 22
2 68004 1 22
2 68005 1 22
2 68006 1 22
2 68007 1 22
2 68008 1 22
2 68009 1 22
2 68010 1 22
2 68011 1 22
2 68012 1 22
2 68013 1 22
2 68014 1 22
2 68015 1 22
2 68016 1 22
2 68017 1 22
2 68018 1 22
2 68019 1 22
2 68020 1 22
2 68021 1 22
2 68022 1 22
2 68023 1 22
2 68024 1 22
2 68025 1 22
2 68026 1 22
2 68027 1 22
2 68028 1 22
2 68029 1 22
2 68030 1 22
2 68031 1 22
2 68032 1 22
2 68033 1 22
2 68034 1 22
2 68035 1 22
2 68036 1 22
2 68037 1 22
2 68038 1 22
2 68039 1 22
2 68040 1 22
2 68041 1 22
2 68042 1 22
2 68043 1 22
2 68044 1 22
2 68045 1 22
2 68046 1 22
2 68047 1 22
2 68048 1 22
2 68049 1 22
2 68050 1 22
2 68051 1 22
2 68052 1 22
2 68053 1 22
2 68054 1 22
2 68055 1 22
2 68056 1 22
2 68057 1 22
2 68058 1 22
2 68059 1 22
2 68060 1 22
2 68061 1 22
2 68062 1 22
2 68063 1 22
2 68064 1 22
2 68065 1 22
2 68066 1 22
2 68067 1 22
2 68068 1 22
2 68069 1 22
2 68070 1 22
2 68071 1 22
2 68072 1 22
2 68073 1 22
2 68074 1 22
2 68075 1 22
2 68076 1 22
2 68077 1 22
2 68078 1 22
2 68079 1 22
2 68080 1 22
2 68081 1 22
2 68082 1 22
2 68083 1 22
2 68084 1 22
2 68085 1 22
2 68086 1 22
2 68087 1 22
2 68088 1 22
2 68089 1 22
2 68090 1 22
2 68091 1 22
2 68092 1 22
2 68093 1 22
2 68094 1 22
2 68095 1 22
2 68096 1 22
2 68097 1 22
2 68098 1 22
2 68099 1 22
2 68100 1 22
2 68101 1 22
2 68102 1 22
2 68103 1 22
2 68104 1 22
2 68105 1 22
2 68106 1 22
2 68107 1 22
2 68108 1 22
2 68109 1 22
2 68110 1 22
2 68111 1 22
2 68112 1 22
2 68113 1 22
2 68114 1 22
2 68115 1 22
2 68116 1 22
2 68117 1 22
2 68118 1 22
2 68119 1 22
2 68120 1 22
2 68121 1 22
2 68122 1 22
2 68123 1 22
2 68124 1 22
2 68125 1 22
2 68126 1 22
2 68127 1 22
2 68128 1 22
2 68129 1 22
2 68130 1 22
2 68131 1 22
2 68132 1 22
2 68133 1 22
2 68134 1 22
2 68135 1 22
2 68136 1 22
2 68137 1 22
2 68138 1 22
2 68139 1 22
2 68140 1 22
2 68141 1 22
2 68142 1 22
2 68143 1 22
2 68144 1 22
2 68145 1 22
2 68146 1 22
2 68147 1 22
2 68148 1 22
2 68149 1 22
2 68150 1 22
2 68151 1 22
2 68152 1 22
2 68153 1 22
2 68154 1 22
2 68155 1 22
2 68156 1 22
2 68157 1 22
2 68158 1 22
2 68159 1 22
2 68160 1 22
2 68161 1 22
2 68162 1 22
2 68163 1 22
2 68164 1 22
2 68165 1 22
2 68166 1 22
2 68167 1 22
2 68168 1 22
2 68169 1 22
2 68170 1 22
2 68171 1 22
2 68172 1 22
2 68173 1 22
2 68174 1 22
2 68175 1 22
2 68176 1 22
2 68177 1 22
2 68178 1 22
2 68179 1 22
2 68180 1 22
2 68181 1 22
2 68182 1 22
2 68183 1 22
2 68184 1 22
2 68185 1 22
2 68186 1 22
2 68187 1 22
2 68188 1 22
2 68189 1 22
2 68190 1 22
2 68191 1 22
2 68192 1 22
2 68193 1 22
2 68194 1 22
2 68195 1 22
2 68196 1 22
2 68197 1 22
2 68198 1 22
2 68199 1 22
2 68200 1 22
2 68201 1 22
2 68202 1 22
2 68203 1 22
2 68204 1 22
2 68205 1 22
2 68206 1 22
2 68207 1 22
2 68208 1 22
2 68209 1 22
2 68210 1 22
2 68211 1 22
2 68212 1 22
2 68213 1 22
2 68214 1 22
2 68215 1 22
2 68216 1 22
2 68217 1 22
2 68218 1 22
2 68219 1 22
2 68220 1 22
2 68221 1 22
2 68222 1 22
2 68223 1 22
2 68224 1 22
2 68225 1 22
2 68226 1 22
2 68227 1 22
2 68228 1 22
2 68229 1 22
2 68230 1 22
1 23 0 310 0
2 68231 1 23
2 68232 1 23
2 68233 1 23
2 68234 1 23
2 68235 1 23
2 68236 1 23
2 68237 1 23
2 68238 1 23
2 68239 1 23
2 68240 1 23
2 68241 1 23
2 68242 1 23
2 68243 1 23
2 68244 1 23
2 68245 1 23
2 68246 1 23
2 68247 1 23
2 68248 1 23
2 68249 1 23
2 68250 1 23
2 68251 1 23
2 68252 1 23
2 68253 1 23
2 68254 1 23
2 68255 1 23
2 68256 1 23
2 68257 1 23
2 68258 1 23
2 68259 1 23
2 68260 1 23
2 68261 1 23
2 68262 1 23
2 68263 1 23
2 68264 1 23
2 68265 1 23
2 68266 1 23
2 68267 1 23
2 68268 1 23
2 68269 1 23
2 68270 1 23
2 68271 1 23
2 68272 1 23
2 68273 1 23
2 68274 1 23
2 68275 1 23
2 68276 1 23
2 68277 1 23
2 68278 1 23
2 68279 1 23
2 68280 1 23
2 68281 1 23
2 68282 1 23
2 68283 1 23
2 68284 1 23
2 68285 1 23
2 68286 1 23
2 68287 1 23
2 68288 1 23
2 68289 1 23
2 68290 1 23
2 68291 1 23
2 68292 1 23
2 68293 1 23
2 68294 1 23
2 68295 1 23
2 68296 1 23
2 68297 1 23
2 68298 1 23
2 68299 1 23
2 68300 1 23
2 68301 1 23
2 68302 1 23
2 68303 1 23
2 68304 1 23
2 68305 1 23
2 68306 1 23
2 68307 1 23
2 68308 1 23
2 68309 1 23
2 68310 1 23
2 68311 1 23
2 68312 1 23
2 68313 1 23
2 68314 1 23
2 68315 1 23
2 68316 1 23
2 68317 1 23
2 68318 1 23
2 68319 1 23
2 68320 1 23
2 68321 1 23
2 68322 1 23
2 68323 1 23
2 68324 1 23
2 68325 1 23
2 68326 1 23
2 68327 1 23
2 68328 1 23
2 68329 1 23
2 68330 1 23
2 68331 1 23
2 68332 1 23
2 68333 1 23
2 68334 1 23
2 68335 1 23
2 68336 1 23
2 68337 1 23
2 68338 1 23
2 68339 1 23
2 68340 1 23
2 68341 1 23
2 68342 1 23
2 68343 1 23
2 68344 1 23
2 68345 1 23
2 68346 1 23
2 68347 1 23
2 68348 1 23
2 68349 1 23
2 68350 1 23
2 68351 1 23
2 68352 1 23
2 68353 1 23
2 68354 1 23
2 68355 1 23
2 68356 1 23
2 68357 1 23
2 68358 1 23
2 68359 1 23
2 68360 1 23
2 68361 1 23
2 68362 1 23
2 68363 1 23
2 68364 1 23
2 68365 1 23
2 68366 1 23
2 68367 1 23
2 68368 1 23
2 68369 1 23
2 68370 1 23
2 68371 1 23
2 68372 1 23
2 68373 1 23
2 68374 1 23
2 68375 1 23
2 68376 1 23
2 68377 1 23
2 68378 1 23
2 68379 1 23
2 68380 1 23
2 68381 1 23
2 68382 1 23
2 68383 1 23
2 68384 1 23
2 68385 1 23
2 68386 1 23
2 68387 1 23
2 68388 1 23
2 68389 1 23
2 68390 1 23
2 68391 1 23
2 68392 1 23
2 68393 1 23
2 68394 1 23
2 68395 1 23
2 68396 1 23
2 68397 1 23
2 68398 1 23
2 68399 1 23
2 68400 1 23
2 68401 1 23
2 68402 1 23
2 68403 1 23
2 68404 1 23
2 68405 1 23
2 68406 1 23
2 68407 1 23
2 68408 1 23
2 68409 1 23
2 68410 1 23
2 68411 1 23
2 68412 1 23
2 68413 1 23
2 68414 1 23
2 68415 1 23
2 68416 1 23
2 68417 1 23
2 68418 1 23
2 68419 1 23
2 68420 1 23
2 68421 1 23
2 68422 1 23
2 68423 1 23
2 68424 1 23
2 68425 1 23
2 68426 1 23
2 68427 1 23
2 68428 1 23
2 68429 1 23
2 68430 1 23
2 68431 1 23
2 68432 1 23
2 68433 1 23
2 68434 1 23
2 68435 1 23
2 68436 1 23
2 68437 1 23
2 68438 1 23
2 68439 1 23
2 68440 1 23
2 68441 1 23
2 68442 1 23
2 68443 1 23
2 68444 1 23
2 68445 1 23
2 68446 1 23
2 68447 1 23
2 68448 1 23
2 68449 1 23
2 68450 1 23
2 68451 1 23
2 68452 1 23
2 68453 1 23
2 68454 1 23
2 68455 1 23
2 68456 1 23
2 68457 1 23
2 68458 1 23
2 68459 1 23
2 68460 1 23
2 68461 1 23
2 68462 1 23
2 68463 1 23
2 68464 1 23
2 68465 1 23
2 68466 1 23
2 68467 1 23
2 68468 1 23
2 68469 1 23
2 68470 1 23
2 68471 1 23
2 68472 1 23
2 68473 1 23
2 68474 1 23
2 68475 1 23
2 68476 1 23
2 68477 1 23
2 68478 1 23
2 68479 1 23
2 68480 1 23
2 68481 1 23
2 68482 1 23
2 68483 1 23
2 68484 1 23
2 68485 1 23
2 68486 1 23
2 68487 1 23
2 68488 1 23
2 68489 1 23
2 68490 1 23
2 68491 1 23
2 68492 1 23
2 68493 1 23
2 68494 1 23
2 68495 1 23
2 68496 1 23
2 68497 1 23
2 68498 1 23
2 68499 1 23
2 68500 1 23
2 68501 1 23
2 68502 1 23
2 68503 1 23
2 68504 1 23
2 68505 1 23
2 68506 1 23
2 68507 1 23
2 68508 1 23
2 68509 1 23
2 68510 1 23
2 68511 1 23
2 68512 1 23
2 68513 1 23
2 68514 1 23
2 68515 1 23
2 68516 1 23
2 68517 1 23
2 68518 1 23
2 68519 1 23
2 68520 1 23
2 68521 1 23
2 68522 1 23
2 68523 1 23
2 68524 1 23
2 68525 1 23
2 68526 1 23
2 68527 1 23
2 68528 1 23
2 68529 1 23
2 68530 1 23
2 68531 1 23
2 68532 1 23
2 68533 1 23
2 68534 1 23
2 68535 1 23
2 68536 1 23
2 68537 1 23
2 68538 1 23
2 68539 1 23
2 68540 1 23
1 24 0 202 0
2 68541 1 24
2 68542 1 24
2 68543 1 24
2 68544 1 24
2 68545 1 24
2 68546 1 24
2 68547 1 24
2 68548 1 24
2 68549 1 24
2 68550 1 24
2 68551 1 24
2 68552 1 24
2 68553 1 24
2 68554 1 24
2 68555 1 24
2 68556 1 24
2 68557 1 24
2 68558 1 24
2 68559 1 24
2 68560 1 24
2 68561 1 24
2 68562 1 24
2 68563 1 24
2 68564 1 24
2 68565 1 24
2 68566 1 24
2 68567 1 24
2 68568 1 24
2 68569 1 24
2 68570 1 24
2 68571 1 24
2 68572 1 24
2 68573 1 24
2 68574 1 24
2 68575 1 24
2 68576 1 24
2 68577 1 24
2 68578 1 24
2 68579 1 24
2 68580 1 24
2 68581 1 24
2 68582 1 24
2 68583 1 24
2 68584 1 24
2 68585 1 24
2 68586 1 24
2 68587 1 24
2 68588 1 24
2 68589 1 24
2 68590 1 24
2 68591 1 24
2 68592 1 24
2 68593 1 24
2 68594 1 24
2 68595 1 24
2 68596 1 24
2 68597 1 24
2 68598 1 24
2 68599 1 24
2 68600 1 24
2 68601 1 24
2 68602 1 24
2 68603 1 24
2 68604 1 24
2 68605 1 24
2 68606 1 24
2 68607 1 24
2 68608 1 24
2 68609 1 24
2 68610 1 24
2 68611 1 24
2 68612 1 24
2 68613 1 24
2 68614 1 24
2 68615 1 24
2 68616 1 24
2 68617 1 24
2 68618 1 24
2 68619 1 24
2 68620 1 24
2 68621 1 24
2 68622 1 24
2 68623 1 24
2 68624 1 24
2 68625 1 24
2 68626 1 24
2 68627 1 24
2 68628 1 24
2 68629 1 24
2 68630 1 24
2 68631 1 24
2 68632 1 24
2 68633 1 24
2 68634 1 24
2 68635 1 24
2 68636 1 24
2 68637 1 24
2 68638 1 24
2 68639 1 24
2 68640 1 24
2 68641 1 24
2 68642 1 24
2 68643 1 24
2 68644 1 24
2 68645 1 24
2 68646 1 24
2 68647 1 24
2 68648 1 24
2 68649 1 24
2 68650 1 24
2 68651 1 24
2 68652 1 24
2 68653 1 24
2 68654 1 24
2 68655 1 24
2 68656 1 24
2 68657 1 24
2 68658 1 24
2 68659 1 24
2 68660 1 24
2 68661 1 24
2 68662 1 24
2 68663 1 24
2 68664 1 24
2 68665 1 24
2 68666 1 24
2 68667 1 24
2 68668 1 24
2 68669 1 24
2 68670 1 24
2 68671 1 24
2 68672 1 24
2 68673 1 24
2 68674 1 24
2 68675 1 24
2 68676 1 24
2 68677 1 24
2 68678 1 24
2 68679 1 24
2 68680 1 24
2 68681 1 24
2 68682 1 24
2 68683 1 24
2 68684 1 24
2 68685 1 24
2 68686 1 24
2 68687 1 24
2 68688 1 24
2 68689 1 24
2 68690 1 24
2 68691 1 24
2 68692 1 24
2 68693 1 24
2 68694 1 24
2 68695 1 24
2 68696 1 24
2 68697 1 24
2 68698 1 24
2 68699 1 24
2 68700 1 24
2 68701 1 24
2 68702 1 24
2 68703 1 24
2 68704 1 24
2 68705 1 24
2 68706 1 24
2 68707 1 24
2 68708 1 24
2 68709 1 24
2 68710 1 24
2 68711 1 24
2 68712 1 24
2 68713 1 24
2 68714 1 24
2 68715 1 24
2 68716 1 24
2 68717 1 24
2 68718 1 24
2 68719 1 24
2 68720 1 24
2 68721 1 24
2 68722 1 24
2 68723 1 24
2 68724 1 24
2 68725 1 24
2 68726 1 24
2 68727 1 24
2 68728 1 24
2 68729 1 24
2 68730 1 24
2 68731 1 24
2 68732 1 24
2 68733 1 24
2 68734 1 24
2 68735 1 24
2 68736 1 24
2 68737 1 24
2 68738 1 24
2 68739 1 24
2 68740 1 24
2 68741 1 24
2 68742 1 24
2 68743 1 27
2 68744 1 27
2 68745 1 27
2 68746 1 27
2 68747 1 27
2 68748 1 27
2 68749 1 27
2 68750 1 27
2 68751 1 27
2 68752 1 27
2 68753 1 27
2 68754 1 27
2 68755 1 27
2 68756 1 27
2 68757 1 27
2 68758 1 27
2 68759 1 27
2 68760 1 27
2 68761 1 27
2 68762 1 27
2 68763 1 27
2 68764 1 27
2 68765 1 27
2 68766 1 27
2 68767 1 27
2 68768 1 27
2 68769 1 27
2 68770 1 27
2 68771 1 27
2 68772 1 27
2 68773 1 27
2 68774 1 27
2 68775 1 27
2 68776 1 27
2 68777 1 27
2 68778 1 27
2 68779 1 27
2 68780 1 27
2 68781 1 27
2 68782 1 27
2 68783 1 27
2 68784 1 27
2 68785 1 27
2 68786 1 27
2 68787 1 27
2 68788 1 27
2 68789 1 27
2 68790 1 27
2 68791 1 27
2 68792 1 27
2 68793 1 27
2 68794 1 27
2 68795 1 27
2 68796 1 27
2 68797 1 27
2 68798 1 27
2 68799 1 27
2 68800 1 27
2 68801 1 27
2 68802 1 27
2 68803 1 27
2 68804 1 27
2 68805 1 27
2 68806 1 27
2 68807 1 27
2 68808 1 27
2 68809 1 27
2 68810 1 27
2 68811 1 27
2 68812 1 27
2 68813 1 27
2 68814 1 27
2 68815 1 27
2 68816 1 27
2 68817 1 27
2 68818 1 27
2 68819 1 27
2 68820 1 27
2 68821 1 27
2 68822 1 27
2 68823 1 27
2 68824 1 27
2 68825 1 27
2 68826 1 27
2 68827 1 27
2 68828 1 27
2 68829 1 27
2 68830 1 27
2 68831 1 27
2 68832 1 27
2 68833 1 27
2 68834 1 27
2 68835 1 27
2 68836 1 27
2 68837 1 27
2 68838 1 27
2 68839 1 27
2 68840 1 27
2 68841 1 27
2 68842 1 27
2 68843 1 27
2 68844 1 27
2 68845 1 27
2 68846 1 27
2 68847 1 27
2 68848 1 27
2 68849 1 27
2 68850 1 27
2 68851 1 27
2 68852 1 27
2 68853 1 27
2 68854 1 27
2 68855 1 27
2 68856 1 27
2 68857 1 27
2 68858 1 27
2 68859 1 27
2 68860 1 27
2 68861 1 27
2 68862 1 27
2 68863 1 27
2 68864 1 27
2 68865 1 27
2 68866 1 27
2 68867 1 27
2 68868 1 27
2 68869 1 27
2 68870 1 27
2 68871 1 27
2 68872 1 27
2 68873 1 27
2 68874 1 27
2 68875 1 27
2 68876 1 27
2 68877 1 27
2 68878 1 27
2 68879 1 27
2 68880 1 27
2 68881 1 27
2 68882 1 27
2 68883 1 27
2 68884 1 27
2 68885 1 27
2 68886 1 27
2 68887 1 27
2 68888 1 27
2 68889 1 27
2 68890 1 27
2 68891 1 27
2 68892 1 27
2 68893 1 27
2 68894 1 27
2 68895 1 27
2 68896 1 27
2 68897 1 27
2 68898 1 27
2 68899 1 27
2 68900 1 27
2 68901 1 27
2 68902 1 27
2 68903 1 27
2 68904 1 27
2 68905 1 27
2 68906 1 27
2 68907 1 27
2 68908 1 28
2 68909 1 28
2 68910 1 28
2 68911 1 28
2 68912 1 28
2 68913 1 28
2 68914 1 28
2 68915 1 28
2 68916 1 28
2 68917 1 28
2 68918 1 28
2 68919 1 28
2 68920 1 28
2 68921 1 28
2 68922 1 28
2 68923 1 28
2 68924 1 28
2 68925 1 28
2 68926 1 28
2 68927 1 28
2 68928 1 28
2 68929 1 28
2 68930 1 28
2 68931 1 28
2 68932 1 28
2 68933 1 28
2 68934 1 28
2 68935 1 28
2 68936 1 28
2 68937 1 28
2 68938 1 28
2 68939 1 28
2 68940 1 28
2 68941 1 28
2 68942 1 28
2 68943 1 28
2 68944 1 28
2 68945 1 28
2 68946 1 28
2 68947 1 28
2 68948 1 28
2 68949 1 28
2 68950 1 28
2 68951 1 28
2 68952 1 28
2 68953 1 28
2 68954 1 28
2 68955 1 28
2 68956 1 28
2 68957 1 28
2 68958 1 28
2 68959 1 28
2 68960 1 28
2 68961 1 28
2 68962 1 28
2 68963 1 28
2 68964 1 28
2 68965 1 28
2 68966 1 28
2 68967 1 28
2 68968 1 28
2 68969 1 28
2 68970 1 28
2 68971 1 28
2 68972 1 28
2 68973 1 28
2 68974 1 28
2 68975 1 28
2 68976 1 28
2 68977 1 28
2 68978 1 28
2 68979 1 28
2 68980 1 28
2 68981 1 28
2 68982 1 28
2 68983 1 28
2 68984 1 28
2 68985 1 28
2 68986 1 28
2 68987 1 28
2 68988 1 28
2 68989 1 28
2 68990 1 28
2 68991 1 28
2 68992 1 28
2 68993 1 28
2 68994 1 28
2 68995 1 28
2 68996 1 28
2 68997 1 28
2 68998 1 28
2 68999 1 28
2 69000 1 28
2 69001 1 28
2 69002 1 28
2 69003 1 28
2 69004 1 28
2 69005 1 28
2 69006 1 28
2 69007 1 28
2 69008 1 28
2 69009 1 28
2 69010 1 28
2 69011 1 28
2 69012 1 28
2 69013 1 28
2 69014 1 28
2 69015 1 28
2 69016 1 28
2 69017 1 28
2 69018 1 28
2 69019 1 28
2 69020 1 28
2 69021 1 28
2 69022 1 28
2 69023 1 28
2 69024 1 28
2 69025 1 28
2 69026 1 28
2 69027 1 28
2 69028 1 28
2 69029 1 28
2 69030 1 28
2 69031 1 28
2 69032 1 28
2 69033 1 28
2 69034 1 28
2 69035 1 28
2 69036 1 28
2 69037 1 28
2 69038 1 28
2 69039 1 28
2 69040 1 29
2 69041 1 29
2 69042 1 29
2 69043 1 29
2 69044 1 29
2 69045 1 29
2 69046 1 29
2 69047 1 29
2 69048 1 29
2 69049 1 29
2 69050 1 29
2 69051 1 29
2 69052 1 29
2 69053 1 29
2 69054 1 29
2 69055 1 29
2 69056 1 29
2 69057 1 29
2 69058 1 29
2 69059 1 29
2 69060 1 29
2 69061 1 29
2 69062 1 29
2 69063 1 29
2 69064 1 29
2 69065 1 29
2 69066 1 29
2 69067 1 29
2 69068 1 29
2 69069 1 29
2 69070 1 29
2 69071 1 29
2 69072 1 29
2 69073 1 29
2 69074 1 29
2 69075 1 29
2 69076 1 29
2 69077 1 29
2 69078 1 29
2 69079 1 29
2 69080 1 29
2 69081 1 29
2 69082 1 29
2 69083 1 29
2 69084 1 29
2 69085 1 29
2 69086 1 29
2 69087 1 29
2 69088 1 29
2 69089 1 29
2 69090 1 29
2 69091 1 30
2 69092 1 30
2 69093 1 30
2 69094 1 30
2 69095 1 30
2 69096 1 30
2 69097 1 30
2 69098 1 30
2 69099 1 30
2 69100 1 30
2 69101 1 30
2 69102 1 30
2 69103 1 30
2 69104 1 30
2 69105 1 30
2 69106 1 30
2 69107 1 30
2 69108 1 30
2 69109 1 30
2 69110 1 30
2 69111 1 30
2 69112 1 30
2 69113 1 30
2 69114 1 30
2 69115 1 30
2 69116 1 30
2 69117 1 30
2 69118 1 30
2 69119 1 30
2 69120 1 30
2 69121 1 30
2 69122 1 30
2 69123 1 30
2 69124 1 30
2 69125 1 30
2 69126 1 30
2 69127 1 30
2 69128 1 30
2 69129 1 30
2 69130 1 30
2 69131 1 30
2 69132 1 30
2 69133 1 30
2 69134 1 30
2 69135 1 30
2 69136 1 30
2 69137 1 30
2 69138 1 30
2 69139 1 30
2 69140 1 30
2 69141 1 30
2 69142 1 30
2 69143 1 30
2 69144 1 30
2 69145 1 30
2 69146 1 30
2 69147 1 30
2 69148 1 30
2 69149 1 30
2 69150 1 30
2 69151 1 30
2 69152 1 30
2 69153 1 30
2 69154 1 30
2 69155 1 30
2 69156 1 30
2 69157 1 30
2 69158 1 30
2 69159 1 30
2 69160 1 30
2 69161 1 30
2 69162 1 30
2 69163 1 30
2 69164 1 30
2 69165 1 30
2 69166 1 30
2 69167 1 30
2 69168 1 30
2 69169 1 30
2 69170 1 30
2 69171 1 30
2 69172 1 30
2 69173 1 30
2 69174 1 30
2 69175 1 30
2 69176 1 30
2 69177 1 30
2 69178 1 30
2 69179 1 30
2 69180 1 30
2 69181 1 30
2 69182 1 30
2 69183 1 30
2 69184 1 30
2 69185 1 30
2 69186 1 30
2 69187 1 30
2 69188 1 30
2 69189 1 30
2 69190 1 30
2 69191 1 30
2 69192 1 30
2 69193 1 30
2 69194 1 30
2 69195 1 30
2 69196 1 30
2 69197 1 30
2 69198 1 30
2 69199 1 30
2 69200 1 30
2 69201 1 30
2 69202 1 30
2 69203 1 30
2 69204 1 30
2 69205 1 30
2 69206 1 30
2 69207 1 30
2 69208 1 30
2 69209 1 30
2 69210 1 30
2 69211 1 30
2 69212 1 30
2 69213 1 30
2 69214 1 30
2 69215 1 30
2 69216 1 30
2 69217 1 30
2 69218 1 30
2 69219 1 30
2 69220 1 30
2 69221 1 30
2 69222 1 30
2 69223 1 30
2 69224 1 30
2 69225 1 30
2 69226 1 30
2 69227 1 30
2 69228 1 30
2 69229 1 30
2 69230 1 30
2 69231 1 30
2 69232 1 30
2 69233 1 30
2 69234 1 30
2 69235 1 30
2 69236 1 30
2 69237 1 30
2 69238 1 30
2 69239 1 30
2 69240 1 30
2 69241 1 30
2 69242 1 30
2 69243 1 30
2 69244 1 30
2 69245 1 30
2 69246 1 30
2 69247 1 30
2 69248 1 30
2 69249 1 30
2 69250 1 30
2 69251 1 30
2 69252 1 30
2 69253 1 30
2 69254 1 30
2 69255 1 30
2 69256 1 30
2 69257 1 30
2 69258 1 30
2 69259 1 30
2 69260 1 30
2 69261 1 30
2 69262 1 30
2 69263 1 30
2 69264 1 30
2 69265 1 30
2 69266 1 30
2 69267 1 30
2 69268 1 30
2 69269 1 30
2 69270 1 30
2 69271 1 30
2 69272 1 30
2 69273 1 30
2 69274 1 30
2 69275 1 30
2 69276 1 30
2 69277 1 30
2 69278 1 30
2 69279 1 30
2 69280 1 30
2 69281 1 30
2 69282 1 30
2 69283 1 30
2 69284 1 30
2 69285 1 30
2 69286 1 30
2 69287 1 30
2 69288 1 30
2 69289 1 30
2 69290 1 30
2 69291 1 30
2 69292 1 30
2 69293 1 30
2 69294 1 30
2 69295 1 30
2 69296 1 30
2 69297 1 30
2 69298 1 30
2 69299 1 30
2 69300 1 30
2 69301 1 30
2 69302 1 30
2 69303 1 30
2 69304 1 30
2 69305 1 30
2 69306 1 30
2 69307 1 30
2 69308 1 30
2 69309 1 30
2 69310 1 30
2 69311 1 30
2 69312 1 30
2 69313 1 30
2 69314 1 30
2 69315 1 30
2 69316 1 30
2 69317 1 30
2 69318 1 30
2 69319 1 30
2 69320 1 30
2 69321 1 30
2 69322 1 30
2 69323 1 30
2 69324 1 30
2 69325 1 30
2 69326 1 30
2 69327 1 30
2 69328 1 30
2 69329 1 30
2 69330 1 30
2 69331 1 30
2 69332 1 30
2 69333 1 31
2 69334 1 31
2 69335 1 31
2 69336 1 31
2 69337 1 31
2 69338 1 31
2 69339 1 31
2 69340 1 31
2 69341 1 31
2 69342 1 31
2 69343 1 31
2 69344 1 31
2 69345 1 31
2 69346 1 31
2 69347 1 31
2 69348 1 31
2 69349 1 31
2 69350 1 31
2 69351 1 31
2 69352 1 31
2 69353 1 31
2 69354 1 31
2 69355 1 31
2 69356 1 31
2 69357 1 31
2 69358 1 31
2 69359 1 31
2 69360 1 31
2 69361 1 31
2 69362 1 31
2 69363 1 31
2 69364 1 31
2 69365 1 31
2 69366 1 31
2 69367 1 31
2 69368 1 31
2 69369 1 31
2 69370 1 31
2 69371 1 31
2 69372 1 31
2 69373 1 31
2 69374 1 31
2 69375 1 31
2 69376 1 31
2 69377 1 31
2 69378 1 31
2 69379 1 31
2 69380 1 31
2 69381 1 31
2 69382 1 31
2 69383 1 31
2 69384 1 31
2 69385 1 31
2 69386 1 31
2 69387 1 31
2 69388 1 31
2 69389 1 31
2 69390 1 31
2 69391 1 31
2 69392 1 31
2 69393 1 31
2 69394 1 31
2 69395 1 31
2 69396 1 31
2 69397 1 31
2 69398 1 31
2 69399 1 31
2 69400 1 31
2 69401 1 31
2 69402 1 31
2 69403 1 31
2 69404 1 31
2 69405 1 31
2 69406 1 31
2 69407 1 31
2 69408 1 31
2 69409 1 31
2 69410 1 31
2 69411 1 31
2 69412 1 31
2 69413 1 31
2 69414 1 31
2 69415 1 31
2 69416 1 31
2 69417 1 31
2 69418 1 31
2 69419 1 31
2 69420 1 31
2 69421 1 31
2 69422 1 31
2 69423 1 31
2 69424 1 31
2 69425 1 31
2 69426 1 31
2 69427 1 31
2 69428 1 31
2 69429 1 31
2 69430 1 31
2 69431 1 31
2 69432 1 31
2 69433 1 31
2 69434 1 31
2 69435 1 31
2 69436 1 31
2 69437 1 31
2 69438 1 31
2 69439 1 31
2 69440 1 31
2 69441 1 31
2 69442 1 31
2 69443 1 31
2 69444 1 31
2 69445 1 31
2 69446 1 31
2 69447 1 31
2 69448 1 31
2 69449 1 31
2 69450 1 31
2 69451 1 31
2 69452 1 31
2 69453 1 31
2 69454 1 31
2 69455 1 31
2 69456 1 31
2 69457 1 31
2 69458 1 31
2 69459 1 31
2 69460 1 31
2 69461 1 31
2 69462 1 31
2 69463 1 31
2 69464 1 31
2 69465 1 31
2 69466 1 31
2 69467 1 31
2 69468 1 31
2 69469 1 31
2 69470 1 31
2 69471 1 31
2 69472 1 31
2 69473 1 31
2 69474 1 31
2 69475 1 31
2 69476 1 31
2 69477 1 31
2 69478 1 31
2 69479 1 31
2 69480 1 31
2 69481 1 31
2 69482 1 31
2 69483 1 31
2 69484 1 31
2 69485 1 31
2 69486 1 31
2 69487 1 31
2 69488 1 31
2 69489 1 31
2 69490 1 31
2 69491 1 31
2 69492 1 31
2 69493 1 31
2 69494 1 31
2 69495 1 31
2 69496 1 31
2 69497 1 31
2 69498 1 31
2 69499 1 31
2 69500 1 31
2 69501 1 31
2 69502 1 31
2 69503 1 31
2 69504 1 31
2 69505 1 31
2 69506 1 31
2 69507 1 31
2 69508 1 31
2 69509 1 31
2 69510 1 31
2 69511 1 31
2 69512 1 31
2 69513 1 31
2 69514 1 31
2 69515 1 31
2 69516 1 31
2 69517 1 31
2 69518 1 31
2 69519 1 31
2 69520 1 31
2 69521 1 31
2 69522 1 31
2 69523 1 31
2 69524 1 31
2 69525 1 31
2 69526 1 31
2 69527 1 31
2 69528 1 31
2 69529 1 31
2 69530 1 31
2 69531 1 31
2 69532 1 31
2 69533 1 31
2 69534 1 31
2 69535 1 31
2 69536 1 31
2 69537 1 31
2 69538 1 31
2 69539 1 31
2 69540 1 31
2 69541 1 31
2 69542 1 31
2 69543 1 31
2 69544 1 31
2 69545 1 31
2 69546 1 31
2 69547 1 31
2 69548 1 31
2 69549 1 31
2 69550 1 31
2 69551 1 31
2 69552 1 31
2 69553 1 31
2 69554 1 31
2 69555 1 31
2 69556 1 31
2 69557 1 31
2 69558 1 31
2 69559 1 31
2 69560 1 31
2 69561 1 31
2 69562 1 31
2 69563 1 31
2 69564 1 31
2 69565 1 31
2 69566 1 31
2 69567 1 31
2 69568 1 31
2 69569 1 31
2 69570 1 31
2 69571 1 31
2 69572 1 31
2 69573 1 31
2 69574 1 31
2 69575 1 31
2 69576 1 31
2 69577 1 31
2 69578 1 31
2 69579 1 31
2 69580 1 31
2 69581 1 31
2 69582 1 31
2 69583 1 31
2 69584 1 31
2 69585 1 31
2 69586 1 31
2 69587 1 31
2 69588 1 31
2 69589 1 31
2 69590 1 31
2 69591 1 31
2 69592 1 31
2 69593 1 31
2 69594 1 31
2 69595 1 31
2 69596 1 31
2 69597 1 31
2 69598 1 31
2 69599 1 31
2 69600 1 31
2 69601 1 31
2 69602 1 31
2 69603 1 31
2 69604 1 31
2 69605 1 31
2 69606 1 31
2 69607 1 31
2 69608 1 31
2 69609 1 31
2 69610 1 31
2 69611 1 31
2 69612 1 31
2 69613 1 31
2 69614 1 31
2 69615 1 31
2 69616 1 31
2 69617 1 31
2 69618 1 31
2 69619 1 31
2 69620 1 31
2 69621 1 31
2 69622 1 31
2 69623 1 31
2 69624 1 31
2 69625 1 31
2 69626 1 31
2 69627 1 31
2 69628 1 31
2 69629 1 31
2 69630 1 31
2 69631 1 31
2 69632 1 31
2 69633 1 31
2 69634 1 31
2 69635 1 31
2 69636 1 31
2 69637 1 31
2 69638 1 31
2 69639 1 31
2 69640 1 31
2 69641 1 31
2 69642 1 31
2 69643 1 31
2 69644 1 31
2 69645 1 31
2 69646 1 31
2 69647 1 31
2 69648 1 31
2 69649 1 31
2 69650 1 31
2 69651 1 31
2 69652 1 31
2 69653 1 31
2 69654 1 31
2 69655 1 31
2 69656 1 31
2 69657 1 31
2 69658 1 31
2 69659 1 31
2 69660 1 31
2 69661 1 31
2 69662 1 31
2 69663 1 31
2 69664 1 31
2 69665 1 31
2 69666 1 31
2 69667 1 31
2 69668 1 31
2 69669 1 31
2 69670 1 31
2 69671 1 31
2 69672 1 31
2 69673 1 31
2 69674 1 31
2 69675 1 31
2 69676 1 31
2 69677 1 32
2 69678 1 32
2 69679 1 32
2 69680 1 32
2 69681 1 32
2 69682 1 32
2 69683 1 32
2 69684 1 32
2 69685 1 32
2 69686 1 32
2 69687 1 32
2 69688 1 32
2 69689 1 32
2 69690 1 32
2 69691 1 32
2 69692 1 32
2 69693 1 32
2 69694 1 32
2 69695 1 32
2 69696 1 32
2 69697 1 32
2 69698 1 32
2 69699 1 32
2 69700 1 32
2 69701 1 32
2 69702 1 32
2 69703 1 32
2 69704 1 32
2 69705 1 32
2 69706 1 32
2 69707 1 32
2 69708 1 32
2 69709 1 32
2 69710 1 32
2 69711 1 32
2 69712 1 32
2 69713 1 32
2 69714 1 32
2 69715 1 32
2 69716 1 32
2 69717 1 32
2 69718 1 32
2 69719 1 32
2 69720 1 32
2 69721 1 32
2 69722 1 32
2 69723 1 32
2 69724 1 32
2 69725 1 32
2 69726 1 32
2 69727 1 32
2 69728 1 32
2 69729 1 32
2 69730 1 32
2 69731 1 32
2 69732 1 32
2 69733 1 32
2 69734 1 32
2 69735 1 32
2 69736 1 32
2 69737 1 32
2 69738 1 32
2 69739 1 32
2 69740 1 32
2 69741 1 32
2 69742 1 32
2 69743 1 32
2 69744 1 32
2 69745 1 32
2 69746 1 32
2 69747 1 32
2 69748 1 32
2 69749 1 32
2 69750 1 32
2 69751 1 32
2 69752 1 32
2 69753 1 32
2 69754 1 32
2 69755 1 32
2 69756 1 32
2 69757 1 32
2 69758 1 32
2 69759 1 32
2 69760 1 32
2 69761 1 32
2 69762 1 32
2 69763 1 32
2 69764 1 32
2 69765 1 32
2 69766 1 32
2 69767 1 32
2 69768 1 32
2 69769 1 32
2 69770 1 32
2 69771 1 32
2 69772 1 32
2 69773 1 32
2 69774 1 32
2 69775 1 32
2 69776 1 32
2 69777 1 32
2 69778 1 32
2 69779 1 32
2 69780 1 32
2 69781 1 32
2 69782 1 32
2 69783 1 32
2 69784 1 32
2 69785 1 32
2 69786 1 32
2 69787 1 32
2 69788 1 32
2 69789 1 32
2 69790 1 32
2 69791 1 32
2 69792 1 32
2 69793 1 32
2 69794 1 32
2 69795 1 32
2 69796 1 32
2 69797 1 32
2 69798 1 32
2 69799 1 32
2 69800 1 32
2 69801 1 32
2 69802 1 32
2 69803 1 32
2 69804 1 32
2 69805 1 32
2 69806 1 32
2 69807 1 32
2 69808 1 32
2 69809 1 32
2 69810 1 32
2 69811 1 32
2 69812 1 32
2 69813 1 32
2 69814 1 32
2 69815 1 32
2 69816 1 32
2 69817 1 32
2 69818 1 32
2 69819 1 32
2 69820 1 32
2 69821 1 32
2 69822 1 32
2 69823 1 32
2 69824 1 32
2 69825 1 32
2 69826 1 32
2 69827 1 32
2 69828 1 32
2 69829 1 32
2 69830 1 32
2 69831 1 32
2 69832 1 32
2 69833 1 32
2 69834 1 32
2 69835 1 32
2 69836 1 32
2 69837 1 32
2 69838 1 32
2 69839 1 32
2 69840 1 32
2 69841 1 32
2 69842 1 32
2 69843 1 32
2 69844 1 32
2 69845 1 32
2 69846 1 32
2 69847 1 32
2 69848 1 32
2 69849 1 32
2 69850 1 32
2 69851 1 32
2 69852 1 32
2 69853 1 32
2 69854 1 32
2 69855 1 32
2 69856 1 32
2 69857 1 32
2 69858 1 32
2 69859 1 32
2 69860 1 32
2 69861 1 32
2 69862 1 32
2 69863 1 32
2 69864 1 32
2 69865 1 32
2 69866 1 32
2 69867 1 32
2 69868 1 32
2 69869 1 32
2 69870 1 32
2 69871 1 32
2 69872 1 32
2 69873 1 32
2 69874 1 32
2 69875 1 32
2 69876 1 32
2 69877 1 32
2 69878 1 32
2 69879 1 32
2 69880 1 32
2 69881 1 32
2 69882 1 32
2 69883 1 32
2 69884 1 32
2 69885 1 32
2 69886 1 32
2 69887 1 32
2 69888 1 32
2 69889 1 32
2 69890 1 32
2 69891 1 32
2 69892 1 32
2 69893 1 32
2 69894 1 32
2 69895 1 32
2 69896 1 32
2 69897 1 32
2 69898 1 32
2 69899 1 32
2 69900 1 32
2 69901 1 32
2 69902 1 32
2 69903 1 32
2 69904 1 32
2 69905 1 32
2 69906 1 32
2 69907 1 32
2 69908 1 32
2 69909 1 32
2 69910 1 32
2 69911 1 32
2 69912 1 32
2 69913 1 32
2 69914 1 32
2 69915 1 32
2 69916 1 32
2 69917 1 32
2 69918 1 32
2 69919 1 32
2 69920 1 32
2 69921 1 32
2 69922 1 32
2 69923 1 32
2 69924 1 32
2 69925 1 32
2 69926 1 32
2 69927 1 32
2 69928 1 32
2 69929 1 32
2 69930 1 32
2 69931 1 32
2 69932 1 32
2 69933 1 32
2 69934 1 32
2 69935 1 32
2 69936 1 32
2 69937 1 32
2 69938 1 32
2 69939 1 32
2 69940 1 32
2 69941 1 32
2 69942 1 32
2 69943 1 32
2 69944 1 32
2 69945 1 32
2 69946 1 32
2 69947 1 32
2 69948 1 32
2 69949 1 32
2 69950 1 32
2 69951 1 32
2 69952 1 32
2 69953 1 32
2 69954 1 32
2 69955 1 32
2 69956 1 32
2 69957 1 32
2 69958 1 32
2 69959 1 32
2 69960 1 32
2 69961 1 32
2 69962 1 32
2 69963 1 32
2 69964 1 32
2 69965 1 32
2 69966 1 32
2 69967 1 32
2 69968 1 32
2 69969 1 32
2 69970 1 32
2 69971 1 32
2 69972 1 32
2 69973 1 32
2 69974 1 32
2 69975 1 32
2 69976 1 32
2 69977 1 32
2 69978 1 32
2 69979 1 32
2 69980 1 32
2 69981 1 32
2 69982 1 32
2 69983 1 32
2 69984 1 32
2 69985 1 32
2 69986 1 32
2 69987 1 32
2 69988 1 32
2 69989 1 32
2 69990 1 32
2 69991 1 32
2 69992 1 32
2 69993 1 32
2 69994 1 32
2 69995 1 32
2 69996 1 32
2 69997 1 32
2 69998 1 32
2 69999 1 32
2 70000 1 32
2 70001 1 32
2 70002 1 32
2 70003 1 32
2 70004 1 32
2 70005 1 32
2 70006 1 32
2 70007 1 32
2 70008 1 32
2 70009 1 32
2 70010 1 32
2 70011 1 32
2 70012 1 32
2 70013 1 32
2 70014 1 32
2 70015 1 32
2 70016 1 32
2 70017 1 32
2 70018 1 32
2 70019 1 32
2 70020 1 32
2 70021 1 32
2 70022 1 32
2 70023 1 32
2 70024 1 32
2 70025 1 32
2 70026 1 32
2 70027 1 32
2 70028 1 32
2 70029 1 32
2 70030 1 32
2 70031 1 32
2 70032 1 32
2 70033 1 32
2 70034 1 32
2 70035 1 32
2 70036 1 32
2 70037 1 32
2 70038 1 33
2 70039 1 33
2 70040 1 33
2 70041 1 33
2 70042 1 33
2 70043 1 33
2 70044 1 33
2 70045 1 33
2 70046 1 33
2 70047 1 33
2 70048 1 33
2 70049 1 33
2 70050 1 33
2 70051 1 33
2 70052 1 33
2 70053 1 33
2 70054 1 33
2 70055 1 33
2 70056 1 33
2 70057 1 33
2 70058 1 33
2 70059 1 33
2 70060 1 33
2 70061 1 33
2 70062 1 33
2 70063 1 33
2 70064 1 33
2 70065 1 33
2 70066 1 33
2 70067 1 33
2 70068 1 33
2 70069 1 33
2 70070 1 33
2 70071 1 33
2 70072 1 33
2 70073 1 33
2 70074 1 33
2 70075 1 33
2 70076 1 33
2 70077 1 33
2 70078 1 33
2 70079 1 33
2 70080 1 33
2 70081 1 33
2 70082 1 33
2 70083 1 33
2 70084 1 33
2 70085 1 33
2 70086 1 33
2 70087 1 33
2 70088 1 33
2 70089 1 33
2 70090 1 33
2 70091 1 33
2 70092 1 33
2 70093 1 33
2 70094 1 33
2 70095 1 33
2 70096 1 33
2 70097 1 33
2 70098 1 33
2 70099 1 33
2 70100 1 33
2 70101 1 33
2 70102 1 33
2 70103 1 33
2 70104 1 33
2 70105 1 33
2 70106 1 33
2 70107 1 33
2 70108 1 33
2 70109 1 33
2 70110 1 33
2 70111 1 33
2 70112 1 33
2 70113 1 33
2 70114 1 33
2 70115 1 33
2 70116 1 33
2 70117 1 33
2 70118 1 33
2 70119 1 33
2 70120 1 33
2 70121 1 33
2 70122 1 33
2 70123 1 33
2 70124 1 33
2 70125 1 33
2 70126 1 33
2 70127 1 33
2 70128 1 33
2 70129 1 33
2 70130 1 33
2 70131 1 33
2 70132 1 33
2 70133 1 33
2 70134 1 33
2 70135 1 33
2 70136 1 33
2 70137 1 33
2 70138 1 33
2 70139 1 33
2 70140 1 33
2 70141 1 33
2 70142 1 33
2 70143 1 33
2 70144 1 33
2 70145 1 33
2 70146 1 33
2 70147 1 33
2 70148 1 33
2 70149 1 33
2 70150 1 33
2 70151 1 33
2 70152 1 33
2 70153 1 33
2 70154 1 33
2 70155 1 33
2 70156 1 33
2 70157 1 33
2 70158 1 33
2 70159 1 33
2 70160 1 33
2 70161 1 33
2 70162 1 33
2 70163 1 33
2 70164 1 33
2 70165 1 33
2 70166 1 33
2 70167 1 33
2 70168 1 33
2 70169 1 33
2 70170 1 33
2 70171 1 33
2 70172 1 33
2 70173 1 33
2 70174 1 33
2 70175 1 33
2 70176 1 33
2 70177 1 33
2 70178 1 33
2 70179 1 33
2 70180 1 33
2 70181 1 33
2 70182 1 33
2 70183 1 33
2 70184 1 33
2 70185 1 33
2 70186 1 33
2 70187 1 33
2 70188 1 33
2 70189 1 33
2 70190 1 33
2 70191 1 33
2 70192 1 33
2 70193 1 33
2 70194 1 33
2 70195 1 33
2 70196 1 33
2 70197 1 33
2 70198 1 33
2 70199 1 33
2 70200 1 33
2 70201 1 33
2 70202 1 33
2 70203 1 33
2 70204 1 33
2 70205 1 33
2 70206 1 33
2 70207 1 33
2 70208 1 33
2 70209 1 33
2 70210 1 33
2 70211 1 33
2 70212 1 33
2 70213 1 33
2 70214 1 33
2 70215 1 33
2 70216 1 33
2 70217 1 33
2 70218 1 33
2 70219 1 33
2 70220 1 33
2 70221 1 33
2 70222 1 33
2 70223 1 33
2 70224 1 33
2 70225 1 33
2 70226 1 33
2 70227 1 33
2 70228 1 33
2 70229 1 33
2 70230 1 33
2 70231 1 33
2 70232 1 33
2 70233 1 33
2 70234 1 33
2 70235 1 33
2 70236 1 33
2 70237 1 33
2 70238 1 33
2 70239 1 33
2 70240 1 33
2 70241 1 33
2 70242 1 33
2 70243 1 33
2 70244 1 33
2 70245 1 33
2 70246 1 33
2 70247 1 33
2 70248 1 33
2 70249 1 33
2 70250 1 33
2 70251 1 33
2 70252 1 33
2 70253 1 33
2 70254 1 33
2 70255 1 33
2 70256 1 33
2 70257 1 33
2 70258 1 33
2 70259 1 33
2 70260 1 33
2 70261 1 33
2 70262 1 33
2 70263 1 33
2 70264 1 33
2 70265 1 33
2 70266 1 33
2 70267 1 33
2 70268 1 33
2 70269 1 33
2 70270 1 33
2 70271 1 33
2 70272 1 33
2 70273 1 33
2 70274 1 33
2 70275 1 33
2 70276 1 33
2 70277 1 33
2 70278 1 33
2 70279 1 33
2 70280 1 33
2 70281 1 33
2 70282 1 33
2 70283 1 33
2 70284 1 33
2 70285 1 33
2 70286 1 33
2 70287 1 33
2 70288 1 33
2 70289 1 33
2 70290 1 33
2 70291 1 33
2 70292 1 33
2 70293 1 33
2 70294 1 33
2 70295 1 33
2 70296 1 33
2 70297 1 33
2 70298 1 33
2 70299 1 33
2 70300 1 33
2 70301 1 33
2 70302 1 33
2 70303 1 33
2 70304 1 33
2 70305 1 33
2 70306 1 33
2 70307 1 33
2 70308 1 33
2 70309 1 34
2 70310 1 34
2 70311 1 34
2 70312 1 34
2 70313 1 34
2 70314 1 34
2 70315 1 34
2 70316 1 34
2 70317 1 34
2 70318 1 34
2 70319 1 34
2 70320 1 34
2 70321 1 34
2 70322 1 34
2 70323 1 34
2 70324 1 34
2 70325 1 34
2 70326 1 34
2 70327 1 34
2 70328 1 34
2 70329 1 34
2 70330 1 34
2 70331 1 34
2 70332 1 34
2 70333 1 34
2 70334 1 34
2 70335 1 34
2 70336 1 34
2 70337 1 34
2 70338 1 34
2 70339 1 34
2 70340 1 34
2 70341 1 34
2 70342 1 34
2 70343 1 34
2 70344 1 34
2 70345 1 34
2 70346 1 34
2 70347 1 34
2 70348 1 34
2 70349 1 34
2 70350 1 34
2 70351 1 34
2 70352 1 34
2 70353 1 34
2 70354 1 34
2 70355 1 34
2 70356 1 34
2 70357 1 34
2 70358 1 34
2 70359 1 34
2 70360 1 34
2 70361 1 34
2 70362 1 34
2 70363 1 34
2 70364 1 34
2 70365 1 34
2 70366 1 34
2 70367 1 34
2 70368 1 34
2 70369 1 34
2 70370 1 34
2 70371 1 34
2 70372 1 34
2 70373 1 34
2 70374 1 34
2 70375 1 34
2 70376 1 34
2 70377 1 34
2 70378 1 34
2 70379 1 34
2 70380 1 34
2 70381 1 34
2 70382 1 34
2 70383 1 34
2 70384 1 34
2 70385 1 34
2 70386 1 34
2 70387 1 34
2 70388 1 34
2 70389 1 34
2 70390 1 34
2 70391 1 34
2 70392 1 34
2 70393 1 34
2 70394 1 34
2 70395 1 34
2 70396 1 34
2 70397 1 34
2 70398 1 34
2 70399 1 34
2 70400 1 34
2 70401 1 34
2 70402 1 34
2 70403 1 34
2 70404 1 34
2 70405 1 34
2 70406 1 34
2 70407 1 34
2 70408 1 34
2 70409 1 34
2 70410 1 34
2 70411 1 34
2 70412 1 34
2 70413 1 34
2 70414 1 34
2 70415 1 34
2 70416 1 34
2 70417 1 34
2 70418 1 34
2 70419 1 34
2 70420 1 34
2 70421 1 34
2 70422 1 34
2 70423 1 34
2 70424 1 34
2 70425 1 34
2 70426 1 34
2 70427 1 34
2 70428 1 34
2 70429 1 34
2 70430 1 34
2 70431 1 34
2 70432 1 34
2 70433 1 34
2 70434 1 34
2 70435 1 34
2 70436 1 34
2 70437 1 34
2 70438 1 34
2 70439 1 34
2 70440 1 34
2 70441 1 34
2 70442 1 34
2 70443 1 34
2 70444 1 34
2 70445 1 34
2 70446 1 34
2 70447 1 34
2 70448 1 34
2 70449 1 34
2 70450 1 34
2 70451 1 34
2 70452 1 34
2 70453 1 34
2 70454 1 34
2 70455 1 34
2 70456 1 34
2 70457 1 34
2 70458 1 34
2 70459 1 34
2 70460 1 34
2 70461 1 34
2 70462 1 34
2 70463 1 34
2 70464 1 34
2 70465 1 34
2 70466 1 34
2 70467 1 34
2 70468 1 34
2 70469 1 34
2 70470 1 34
2 70471 1 34
2 70472 1 34
2 70473 1 34
2 70474 1 34
2 70475 1 34
2 70476 1 34
2 70477 1 34
2 70478 1 34
2 70479 1 34
2 70480 1 34
2 70481 1 34
2 70482 1 34
2 70483 1 34
2 70484 1 34
2 70485 1 34
2 70486 1 34
2 70487 1 34
2 70488 1 34
2 70489 1 34
2 70490 1 34
2 70491 1 34
2 70492 1 34
2 70493 1 34
2 70494 1 34
2 70495 1 34
2 70496 1 34
2 70497 1 34
2 70498 1 34
2 70499 1 34
2 70500 1 34
2 70501 1 34
2 70502 1 34
2 70503 1 34
2 70504 1 34
2 70505 1 34
2 70506 1 34
2 70507 1 34
2 70508 1 34
2 70509 1 34
2 70510 1 34
2 70511 1 34
2 70512 1 34
2 70513 1 34
2 70514 1 34
2 70515 1 34
2 70516 1 34
2 70517 1 34
2 70518 1 34
2 70519 1 34
2 70520 1 34
2 70521 1 34
2 70522 1 34
2 70523 1 34
2 70524 1 34
2 70525 1 34
2 70526 1 34
2 70527 1 34
2 70528 1 34
2 70529 1 34
2 70530 1 34
2 70531 1 34
2 70532 1 34
2 70533 1 34
2 70534 1 34
2 70535 1 34
2 70536 1 34
2 70537 1 34
2 70538 1 34
2 70539 1 34
2 70540 1 34
2 70541 1 34
2 70542 1 34
2 70543 1 34
2 70544 1 34
2 70545 1 34
2 70546 1 34
2 70547 1 34
2 70548 1 34
2 70549 1 34
2 70550 1 34
2 70551 1 34
2 70552 1 34
2 70553 1 34
2 70554 1 34
2 70555 1 34
2 70556 1 34
2 70557 1 34
2 70558 1 34
2 70559 1 34
2 70560 1 34
2 70561 1 34
2 70562 1 34
2 70563 1 34
2 70564 1 34
2 70565 1 34
2 70566 1 34
2 70567 1 34
2 70568 1 34
2 70569 1 34
2 70570 1 34
2 70571 1 34
2 70572 1 34
2 70573 1 34
2 70574 1 34
2 70575 1 34
2 70576 1 34
2 70577 1 34
2 70578 1 34
2 70579 1 34
2 70580 1 34
2 70581 1 34
2 70582 1 34
2 70583 1 34
2 70584 1 34
2 70585 1 34
2 70586 1 34
2 70587 1 35
2 70588 1 35
2 70589 1 35
2 70590 1 35
2 70591 1 35
2 70592 1 35
2 70593 1 35
2 70594 1 35
2 70595 1 35
2 70596 1 35
2 70597 1 35
2 70598 1 35
2 70599 1 35
2 70600 1 35
2 70601 1 35
2 70602 1 35
2 70603 1 35
2 70604 1 35
2 70605 1 35
2 70606 1 35
2 70607 1 35
2 70608 1 35
2 70609 1 35
2 70610 1 35
2 70611 1 35
2 70612 1 35
2 70613 1 35
2 70614 1 35
2 70615 1 35
2 70616 1 35
2 70617 1 35
2 70618 1 35
2 70619 1 35
2 70620 1 35
2 70621 1 35
2 70622 1 35
2 70623 1 35
2 70624 1 35
2 70625 1 35
2 70626 1 35
2 70627 1 35
2 70628 1 35
2 70629 1 35
2 70630 1 35
2 70631 1 35
2 70632 1 35
2 70633 1 35
2 70634 1 35
2 70635 1 35
2 70636 1 35
2 70637 1 35
2 70638 1 35
2 70639 1 35
2 70640 1 35
2 70641 1 35
2 70642 1 35
2 70643 1 35
2 70644 1 35
2 70645 1 35
2 70646 1 35
2 70647 1 35
2 70648 1 35
2 70649 1 35
2 70650 1 36
2 70651 1 36
2 70652 1 36
2 70653 1 36
2 70654 1 36
2 70655 1 36
2 70656 1 36
2 70657 1 36
2 70658 1 36
2 70659 1 36
2 70660 1 36
2 70661 1 36
2 70662 1 36
2 70663 1 36
2 70664 1 36
2 70665 1 36
2 70666 1 36
2 70667 1 36
2 70668 1 36
2 70669 1 36
2 70670 1 36
2 70671 1 36
2 70672 1 36
2 70673 1 36
2 70674 1 36
2 70675 1 36
2 70676 1 36
2 70677 1 36
2 70678 1 36
2 70679 1 36
2 70680 1 36
2 70681 1 36
2 70682 1 36
2 70683 1 36
2 70684 1 36
2 70685 1 36
2 70686 1 36
2 70687 1 36
2 70688 1 36
2 70689 1 36
2 70690 1 36
2 70691 1 36
2 70692 1 36
2 70693 1 36
2 70694 1 36
2 70695 1 36
2 70696 1 36
2 70697 1 36
2 70698 1 36
2 70699 1 36
2 70700 1 36
2 70701 1 37
2 70702 1 37
2 70703 1 37
2 70704 1 37
2 70705 1 37
2 70706 1 37
2 70707 1 37
2 70708 1 37
2 70709 1 37
2 70710 1 37
2 70711 1 37
2 70712 1 37
2 70713 1 37
2 70714 1 37
2 70715 1 37
2 70716 1 37
2 70717 1 37
2 70718 1 37
2 70719 1 37
2 70720 1 37
2 70721 1 37
2 70722 1 37
2 70723 1 37
2 70724 1 37
2 70725 1 37
2 70726 1 37
2 70727 1 37
2 70728 1 37
2 70729 1 37
2 70730 1 37
2 70731 1 37
2 70732 1 37
2 70733 1 37
2 70734 1 37
2 70735 1 37
2 70736 1 37
2 70737 1 37
2 70738 1 37
2 70739 1 37
2 70740 1 37
2 70741 1 37
2 70742 1 37
2 70743 1 37
2 70744 1 37
2 70745 1 37
2 70746 1 37
2 70747 1 37
2 70748 1 37
2 70749 1 37
2 70750 1 37
2 70751 1 37
2 70752 1 37
2 70753 1 37
2 70754 1 37
2 70755 1 37
2 70756 1 38
2 70757 1 38
2 70758 1 38
2 70759 1 38
2 70760 1 38
2 70761 1 38
2 70762 1 38
2 70763 1 38
2 70764 1 38
2 70765 1 38
2 70766 1 38
2 70767 1 38
2 70768 1 38
2 70769 1 38
2 70770 1 38
2 70771 1 38
2 70772 1 38
2 70773 1 38
2 70774 1 38
2 70775 1 38
2 70776 1 38
2 70777 1 38
2 70778 1 38
2 70779 1 38
2 70780 1 38
2 70781 1 38
2 70782 1 38
2 70783 1 38
2 70784 1 38
2 70785 1 38
2 70786 1 38
2 70787 1 38
2 70788 1 38
2 70789 1 38
2 70790 1 38
2 70791 1 38
2 70792 1 38
2 70793 1 38
2 70794 1 38
2 70795 1 38
2 70796 1 38
2 70797 1 38
2 70798 1 38
2 70799 1 38
2 70800 1 38
2 70801 1 38
2 70802 1 38
2 70803 1 38
2 70804 1 38
2 70805 1 38
2 70806 1 38
2 70807 1 38
2 70808 1 38
2 70809 1 38
2 70810 1 38
2 70811 1 38
2 70812 1 38
2 70813 1 38
2 70814 1 38
2 70815 1 38
2 70816 1 38
2 70817 1 38
2 70818 1 38
2 70819 1 38
2 70820 1 38
2 70821 1 38
2 70822 1 38
2 70823 1 38
2 70824 1 38
2 70825 1 38
2 70826 1 38
2 70827 1 38
2 70828 1 38
2 70829 1 38
2 70830 1 38
2 70831 1 38
2 70832 1 38
2 70833 1 38
2 70834 1 38
2 70835 1 38
2 70836 1 38
2 70837 1 38
2 70838 1 38
2 70839 1 38
2 70840 1 38
2 70841 1 38
2 70842 1 38
2 70843 1 38
2 70844 1 38
2 70845 1 38
2 70846 1 38
2 70847 1 38
2 70848 1 38
2 70849 1 38
2 70850 1 38
2 70851 1 38
2 70852 1 38
2 70853 1 38
2 70854 1 38
2 70855 1 38
2 70856 1 38
2 70857 1 38
2 70858 1 38
2 70859 1 38
2 70860 1 38
2 70861 1 38
2 70862 1 38
2 70863 1 38
2 70864 1 38
2 70865 1 38
2 70866 1 38
2 70867 1 38
2 70868 1 38
2 70869 1 38
2 70870 1 38
2 70871 1 38
2 70872 1 38
2 70873 1 38
2 70874 1 38
2 70875 1 38
2 70876 1 38
2 70877 1 38
2 70878 1 38
2 70879 1 38
2 70880 1 38
2 70881 1 38
2 70882 1 38
2 70883 1 38
2 70884 1 38
2 70885 1 38
2 70886 1 38
2 70887 1 38
2 70888 1 38
2 70889 1 38
2 70890 1 38
2 70891 1 38
2 70892 1 38
2 70893 1 38
2 70894 1 38
2 70895 1 38
2 70896 1 38
2 70897 1 38
2 70898 1 38
2 70899 1 38
2 70900 1 38
2 70901 1 38
2 70902 1 38
2 70903 1 38
2 70904 1 38
2 70905 1 38
2 70906 1 38
2 70907 1 38
2 70908 1 38
2 70909 1 38
2 70910 1 38
2 70911 1 38
2 70912 1 38
2 70913 1 38
2 70914 1 38
2 70915 1 38
2 70916 1 38
2 70917 1 38
2 70918 1 38
2 70919 1 38
2 70920 1 38
2 70921 1 38
2 70922 1 38
2 70923 1 38
2 70924 1 38
2 70925 1 38
2 70926 1 38
2 70927 1 38
2 70928 1 38
2 70929 1 38
2 70930 1 38
2 70931 1 38
2 70932 1 38
2 70933 1 38
2 70934 1 38
2 70935 1 38
2 70936 1 39
2 70937 1 39
2 70938 1 39
2 70939 1 39
2 70940 1 39
2 70941 1 39
2 70942 1 39
2 70943 1 39
2 70944 1 39
2 70945 1 39
2 70946 1 39
2 70947 1 39
2 70948 1 39
2 70949 1 39
2 70950 1 39
2 70951 1 39
2 70952 1 39
2 70953 1 39
2 70954 1 39
2 70955 1 39
2 70956 1 39
2 70957 1 39
2 70958 1 39
2 70959 1 39
2 70960 1 39
2 70961 1 39
2 70962 1 39
2 70963 1 39
2 70964 1 39
2 70965 1 39
2 70966 1 39
2 70967 1 39
2 70968 1 39
2 70969 1 39
2 70970 1 39
2 70971 1 39
2 70972 1 39
2 70973 1 39
2 70974 1 39
2 70975 1 39
2 70976 1 39
2 70977 1 39
2 70978 1 39
2 70979 1 39
2 70980 1 39
2 70981 1 39
2 70982 1 39
2 70983 1 39
2 70984 1 39
2 70985 1 39
2 70986 1 39
2 70987 1 39
2 70988 1 39
2 70989 1 39
2 70990 1 39
2 70991 1 39
2 70992 1 39
2 70993 1 39
2 70994 1 39
2 70995 1 39
2 70996 1 39
2 70997 1 39
2 70998 1 39
2 70999 1 39
2 71000 1 39
2 71001 1 39
2 71002 1 39
2 71003 1 39
2 71004 1 39
2 71005 1 39
2 71006 1 39
2 71007 1 39
2 71008 1 39
2 71009 1 39
2 71010 1 39
2 71011 1 39
2 71012 1 39
2 71013 1 39
2 71014 1 39
2 71015 1 39
2 71016 1 39
2 71017 1 39
2 71018 1 39
2 71019 1 39
2 71020 1 39
2 71021 1 39
2 71022 1 39
2 71023 1 39
2 71024 1 39
2 71025 1 39
2 71026 1 39
2 71027 1 39
2 71028 1 39
2 71029 1 39
2 71030 1 39
2 71031 1 39
2 71032 1 39
2 71033 1 39
2 71034 1 39
2 71035 1 39
2 71036 1 39
2 71037 1 39
2 71038 1 39
2 71039 1 39
2 71040 1 39
2 71041 1 39
2 71042 1 39
2 71043 1 39
2 71044 1 39
2 71045 1 39
2 71046 1 39
2 71047 1 39
2 71048 1 39
2 71049 1 39
2 71050 1 39
2 71051 1 39
2 71052 1 39
2 71053 1 39
2 71054 1 39
2 71055 1 39
2 71056 1 39
2 71057 1 39
2 71058 1 39
2 71059 1 39
2 71060 1 39
2 71061 1 39
2 71062 1 39
2 71063 1 39
2 71064 1 39
2 71065 1 39
2 71066 1 39
2 71067 1 39
2 71068 1 39
2 71069 1 39
2 71070 1 39
2 71071 1 39
2 71072 1 39
2 71073 1 39
2 71074 1 39
2 71075 1 39
2 71076 1 39
2 71077 1 39
2 71078 1 39
2 71079 1 39
2 71080 1 39
2 71081 1 39
2 71082 1 39
2 71083 1 39
2 71084 1 39
2 71085 1 39
2 71086 1 39
2 71087 1 39
2 71088 1 39
2 71089 1 39
2 71090 1 39
2 71091 1 39
2 71092 1 39
2 71093 1 39
2 71094 1 39
2 71095 1 39
2 71096 1 39
2 71097 1 39
2 71098 1 39
2 71099 1 39
2 71100 1 39
2 71101 1 39
2 71102 1 39
2 71103 1 39
2 71104 1 39
2 71105 1 39
2 71106 1 39
2 71107 1 39
2 71108 1 39
2 71109 1 39
2 71110 1 39
2 71111 1 39
2 71112 1 39
2 71113 1 39
2 71114 1 39
2 71115 1 39
2 71116 1 39
2 71117 1 39
2 71118 1 39
2 71119 1 39
2 71120 1 39
2 71121 1 39
2 71122 1 39
2 71123 1 39
2 71124 1 39
2 71125 1 39
2 71126 1 39
2 71127 1 39
2 71128 1 39
2 71129 1 39
2 71130 1 39
2 71131 1 39
2 71132 1 39
2 71133 1 39
2 71134 1 39
2 71135 1 39
2 71136 1 39
2 71137 1 39
2 71138 1 39
2 71139 1 39
2 71140 1 39
2 71141 1 39
2 71142 1 39
2 71143 1 39
2 71144 1 39
2 71145 1 39
2 71146 1 39
2 71147 1 39
2 71148 1 39
2 71149 1 39
2 71150 1 39
2 71151 1 39
2 71152 1 39
2 71153 1 39
2 71154 1 39
2 71155 1 39
2 71156 1 39
2 71157 1 39
2 71158 1 39
2 71159 1 39
2 71160 1 39
2 71161 1 39
2 71162 1 39
2 71163 1 39
2 71164 1 39
2 71165 1 39
2 71166 1 39
2 71167 1 39
2 71168 1 39
2 71169 1 39
2 71170 1 39
2 71171 1 39
2 71172 1 39
2 71173 1 39
2 71174 1 39
2 71175 1 39
2 71176 1 39
2 71177 1 39
2 71178 1 39
2 71179 1 39
2 71180 1 39
2 71181 1 39
2 71182 1 39
2 71183 1 39
2 71184 1 39
2 71185 1 39
2 71186 1 39
2 71187 1 39
2 71188 1 39
2 71189 1 39
2 71190 1 39
2 71191 1 39
2 71192 1 39
2 71193 1 39
2 71194 1 39
2 71195 1 39
2 71196 1 39
2 71197 1 39
2 71198 1 39
2 71199 1 39
2 71200 1 39
2 71201 1 39
2 71202 1 39
2 71203 1 39
2 71204 1 39
2 71205 1 39
2 71206 1 39
2 71207 1 39
2 71208 1 39
2 71209 1 39
2 71210 1 39
2 71211 1 39
2 71212 1 39
2 71213 1 39
2 71214 1 39
2 71215 1 39
2 71216 1 39
2 71217 1 39
2 71218 1 39
2 71219 1 39
2 71220 1 40
2 71221 1 40
2 71222 1 40
2 71223 1 40
2 71224 1 40
2 71225 1 40
2 71226 1 40
2 71227 1 40
2 71228 1 40
2 71229 1 40
2 71230 1 40
2 71231 1 40
2 71232 1 40
2 71233 1 40
2 71234 1 40
2 71235 1 40
2 71236 1 40
2 71237 1 40
2 71238 1 40
2 71239 1 40
2 71240 1 40
2 71241 1 40
2 71242 1 40
2 71243 1 40
2 71244 1 40
2 71245 1 40
2 71246 1 40
2 71247 1 40
2 71248 1 40
2 71249 1 40
2 71250 1 40
2 71251 1 40
2 71252 1 40
2 71253 1 40
2 71254 1 40
2 71255 1 40
2 71256 1 40
2 71257 1 40
2 71258 1 40
2 71259 1 40
2 71260 1 40
2 71261 1 40
2 71262 1 40
2 71263 1 40
2 71264 1 40
2 71265 1 40
2 71266 1 40
2 71267 1 40
2 71268 1 40
2 71269 1 40
2 71270 1 40
2 71271 1 40
2 71272 1 40
2 71273 1 40
2 71274 1 40
2 71275 1 40
2 71276 1 40
2 71277 1 40
2 71278 1 40
2 71279 1 40
2 71280 1 40
2 71281 1 40
2 71282 1 40
2 71283 1 40
2 71284 1 40
2 71285 1 40
2 71286 1 40
2 71287 1 40
2 71288 1 40
2 71289 1 40
2 71290 1 40
2 71291 1 40
2 71292 1 40
2 71293 1 40
2 71294 1 40
2 71295 1 40
2 71296 1 40
2 71297 1 40
2 71298 1 40
2 71299 1 40
2 71300 1 40
2 71301 1 40
2 71302 1 40
2 71303 1 40
2 71304 1 40
2 71305 1 40
2 71306 1 40
2 71307 1 40
2 71308 1 40
2 71309 1 40
2 71310 1 40
2 71311 1 40
2 71312 1 40
2 71313 1 40
2 71314 1 40
2 71315 1 40
2 71316 1 40
2 71317 1 40
2 71318 1 40
2 71319 1 40
2 71320 1 40
2 71321 1 40
2 71322 1 40
2 71323 1 40
2 71324 1 40
2 71325 1 40
2 71326 1 40
2 71327 1 40
2 71328 1 40
2 71329 1 40
2 71330 1 40
2 71331 1 40
2 71332 1 40
2 71333 1 40
2 71334 1 40
2 71335 1 40
2 71336 1 40
2 71337 1 40
2 71338 1 40
2 71339 1 40
2 71340 1 40
2 71341 1 40
2 71342 1 40
2 71343 1 40
2 71344 1 40
2 71345 1 40
2 71346 1 40
2 71347 1 40
2 71348 1 40
2 71349 1 40
2 71350 1 40
2 71351 1 40
2 71352 1 40
2 71353 1 40
2 71354 1 40
2 71355 1 40
2 71356 1 40
2 71357 1 40
2 71358 1 40
2 71359 1 40
2 71360 1 40
2 71361 1 40
2 71362 1 40
2 71363 1 40
2 71364 1 40
2 71365 1 40
2 71366 1 40
2 71367 1 40
2 71368 1 40
2 71369 1 40
2 71370 1 40
2 71371 1 40
2 71372 1 40
2 71373 1 40
2 71374 1 40
2 71375 1 40
2 71376 1 40
2 71377 1 40
2 71378 1 40
2 71379 1 40
2 71380 1 40
2 71381 1 40
2 71382 1 40
2 71383 1 40
2 71384 1 40
2 71385 1 40
2 71386 1 40
2 71387 1 40
2 71388 1 40
2 71389 1 40
2 71390 1 40
2 71391 1 40
2 71392 1 40
2 71393 1 40
2 71394 1 40
2 71395 1 40
2 71396 1 40
2 71397 1 40
2 71398 1 40
2 71399 1 40
2 71400 1 40
2 71401 1 40
2 71402 1 40
2 71403 1 40
2 71404 1 40
2 71405 1 40
2 71406 1 40
2 71407 1 40
2 71408 1 40
2 71409 1 40
2 71410 1 40
2 71411 1 40
2 71412 1 40
2 71413 1 40
2 71414 1 40
2 71415 1 40
2 71416 1 40
2 71417 1 40
2 71418 1 40
2 71419 1 40
2 71420 1 40
2 71421 1 40
2 71422 1 40
2 71423 1 40
2 71424 1 40
2 71425 1 40
2 71426 1 40
2 71427 1 40
2 71428 1 40
2 71429 1 40
2 71430 1 40
2 71431 1 40
2 71432 1 40
2 71433 1 40
2 71434 1 40
2 71435 1 40
2 71436 1 40
2 71437 1 40
2 71438 1 40
2 71439 1 40
2 71440 1 40
2 71441 1 40
2 71442 1 40
2 71443 1 40
2 71444 1 40
2 71445 1 40
2 71446 1 40
2 71447 1 40
2 71448 1 40
2 71449 1 40
2 71450 1 40
2 71451 1 40
2 71452 1 40
2 71453 1 40
2 71454 1 40
2 71455 1 40
2 71456 1 40
2 71457 1 40
2 71458 1 40
2 71459 1 40
2 71460 1 40
2 71461 1 40
2 71462 1 40
2 71463 1 40
2 71464 1 40
2 71465 1 40
2 71466 1 40
2 71467 1 40
2 71468 1 40
2 71469 1 40
2 71470 1 40
2 71471 1 40
2 71472 1 40
2 71473 1 40
2 71474 1 40
2 71475 1 40
2 71476 1 40
2 71477 1 40
2 71478 1 40
2 71479 1 40
2 71480 1 40
2 71481 1 40
2 71482 1 40
2 71483 1 40
2 71484 1 40
2 71485 1 40
2 71486 1 40
2 71487 1 40
2 71488 1 40
2 71489 1 40
2 71490 1 40
2 71491 1 40
2 71492 1 40
2 71493 1 40
2 71494 1 40
2 71495 1 40
2 71496 1 40
2 71497 1 40
2 71498 1 40
2 71499 1 40
2 71500 1 40
2 71501 1 40
2 71502 1 40
2 71503 1 40
2 71504 1 40
2 71505 1 40
2 71506 1 40
2 71507 1 40
2 71508 1 40
2 71509 1 40
2 71510 1 40
2 71511 1 40
2 71512 1 40
2 71513 1 40
2 71514 1 40
2 71515 1 40
2 71516 1 40
2 71517 1 40
2 71518 1 40
2 71519 1 40
2 71520 1 40
2 71521 1 41
2 71522 1 41
2 71523 1 41
2 71524 1 41
2 71525 1 41
2 71526 1 41
2 71527 1 41
2 71528 1 41
2 71529 1 41
2 71530 1 41
2 71531 1 41
2 71532 1 41
2 71533 1 41
2 71534 1 41
2 71535 1 41
2 71536 1 41
2 71537 1 41
2 71538 1 41
2 71539 1 41
2 71540 1 41
2 71541 1 41
2 71542 1 41
2 71543 1 41
2 71544 1 41
2 71545 1 41
2 71546 1 41
2 71547 1 41
2 71548 1 41
2 71549 1 41
2 71550 1 41
2 71551 1 41
2 71552 1 41
2 71553 1 41
2 71554 1 41
2 71555 1 41
2 71556 1 41
2 71557 1 41
2 71558 1 41
2 71559 1 41
2 71560 1 41
2 71561 1 41
2 71562 1 41
2 71563 1 41
2 71564 1 41
2 71565 1 41
2 71566 1 41
2 71567 1 41
2 71568 1 41
2 71569 1 41
2 71570 1 41
2 71571 1 41
2 71572 1 41
2 71573 1 41
2 71574 1 41
2 71575 1 41
2 71576 1 41
2 71577 1 41
2 71578 1 41
2 71579 1 41
2 71580 1 41
2 71581 1 41
2 71582 1 41
2 71583 1 41
2 71584 1 41
2 71585 1 41
2 71586 1 41
2 71587 1 41
2 71588 1 41
2 71589 1 41
2 71590 1 41
2 71591 1 41
2 71592 1 41
2 71593 1 41
2 71594 1 41
2 71595 1 41
2 71596 1 41
2 71597 1 41
2 71598 1 41
2 71599 1 41
2 71600 1 41
2 71601 1 41
2 71602 1 41
2 71603 1 41
2 71604 1 41
2 71605 1 41
2 71606 1 41
2 71607 1 41
2 71608 1 41
2 71609 1 41
2 71610 1 41
2 71611 1 41
2 71612 1 41
2 71613 1 41
2 71614 1 41
2 71615 1 41
2 71616 1 41
2 71617 1 41
2 71618 1 41
2 71619 1 41
2 71620 1 41
2 71621 1 41
2 71622 1 41
2 71623 1 41
2 71624 1 41
2 71625 1 41
2 71626 1 41
2 71627 1 41
2 71628 1 41
2 71629 1 41
2 71630 1 41
2 71631 1 41
2 71632 1 41
2 71633 1 41
2 71634 1 41
2 71635 1 41
2 71636 1 41
2 71637 1 41
2 71638 1 41
2 71639 1 41
2 71640 1 41
2 71641 1 41
2 71642 1 41
2 71643 1 41
2 71644 1 41
2 71645 1 41
2 71646 1 41
2 71647 1 41
2 71648 1 41
2 71649 1 41
2 71650 1 41
2 71651 1 41
2 71652 1 41
2 71653 1 41
2 71654 1 41
2 71655 1 41
2 71656 1 41
2 71657 1 41
2 71658 1 41
2 71659 1 41
2 71660 1 41
2 71661 1 41
2 71662 1 41
2 71663 1 41
2 71664 1 41
2 71665 1 41
2 71666 1 41
2 71667 1 41
2 71668 1 41
2 71669 1 41
2 71670 1 41
2 71671 1 41
2 71672 1 41
2 71673 1 41
2 71674 1 41
2 71675 1 41
2 71676 1 41
2 71677 1 41
2 71678 1 41
2 71679 1 41
2 71680 1 41
2 71681 1 41
2 71682 1 41
2 71683 1 41
2 71684 1 41
2 71685 1 41
2 71686 1 41
2 71687 1 41
2 71688 1 41
2 71689 1 41
2 71690 1 41
2 71691 1 41
2 71692 1 41
2 71693 1 41
2 71694 1 41
2 71695 1 41
2 71696 1 41
2 71697 1 41
2 71698 1 41
2 71699 1 41
2 71700 1 41
2 71701 1 41
2 71702 1 41
2 71703 1 41
2 71704 1 41
2 71705 1 41
2 71706 1 41
2 71707 1 41
2 71708 1 41
2 71709 1 41
2 71710 1 41
2 71711 1 41
2 71712 1 41
2 71713 1 42
2 71714 1 42
2 71715 1 42
2 71716 1 42
2 71717 1 42
2 71718 1 42
2 71719 1 42
2 71720 1 42
2 71721 1 42
2 71722 1 42
2 71723 1 42
2 71724 1 42
2 71725 1 42
2 71726 1 42
2 71727 1 42
2 71728 1 42
2 71729 1 42
2 71730 1 42
2 71731 1 42
2 71732 1 42
2 71733 1 42
2 71734 1 42
2 71735 1 42
2 71736 1 42
2 71737 1 42
2 71738 1 42
2 71739 1 42
2 71740 1 42
2 71741 1 42
2 71742 1 42
2 71743 1 42
2 71744 1 42
2 71745 1 42
2 71746 1 42
2 71747 1 42
2 71748 1 42
2 71749 1 42
2 71750 1 42
2 71751 1 42
2 71752 1 42
2 71753 1 42
2 71754 1 42
2 71755 1 42
2 71756 1 42
2 71757 1 42
2 71758 1 42
2 71759 1 42
2 71760 1 42
2 71761 1 42
2 71762 1 42
2 71763 1 42
2 71764 1 42
2 71765 1 42
2 71766 1 42
2 71767 1 42
2 71768 1 42
2 71769 1 42
2 71770 1 42
2 71771 1 42
2 71772 1 42
2 71773 1 42
2 71774 1 42
2 71775 1 42
2 71776 1 42
2 71777 1 42
2 71778 1 42
2 71779 1 42
2 71780 1 42
2 71781 1 42
2 71782 1 42
2 71783 1 42
2 71784 1 42
2 71785 1 42
2 71786 1 42
2 71787 1 42
2 71788 1 42
2 71789 1 42
2 71790 1 42
2 71791 1 42
2 71792 1 42
2 71793 1 42
2 71794 1 42
2 71795 1 42
2 71796 1 42
2 71797 1 42
2 71798 1 42
2 71799 1 42
2 71800 1 42
2 71801 1 42
2 71802 1 42
2 71803 1 42
2 71804 1 42
2 71805 1 42
2 71806 1 42
2 71807 1 42
2 71808 1 42
2 71809 1 42
2 71810 1 42
2 71811 1 42
2 71812 1 42
2 71813 1 42
2 71814 1 42
2 71815 1 42
2 71816 1 42
2 71817 1 42
2 71818 1 42
2 71819 1 42
2 71820 1 42
2 71821 1 42
2 71822 1 42
2 71823 1 42
2 71824 1 42
2 71825 1 42
2 71826 1 42
2 71827 1 42
2 71828 1 42
2 71829 1 42
2 71830 1 42
2 71831 1 42
2 71832 1 42
2 71833 1 42
2 71834 1 42
2 71835 1 42
2 71836 1 42
2 71837 1 42
2 71838 1 42
2 71839 1 42
2 71840 1 42
2 71841 1 42
2 71842 1 42
2 71843 1 42
2 71844 1 42
2 71845 1 42
2 71846 1 42
2 71847 1 42
2 71848 1 42
2 71849 1 42
2 71850 1 42
2 71851 1 42
2 71852 1 42
2 71853 1 42
2 71854 1 42
2 71855 1 42
2 71856 1 42
2 71857 1 42
2 71858 1 42
2 71859 1 42
2 71860 1 42
2 71861 1 42
2 71862 1 42
2 71863 1 42
2 71864 1 42
2 71865 1 42
2 71866 1 42
2 71867 1 42
2 71868 1 42
2 71869 1 42
2 71870 1 42
2 71871 1 42
2 71872 1 42
2 71873 1 42
2 71874 1 42
2 71875 1 42
2 71876 1 42
2 71877 1 42
2 71878 1 42
2 71879 1 43
2 71880 1 43
2 71881 1 43
2 71882 1 43
2 71883 1 43
2 71884 1 43
2 71885 1 43
2 71886 1 43
2 71887 1 43
2 71888 1 43
2 71889 1 43
2 71890 1 43
2 71891 1 43
2 71892 1 43
2 71893 1 43
2 71894 1 43
2 71895 1 43
2 71896 1 43
2 71897 1 43
2 71898 1 43
2 71899 1 43
2 71900 1 43
2 71901 1 43
2 71902 1 43
2 71903 1 43
2 71904 1 43
2 71905 1 43
2 71906 1 43
2 71907 1 43
2 71908 1 43
2 71909 1 43
2 71910 1 43
2 71911 1 43
2 71912 1 43
2 71913 1 43
2 71914 1 43
2 71915 1 43
2 71916 1 43
2 71917 1 43
2 71918 1 43
2 71919 1 43
2 71920 1 43
2 71921 1 43
2 71922 1 43
2 71923 1 43
2 71924 1 43
2 71925 1 43
2 71926 1 43
2 71927 1 43
2 71928 1 43
2 71929 1 43
2 71930 1 43
2 71931 1 43
2 71932 1 43
2 71933 1 43
2 71934 1 43
2 71935 1 43
2 71936 1 43
2 71937 1 43
2 71938 1 43
2 71939 1 43
2 71940 1 43
2 71941 1 43
2 71942 1 43
2 71943 1 43
2 71944 1 43
2 71945 1 43
2 71946 1 43
2 71947 1 43
2 71948 1 43
2 71949 1 43
2 71950 1 43
2 71951 1 43
2 71952 1 43
2 71953 1 43
2 71954 1 43
2 71955 1 43
2 71956 1 43
2 71957 1 43
2 71958 1 43
2 71959 1 43
2 71960 1 43
2 71961 1 43
2 71962 1 43
2 71963 1 43
2 71964 1 43
2 71965 1 43
2 71966 1 43
2 71967 1 43
2 71968 1 43
2 71969 1 43
2 71970 1 43
2 71971 1 43
2 71972 1 43
2 71973 1 43
2 71974 1 43
2 71975 1 43
2 71976 1 43
2 71977 1 44
2 71978 1 44
2 71979 1 44
2 71980 1 44
2 71981 1 44
2 71982 1 44
2 71983 1 44
2 71984 1 44
2 71985 1 44
2 71986 1 44
2 71987 1 44
2 71988 1 44
2 71989 1 44
2 71990 1 44
2 71991 1 44
2 71992 1 44
2 71993 1 44
2 71994 1 44
2 71995 1 44
2 71996 1 44
2 71997 1 44
2 71998 1 44
2 71999 1 44
2 72000 1 44
2 72001 1 44
2 72002 1 44
2 72003 1 44
2 72004 1 44
2 72005 1 44
2 72006 1 44
2 72007 1 44
2 72008 1 44
2 72009 1 44
2 72010 1 44
2 72011 1 44
2 72012 1 44
2 72013 1 44
2 72014 1 44
2 72015 1 44
2 72016 1 44
2 72017 1 44
2 72018 1 44
2 72019 1 44
2 72020 1 44
2 72021 1 44
2 72022 1 44
2 72023 1 44
2 72024 1 44
2 72025 1 44
2 72026 1 44
2 72027 1 44
2 72028 1 44
2 72029 1 44
2 72030 1 44
2 72031 1 44
2 72032 1 44
2 72033 1 44
2 72034 1 44
2 72035 1 44
2 72036 1 44
2 72037 1 44
2 72038 1 44
2 72039 1 44
2 72040 1 44
2 72041 1 44
2 72042 1 44
2 72043 1 44
2 72044 1 44
2 72045 1 44
2 72046 1 44
2 72047 1 44
2 72048 1 44
2 72049 1 44
2 72050 1 44
2 72051 1 44
2 72052 1 44
2 72053 1 44
2 72054 1 44
2 72055 1 44
2 72056 1 44
2 72057 1 44
2 72058 1 44
2 72059 1 44
2 72060 1 44
2 72061 1 44
2 72062 1 44
2 72063 1 44
2 72064 1 44
2 72065 1 44
2 72066 1 44
2 72067 1 44
2 72068 1 44
2 72069 1 44
2 72070 1 44
2 72071 1 44
2 72072 1 44
2 72073 1 44
2 72074 1 44
2 72075 1 44
2 72076 1 44
2 72077 1 44
2 72078 1 44
2 72079 1 44
2 72080 1 45
2 72081 1 45
2 72082 1 45
2 72083 1 45
2 72084 1 45
2 72085 1 45
2 72086 1 45
2 72087 1 45
2 72088 1 45
2 72089 1 45
2 72090 1 45
2 72091 1 45
2 72092 1 45
2 72093 1 45
2 72094 1 45
2 72095 1 45
2 72096 1 45
2 72097 1 45
2 72098 1 45
2 72099 1 45
2 72100 1 45
2 72101 1 45
2 72102 1 45
2 72103 1 45
2 72104 1 45
2 72105 1 45
2 72106 1 45
2 72107 1 45
2 72108 1 45
2 72109 1 45
2 72110 1 45
2 72111 1 45
2 72112 1 45
2 72113 1 45
2 72114 1 45
2 72115 1 45
2 72116 1 45
2 72117 1 45
2 72118 1 45
2 72119 1 45
2 72120 1 45
2 72121 1 45
2 72122 1 45
2 72123 1 45
2 72124 1 45
2 72125 1 45
2 72126 1 45
2 72127 1 45
2 72128 1 45
2 72129 1 45
2 72130 1 45
2 72131 1 45
2 72132 1 45
2 72133 1 45
2 72134 1 45
2 72135 1 45
2 72136 1 45
2 72137 1 45
2 72138 1 45
2 72139 1 45
2 72140 1 45
2 72141 1 45
2 72142 1 45
2 72143 1 45
2 72144 1 45
2 72145 1 45
2 72146 1 45
2 72147 1 45
2 72148 1 45
2 72149 1 45
2 72150 1 45
2 72151 1 45
2 72152 1 45
2 72153 1 45
2 72154 1 45
2 72155 1 45
2 72156 1 45
2 72157 1 45
2 72158 1 45
2 72159 1 45
2 72160 1 45
2 72161 1 45
2 72162 1 45
2 72163 1 45
2 72164 1 45
2 72165 1 45
2 72166 1 45
2 72167 1 45
2 72168 1 45
2 72169 1 45
2 72170 1 45
2 72171 1 45
2 72172 1 45
2 72173 1 45
2 72174 1 45
2 72175 1 45
2 72176 1 45
2 72177 1 45
2 72178 1 45
2 72179 1 45
2 72180 1 45
2 72181 1 45
2 72182 1 45
2 72183 1 45
2 72184 1 45
2 72185 1 45
2 72186 1 45
2 72187 1 45
2 72188 1 45
2 72189 1 45
2 72190 1 45
2 72191 1 45
2 72192 1 45
2 72193 1 45
2 72194 1 45
2 72195 1 45
2 72196 1 45
2 72197 1 45
2 72198 1 45
2 72199 1 45
2 72200 1 45
2 72201 1 45
2 72202 1 45
2 72203 1 45
2 72204 1 45
2 72205 1 45
2 72206 1 45
2 72207 1 45
2 72208 1 45
2 72209 1 45
2 72210 1 46
2 72211 1 46
2 72212 1 46
2 72213 1 46
2 72214 1 46
2 72215 1 46
2 72216 1 46
2 72217 1 46
2 72218 1 46
2 72219 1 46
2 72220 1 46
2 72221 1 46
2 72222 1 46
2 72223 1 46
2 72224 1 46
2 72225 1 46
2 72226 1 46
2 72227 1 46
2 72228 1 46
2 72229 1 46
2 72230 1 46
2 72231 1 46
2 72232 1 46
2 72233 1 46
2 72234 1 46
2 72235 1 46
2 72236 1 46
2 72237 1 46
2 72238 1 46
2 72239 1 46
2 72240 1 46
2 72241 1 46
2 72242 1 46
2 72243 1 46
2 72244 1 46
2 72245 1 46
2 72246 1 46
2 72247 1 46
2 72248 1 46
2 72249 1 46
2 72250 1 46
2 72251 1 46
2 72252 1 46
2 72253 1 46
2 72254 1 46
2 72255 1 46
2 72256 1 46
2 72257 1 46
2 72258 1 46
2 72259 1 46
2 72260 1 46
2 72261 1 46
2 72262 1 46
2 72263 1 46
2 72264 1 46
2 72265 1 46
2 72266 1 46
2 72267 1 46
2 72268 1 46
2 72269 1 46
2 72270 1 46
2 72271 1 46
2 72272 1 46
2 72273 1 46
2 72274 1 46
2 72275 1 46
2 72276 1 46
2 72277 1 46
2 72278 1 46
2 72279 1 46
2 72280 1 46
2 72281 1 46
2 72282 1 46
2 72283 1 46
2 72284 1 46
2 72285 1 46
2 72286 1 46
2 72287 1 46
2 72288 1 46
2 72289 1 46
2 72290 1 46
2 72291 1 46
2 72292 1 46
2 72293 1 46
2 72294 1 46
2 72295 1 46
2 72296 1 46
2 72297 1 47
2 72298 1 47
2 72299 1 47
2 72300 1 47
2 72301 1 47
2 72302 1 47
2 72303 1 47
2 72304 1 47
2 72305 1 47
2 72306 1 47
2 72307 1 47
2 72308 1 47
2 72309 1 47
2 72310 1 47
2 72311 1 47
2 72312 1 47
2 72313 1 47
2 72314 1 47
2 72315 1 47
2 72316 1 47
2 72317 1 47
2 72318 1 47
2 72319 1 47
2 72320 1 47
2 72321 1 47
2 72322 1 47
2 72323 1 47
2 72324 1 47
2 72325 1 47
2 72326 1 47
2 72327 1 47
2 72328 1 47
2 72329 1 47
2 72330 1 47
2 72331 1 47
2 72332 1 47
2 72333 1 47
2 72334 1 47
2 72335 1 47
2 72336 1 47
2 72337 1 47
2 72338 1 47
2 72339 1 47
2 72340 1 47
2 72341 1 47
2 72342 1 47
2 72343 1 47
2 72344 1 47
2 72345 1 47
2 72346 1 47
2 72347 1 47
2 72348 1 47
2 72349 1 47
2 72350 1 47
2 72351 1 47
2 72352 1 47
2 72353 1 47
2 72354 1 47
2 72355 1 47
2 72356 1 47
2 72357 1 47
2 72358 1 47
2 72359 1 47
2 72360 1 47
2 72361 1 47
2 72362 1 47
2 72363 1 47
2 72364 1 47
2 72365 1 47
2 72366 1 47
2 72367 1 47
2 72368 1 47
2 72369 1 47
2 72370 1 47
2 72371 1 47
2 72372 1 47
2 72373 1 47
2 72374 1 47
2 72375 1 47
2 72376 1 47
2 72377 1 47
2 72378 1 47
2 72379 1 47
2 72380 1 47
2 72381 1 47
2 72382 1 47
2 72383 1 47
2 72384 1 47
2 72385 1 47
2 72386 1 47
2 72387 1 47
2 72388 1 47
2 72389 1 47
2 72390 1 47
2 72391 1 47
2 72392 1 47
2 72393 1 47
2 72394 1 47
2 72395 1 47
2 72396 1 47
2 72397 1 47
2 72398 1 47
2 72399 1 47
2 72400 1 47
2 72401 1 47
2 72402 1 47
2 72403 1 47
2 72404 1 47
2 72405 1 47
2 72406 1 47
2 72407 1 47
2 72408 1 47
2 72409 1 47
2 72410 1 47
2 72411 1 47
2 72412 1 47
2 72413 1 47
2 72414 1 47
2 72415 1 47
2 72416 1 47
2 72417 1 47
2 72418 1 47
2 72419 1 47
2 72420 1 47
2 72421 1 47
2 72422 1 47
2 72423 1 47
2 72424 1 47
2 72425 1 47
2 72426 1 47
2 72427 1 47
2 72428 1 47
2 72429 1 47
2 72430 1 47
2 72431 1 47
2 72432 1 47
2 72433 1 47
2 72434 1 47
2 72435 1 47
2 72436 1 47
2 72437 1 47
2 72438 1 47
2 72439 1 47
2 72440 1 47
2 72441 1 47
2 72442 1 47
2 72443 1 47
2 72444 1 47
2 72445 1 47
2 72446 1 47
2 72447 1 47
2 72448 1 47
2 72449 1 47
2 72450 1 47
2 72451 1 47
2 72452 1 47
2 72453 1 47
2 72454 1 47
2 72455 1 47
2 72456 1 47
2 72457 1 47
2 72458 1 47
2 72459 1 47
2 72460 1 47
2 72461 1 47
2 72462 1 47
2 72463 1 47
2 72464 1 47
2 72465 1 47
2 72466 1 47
2 72467 1 47
2 72468 1 47
2 72469 1 47
2 72470 1 47
2 72471 1 47
2 72472 1 47
2 72473 1 47
2 72474 1 47
2 72475 1 47
2 72476 1 47
2 72477 1 47
2 72478 1 47
2 72479 1 47
2 72480 1 47
2 72481 1 47
2 72482 1 47
2 72483 1 47
2 72484 1 47
2 72485 1 47
2 72486 1 47
2 72487 1 47
2 72488 1 47
2 72489 1 47
2 72490 1 47
2 72491 1 47
2 72492 1 47
2 72493 1 47
2 72494 1 47
2 72495 1 47
2 72496 1 47
2 72497 1 47
2 72498 1 47
2 72499 1 47
2 72500 1 47
2 72501 1 47
2 72502 1 47
2 72503 1 47
2 72504 1 47
2 72505 1 48
2 72506 1 48
2 72507 1 48
2 72508 1 48
2 72509 1 48
2 72510 1 48
2 72511 1 48
2 72512 1 48
2 72513 1 48
2 72514 1 48
2 72515 1 48
2 72516 1 48
2 72517 1 48
2 72518 1 48
2 72519 1 48
2 72520 1 48
2 72521 1 48
2 72522 1 48
2 72523 1 48
2 72524 1 48
2 72525 1 48
2 72526 1 48
2 72527 1 48
2 72528 1 48
2 72529 1 48
2 72530 1 48
2 72531 1 48
2 72532 1 48
2 72533 1 48
2 72534 1 48
2 72535 1 48
2 72536 1 48
2 72537 1 48
2 72538 1 48
2 72539 1 48
2 72540 1 48
2 72541 1 48
2 72542 1 48
2 72543 1 48
2 72544 1 48
2 72545 1 48
2 72546 1 48
2 72547 1 48
2 72548 1 48
2 72549 1 48
2 72550 1 48
2 72551 1 48
2 72552 1 48
2 72553 1 48
2 72554 1 48
2 72555 1 48
2 72556 1 48
2 72557 1 48
2 72558 1 48
2 72559 1 48
2 72560 1 48
2 72561 1 48
2 72562 1 48
2 72563 1 48
2 72564 1 48
2 72565 1 48
2 72566 1 48
2 72567 1 48
2 72568 1 48
2 72569 1 48
2 72570 1 48
2 72571 1 48
2 72572 1 48
2 72573 1 48
2 72574 1 48
2 72575 1 48
2 72576 1 48
2 72577 1 48
2 72578 1 48
2 72579 1 48
2 72580 1 48
2 72581 1 48
2 72582 1 48
2 72583 1 48
2 72584 1 48
2 72585 1 48
2 72586 1 48
2 72587 1 48
2 72588 1 48
2 72589 1 48
2 72590 1 48
2 72591 1 48
2 72592 1 48
2 72593 1 48
2 72594 1 48
2 72595 1 48
2 72596 1 48
2 72597 1 48
2 72598 1 48
2 72599 1 48
2 72600 1 48
2 72601 1 48
2 72602 1 48
2 72603 1 48
2 72604 1 48
2 72605 1 48
2 72606 1 48
2 72607 1 48
2 72608 1 48
2 72609 1 48
2 72610 1 48
2 72611 1 48
2 72612 1 48
2 72613 1 48
2 72614 1 48
2 72615 1 48
2 72616 1 48
2 72617 1 48
2 72618 1 48
2 72619 1 48
2 72620 1 48
2 72621 1 48
2 72622 1 48
2 72623 1 48
2 72624 1 48
2 72625 1 48
2 72626 1 48
2 72627 1 48
2 72628 1 48
2 72629 1 48
2 72630 1 48
2 72631 1 48
2 72632 1 48
2 72633 1 48
2 72634 1 48
2 72635 1 48
2 72636 1 48
2 72637 1 48
2 72638 1 48
2 72639 1 48
2 72640 1 48
2 72641 1 48
2 72642 1 48
2 72643 1 48
2 72644 1 48
2 72645 1 48
2 72646 1 48
2 72647 1 48
2 72648 1 48
2 72649 1 48
2 72650 1 48
2 72651 1 48
2 72652 1 48
2 72653 1 48
2 72654 1 48
2 72655 1 48
2 72656 1 48
2 72657 1 48
2 72658 1 48
2 72659 1 48
2 72660 1 48
2 72661 1 48
2 72662 1 48
2 72663 1 48
2 72664 1 48
2 72665 1 48
2 72666 1 48
2 72667 1 48
2 72668 1 48
2 72669 1 48
2 72670 1 48
2 72671 1 48
2 72672 1 48
2 72673 1 48
2 72674 1 48
2 72675 1 48
2 72676 1 48
2 72677 1 48
2 72678 1 48
2 72679 1 48
2 72680 1 48
2 72681 1 48
2 72682 1 48
2 72683 1 48
2 72684 1 48
2 72685 1 48
2 72686 1 48
2 72687 1 48
2 72688 1 48
2 72689 1 48
2 72690 1 48
2 72691 1 48
2 72692 1 48
2 72693 1 48
2 72694 1 48
2 72695 1 48
2 72696 1 48
2 72697 1 48
2 72698 1 48
2 72699 1 48
2 72700 1 48
2 72701 1 48
2 72702 1 48
2 72703 1 48
2 72704 1 48
2 72705 1 48
2 72706 1 48
2 72707 1 48
2 72708 1 48
2 72709 1 48
2 72710 1 48
2 72711 1 48
2 72712 1 48
2 72713 1 48
2 72714 1 48
2 72715 1 48
2 72716 1 48
2 72717 1 48
2 72718 1 48
2 72719 1 48
2 72720 1 48
2 72721 1 48
2 72722 1 48
2 72723 1 48
2 72724 1 48
2 72725 1 48
2 72726 1 48
2 72727 1 48
2 72728 1 48
2 72729 1 48
2 72730 1 48
2 72731 1 48
2 72732 1 48
2 72733 1 48
2 72734 1 48
2 72735 1 48
2 72736 1 48
2 72737 1 48
2 72738 1 48
2 72739 1 48
2 72740 1 48
2 72741 1 48
2 72742 1 48
2 72743 1 48
2 72744 1 48
2 72745 1 48
2 72746 1 48
2 72747 1 48
2 72748 1 48
2 72749 1 48
2 72750 1 48
2 72751 1 48
2 72752 1 48
2 72753 1 48
2 72754 1 48
2 72755 1 48
2 72756 1 48
2 72757 1 48
2 72758 1 48
2 72759 1 48
2 72760 1 48
2 72761 1 48
2 72762 1 48
2 72763 1 48
2 72764 1 48
2 72765 1 48
2 72766 1 48
2 72767 1 48
2 72768 1 48
2 72769 1 48
2 72770 1 48
2 72771 1 48
2 72772 1 48
2 72773 1 48
2 72774 1 48
2 72775 1 48
2 72776 1 48
2 72777 1 48
2 72778 1 48
2 72779 1 48
2 72780 1 48
2 72781 1 48
2 72782 1 48
2 72783 1 48
2 72784 1 48
2 72785 1 48
2 72786 1 48
2 72787 1 48
2 72788 1 48
2 72789 1 48
2 72790 1 48
2 72791 1 48
2 72792 1 48
2 72793 1 48
2 72794 1 48
2 72795 1 48
2 72796 1 48
2 72797 1 48
2 72798 1 48
2 72799 1 48
2 72800 1 48
2 72801 1 48
2 72802 1 48
2 72803 1 48
2 72804 1 48
2 72805 1 48
2 72806 1 48
2 72807 1 48
2 72808 1 48
2 72809 1 48
2 72810 1 48
2 72811 1 48
2 72812 1 48
2 72813 1 48
2 72814 1 48
2 72815 1 48
2 72816 1 48
2 72817 1 48
2 72818 1 48
2 72819 1 48
2 72820 1 48
2 72821 1 48
2 72822 1 48
2 72823 1 48
2 72824 1 48
2 72825 1 48
2 72826 1 48
2 72827 1 48
2 72828 1 48
2 72829 1 48
2 72830 1 48
2 72831 1 48
2 72832 1 48
2 72833 1 48
2 72834 1 48
2 72835 1 48
2 72836 1 48
2 72837 1 48
2 72838 1 48
2 72839 1 48
2 72840 1 48
2 72841 1 48
2 72842 1 48
2 72843 1 48
2 72844 1 48
2 72845 1 48
2 72846 1 48
2 72847 1 48
2 72848 1 48
2 72849 1 48
2 72850 1 48
2 72851 1 48
2 72852 1 49
2 72853 1 49
2 72854 1 49
2 72855 1 49
2 72856 1 49
2 72857 1 49
2 72858 1 49
2 72859 1 49
2 72860 1 49
2 72861 1 49
2 72862 1 49
2 72863 1 49
2 72864 1 49
2 72865 1 49
2 72866 1 49
2 72867 1 49
2 72868 1 49
2 72869 1 49
2 72870 1 49
2 72871 1 49
2 72872 1 49
2 72873 1 49
2 72874 1 49
2 72875 1 49
2 72876 1 49
2 72877 1 49
2 72878 1 49
2 72879 1 49
2 72880 1 49
2 72881 1 49
2 72882 1 49
2 72883 1 49
2 72884 1 49
2 72885 1 49
2 72886 1 49
2 72887 1 49
2 72888 1 49
2 72889 1 49
2 72890 1 49
2 72891 1 49
2 72892 1 49
2 72893 1 49
2 72894 1 49
2 72895 1 49
2 72896 1 49
2 72897 1 49
2 72898 1 49
2 72899 1 49
2 72900 1 49
2 72901 1 49
2 72902 1 49
2 72903 1 49
2 72904 1 49
2 72905 1 49
2 72906 1 49
2 72907 1 49
2 72908 1 49
2 72909 1 49
2 72910 1 49
2 72911 1 49
2 72912 1 49
2 72913 1 49
2 72914 1 49
2 72915 1 49
2 72916 1 49
2 72917 1 49
2 72918 1 49
2 72919 1 49
2 72920 1 49
2 72921 1 49
2 72922 1 49
2 72923 1 49
2 72924 1 49
2 72925 1 49
2 72926 1 49
2 72927 1 49
2 72928 1 49
2 72929 1 49
2 72930 1 49
2 72931 1 49
2 72932 1 49
2 72933 1 49
2 72934 1 49
2 72935 1 49
2 72936 1 49
2 72937 1 49
2 72938 1 49
2 72939 1 49
2 72940 1 49
2 72941 1 49
2 72942 1 49
2 72943 1 49
2 72944 1 49
2 72945 1 49
2 72946 1 49
2 72947 1 49
2 72948 1 49
2 72949 1 49
2 72950 1 49
2 72951 1 49
2 72952 1 49
2 72953 1 49
2 72954 1 49
2 72955 1 49
2 72956 1 49
2 72957 1 49
2 72958 1 49
2 72959 1 49
2 72960 1 49
2 72961 1 49
2 72962 1 49
2 72963 1 49
2 72964 1 49
2 72965 1 49
2 72966 1 49
2 72967 1 49
2 72968 1 49
2 72969 1 49
2 72970 1 49
2 72971 1 49
2 72972 1 49
2 72973 1 49
2 72974 1 49
2 72975 1 49
2 72976 1 49
2 72977 1 49
2 72978 1 49
2 72979 1 49
2 72980 1 49
2 72981 1 49
2 72982 1 49
2 72983 1 49
2 72984 1 49
2 72985 1 49
2 72986 1 49
2 72987 1 49
2 72988 1 49
2 72989 1 49
2 72990 1 49
2 72991 1 49
2 72992 1 49
2 72993 1 49
2 72994 1 49
2 72995 1 49
2 72996 1 49
2 72997 1 49
2 72998 1 49
2 72999 1 49
2 73000 1 49
2 73001 1 49
2 73002 1 49
2 73003 1 49
2 73004 1 49
2 73005 1 49
2 73006 1 49
2 73007 1 49
2 73008 1 49
2 73009 1 49
2 73010 1 49
2 73011 1 49
2 73012 1 49
2 73013 1 49
2 73014 1 49
2 73015 1 49
2 73016 1 49
2 73017 1 49
2 73018 1 49
2 73019 1 49
2 73020 1 49
2 73021 1 49
2 73022 1 49
2 73023 1 49
2 73024 1 49
2 73025 1 49
2 73026 1 49
2 73027 1 49
2 73028 1 49
2 73029 1 49
2 73030 1 49
2 73031 1 49
2 73032 1 49
2 73033 1 49
2 73034 1 49
2 73035 1 49
2 73036 1 49
2 73037 1 49
2 73038 1 49
2 73039 1 49
2 73040 1 49
2 73041 1 49
2 73042 1 49
2 73043 1 49
2 73044 1 49
2 73045 1 49
2 73046 1 49
2 73047 1 49
2 73048 1 49
2 73049 1 49
2 73050 1 49
2 73051 1 49
2 73052 1 49
2 73053 1 49
2 73054 1 49
2 73055 1 49
2 73056 1 49
2 73057 1 49
2 73058 1 49
2 73059 1 49
2 73060 1 49
2 73061 1 49
2 73062 1 49
2 73063 1 49
2 73064 1 49
2 73065 1 49
2 73066 1 49
2 73067 1 49
2 73068 1 49
2 73069 1 49
2 73070 1 49
2 73071 1 49
2 73072 1 49
2 73073 1 49
2 73074 1 49
2 73075 1 49
2 73076 1 49
2 73077 1 49
2 73078 1 49
2 73079 1 49
2 73080 1 49
2 73081 1 49
2 73082 1 49
2 73083 1 49
2 73084 1 49
2 73085 1 49
2 73086 1 49
2 73087 1 49
2 73088 1 49
2 73089 1 49
2 73090 1 49
2 73091 1 49
2 73092 1 49
2 73093 1 49
2 73094 1 49
2 73095 1 49
2 73096 1 49
2 73097 1 49
2 73098 1 49
2 73099 1 49
2 73100 1 49
2 73101 1 49
2 73102 1 49
2 73103 1 49
2 73104 1 49
2 73105 1 49
2 73106 1 49
2 73107 1 49
2 73108 1 49
2 73109 1 49
2 73110 1 49
2 73111 1 49
2 73112 1 49
2 73113 1 49
2 73114 1 49
2 73115 1 49
2 73116 1 49
2 73117 1 49
2 73118 1 49
2 73119 1 49
2 73120 1 49
2 73121 1 49
2 73122 1 49
2 73123 1 49
2 73124 1 49
2 73125 1 49
2 73126 1 49
2 73127 1 49
2 73128 1 49
2 73129 1 49
2 73130 1 49
2 73131 1 49
2 73132 1 49
2 73133 1 49
2 73134 1 49
2 73135 1 49
2 73136 1 49
2 73137 1 49
2 73138 1 49
2 73139 1 49
2 73140 1 49
2 73141 1 49
2 73142 1 49
2 73143 1 49
2 73144 1 49
2 73145 1 49
2 73146 1 49
2 73147 1 49
2 73148 1 49
2 73149 1 49
2 73150 1 49
2 73151 1 49
2 73152 1 49
2 73153 1 49
2 73154 1 49
2 73155 1 49
2 73156 1 49
2 73157 1 49
2 73158 1 49
2 73159 1 49
2 73160 1 49
2 73161 1 49
2 73162 1 49
2 73163 1 49
2 73164 1 49
2 73165 1 49
2 73166 1 49
2 73167 1 49
2 73168 1 49
2 73169 1 49
2 73170 1 49
2 73171 1 49
2 73172 1 49
2 73173 1 49
2 73174 1 49
2 73175 1 49
2 73176 1 49
2 73177 1 49
2 73178 1 49
2 73179 1 49
2 73180 1 49
2 73181 1 49
2 73182 1 49
2 73183 1 49
2 73184 1 49
2 73185 1 49
2 73186 1 49
2 73187 1 49
2 73188 1 49
2 73189 1 49
2 73190 1 49
2 73191 1 49
2 73192 1 49
2 73193 1 49
2 73194 1 49
2 73195 1 49
2 73196 1 49
2 73197 1 49
2 73198 1 49
2 73199 1 49
2 73200 1 49
2 73201 1 49
2 73202 1 49
2 73203 1 49
2 73204 1 49
2 73205 1 49
2 73206 1 49
2 73207 1 49
2 73208 1 49
2 73209 1 49
2 73210 1 49
2 73211 1 49
2 73212 1 49
2 73213 1 49
2 73214 1 49
2 73215 1 49
2 73216 1 49
2 73217 1 49
2 73218 1 49
2 73219 1 49
2 73220 1 49
2 73221 1 49
2 73222 1 49
2 73223 1 49
2 73224 1 49
2 73225 1 49
2 73226 1 49
2 73227 1 49
2 73228 1 49
2 73229 1 49
2 73230 1 49
2 73231 1 49
2 73232 1 49
2 73233 1 49
2 73234 1 49
2 73235 1 49
2 73236 1 49
2 73237 1 49
2 73238 1 49
2 73239 1 49
2 73240 1 49
2 73241 1 49
2 73242 1 49
2 73243 1 49
2 73244 1 49
2 73245 1 49
2 73246 1 49
2 73247 1 49
2 73248 1 49
2 73249 1 49
2 73250 1 49
2 73251 1 49
2 73252 1 49
2 73253 1 49
2 73254 1 49
2 73255 1 49
2 73256 1 49
2 73257 1 49
2 73258 1 49
2 73259 1 49
2 73260 1 49
2 73261 1 49
2 73262 1 49
2 73263 1 49
2 73264 1 49
2 73265 1 49
2 73266 1 49
2 73267 1 49
2 73268 1 49
2 73269 1 49
2 73270 1 49
2 73271 1 49
2 73272 1 49
2 73273 1 49
2 73274 1 49
2 73275 1 49
2 73276 1 49
2 73277 1 49
2 73278 1 49
2 73279 1 49
2 73280 1 49
2 73281 1 49
2 73282 1 49
2 73283 1 49
2 73284 1 49
2 73285 1 49
2 73286 1 49
2 73287 1 49
2 73288 1 49
2 73289 1 49
2 73290 1 49
2 73291 1 49
2 73292 1 49
2 73293 1 49
2 73294 1 49
2 73295 1 49
2 73296 1 49
2 73297 1 49
2 73298 1 49
2 73299 1 49
2 73300 1 49
2 73301 1 49
2 73302 1 49
2 73303 1 49
2 73304 1 49
2 73305 1 49
2 73306 1 49
2 73307 1 50
2 73308 1 50
2 73309 1 50
2 73310 1 50
2 73311 1 50
2 73312 1 50
2 73313 1 50
2 73314 1 50
2 73315 1 50
2 73316 1 50
2 73317 1 50
2 73318 1 50
2 73319 1 50
2 73320 1 50
2 73321 1 50
2 73322 1 50
2 73323 1 50
2 73324 1 50
2 73325 1 50
2 73326 1 50
2 73327 1 50
2 73328 1 50
2 73329 1 50
2 73330 1 50
2 73331 1 50
2 73332 1 50
2 73333 1 50
2 73334 1 50
2 73335 1 50
2 73336 1 50
2 73337 1 50
2 73338 1 50
2 73339 1 50
2 73340 1 50
2 73341 1 50
2 73342 1 50
2 73343 1 50
2 73344 1 50
2 73345 1 50
2 73346 1 50
2 73347 1 50
2 73348 1 50
2 73349 1 50
2 73350 1 50
2 73351 1 50
2 73352 1 50
2 73353 1 50
2 73354 1 50
2 73355 1 50
2 73356 1 50
2 73357 1 50
2 73358 1 50
2 73359 1 50
2 73360 1 50
2 73361 1 50
2 73362 1 50
2 73363 1 50
2 73364 1 50
2 73365 1 50
2 73366 1 50
2 73367 1 50
2 73368 1 50
2 73369 1 50
2 73370 1 50
2 73371 1 50
2 73372 1 50
2 73373 1 50
2 73374 1 50
2 73375 1 50
2 73376 1 50
2 73377 1 50
2 73378 1 50
2 73379 1 50
2 73380 1 50
2 73381 1 50
2 73382 1 50
2 73383 1 50
2 73384 1 50
2 73385 1 50
2 73386 1 50
2 73387 1 50
2 73388 1 50
2 73389 1 50
2 73390 1 50
2 73391 1 50
2 73392 1 50
2 73393 1 50
2 73394 1 50
2 73395 1 50
2 73396 1 50
2 73397 1 50
2 73398 1 50
2 73399 1 50
2 73400 1 50
2 73401 1 50
2 73402 1 50
2 73403 1 50
2 73404 1 50
2 73405 1 50
2 73406 1 50
2 73407 1 50
2 73408 1 50
2 73409 1 50
2 73410 1 50
2 73411 1 50
2 73412 1 50
2 73413 1 50
2 73414 1 50
2 73415 1 50
2 73416 1 50
2 73417 1 50
2 73418 1 50
2 73419 1 50
2 73420 1 50
2 73421 1 50
2 73422 1 50
2 73423 1 50
2 73424 1 50
2 73425 1 50
2 73426 1 50
2 73427 1 50
2 73428 1 50
2 73429 1 50
2 73430 1 50
2 73431 1 50
2 73432 1 50
2 73433 1 50
2 73434 1 50
2 73435 1 50
2 73436 1 50
2 73437 1 50
2 73438 1 50
2 73439 1 50
2 73440 1 50
2 73441 1 50
2 73442 1 50
2 73443 1 50
2 73444 1 50
2 73445 1 50
2 73446 1 50
2 73447 1 50
2 73448 1 50
2 73449 1 50
2 73450 1 50
2 73451 1 50
2 73452 1 50
2 73453 1 50
2 73454 1 50
2 73455 1 50
2 73456 1 50
2 73457 1 50
2 73458 1 50
2 73459 1 50
2 73460 1 50
2 73461 1 50
2 73462 1 50
2 73463 1 50
2 73464 1 50
2 73465 1 50
2 73466 1 50
2 73467 1 50
2 73468 1 50
2 73469 1 50
2 73470 1 50
2 73471 1 50
2 73472 1 50
2 73473 1 50
2 73474 1 50
2 73475 1 50
2 73476 1 50
2 73477 1 50
2 73478 1 50
2 73479 1 50
2 73480 1 50
2 73481 1 50
2 73482 1 50
2 73483 1 50
2 73484 1 50
2 73485 1 50
2 73486 1 50
2 73487 1 50
2 73488 1 50
2 73489 1 50
2 73490 1 50
2 73491 1 50
2 73492 1 50
2 73493 1 50
2 73494 1 50
2 73495 1 50
2 73496 1 50
2 73497 1 50
2 73498 1 50
2 73499 1 50
2 73500 1 50
2 73501 1 50
2 73502 1 50
2 73503 1 50
2 73504 1 50
2 73505 1 50
2 73506 1 50
2 73507 1 50
2 73508 1 50
2 73509 1 50
2 73510 1 50
2 73511 1 50
2 73512 1 50
2 73513 1 50
2 73514 1 50
2 73515 1 50
2 73516 1 50
2 73517 1 50
2 73518 1 50
2 73519 1 50
2 73520 1 50
2 73521 1 50
2 73522 1 50
2 73523 1 50
2 73524 1 50
2 73525 1 50
2 73526 1 50
2 73527 1 50
2 73528 1 50
2 73529 1 50
2 73530 1 50
2 73531 1 50
2 73532 1 50
2 73533 1 50
2 73534 1 50
2 73535 1 50
2 73536 1 50
2 73537 1 50
2 73538 1 50
2 73539 1 50
2 73540 1 50
2 73541 1 50
2 73542 1 50
2 73543 1 50
2 73544 1 50
2 73545 1 50
2 73546 1 50
2 73547 1 50
2 73548 1 50
2 73549 1 50
2 73550 1 50
2 73551 1 50
2 73552 1 50
2 73553 1 50
2 73554 1 50
2 73555 1 50
2 73556 1 50
2 73557 1 50
2 73558 1 50
2 73559 1 50
2 73560 1 50
2 73561 1 50
2 73562 1 50
2 73563 1 50
2 73564 1 50
2 73565 1 50
2 73566 1 50
2 73567 1 50
2 73568 1 50
2 73569 1 50
2 73570 1 50
2 73571 1 50
2 73572 1 50
2 73573 1 50
2 73574 1 50
2 73575 1 50
2 73576 1 50
2 73577 1 50
2 73578 1 50
2 73579 1 50
2 73580 1 50
2 73581 1 50
2 73582 1 50
2 73583 1 50
2 73584 1 50
2 73585 1 50
2 73586 1 50
2 73587 1 50
2 73588 1 50
2 73589 1 50
2 73590 1 50
2 73591 1 50
2 73592 1 50
2 73593 1 50
2 73594 1 50
2 73595 1 50
2 73596 1 50
2 73597 1 50
2 73598 1 50
2 73599 1 50
2 73600 1 50
2 73601 1 50
2 73602 1 50
2 73603 1 50
2 73604 1 50
2 73605 1 50
2 73606 1 50
2 73607 1 50
2 73608 1 50
2 73609 1 50
2 73610 1 50
2 73611 1 50
2 73612 1 50
2 73613 1 50
2 73614 1 50
2 73615 1 50
2 73616 1 50
2 73617 1 50
2 73618 1 50
2 73619 1 50
2 73620 1 50
2 73621 1 50
2 73622 1 50
2 73623 1 51
2 73624 1 51
2 73625 1 51
2 73626 1 51
2 73627 1 51
2 73628 1 51
2 73629 1 51
2 73630 1 51
2 73631 1 51
2 73632 1 51
2 73633 1 51
2 73634 1 51
2 73635 1 51
2 73636 1 51
2 73637 1 51
2 73638 1 51
2 73639 1 51
2 73640 1 51
2 73641 1 51
2 73642 1 51
2 73643 1 51
2 73644 1 51
2 73645 1 51
2 73646 1 51
2 73647 1 51
2 73648 1 51
2 73649 1 51
2 73650 1 51
2 73651 1 51
2 73652 1 51
2 73653 1 51
2 73654 1 51
2 73655 1 51
2 73656 1 51
2 73657 1 51
2 73658 1 51
2 73659 1 51
2 73660 1 51
2 73661 1 51
2 73662 1 51
2 73663 1 51
2 73664 1 51
2 73665 1 51
2 73666 1 51
2 73667 1 51
2 73668 1 51
2 73669 1 51
2 73670 1 51
2 73671 1 51
2 73672 1 51
2 73673 1 51
2 73674 1 51
2 73675 1 51
2 73676 1 51
2 73677 1 51
2 73678 1 51
2 73679 1 51
2 73680 1 51
2 73681 1 51
2 73682 1 51
2 73683 1 51
2 73684 1 51
2 73685 1 51
2 73686 1 51
2 73687 1 51
2 73688 1 51
2 73689 1 51
2 73690 1 51
2 73691 1 51
2 73692 1 51
2 73693 1 51
2 73694 1 51
2 73695 1 51
2 73696 1 51
2 73697 1 51
2 73698 1 51
2 73699 1 51
2 73700 1 51
2 73701 1 51
2 73702 1 51
2 73703 1 51
2 73704 1 51
2 73705 1 51
2 73706 1 51
2 73707 1 51
2 73708 1 51
2 73709 1 51
2 73710 1 51
2 73711 1 51
2 73712 1 51
2 73713 1 51
2 73714 1 51
2 73715 1 51
2 73716 1 51
2 73717 1 51
2 73718 1 51
2 73719 1 51
2 73720 1 51
2 73721 1 51
2 73722 1 51
2 73723 1 51
2 73724 1 51
2 73725 1 51
2 73726 1 51
2 73727 1 51
2 73728 1 51
2 73729 1 51
2 73730 1 51
2 73731 1 51
2 73732 1 51
2 73733 1 51
2 73734 1 51
2 73735 1 51
2 73736 1 51
2 73737 1 51
2 73738 1 51
2 73739 1 51
2 73740 1 51
2 73741 1 51
2 73742 1 51
2 73743 1 51
2 73744 1 51
2 73745 1 51
2 73746 1 51
2 73747 1 51
2 73748 1 51
2 73749 1 51
2 73750 1 51
2 73751 1 51
2 73752 1 51
2 73753 1 51
2 73754 1 51
2 73755 1 51
2 73756 1 51
2 73757 1 51
2 73758 1 51
2 73759 1 51
2 73760 1 51
2 73761 1 51
2 73762 1 51
2 73763 1 51
2 73764 1 51
2 73765 1 51
2 73766 1 51
2 73767 1 51
2 73768 1 51
2 73769 1 51
2 73770 1 51
2 73771 1 51
2 73772 1 51
2 73773 1 51
2 73774 1 51
2 73775 1 51
2 73776 1 51
2 73777 1 51
2 73778 1 51
2 73779 1 51
2 73780 1 51
2 73781 1 51
2 73782 1 51
2 73783 1 51
2 73784 1 51
2 73785 1 51
2 73786 1 51
2 73787 1 51
2 73788 1 51
2 73789 1 51
2 73790 1 51
2 73791 1 51
2 73792 1 51
2 73793 1 51
2 73794 1 51
2 73795 1 51
2 73796 1 51
2 73797 1 51
2 73798 1 51
2 73799 1 51
2 73800 1 51
2 73801 1 51
2 73802 1 51
2 73803 1 51
2 73804 1 51
2 73805 1 51
2 73806 1 51
2 73807 1 52
2 73808 1 52
2 73809 1 52
2 73810 1 52
2 73811 1 52
2 73812 1 52
2 73813 1 52
2 73814 1 52
2 73815 1 52
2 73816 1 53
2 73817 1 53
2 73818 1 53
2 73819 1 53
2 73820 1 53
2 73821 1 53
2 73822 1 53
2 73823 1 53
2 73824 1 55
2 73825 1 55
2 73826 1 55
2 73827 1 55
2 73828 1 55
2 73829 1 56
2 73830 1 56
2 73831 1 56
2 73832 1 56
2 73833 1 56
2 73834 1 56
2 73835 1 59
2 73836 1 59
2 73837 1 59
2 73838 1 59
2 73839 1 59
2 73840 1 59
2 73841 1 59
2 73842 1 59
2 73843 1 59
2 73844 1 59
2 73845 1 59
2 73846 1 59
2 73847 1 59
2 73848 1 59
2 73849 1 59
2 73850 1 59
2 73851 1 59
2 73852 1 59
2 73853 1 59
2 73854 1 59
2 73855 1 59
2 73856 1 59
2 73857 1 59
2 73858 1 59
2 73859 1 59
2 73860 1 59
2 73861 1 59
2 73862 1 59
2 73863 1 59
2 73864 1 59
2 73865 1 59
2 73866 1 59
2 73867 1 59
2 73868 1 59
2 73869 1 59
2 73870 1 59
2 73871 1 59
2 73872 1 59
2 73873 1 59
2 73874 1 59
2 73875 1 59
2 73876 1 59
2 73877 1 59
2 73878 1 59
2 73879 1 59
2 73880 1 59
2 73881 1 59
2 73882 1 59
2 73883 1 59
2 73884 1 59
2 73885 1 60
2 73886 1 60
2 73887 1 60
2 73888 1 60
2 73889 1 60
2 73890 1 60
2 73891 1 60
2 73892 1 60
2 73893 1 60
2 73894 1 60
2 73895 1 60
2 73896 1 60
2 73897 1 60
2 73898 1 60
2 73899 1 60
2 73900 1 60
2 73901 1 60
2 73902 1 60
2 73903 1 60
2 73904 1 60
2 73905 1 60
2 73906 1 60
2 73907 1 60
2 73908 1 60
2 73909 1 60
2 73910 1 60
2 73911 1 60
2 73912 1 60
2 73913 1 60
2 73914 1 60
2 73915 1 60
2 73916 1 60
2 73917 1 60
2 73918 1 60
2 73919 1 60
2 73920 1 60
2 73921 1 60
2 73922 1 60
2 73923 1 60
2 73924 1 60
2 73925 1 60
2 73926 1 60
2 73927 1 60
2 73928 1 60
2 73929 1 60
2 73930 1 60
2 73931 1 61
2 73932 1 61
2 73933 1 61
2 73934 1 61
2 73935 1 61
2 73936 1 61
2 73937 1 61
2 73938 1 61
2 73939 1 61
2 73940 1 61
2 73941 1 61
2 73942 1 61
2 73943 1 61
2 73944 1 61
2 73945 1 61
2 73946 1 61
2 73947 1 61
2 73948 1 61
2 73949 1 61
2 73950 1 61
2 73951 1 61
2 73952 1 61
2 73953 1 61
2 73954 1 61
2 73955 1 61
2 73956 1 61
2 73957 1 61
2 73958 1 61
2 73959 1 61
2 73960 1 61
2 73961 1 61
2 73962 1 61
2 73963 1 61
2 73964 1 61
2 73965 1 61
2 73966 1 61
2 73967 1 61
2 73968 1 61
2 73969 1 61
2 73970 1 61
2 73971 1 61
2 73972 1 61
2 73973 1 61
2 73974 1 61
2 73975 1 61
2 73976 1 61
2 73977 1 61
2 73978 1 61
2 73979 1 61
2 73980 1 61
2 73981 1 61
2 73982 1 61
2 73983 1 61
2 73984 1 61
2 73985 1 61
2 73986 1 61
2 73987 1 61
2 73988 1 61
2 73989 1 61
2 73990 1 61
2 73991 1 61
2 73992 1 61
2 73993 1 61
2 73994 1 61
2 73995 1 61
2 73996 1 61
2 73997 1 62
2 73998 1 62
2 73999 1 62
2 74000 1 62
2 74001 1 62
2 74002 1 64
2 74003 1 64
2 74004 1 64
2 74005 1 64
2 74006 1 64
2 74007 1 64
2 74008 1 64
2 74009 1 64
2 74010 1 66
2 74011 1 66
2 74012 1 66
2 74013 1 66
2 74014 1 66
2 74015 1 67
2 74016 1 67
2 74017 1 67
2 74018 1 67
2 74019 1 67
2 74020 1 67
2 74021 1 67
2 74022 1 67
2 74023 1 67
2 74024 1 67
2 74025 1 67
2 74026 1 67
2 74027 1 67
2 74028 1 67
2 74029 1 67
2 74030 1 67
2 74031 1 67
2 74032 1 67
2 74033 1 67
2 74034 1 67
2 74035 1 67
2 74036 1 67
2 74037 1 67
2 74038 1 67
2 74039 1 67
2 74040 1 67
2 74041 1 67
2 74042 1 67
2 74043 1 67
2 74044 1 67
2 74045 1 67
2 74046 1 67
2 74047 1 67
2 74048 1 67
2 74049 1 68
2 74050 1 68
2 74051 1 68
2 74052 1 68
2 74053 1 68
2 74054 1 68
2 74055 1 68
2 74056 1 68
2 74057 1 68
2 74058 1 68
2 74059 1 68
2 74060 1 68
2 74061 1 68
2 74062 1 68
2 74063 1 68
2 74064 1 68
2 74065 1 68
2 74066 1 68
2 74067 1 68
2 74068 1 68
2 74069 1 68
2 74070 1 68
2 74071 1 68
2 74072 1 68
2 74073 1 68
2 74074 1 68
2 74075 1 68
2 74076 1 68
2 74077 1 68
2 74078 1 68
2 74079 1 68
2 74080 1 68
2 74081 1 70
2 74082 1 70
2 74083 1 71
2 74084 1 71
2 74085 1 71
2 74086 1 71
2 74087 1 71
2 74088 1 71
2 74089 1 71
2 74090 1 71
2 74091 1 72
2 74092 1 72
2 74093 1 72
2 74094 1 72
2 74095 1 72
2 74096 1 72
2 74097 1 72
2 74098 1 72
2 74099 1 72
2 74100 1 72
2 74101 1 72
2 74102 1 72
2 74103 1 72
2 74104 1 72
2 74105 1 72
2 74106 1 72
2 74107 1 72
2 74108 1 73
2 74109 1 73
2 74110 1 73
2 74111 1 73
2 74112 1 73
2 74113 1 73
2 74114 1 73
2 74115 1 73
2 74116 1 73
2 74117 1 73
2 74118 1 73
2 74119 1 73
2 74120 1 73
2 74121 1 73
2 74122 1 73
2 74123 1 73
2 74124 1 73
2 74125 1 74
2 74126 1 74
2 74127 1 74
2 74128 1 74
2 74129 1 74
2 74130 1 74
2 74131 1 75
2 74132 1 75
2 74133 1 76
2 74134 1 76
2 74135 1 76
2 74136 1 76
2 74137 1 76
2 74138 1 81
2 74139 1 81
2 74140 1 81
2 74141 1 81
2 74142 1 81
2 74143 1 81
2 74144 1 81
2 74145 1 81
2 74146 1 81
2 74147 1 81
2 74148 1 81
2 74149 1 81
2 74150 1 81
2 74151 1 81
2 74152 1 81
2 74153 1 81
2 74154 1 81
2 74155 1 81
2 74156 1 82
2 74157 1 82
2 74158 1 83
2 74159 1 83
2 74160 1 83
2 74161 1 83
2 74162 1 84
2 74163 1 84
2 74164 1 84
2 74165 1 84
2 74166 1 84
2 74167 1 84
2 74168 1 84
2 74169 1 84
2 74170 1 84
2 74171 1 84
2 74172 1 84
2 74173 1 84
2 74174 1 84
2 74175 1 84
2 74176 1 84
2 74177 1 84
2 74178 1 87
2 74179 1 87
2 74180 1 88
2 74181 1 88
2 74182 1 88
2 74183 1 88
2 74184 1 88
2 74185 1 88
2 74186 1 88
2 74187 1 88
2 74188 1 88
2 74189 1 88
2 74190 1 88
2 74191 1 88
2 74192 1 88
2 74193 1 88
2 74194 1 88
2 74195 1 88
2 74196 1 88
2 74197 1 88
2 74198 1 88
2 74199 1 88
2 74200 1 88
2 74201 1 88
2 74202 1 89
2 74203 1 89
2 74204 1 90
2 74205 1 90
2 74206 1 90
2 74207 1 90
2 74208 1 90
2 74209 1 90
2 74210 1 90
2 74211 1 91
2 74212 1 91
2 74213 1 91
2 74214 1 91
2 74215 1 91
2 74216 1 91
2 74217 1 91
2 74218 1 91
2 74219 1 91
2 74220 1 91
2 74221 1 91
2 74222 1 91
2 74223 1 91
2 74224 1 91
2 74225 1 91
2 74226 1 91
2 74227 1 91
2 74228 1 101
2 74229 1 101
2 74230 1 101
2 74231 1 101
2 74232 1 101
2 74233 1 101
2 74234 1 101
2 74235 1 101
2 74236 1 101
2 74237 1 101
2 74238 1 101
2 74239 1 101
2 74240 1 101
2 74241 1 101
2 74242 1 101
2 74243 1 101
2 74244 1 101
2 74245 1 101
2 74246 1 101
2 74247 1 101
2 74248 1 101
2 74249 1 101
2 74250 1 101
2 74251 1 101
2 74252 1 101
2 74253 1 101
2 74254 1 101
2 74255 1 101
2 74256 1 101
2 74257 1 101
2 74258 1 102
2 74259 1 102
2 74260 1 102
2 74261 1 102
2 74262 1 102
2 74263 1 102
2 74264 1 102
2 74265 1 102
2 74266 1 102
2 74267 1 102
2 74268 1 102
2 74269 1 102
2 74270 1 103
2 74271 1 103
2 74272 1 103
2 74273 1 103
2 74274 1 103
2 74275 1 103
2 74276 1 103
2 74277 1 104
2 74278 1 104
2 74279 1 104
2 74280 1 104
2 74281 1 104
2 74282 1 104
2 74283 1 104
2 74284 1 104
2 74285 1 104
2 74286 1 104
2 74287 1 104
2 74288 1 104
2 74289 1 104
2 74290 1 104
2 74291 1 105
2 74292 1 105
2 74293 1 105
2 74294 1 105
2 74295 1 105
2 74296 1 105
2 74297 1 105
2 74298 1 105
2 74299 1 105
2 74300 1 105
2 74301 1 106
2 74302 1 106
2 74303 1 109
2 74304 1 109
2 74305 1 109
2 74306 1 110
2 74307 1 110
2 74308 1 111
2 74309 1 111
2 74310 1 111
2 74311 1 111
2 74312 1 111
2 74313 1 111
2 74314 1 111
2 74315 1 111
2 74316 1 111
2 74317 1 111
2 74318 1 111
2 74319 1 111
2 74320 1 111
2 74321 1 111
2 74322 1 112
2 74323 1 112
2 74324 1 112
2 74325 1 114
2 74326 1 114
2 74327 1 114
2 74328 1 114
2 74329 1 114
2 74330 1 114
2 74331 1 114
2 74332 1 114
2 74333 1 114
2 74334 1 114
2 74335 1 114
2 74336 1 114
2 74337 1 114
2 74338 1 114
2 74339 1 116
2 74340 1 116
2 74341 1 116
2 74342 1 116
2 74343 1 116
2 74344 1 116
2 74345 1 116
2 74346 1 116
2 74347 1 116
2 74348 1 118
2 74349 1 118
2 74350 1 118
2 74351 1 118
2 74352 1 118
2 74353 1 118
2 74354 1 118
2 74355 1 118
2 74356 1 118
2 74357 1 118
2 74358 1 118
2 74359 1 118
2 74360 1 118
2 74361 1 119
2 74362 1 119
2 74363 1 128
2 74364 1 128
2 74365 1 128
2 74366 1 128
2 74367 1 128
2 74368 1 128
2 74369 1 128
2 74370 1 128
2 74371 1 128
2 74372 1 128
2 74373 1 128
2 74374 1 128
2 74375 1 128
2 74376 1 128
2 74377 1 128
2 74378 1 128
2 74379 1 128
2 74380 1 128
2 74381 1 128
2 74382 1 128
2 74383 1 128
2 74384 1 128
2 74385 1 128
2 74386 1 128
2 74387 1 128
2 74388 1 128
2 74389 1 128
2 74390 1 128
2 74391 1 128
2 74392 1 128
2 74393 1 128
2 74394 1 128
2 74395 1 128
2 74396 1 128
2 74397 1 128
2 74398 1 128
2 74399 1 128
2 74400 1 128
2 74401 1 128
2 74402 1 128
2 74403 1 128
2 74404 1 128
2 74405 1 128
2 74406 1 128
2 74407 1 128
2 74408 1 128
2 74409 1 128
2 74410 1 128
2 74411 1 128
2 74412 1 128
2 74413 1 128
2 74414 1 128
2 74415 1 128
2 74416 1 129
2 74417 1 129
2 74418 1 129
2 74419 1 129
2 74420 1 129
2 74421 1 129
2 74422 1 129
2 74423 1 129
2 74424 1 129
2 74425 1 129
2 74426 1 129
2 74427 1 129
2 74428 1 129
2 74429 1 129
2 74430 1 129
2 74431 1 129
2 74432 1 129
2 74433 1 129
2 74434 1 129
2 74435 1 129
2 74436 1 129
2 74437 1 129
2 74438 1 129
2 74439 1 129
2 74440 1 129
2 74441 1 129
2 74442 1 129
2 74443 1 129
2 74444 1 129
2 74445 1 129
2 74446 1 130
2 74447 1 130
2 74448 1 130
2 74449 1 130
2 74450 1 130
2 74451 1 130
2 74452 1 130
2 74453 1 130
2 74454 1 130
2 74455 1 130
2 74456 1 130
2 74457 1 131
2 74458 1 131
2 74459 1 131
2 74460 1 131
2 74461 1 131
2 74462 1 131
2 74463 1 131
2 74464 1 131
2 74465 1 131
2 74466 1 131
2 74467 1 131
2 74468 1 131
2 74469 1 131
2 74470 1 131
2 74471 1 131
2 74472 1 131
2 74473 1 131
2 74474 1 131
2 74475 1 131
2 74476 1 131
2 74477 1 131
2 74478 1 131
2 74479 1 131
2 74480 1 131
2 74481 1 131
2 74482 1 131
2 74483 1 131
2 74484 1 132
2 74485 1 132
2 74486 1 132
2 74487 1 132
2 74488 1 132
2 74489 1 132
2 74490 1 132
2 74491 1 132
2 74492 1 133
2 74493 1 133
2 74494 1 133
2 74495 1 134
2 74496 1 134
2 74497 1 134
2 74498 1 134
2 74499 1 135
2 74500 1 135
2 74501 1 135
2 74502 1 135
2 74503 1 135
2 74504 1 135
2 74505 1 135
2 74506 1 135
2 74507 1 135
2 74508 1 135
2 74509 1 135
2 74510 1 135
2 74511 1 135
2 74512 1 135
2 74513 1 135
2 74514 1 135
2 74515 1 135
2 74516 1 135
2 74517 1 135
2 74518 1 135
2 74519 1 135
2 74520 1 135
2 74521 1 135
2 74522 1 135
2 74523 1 135
2 74524 1 135
2 74525 1 135
2 74526 1 135
2 74527 1 135
2 74528 1 135
2 74529 1 135
2 74530 1 135
2 74531 1 135
2 74532 1 135
2 74533 1 135
2 74534 1 135
2 74535 1 135
2 74536 1 135
2 74537 1 135
2 74538 1 135
2 74539 1 135
2 74540 1 135
2 74541 1 135
2 74542 1 135
2 74543 1 135
2 74544 1 135
2 74545 1 135
2 74546 1 135
2 74547 1 135
2 74548 1 135
2 74549 1 135
2 74550 1 135
2 74551 1 135
2 74552 1 135
2 74553 1 135
2 74554 1 135
2 74555 1 135
2 74556 1 135
2 74557 1 135
2 74558 1 135
2 74559 1 135
2 74560 1 135
2 74561 1 135
2 74562 1 135
2 74563 1 135
2 74564 1 135
2 74565 1 135
2 74566 1 135
2 74567 1 135
2 74568 1 135
2 74569 1 135
2 74570 1 135
2 74571 1 135
2 74572 1 135
2 74573 1 135
2 74574 1 135
2 74575 1 135
2 74576 1 135
2 74577 1 135
2 74578 1 135
2 74579 1 135
2 74580 1 135
2 74581 1 136
2 74582 1 136
2 74583 1 136
2 74584 1 136
2 74585 1 136
2 74586 1 136
2 74587 1 136
2 74588 1 136
2 74589 1 136
2 74590 1 136
2 74591 1 136
2 74592 1 136
2 74593 1 136
2 74594 1 136
2 74595 1 136
2 74596 1 136
2 74597 1 136
2 74598 1 136
2 74599 1 136
2 74600 1 136
2 74601 1 136
2 74602 1 136
2 74603 1 136
2 74604 1 136
2 74605 1 136
2 74606 1 136
2 74607 1 136
2 74608 1 136
2 74609 1 136
2 74610 1 136
2 74611 1 136
2 74612 1 136
2 74613 1 136
2 74614 1 136
2 74615 1 136
2 74616 1 136
2 74617 1 136
2 74618 1 136
2 74619 1 136
2 74620 1 136
2 74621 1 136
2 74622 1 136
2 74623 1 136
2 74624 1 136
2 74625 1 136
2 74626 1 136
2 74627 1 136
2 74628 1 136
2 74629 1 136
2 74630 1 136
2 74631 1 136
2 74632 1 136
2 74633 1 136
2 74634 1 136
2 74635 1 136
2 74636 1 136
2 74637 1 136
2 74638 1 136
2 74639 1 136
2 74640 1 136
2 74641 1 136
2 74642 1 136
2 74643 1 136
2 74644 1 136
2 74645 1 136
2 74646 1 136
2 74647 1 136
2 74648 1 136
2 74649 1 136
2 74650 1 136
2 74651 1 136
2 74652 1 136
2 74653 1 136
2 74654 1 136
2 74655 1 136
2 74656 1 136
2 74657 1 136
2 74658 1 136
2 74659 1 136
2 74660 1 136
2 74661 1 136
2 74662 1 136
2 74663 1 136
2 74664 1 136
2 74665 1 136
2 74666 1 136
2 74667 1 136
2 74668 1 136
2 74669 1 136
2 74670 1 136
2 74671 1 136
2 74672 1 136
2 74673 1 136
2 74674 1 136
2 74675 1 136
2 74676 1 136
2 74677 1 136
2 74678 1 136
2 74679 1 136
2 74680 1 136
2 74681 1 136
2 74682 1 136
2 74683 1 136
2 74684 1 136
2 74685 1 136
2 74686 1 136
2 74687 1 136
2 74688 1 136
2 74689 1 136
2 74690 1 136
2 74691 1 136
2 74692 1 136
2 74693 1 136
2 74694 1 136
2 74695 1 136
2 74696 1 136
2 74697 1 136
2 74698 1 136
2 74699 1 136
2 74700 1 136
2 74701 1 136
2 74702 1 136
2 74703 1 136
2 74704 1 136
2 74705 1 136
2 74706 1 136
2 74707 1 136
2 74708 1 136
2 74709 1 136
2 74710 1 136
2 74711 1 136
2 74712 1 136
2 74713 1 136
2 74714 1 136
2 74715 1 136
2 74716 1 137
2 74717 1 137
2 74718 1 137
2 74719 1 137
2 74720 1 137
2 74721 1 137
2 74722 1 137
2 74723 1 137
2 74724 1 137
2 74725 1 137
2 74726 1 137
2 74727 1 137
2 74728 1 137
2 74729 1 137
2 74730 1 137
2 74731 1 137
2 74732 1 137
2 74733 1 137
2 74734 1 137
2 74735 1 137
2 74736 1 137
2 74737 1 137
2 74738 1 137
2 74739 1 137
2 74740 1 137
2 74741 1 137
2 74742 1 137
2 74743 1 137
2 74744 1 137
2 74745 1 137
2 74746 1 137
2 74747 1 137
2 74748 1 137
2 74749 1 138
2 74750 1 138
2 74751 1 138
2 74752 1 138
2 74753 1 138
2 74754 1 138
2 74755 1 138
2 74756 1 139
2 74757 1 139
2 74758 1 139
2 74759 1 140
2 74760 1 140
2 74761 1 140
2 74762 1 141
2 74763 1 141
2 74764 1 145
2 74765 1 145
2 74766 1 145
2 74767 1 145
2 74768 1 145
2 74769 1 145
2 74770 1 145
2 74771 1 145
2 74772 1 145
2 74773 1 145
2 74774 1 145
2 74775 1 145
2 74776 1 145
2 74777 1 145
2 74778 1 145
2 74779 1 145
2 74780 1 145
2 74781 1 145
2 74782 1 145
2 74783 1 145
2 74784 1 145
2 74785 1 145
2 74786 1 145
2 74787 1 145
2 74788 1 145
2 74789 1 145
2 74790 1 145
2 74791 1 145
2 74792 1 145
2 74793 1 145
2 74794 1 145
2 74795 1 145
2 74796 1 145
2 74797 1 145
2 74798 1 145
2 74799 1 145
2 74800 1 145
2 74801 1 145
2 74802 1 145
2 74803 1 145
2 74804 1 145
2 74805 1 146
2 74806 1 146
2 74807 1 146
2 74808 1 146
2 74809 1 146
2 74810 1 147
2 74811 1 147
2 74812 1 147
2 74813 1 147
2 74814 1 147
2 74815 1 148
2 74816 1 148
2 74817 1 148
2 74818 1 149
2 74819 1 149
2 74820 1 149
2 74821 1 149
2 74822 1 149
2 74823 1 149
2 74824 1 149
2 74825 1 150
2 74826 1 150
2 74827 1 150
2 74828 1 161
2 74829 1 161
2 74830 1 161
2 74831 1 161
2 74832 1 161
2 74833 1 161
2 74834 1 161
2 74835 1 161
2 74836 1 161
2 74837 1 161
2 74838 1 161
2 74839 1 161
2 74840 1 161
2 74841 1 161
2 74842 1 161
2 74843 1 161
2 74844 1 161
2 74845 1 161
2 74846 1 161
2 74847 1 161
2 74848 1 161
2 74849 1 161
2 74850 1 161
2 74851 1 161
2 74852 1 161
2 74853 1 161
2 74854 1 161
2 74855 1 161
2 74856 1 161
2 74857 1 161
2 74858 1 161
2 74859 1 161
2 74860 1 161
2 74861 1 161
2 74862 1 161
2 74863 1 161
2 74864 1 161
2 74865 1 162
2 74866 1 162
2 74867 1 162
2 74868 1 162
2 74869 1 162
2 74870 1 162
2 74871 1 162
2 74872 1 162
2 74873 1 162
2 74874 1 162
2 74875 1 162
2 74876 1 162
2 74877 1 162
2 74878 1 162
2 74879 1 162
2 74880 1 162
2 74881 1 162
2 74882 1 162
2 74883 1 162
2 74884 1 163
2 74885 1 163
2 74886 1 163
2 74887 1 164
2 74888 1 164
2 74889 1 164
2 74890 1 164
2 74891 1 164
2 74892 1 165
2 74893 1 165
2 74894 1 165
2 74895 1 165
2 74896 1 165
2 74897 1 165
2 74898 1 165
2 74899 1 165
2 74900 1 165
2 74901 1 165
2 74902 1 165
2 74903 1 165
2 74904 1 165
2 74905 1 165
2 74906 1 165
2 74907 1 165
2 74908 1 165
2 74909 1 165
2 74910 1 165
2 74911 1 165
2 74912 1 165
2 74913 1 165
2 74914 1 167
2 74915 1 167
2 74916 1 174
2 74917 1 174
2 74918 1 174
2 74919 1 174
2 74920 1 174
2 74921 1 174
2 74922 1 174
2 74923 1 175
2 74924 1 175
2 74925 1 175
2 74926 1 175
2 74927 1 175
2 74928 1 176
2 74929 1 176
2 74930 1 177
2 74931 1 177
2 74932 1 177
2 74933 1 177
2 74934 1 177
2 74935 1 177
2 74936 1 177
2 74937 1 177
2 74938 1 177
2 74939 1 177
2 74940 1 177
2 74941 1 177
2 74942 1 177
2 74943 1 177
2 74944 1 177
2 74945 1 177
2 74946 1 177
2 74947 1 177
2 74948 1 177
2 74949 1 177
2 74950 1 177
2 74951 1 177
2 74952 1 177
2 74953 1 177
2 74954 1 177
2 74955 1 177
2 74956 1 177
2 74957 1 177
2 74958 1 177
2 74959 1 177
2 74960 1 177
2 74961 1 177
2 74962 1 177
2 74963 1 177
2 74964 1 177
2 74965 1 177
2 74966 1 177
2 74967 1 177
2 74968 1 177
2 74969 1 177
2 74970 1 177
2 74971 1 177
2 74972 1 177
2 74973 1 177
2 74974 1 177
2 74975 1 177
2 74976 1 177
2 74977 1 177
2 74978 1 177
2 74979 1 177
2 74980 1 177
2 74981 1 177
2 74982 1 177
2 74983 1 177
2 74984 1 177
2 74985 1 177
2 74986 1 178
2 74987 1 178
2 74988 1 178
2 74989 1 178
2 74990 1 178
2 74991 1 178
2 74992 1 178
2 74993 1 178
2 74994 1 178
2 74995 1 178
2 74996 1 178
2 74997 1 178
2 74998 1 178
2 74999 1 178
2 75000 1 178
2 75001 1 178
2 75002 1 178
2 75003 1 178
2 75004 1 178
2 75005 1 178
2 75006 1 178
2 75007 1 178
2 75008 1 178
2 75009 1 178
2 75010 1 178
2 75011 1 178
2 75012 1 178
2 75013 1 178
2 75014 1 178
2 75015 1 178
2 75016 1 178
2 75017 1 178
2 75018 1 178
2 75019 1 178
2 75020 1 178
2 75021 1 178
2 75022 1 178
2 75023 1 178
2 75024 1 178
2 75025 1 178
2 75026 1 179
2 75027 1 179
2 75028 1 179
2 75029 1 179
2 75030 1 179
2 75031 1 179
2 75032 1 179
2 75033 1 179
2 75034 1 179
2 75035 1 180
2 75036 1 180
2 75037 1 180
2 75038 1 180
2 75039 1 180
2 75040 1 180
2 75041 1 180
2 75042 1 180
2 75043 1 180
2 75044 1 180
2 75045 1 180
2 75046 1 180
2 75047 1 180
2 75048 1 180
2 75049 1 180
2 75050 1 180
2 75051 1 180
2 75052 1 180
2 75053 1 180
2 75054 1 189
2 75055 1 189
2 75056 1 189
2 75057 1 189
2 75058 1 189
2 75059 1 189
2 75060 1 189
2 75061 1 189
2 75062 1 189
2 75063 1 189
2 75064 1 190
2 75065 1 190
2 75066 1 190
2 75067 1 190
2 75068 1 190
2 75069 1 190
2 75070 1 191
2 75071 1 191
2 75072 1 191
2 75073 1 191
2 75074 1 191
2 75075 1 191
2 75076 1 191
2 75077 1 191
2 75078 1 191
2 75079 1 191
2 75080 1 191
2 75081 1 191
2 75082 1 191
2 75083 1 191
2 75084 1 191
2 75085 1 191
2 75086 1 191
2 75087 1 191
2 75088 1 192
2 75089 1 192
2 75090 1 192
2 75091 1 192
2 75092 1 192
2 75093 1 193
2 75094 1 193
2 75095 1 193
2 75096 1 193
2 75097 1 193
2 75098 1 193
2 75099 1 193
2 75100 1 193
2 75101 1 193
2 75102 1 193
2 75103 1 193
2 75104 1 193
2 75105 1 193
2 75106 1 193
2 75107 1 193
2 75108 1 193
2 75109 1 193
2 75110 1 193
2 75111 1 194
2 75112 1 194
2 75113 1 194
2 75114 1 194
2 75115 1 194
2 75116 1 194
2 75117 1 194
2 75118 1 194
2 75119 1 194
2 75120 1 194
2 75121 1 194
2 75122 1 194
2 75123 1 194
2 75124 1 194
2 75125 1 194
2 75126 1 194
2 75127 1 194
2 75128 1 194
2 75129 1 194
2 75130 1 194
2 75131 1 194
2 75132 1 194
2 75133 1 194
2 75134 1 194
2 75135 1 194
2 75136 1 195
2 75137 1 195
2 75138 1 196
2 75139 1 196
2 75140 1 196
2 75141 1 196
2 75142 1 201
2 75143 1 201
2 75144 1 201
2 75145 1 201
2 75146 1 201
2 75147 1 201
2 75148 1 201
2 75149 1 202
2 75150 1 202
2 75151 1 202
2 75152 1 202
2 75153 1 202
2 75154 1 202
2 75155 1 202
2 75156 1 202
2 75157 1 202
2 75158 1 202
2 75159 1 202
2 75160 1 202
2 75161 1 202
2 75162 1 202
2 75163 1 202
2 75164 1 202
2 75165 1 202
2 75166 1 202
2 75167 1 202
2 75168 1 202
2 75169 1 202
2 75170 1 202
2 75171 1 203
2 75172 1 203
2 75173 1 203
2 75174 1 203
2 75175 1 203
2 75176 1 203
2 75177 1 203
2 75178 1 203
2 75179 1 203
2 75180 1 203
2 75181 1 203
2 75182 1 203
2 75183 1 203
2 75184 1 203
2 75185 1 203
2 75186 1 203
2 75187 1 203
2 75188 1 203
2 75189 1 211
2 75190 1 211
2 75191 1 211
2 75192 1 211
2 75193 1 211
2 75194 1 211
2 75195 1 211
2 75196 1 211
2 75197 1 211
2 75198 1 211
2 75199 1 211
2 75200 1 212
2 75201 1 212
2 75202 1 212
2 75203 1 212
2 75204 1 212
2 75205 1 212
2 75206 1 212
2 75207 1 212
2 75208 1 212
2 75209 1 212
2 75210 1 212
2 75211 1 212
2 75212 1 212
2 75213 1 212
2 75214 1 212
2 75215 1 212
2 75216 1 212
2 75217 1 212
2 75218 1 212
2 75219 1 212
2 75220 1 212
2 75221 1 212
2 75222 1 212
2 75223 1 212
2 75224 1 212
2 75225 1 212
2 75226 1 212
2 75227 1 212
2 75228 1 212
2 75229 1 212
2 75230 1 212
2 75231 1 212
2 75232 1 212
2 75233 1 212
2 75234 1 212
2 75235 1 212
2 75236 1 212
2 75237 1 212
2 75238 1 212
2 75239 1 213
2 75240 1 213
2 75241 1 214
2 75242 1 214
2 75243 1 214
2 75244 1 214
2 75245 1 214
2 75246 1 214
2 75247 1 214
2 75248 1 214
2 75249 1 214
2 75250 1 214
2 75251 1 214
2 75252 1 214
2 75253 1 214
2 75254 1 214
2 75255 1 214
2 75256 1 214
2 75257 1 214
2 75258 1 214
2 75259 1 214
2 75260 1 214
2 75261 1 214
2 75262 1 214
2 75263 1 214
2 75264 1 214
2 75265 1 214
2 75266 1 214
2 75267 1 214
2 75268 1 214
2 75269 1 214
2 75270 1 214
2 75271 1 214
2 75272 1 214
2 75273 1 214
2 75274 1 214
2 75275 1 214
2 75276 1 214
2 75277 1 214
2 75278 1 214
2 75279 1 214
2 75280 1 214
2 75281 1 214
2 75282 1 214
2 75283 1 214
2 75284 1 214
2 75285 1 214
2 75286 1 214
2 75287 1 214
2 75288 1 214
2 75289 1 214
2 75290 1 214
2 75291 1 214
2 75292 1 214
2 75293 1 214
2 75294 1 214
2 75295 1 214
2 75296 1 214
2 75297 1 214
2 75298 1 214
2 75299 1 214
2 75300 1 214
2 75301 1 214
2 75302 1 214
2 75303 1 215
2 75304 1 215
2 75305 1 215
2 75306 1 215
2 75307 1 215
2 75308 1 215
2 75309 1 215
2 75310 1 215
2 75311 1 215
2 75312 1 215
2 75313 1 215
2 75314 1 215
2 75315 1 215
2 75316 1 215
2 75317 1 215
2 75318 1 215
2 75319 1 215
2 75320 1 215
2 75321 1 215
2 75322 1 215
2 75323 1 215
2 75324 1 215
2 75325 1 215
2 75326 1 215
2 75327 1 215
2 75328 1 215
2 75329 1 215
2 75330 1 215
2 75331 1 215
2 75332 1 215
2 75333 1 215
2 75334 1 215
2 75335 1 215
2 75336 1 215
2 75337 1 215
2 75338 1 215
2 75339 1 215
2 75340 1 215
2 75341 1 215
2 75342 1 215
2 75343 1 215
2 75344 1 215
2 75345 1 215
2 75346 1 215
2 75347 1 215
2 75348 1 215
2 75349 1 215
2 75350 1 215
2 75351 1 215
2 75352 1 215
2 75353 1 215
2 75354 1 215
2 75355 1 215
2 75356 1 215
2 75357 1 215
2 75358 1 215
2 75359 1 215
2 75360 1 215
2 75361 1 215
2 75362 1 215
2 75363 1 215
2 75364 1 215
2 75365 1 215
2 75366 1 215
2 75367 1 215
2 75368 1 215
2 75369 1 215
2 75370 1 215
2 75371 1 215
2 75372 1 215
2 75373 1 215
2 75374 1 215
2 75375 1 215
2 75376 1 215
2 75377 1 215
2 75378 1 215
2 75379 1 215
2 75380 1 215
2 75381 1 215
2 75382 1 215
2 75383 1 215
2 75384 1 215
2 75385 1 215
2 75386 1 215
2 75387 1 215
2 75388 1 215
2 75389 1 215
2 75390 1 215
2 75391 1 215
2 75392 1 215
2 75393 1 215
2 75394 1 215
2 75395 1 215
2 75396 1 215
2 75397 1 215
2 75398 1 215
2 75399 1 215
2 75400 1 215
2 75401 1 215
2 75402 1 215
2 75403 1 215
2 75404 1 215
2 75405 1 215
2 75406 1 215
2 75407 1 215
2 75408 1 215
2 75409 1 215
2 75410 1 215
2 75411 1 215
2 75412 1 215
2 75413 1 215
2 75414 1 215
2 75415 1 215
2 75416 1 215
2 75417 1 215
2 75418 1 215
2 75419 1 215
2 75420 1 215
2 75421 1 215
2 75422 1 215
2 75423 1 215
2 75424 1 215
2 75425 1 215
2 75426 1 215
2 75427 1 215
2 75428 1 215
2 75429 1 215
2 75430 1 215
2 75431 1 215
2 75432 1 215
2 75433 1 215
2 75434 1 215
2 75435 1 215
2 75436 1 215
2 75437 1 215
2 75438 1 215
2 75439 1 215
2 75440 1 215
2 75441 1 215
2 75442 1 215
2 75443 1 215
2 75444 1 215
2 75445 1 215
2 75446 1 215
2 75447 1 215
2 75448 1 215
2 75449 1 215
2 75450 1 215
2 75451 1 215
2 75452 1 215
2 75453 1 215
2 75454 1 215
2 75455 1 215
2 75456 1 215
2 75457 1 215
2 75458 1 215
2 75459 1 215
2 75460 1 215
2 75461 1 215
2 75462 1 215
2 75463 1 215
2 75464 1 215
2 75465 1 215
2 75466 1 215
2 75467 1 215
2 75468 1 215
2 75469 1 216
2 75470 1 216
2 75471 1 216
2 75472 1 216
2 75473 1 216
2 75474 1 216
2 75475 1 216
2 75476 1 216
2 75477 1 217
2 75478 1 217
2 75479 1 218
2 75480 1 218
2 75481 1 218
2 75482 1 218
2 75483 1 220
2 75484 1 220
2 75485 1 220
2 75486 1 220
2 75487 1 220
2 75488 1 220
2 75489 1 220
2 75490 1 221
2 75491 1 221
2 75492 1 222
2 75493 1 222
2 75494 1 222
2 75495 1 225
2 75496 1 225
2 75497 1 225
2 75498 1 225
2 75499 1 225
2 75500 1 225
2 75501 1 225
2 75502 1 225
2 75503 1 225
2 75504 1 225
2 75505 1 225
2 75506 1 225
2 75507 1 225
2 75508 1 225
2 75509 1 225
2 75510 1 225
2 75511 1 225
2 75512 1 225
2 75513 1 225
2 75514 1 226
2 75515 1 226
2 75516 1 226
2 75517 1 227
2 75518 1 227
2 75519 1 227
2 75520 1 227
2 75521 1 228
2 75522 1 228
2 75523 1 228
2 75524 1 228
2 75525 1 228
2 75526 1 228
2 75527 1 228
2 75528 1 229
2 75529 1 229
2 75530 1 229
2 75531 1 229
2 75532 1 229
2 75533 1 229
2 75534 1 229
2 75535 1 229
2 75536 1 229
2 75537 1 229
2 75538 1 235
2 75539 1 235
2 75540 1 235
2 75541 1 235
2 75542 1 235
2 75543 1 235
2 75544 1 235
2 75545 1 235
2 75546 1 235
2 75547 1 235
2 75548 1 235
2 75549 1 235
2 75550 1 235
2 75551 1 235
2 75552 1 235
2 75553 1 235
2 75554 1 235
2 75555 1 235
2 75556 1 235
2 75557 1 235
2 75558 1 235
2 75559 1 235
2 75560 1 235
2 75561 1 235
2 75562 1 235
2 75563 1 235
2 75564 1 235
2 75565 1 235
2 75566 1 235
2 75567 1 235
2 75568 1 235
2 75569 1 235
2 75570 1 235
2 75571 1 235
2 75572 1 235
2 75573 1 235
2 75574 1 235
2 75575 1 235
2 75576 1 235
2 75577 1 235
2 75578 1 235
2 75579 1 235
2 75580 1 235
2 75581 1 235
2 75582 1 235
2 75583 1 235
2 75584 1 235
2 75585 1 236
2 75586 1 236
2 75587 1 236
2 75588 1 236
2 75589 1 237
2 75590 1 237
2 75591 1 237
2 75592 1 237
2 75593 1 237
2 75594 1 237
2 75595 1 245
2 75596 1 245
2 75597 1 245
2 75598 1 245
2 75599 1 245
2 75600 1 245
2 75601 1 245
2 75602 1 245
2 75603 1 245
2 75604 1 245
2 75605 1 245
2 75606 1 245
2 75607 1 245
2 75608 1 245
2 75609 1 245
2 75610 1 245
2 75611 1 245
2 75612 1 245
2 75613 1 246
2 75614 1 246
2 75615 1 246
2 75616 1 246
2 75617 1 246
2 75618 1 246
2 75619 1 246
2 75620 1 246
2 75621 1 246
2 75622 1 246
2 75623 1 246
2 75624 1 246
2 75625 1 246
2 75626 1 246
2 75627 1 246
2 75628 1 246
2 75629 1 246
2 75630 1 246
2 75631 1 246
2 75632 1 247
2 75633 1 247
2 75634 1 247
2 75635 1 247
2 75636 1 248
2 75637 1 248
2 75638 1 249
2 75639 1 249
2 75640 1 252
2 75641 1 252
2 75642 1 252
2 75643 1 252
2 75644 1 252
2 75645 1 252
2 75646 1 252
2 75647 1 252
2 75648 1 252
2 75649 1 252
2 75650 1 252
2 75651 1 253
2 75652 1 253
2 75653 1 253
2 75654 1 253
2 75655 1 254
2 75656 1 254
2 75657 1 255
2 75658 1 255
2 75659 1 262
2 75660 1 262
2 75661 1 262
2 75662 1 262
2 75663 1 262
2 75664 1 262
2 75665 1 262
2 75666 1 262
2 75667 1 262
2 75668 1 262
2 75669 1 262
2 75670 1 262
2 75671 1 262
2 75672 1 263
2 75673 1 263
2 75674 1 263
2 75675 1 263
2 75676 1 264
2 75677 1 264
2 75678 1 264
2 75679 1 264
2 75680 1 264
2 75681 1 264
2 75682 1 264
2 75683 1 264
2 75684 1 265
2 75685 1 265
2 75686 1 272
2 75687 1 272
2 75688 1 272
2 75689 1 272
2 75690 1 272
2 75691 1 272
2 75692 1 272
2 75693 1 272
2 75694 1 272
2 75695 1 272
2 75696 1 272
2 75697 1 273
2 75698 1 273
2 75699 1 273
2 75700 1 274
2 75701 1 274
2 75702 1 275
2 75703 1 275
2 75704 1 276
2 75705 1 276
2 75706 1 276
2 75707 1 276
2 75708 1 276
2 75709 1 276
2 75710 1 276
2 75711 1 276
2 75712 1 277
2 75713 1 277
2 75714 1 277
2 75715 1 277
2 75716 1 277
2 75717 1 277
2 75718 1 277
2 75719 1 277
2 75720 1 277
2 75721 1 277
2 75722 1 277
2 75723 1 277
2 75724 1 277
2 75725 1 277
2 75726 1 277
2 75727 1 277
2 75728 1 277
2 75729 1 277
2 75730 1 277
2 75731 1 277
2 75732 1 277
2 75733 1 277
2 75734 1 277
2 75735 1 277
2 75736 1 277
2 75737 1 277
2 75738 1 277
2 75739 1 277
2 75740 1 277
2 75741 1 277
2 75742 1 277
2 75743 1 277
2 75744 1 277
2 75745 1 277
2 75746 1 277
2 75747 1 277
2 75748 1 277
2 75749 1 277
2 75750 1 277
2 75751 1 277
2 75752 1 277
2 75753 1 277
2 75754 1 277
2 75755 1 277
2 75756 1 277
2 75757 1 277
2 75758 1 277
2 75759 1 277
2 75760 1 277
2 75761 1 277
2 75762 1 277
2 75763 1 277
2 75764 1 277
2 75765 1 278
2 75766 1 278
2 75767 1 278
2 75768 1 278
2 75769 1 278
2 75770 1 278
2 75771 1 278
2 75772 1 278
2 75773 1 278
2 75774 1 278
2 75775 1 278
2 75776 1 282
2 75777 1 282
2 75778 1 282
2 75779 1 282
2 75780 1 282
2 75781 1 282
2 75782 1 282
2 75783 1 282
2 75784 1 282
2 75785 1 282
2 75786 1 282
2 75787 1 282
2 75788 1 283
2 75789 1 283
2 75790 1 283
2 75791 1 283
2 75792 1 284
2 75793 1 284
2 75794 1 287
2 75795 1 287
2 75796 1 288
2 75797 1 288
2 75798 1 288
2 75799 1 288
2 75800 1 288
2 75801 1 288
2 75802 1 288
2 75803 1 288
2 75804 1 288
2 75805 1 288
2 75806 1 288
2 75807 1 288
2 75808 1 288
2 75809 1 288
2 75810 1 288
2 75811 1 289
2 75812 1 289
2 75813 1 289
2 75814 1 289
2 75815 1 289
2 75816 1 289
2 75817 1 289
2 75818 1 289
2 75819 1 289
2 75820 1 289
2 75821 1 289
2 75822 1 289
2 75823 1 289
2 75824 1 289
2 75825 1 289
2 75826 1 289
2 75827 1 289
2 75828 1 290
2 75829 1 290
2 75830 1 290
2 75831 1 290
2 75832 1 290
2 75833 1 290
2 75834 1 290
2 75835 1 290
2 75836 1 290
2 75837 1 290
2 75838 1 290
2 75839 1 290
2 75840 1 290
2 75841 1 296
2 75842 1 296
2 75843 1 296
2 75844 1 296
2 75845 1 296
2 75846 1 296
2 75847 1 296
2 75848 1 296
2 75849 1 296
2 75850 1 296
2 75851 1 296
2 75852 1 296
2 75853 1 296
2 75854 1 297
2 75855 1 297
2 75856 1 297
2 75857 1 298
2 75858 1 298
2 75859 1 298
2 75860 1 298
2 75861 1 298
2 75862 1 306
2 75863 1 306
2 75864 1 306
2 75865 1 306
2 75866 1 307
2 75867 1 307
2 75868 1 307
2 75869 1 307
2 75870 1 307
2 75871 1 307
2 75872 1 307
2 75873 1 307
2 75874 1 307
2 75875 1 307
2 75876 1 307
2 75877 1 307
2 75878 1 307
2 75879 1 307
2 75880 1 307
2 75881 1 307
2 75882 1 307
2 75883 1 307
2 75884 1 307
2 75885 1 309
2 75886 1 309
2 75887 1 309
2 75888 1 310
2 75889 1 310
2 75890 1 310
2 75891 1 310
2 75892 1 313
2 75893 1 313
2 75894 1 316
2 75895 1 316
2 75896 1 316
2 75897 1 316
2 75898 1 316
2 75899 1 316
2 75900 1 316
2 75901 1 316
2 75902 1 316
2 75903 1 316
2 75904 1 316
2 75905 1 316
2 75906 1 316
2 75907 1 316
2 75908 1 316
2 75909 1 316
2 75910 1 316
2 75911 1 316
2 75912 1 316
2 75913 1 316
2 75914 1 316
2 75915 1 316
2 75916 1 316
2 75917 1 316
2 75918 1 316
2 75919 1 316
2 75920 1 316
2 75921 1 316
2 75922 1 316
2 75923 1 316
2 75924 1 316
2 75925 1 316
2 75926 1 316
2 75927 1 316
2 75928 1 316
2 75929 1 316
2 75930 1 316
2 75931 1 316
2 75932 1 316
2 75933 1 316
2 75934 1 316
2 75935 1 316
2 75936 1 316
2 75937 1 316
2 75938 1 316
2 75939 1 316
2 75940 1 316
2 75941 1 316
2 75942 1 316
2 75943 1 316
2 75944 1 316
2 75945 1 316
2 75946 1 317
2 75947 1 317
2 75948 1 317
2 75949 1 317
2 75950 1 317
2 75951 1 317
2 75952 1 317
2 75953 1 317
2 75954 1 317
2 75955 1 317
2 75956 1 317
2 75957 1 317
2 75958 1 317
2 75959 1 317
2 75960 1 317
2 75961 1 317
2 75962 1 317
2 75963 1 317
2 75964 1 317
2 75965 1 317
2 75966 1 317
2 75967 1 317
2 75968 1 317
2 75969 1 317
2 75970 1 317
2 75971 1 317
2 75972 1 317
2 75973 1 317
2 75974 1 317
2 75975 1 317
2 75976 1 317
2 75977 1 317
2 75978 1 317
2 75979 1 317
2 75980 1 317
2 75981 1 317
2 75982 1 317
2 75983 1 317
2 75984 1 317
2 75985 1 317
2 75986 1 317
2 75987 1 317
2 75988 1 317
2 75989 1 317
2 75990 1 317
2 75991 1 317
2 75992 1 317
2 75993 1 318
2 75994 1 318
2 75995 1 320
2 75996 1 320
2 75997 1 320
2 75998 1 320
2 75999 1 320
2 76000 1 320
2 76001 1 320
2 76002 1 320
2 76003 1 320
2 76004 1 320
2 76005 1 320
2 76006 1 320
2 76007 1 322
2 76008 1 322
2 76009 1 322
2 76010 1 322
2 76011 1 322
2 76012 1 322
2 76013 1 323
2 76014 1 323
2 76015 1 323
2 76016 1 330
2 76017 1 330
2 76018 1 330
2 76019 1 330
2 76020 1 330
2 76021 1 330
2 76022 1 330
2 76023 1 330
2 76024 1 330
2 76025 1 330
2 76026 1 330
2 76027 1 330
2 76028 1 330
2 76029 1 330
2 76030 1 330
2 76031 1 330
2 76032 1 330
2 76033 1 330
2 76034 1 330
2 76035 1 331
2 76036 1 331
2 76037 1 331
2 76038 1 331
2 76039 1 331
2 76040 1 331
2 76041 1 332
2 76042 1 332
2 76043 1 332
2 76044 1 332
2 76045 1 332
2 76046 1 332
2 76047 1 332
2 76048 1 332
2 76049 1 332
2 76050 1 332
2 76051 1 332
2 76052 1 332
2 76053 1 332
2 76054 1 332
2 76055 1 333
2 76056 1 333
2 76057 1 333
2 76058 1 333
2 76059 1 334
2 76060 1 334
2 76061 1 334
2 76062 1 335
2 76063 1 335
2 76064 1 335
2 76065 1 335
2 76066 1 335
2 76067 1 335
2 76068 1 335
2 76069 1 335
2 76070 1 335
2 76071 1 335
2 76072 1 335
2 76073 1 335
2 76074 1 335
2 76075 1 335
2 76076 1 335
2 76077 1 335
2 76078 1 335
2 76079 1 335
2 76080 1 335
2 76081 1 335
2 76082 1 335
2 76083 1 335
2 76084 1 335
2 76085 1 335
2 76086 1 335
2 76087 1 335
2 76088 1 335
2 76089 1 335
2 76090 1 335
2 76091 1 335
2 76092 1 335
2 76093 1 335
2 76094 1 335
2 76095 1 335
2 76096 1 335
2 76097 1 335
2 76098 1 335
2 76099 1 335
2 76100 1 335
2 76101 1 335
2 76102 1 335
2 76103 1 335
2 76104 1 335
2 76105 1 335
2 76106 1 335
2 76107 1 335
2 76108 1 335
2 76109 1 335
2 76110 1 335
2 76111 1 335
2 76112 1 335
2 76113 1 335
2 76114 1 336
2 76115 1 336
2 76116 1 336
2 76117 1 336
2 76118 1 336
2 76119 1 336
2 76120 1 337
2 76121 1 337
2 76122 1 337
2 76123 1 337
2 76124 1 338
2 76125 1 338
2 76126 1 338
2 76127 1 342
2 76128 1 342
2 76129 1 342
2 76130 1 342
2 76131 1 342
2 76132 1 342
2 76133 1 342
2 76134 1 342
2 76135 1 342
2 76136 1 342
2 76137 1 343
2 76138 1 343
2 76139 1 344
2 76140 1 344
2 76141 1 344
2 76142 1 344
2 76143 1 344
2 76144 1 344
2 76145 1 344
2 76146 1 344
2 76147 1 344
2 76148 1 344
2 76149 1 344
2 76150 1 344
2 76151 1 344
2 76152 1 344
2 76153 1 344
2 76154 1 344
2 76155 1 344
2 76156 1 344
2 76157 1 344
2 76158 1 344
2 76159 1 344
2 76160 1 344
2 76161 1 344
2 76162 1 344
2 76163 1 344
2 76164 1 344
2 76165 1 344
2 76166 1 344
2 76167 1 344
2 76168 1 346
2 76169 1 346
2 76170 1 346
2 76171 1 346
2 76172 1 355
2 76173 1 355
2 76174 1 355
2 76175 1 355
2 76176 1 355
2 76177 1 355
2 76178 1 355
2 76179 1 355
2 76180 1 355
2 76181 1 355
2 76182 1 355
2 76183 1 355
2 76184 1 355
2 76185 1 355
2 76186 1 355
2 76187 1 355
2 76188 1 355
2 76189 1 355
2 76190 1 355
2 76191 1 355
2 76192 1 355
2 76193 1 355
2 76194 1 355
2 76195 1 355
2 76196 1 355
2 76197 1 355
2 76198 1 355
2 76199 1 355
2 76200 1 355
2 76201 1 355
2 76202 1 355
2 76203 1 355
2 76204 1 355
2 76205 1 355
2 76206 1 355
2 76207 1 355
2 76208 1 355
2 76209 1 355
2 76210 1 355
2 76211 1 355
2 76212 1 355
2 76213 1 355
2 76214 1 355
2 76215 1 355
2 76216 1 355
2 76217 1 355
2 76218 1 355
2 76219 1 355
2 76220 1 355
2 76221 1 355
2 76222 1 355
2 76223 1 355
2 76224 1 355
2 76225 1 355
2 76226 1 355
2 76227 1 355
2 76228 1 355
2 76229 1 355
2 76230 1 355
2 76231 1 355
2 76232 1 355
2 76233 1 355
2 76234 1 355
2 76235 1 355
2 76236 1 355
2 76237 1 355
2 76238 1 355
2 76239 1 355
2 76240 1 355
2 76241 1 355
2 76242 1 355
2 76243 1 355
2 76244 1 355
2 76245 1 355
2 76246 1 355
2 76247 1 355
2 76248 1 355
2 76249 1 355
2 76250 1 355
2 76251 1 355
2 76252 1 355
2 76253 1 355
2 76254 1 355
2 76255 1 355
2 76256 1 356
2 76257 1 356
2 76258 1 356
2 76259 1 356
2 76260 1 356
2 76261 1 356
2 76262 1 356
2 76263 1 356
2 76264 1 356
2 76265 1 356
2 76266 1 356
2 76267 1 356
2 76268 1 356
2 76269 1 356
2 76270 1 356
2 76271 1 356
2 76272 1 356
2 76273 1 356
2 76274 1 356
2 76275 1 356
2 76276 1 356
2 76277 1 356
2 76278 1 356
2 76279 1 356
2 76280 1 356
2 76281 1 356
2 76282 1 356
2 76283 1 356
2 76284 1 356
2 76285 1 356
2 76286 1 356
2 76287 1 356
2 76288 1 356
2 76289 1 356
2 76290 1 356
2 76291 1 356
2 76292 1 356
2 76293 1 356
2 76294 1 356
2 76295 1 356
2 76296 1 356
2 76297 1 356
2 76298 1 356
2 76299 1 356
2 76300 1 356
2 76301 1 356
2 76302 1 356
2 76303 1 356
2 76304 1 356
2 76305 1 356
2 76306 1 356
2 76307 1 356
2 76308 1 356
2 76309 1 356
2 76310 1 356
2 76311 1 356
2 76312 1 356
2 76313 1 356
2 76314 1 356
2 76315 1 356
2 76316 1 356
2 76317 1 356
2 76318 1 356
2 76319 1 356
2 76320 1 356
2 76321 1 356
2 76322 1 356
2 76323 1 356
2 76324 1 356
2 76325 1 356
2 76326 1 356
2 76327 1 356
2 76328 1 356
2 76329 1 356
2 76330 1 356
2 76331 1 356
2 76332 1 356
2 76333 1 356
2 76334 1 356
2 76335 1 356
2 76336 1 356
2 76337 1 356
2 76338 1 356
2 76339 1 356
2 76340 1 356
2 76341 1 356
2 76342 1 356
2 76343 1 356
2 76344 1 356
2 76345 1 356
2 76346 1 356
2 76347 1 357
2 76348 1 357
2 76349 1 361
2 76350 1 361
2 76351 1 361
2 76352 1 361
2 76353 1 361
2 76354 1 361
2 76355 1 361
2 76356 1 361
2 76357 1 361
2 76358 1 361
2 76359 1 369
2 76360 1 369
2 76361 1 369
2 76362 1 369
2 76363 1 369
2 76364 1 369
2 76365 1 369
2 76366 1 369
2 76367 1 369
2 76368 1 369
2 76369 1 369
2 76370 1 369
2 76371 1 369
2 76372 1 369
2 76373 1 369
2 76374 1 369
2 76375 1 369
2 76376 1 369
2 76377 1 369
2 76378 1 369
2 76379 1 369
2 76380 1 369
2 76381 1 369
2 76382 1 369
2 76383 1 369
2 76384 1 369
2 76385 1 369
2 76386 1 369
2 76387 1 369
2 76388 1 369
2 76389 1 369
2 76390 1 369
2 76391 1 369
2 76392 1 369
2 76393 1 369
2 76394 1 369
2 76395 1 369
2 76396 1 369
2 76397 1 369
2 76398 1 369
2 76399 1 369
2 76400 1 370
2 76401 1 370
2 76402 1 371
2 76403 1 371
2 76404 1 371
2 76405 1 371
2 76406 1 371
2 76407 1 371
2 76408 1 371
2 76409 1 371
2 76410 1 371
2 76411 1 371
2 76412 1 371
2 76413 1 371
2 76414 1 371
2 76415 1 371
2 76416 1 371
2 76417 1 371
2 76418 1 371
2 76419 1 371
2 76420 1 371
2 76421 1 371
2 76422 1 371
2 76423 1 371
2 76424 1 371
2 76425 1 371
2 76426 1 381
2 76427 1 381
2 76428 1 381
2 76429 1 381
2 76430 1 381
2 76431 1 382
2 76432 1 382
2 76433 1 382
2 76434 1 382
2 76435 1 382
2 76436 1 382
2 76437 1 382
2 76438 1 382
2 76439 1 382
2 76440 1 382
2 76441 1 382
2 76442 1 382
2 76443 1 382
2 76444 1 382
2 76445 1 382
2 76446 1 382
2 76447 1 382
2 76448 1 382
2 76449 1 382
2 76450 1 382
2 76451 1 382
2 76452 1 382
2 76453 1 382
2 76454 1 382
2 76455 1 382
2 76456 1 382
2 76457 1 382
2 76458 1 382
2 76459 1 382
2 76460 1 382
2 76461 1 382
2 76462 1 382
2 76463 1 382
2 76464 1 382
2 76465 1 382
2 76466 1 382
2 76467 1 382
2 76468 1 382
2 76469 1 382
2 76470 1 382
2 76471 1 382
2 76472 1 382
2 76473 1 382
2 76474 1 382
2 76475 1 382
2 76476 1 382
2 76477 1 382
2 76478 1 382
2 76479 1 382
2 76480 1 382
2 76481 1 382
2 76482 1 382
2 76483 1 382
2 76484 1 382
2 76485 1 382
2 76486 1 382
2 76487 1 382
2 76488 1 382
2 76489 1 382
2 76490 1 382
2 76491 1 382
2 76492 1 382
2 76493 1 382
2 76494 1 382
2 76495 1 382
2 76496 1 382
2 76497 1 382
2 76498 1 382
2 76499 1 382
2 76500 1 382
2 76501 1 382
2 76502 1 382
2 76503 1 382
2 76504 1 382
2 76505 1 382
2 76506 1 382
2 76507 1 382
2 76508 1 382
2 76509 1 382
2 76510 1 382
2 76511 1 382
2 76512 1 382
2 76513 1 382
2 76514 1 382
2 76515 1 382
2 76516 1 382
2 76517 1 382
2 76518 1 382
2 76519 1 382
2 76520 1 382
2 76521 1 382
2 76522 1 382
2 76523 1 382
2 76524 1 382
2 76525 1 382
2 76526 1 383
2 76527 1 383
2 76528 1 383
2 76529 1 383
2 76530 1 383
2 76531 1 383
2 76532 1 383
2 76533 1 383
2 76534 1 383
2 76535 1 383
2 76536 1 383
2 76537 1 383
2 76538 1 383
2 76539 1 383
2 76540 1 383
2 76541 1 383
2 76542 1 383
2 76543 1 383
2 76544 1 383
2 76545 1 383
2 76546 1 383
2 76547 1 383
2 76548 1 383
2 76549 1 383
2 76550 1 383
2 76551 1 383
2 76552 1 383
2 76553 1 383
2 76554 1 383
2 76555 1 383
2 76556 1 383
2 76557 1 383
2 76558 1 383
2 76559 1 383
2 76560 1 383
2 76561 1 383
2 76562 1 383
2 76563 1 383
2 76564 1 383
2 76565 1 383
2 76566 1 383
2 76567 1 383
2 76568 1 383
2 76569 1 383
2 76570 1 383
2 76571 1 383
2 76572 1 383
2 76573 1 383
2 76574 1 383
2 76575 1 383
2 76576 1 383
2 76577 1 383
2 76578 1 383
2 76579 1 383
2 76580 1 383
2 76581 1 383
2 76582 1 383
2 76583 1 383
2 76584 1 383
2 76585 1 383
2 76586 1 383
2 76587 1 383
2 76588 1 383
2 76589 1 383
2 76590 1 383
2 76591 1 383
2 76592 1 383
2 76593 1 383
2 76594 1 383
2 76595 1 383
2 76596 1 383
2 76597 1 383
2 76598 1 383
2 76599 1 383
2 76600 1 383
2 76601 1 383
2 76602 1 383
2 76603 1 383
2 76604 1 383
2 76605 1 383
2 76606 1 383
2 76607 1 383
2 76608 1 383
2 76609 1 383
2 76610 1 383
2 76611 1 383
2 76612 1 383
2 76613 1 383
2 76614 1 383
2 76615 1 383
2 76616 1 383
2 76617 1 384
2 76618 1 384
2 76619 1 384
2 76620 1 384
2 76621 1 384
2 76622 1 384
2 76623 1 384
2 76624 1 384
2 76625 1 385
2 76626 1 385
2 76627 1 386
2 76628 1 386
2 76629 1 386
2 76630 1 395
2 76631 1 395
2 76632 1 395
2 76633 1 395
2 76634 1 396
2 76635 1 396
2 76636 1 396
2 76637 1 396
2 76638 1 396
2 76639 1 396
2 76640 1 396
2 76641 1 396
2 76642 1 396
2 76643 1 396
2 76644 1 396
2 76645 1 396
2 76646 1 396
2 76647 1 396
2 76648 1 396
2 76649 1 396
2 76650 1 396
2 76651 1 396
2 76652 1 396
2 76653 1 396
2 76654 1 396
2 76655 1 396
2 76656 1 396
2 76657 1 396
2 76658 1 396
2 76659 1 396
2 76660 1 396
2 76661 1 396
2 76662 1 396
2 76663 1 396
2 76664 1 396
2 76665 1 396
2 76666 1 396
2 76667 1 396
2 76668 1 397
2 76669 1 397
2 76670 1 397
2 76671 1 397
2 76672 1 397
2 76673 1 397
2 76674 1 397
2 76675 1 397
2 76676 1 397
2 76677 1 397
2 76678 1 397
2 76679 1 397
2 76680 1 397
2 76681 1 397
2 76682 1 397
2 76683 1 397
2 76684 1 397
2 76685 1 397
2 76686 1 397
2 76687 1 397
2 76688 1 397
2 76689 1 397
2 76690 1 397
2 76691 1 397
2 76692 1 397
2 76693 1 397
2 76694 1 397
2 76695 1 398
2 76696 1 398
2 76697 1 398
2 76698 1 399
2 76699 1 399
2 76700 1 399
2 76701 1 399
2 76702 1 399
2 76703 1 399
2 76704 1 399
2 76705 1 399
2 76706 1 399
2 76707 1 399
2 76708 1 399
2 76709 1 399
2 76710 1 399
2 76711 1 399
2 76712 1 399
2 76713 1 399
2 76714 1 399
2 76715 1 399
2 76716 1 400
2 76717 1 400
2 76718 1 403
2 76719 1 403
2 76720 1 403
2 76721 1 403
2 76722 1 403
2 76723 1 403
2 76724 1 403
2 76725 1 403
2 76726 1 403
2 76727 1 403
2 76728 1 403
2 76729 1 403
2 76730 1 403
2 76731 1 403
2 76732 1 403
2 76733 1 403
2 76734 1 403
2 76735 1 403
2 76736 1 403
2 76737 1 403
2 76738 1 403
2 76739 1 404
2 76740 1 404
2 76741 1 404
2 76742 1 404
2 76743 1 404
2 76744 1 405
2 76745 1 405
2 76746 1 405
2 76747 1 405
2 76748 1 407
2 76749 1 407
2 76750 1 407
2 76751 1 407
2 76752 1 407
2 76753 1 407
2 76754 1 407
2 76755 1 407
2 76756 1 418
2 76757 1 418
2 76758 1 418
2 76759 1 418
2 76760 1 418
2 76761 1 418
2 76762 1 418
2 76763 1 418
2 76764 1 418
2 76765 1 418
2 76766 1 418
2 76767 1 418
2 76768 1 418
2 76769 1 418
2 76770 1 418
2 76771 1 418
2 76772 1 418
2 76773 1 418
2 76774 1 418
2 76775 1 418
2 76776 1 418
2 76777 1 418
2 76778 1 418
2 76779 1 418
2 76780 1 420
2 76781 1 420
2 76782 1 420
2 76783 1 420
2 76784 1 420
2 76785 1 420
2 76786 1 420
2 76787 1 420
2 76788 1 420
2 76789 1 420
2 76790 1 420
2 76791 1 420
2 76792 1 422
2 76793 1 422
2 76794 1 422
2 76795 1 422
2 76796 1 422
2 76797 1 422
2 76798 1 422
2 76799 1 422
2 76800 1 422
2 76801 1 422
2 76802 1 422
2 76803 1 422
2 76804 1 422
2 76805 1 422
2 76806 1 422
2 76807 1 422
2 76808 1 422
2 76809 1 422
2 76810 1 422
2 76811 1 422
2 76812 1 422
2 76813 1 422
2 76814 1 422
2 76815 1 422
2 76816 1 422
2 76817 1 431
2 76818 1 431
2 76819 1 431
2 76820 1 431
2 76821 1 431
2 76822 1 431
2 76823 1 431
2 76824 1 431
2 76825 1 431
2 76826 1 431
2 76827 1 431
2 76828 1 431
2 76829 1 434
2 76830 1 434
2 76831 1 434
2 76832 1 434
2 76833 1 434
2 76834 1 434
2 76835 1 434
2 76836 1 434
2 76837 1 434
2 76838 1 434
2 76839 1 434
2 76840 1 434
2 76841 1 434
2 76842 1 434
2 76843 1 434
2 76844 1 434
2 76845 1 434
2 76846 1 434
2 76847 1 434
2 76848 1 434
2 76849 1 434
2 76850 1 434
2 76851 1 434
2 76852 1 434
2 76853 1 434
2 76854 1 434
2 76855 1 434
2 76856 1 434
2 76857 1 434
2 76858 1 434
2 76859 1 434
2 76860 1 434
2 76861 1 434
2 76862 1 435
2 76863 1 435
2 76864 1 435
2 76865 1 435
2 76866 1 436
2 76867 1 436
2 76868 1 436
2 76869 1 436
2 76870 1 436
2 76871 1 436
2 76872 1 436
2 76873 1 436
2 76874 1 436
2 76875 1 436
2 76876 1 436
2 76877 1 437
2 76878 1 437
2 76879 1 437
2 76880 1 437
2 76881 1 437
2 76882 1 437
2 76883 1 437
2 76884 1 437
2 76885 1 437
2 76886 1 437
2 76887 1 437
2 76888 1 437
2 76889 1 437
2 76890 1 437
2 76891 1 437
2 76892 1 437
2 76893 1 437
2 76894 1 438
2 76895 1 438
2 76896 1 446
2 76897 1 446
2 76898 1 446
2 76899 1 446
2 76900 1 446
2 76901 1 446
2 76902 1 446
2 76903 1 446
2 76904 1 446
2 76905 1 446
2 76906 1 446
2 76907 1 446
2 76908 1 447
2 76909 1 447
2 76910 1 448
2 76911 1 448
2 76912 1 448
2 76913 1 448
2 76914 1 448
2 76915 1 448
2 76916 1 448
2 76917 1 448
2 76918 1 448
2 76919 1 448
2 76920 1 448
2 76921 1 448
2 76922 1 448
2 76923 1 448
2 76924 1 448
2 76925 1 449
2 76926 1 449
2 76927 1 449
2 76928 1 449
2 76929 1 449
2 76930 1 449
2 76931 1 449
2 76932 1 449
2 76933 1 449
2 76934 1 449
2 76935 1 449
2 76936 1 449
2 76937 1 449
2 76938 1 449
2 76939 1 449
2 76940 1 449
2 76941 1 449
2 76942 1 449
2 76943 1 449
2 76944 1 451
2 76945 1 451
2 76946 1 459
2 76947 1 459
2 76948 1 459
2 76949 1 459
2 76950 1 459
2 76951 1 459
2 76952 1 459
2 76953 1 459
2 76954 1 459
2 76955 1 459
2 76956 1 459
2 76957 1 459
2 76958 1 459
2 76959 1 459
2 76960 1 459
2 76961 1 459
2 76962 1 459
2 76963 1 459
2 76964 1 459
2 76965 1 459
2 76966 1 459
2 76967 1 459
2 76968 1 459
2 76969 1 460
2 76970 1 460
2 76971 1 461
2 76972 1 461
2 76973 1 461
2 76974 1 462
2 76975 1 462
2 76976 1 462
2 76977 1 462
2 76978 1 462
2 76979 1 462
2 76980 1 463
2 76981 1 463
2 76982 1 474
2 76983 1 474
2 76984 1 474
2 76985 1 474
2 76986 1 474
2 76987 1 474
2 76988 1 474
2 76989 1 474
2 76990 1 474
2 76991 1 474
2 76992 1 474
2 76993 1 474
2 76994 1 474
2 76995 1 474
2 76996 1 474
2 76997 1 474
2 76998 1 474
2 76999 1 474
2 77000 1 474
2 77001 1 474
2 77002 1 474
2 77003 1 474
2 77004 1 474
2 77005 1 474
2 77006 1 474
2 77007 1 475
2 77008 1 475
2 77009 1 475
2 77010 1 476
2 77011 1 476
2 77012 1 476
2 77013 1 476
2 77014 1 476
2 77015 1 476
2 77016 1 476
2 77017 1 476
2 77018 1 476
2 77019 1 476
2 77020 1 476
2 77021 1 476
2 77022 1 476
2 77023 1 477
2 77024 1 477
2 77025 1 477
2 77026 1 478
2 77027 1 478
2 77028 1 478
2 77029 1 478
2 77030 1 478
2 77031 1 481
2 77032 1 481
2 77033 1 481
2 77034 1 481
2 77035 1 481
2 77036 1 481
2 77037 1 482
2 77038 1 482
2 77039 1 482
2 77040 1 482
2 77041 1 482
2 77042 1 482
2 77043 1 482
2 77044 1 482
2 77045 1 482
2 77046 1 482
2 77047 1 482
2 77048 1 482
2 77049 1 482
2 77050 1 482
2 77051 1 482
2 77052 1 482
2 77053 1 482
2 77054 1 483
2 77055 1 483
2 77056 1 483
2 77057 1 484
2 77058 1 484
2 77059 1 484
2 77060 1 484
2 77061 1 484
2 77062 1 484
2 77063 1 484
2 77064 1 484
2 77065 1 484
2 77066 1 484
2 77067 1 484
2 77068 1 484
2 77069 1 484
2 77070 1 484
2 77071 1 484
2 77072 1 484
2 77073 1 484
2 77074 1 484
2 77075 1 484
2 77076 1 485
2 77077 1 485
2 77078 1 492
2 77079 1 492
2 77080 1 492
2 77081 1 492
2 77082 1 492
2 77083 1 492
2 77084 1 492
2 77085 1 492
2 77086 1 492
2 77087 1 492
2 77088 1 492
2 77089 1 492
2 77090 1 492
2 77091 1 492
2 77092 1 493
2 77093 1 493
2 77094 1 493
2 77095 1 493
2 77096 1 493
2 77097 1 493
2 77098 1 493
2 77099 1 493
2 77100 1 493
2 77101 1 493
2 77102 1 493
2 77103 1 493
2 77104 1 493
2 77105 1 493
2 77106 1 493
2 77107 1 494
2 77108 1 494
2 77109 1 494
2 77110 1 494
2 77111 1 494
2 77112 1 494
2 77113 1 494
2 77114 1 494
2 77115 1 494
2 77116 1 494
2 77117 1 495
2 77118 1 495
2 77119 1 495
2 77120 1 495
2 77121 1 495
2 77122 1 495
2 77123 1 495
2 77124 1 495
2 77125 1 495
2 77126 1 495
2 77127 1 495
2 77128 1 495
2 77129 1 495
2 77130 1 496
2 77131 1 496
2 77132 1 497
2 77133 1 497
2 77134 1 498
2 77135 1 498
2 77136 1 498
2 77137 1 498
2 77138 1 498
2 77139 1 498
2 77140 1 498
2 77141 1 498
2 77142 1 498
2 77143 1 498
2 77144 1 498
2 77145 1 498
2 77146 1 498
2 77147 1 498
2 77148 1 498
2 77149 1 498
2 77150 1 498
2 77151 1 498
2 77152 1 498
2 77153 1 498
2 77154 1 498
2 77155 1 498
2 77156 1 498
2 77157 1 498
2 77158 1 498
2 77159 1 498
2 77160 1 498
2 77161 1 498
2 77162 1 498
2 77163 1 498
2 77164 1 498
2 77165 1 498
2 77166 1 498
2 77167 1 498
2 77168 1 498
2 77169 1 498
2 77170 1 498
2 77171 1 498
2 77172 1 498
2 77173 1 498
2 77174 1 498
2 77175 1 498
2 77176 1 498
2 77177 1 498
2 77178 1 498
2 77179 1 498
2 77180 1 498
2 77181 1 498
2 77182 1 498
2 77183 1 498
2 77184 1 498
2 77185 1 498
2 77186 1 498
2 77187 1 498
2 77188 1 498
2 77189 1 498
2 77190 1 498
2 77191 1 498
2 77192 1 498
2 77193 1 498
2 77194 1 498
2 77195 1 498
2 77196 1 498
2 77197 1 498
2 77198 1 499
2 77199 1 499
2 77200 1 499
2 77201 1 499
2 77202 1 499
2 77203 1 499
2 77204 1 499
2 77205 1 499
2 77206 1 499
2 77207 1 499
2 77208 1 499
2 77209 1 499
2 77210 1 499
2 77211 1 499
2 77212 1 499
2 77213 1 499
2 77214 1 499
2 77215 1 499
2 77216 1 499
2 77217 1 499
2 77218 1 499
2 77219 1 499
2 77220 1 499
2 77221 1 499
2 77222 1 499
2 77223 1 499
2 77224 1 499
2 77225 1 499
2 77226 1 499
2 77227 1 499
2 77228 1 499
2 77229 1 499
2 77230 1 499
2 77231 1 499
2 77232 1 499
2 77233 1 499
2 77234 1 499
2 77235 1 499
2 77236 1 499
2 77237 1 499
2 77238 1 499
2 77239 1 499
2 77240 1 499
2 77241 1 499
2 77242 1 499
2 77243 1 499
2 77244 1 499
2 77245 1 499
2 77246 1 499
2 77247 1 499
2 77248 1 499
2 77249 1 499
2 77250 1 499
2 77251 1 499
2 77252 1 499
2 77253 1 499
2 77254 1 499
2 77255 1 499
2 77256 1 499
2 77257 1 499
2 77258 1 499
2 77259 1 499
2 77260 1 499
2 77261 1 499
2 77262 1 499
2 77263 1 499
2 77264 1 499
2 77265 1 499
2 77266 1 499
2 77267 1 499
2 77268 1 499
2 77269 1 499
2 77270 1 499
2 77271 1 499
2 77272 1 499
2 77273 1 499
2 77274 1 499
2 77275 1 499
2 77276 1 499
2 77277 1 503
2 77278 1 503
2 77279 1 503
2 77280 1 503
2 77281 1 503
2 77282 1 503
2 77283 1 503
2 77284 1 503
2 77285 1 503
2 77286 1 503
2 77287 1 503
2 77288 1 503
2 77289 1 504
2 77290 1 504
2 77291 1 504
2 77292 1 504
2 77293 1 504
2 77294 1 504
2 77295 1 504
2 77296 1 505
2 77297 1 505
2 77298 1 505
2 77299 1 505
2 77300 1 505
2 77301 1 506
2 77302 1 506
2 77303 1 506
2 77304 1 506
2 77305 1 506
2 77306 1 506
2 77307 1 506
2 77308 1 506
2 77309 1 506
2 77310 1 506
2 77311 1 506
2 77312 1 506
2 77313 1 506
2 77314 1 507
2 77315 1 507
2 77316 1 507
2 77317 1 507
2 77318 1 507
2 77319 1 507
2 77320 1 507
2 77321 1 507
2 77322 1 507
2 77323 1 507
2 77324 1 507
2 77325 1 507
2 77326 1 507
2 77327 1 507
2 77328 1 507
2 77329 1 507
2 77330 1 507
2 77331 1 507
2 77332 1 507
2 77333 1 507
2 77334 1 507
2 77335 1 507
2 77336 1 507
2 77337 1 507
2 77338 1 507
2 77339 1 507
2 77340 1 507
2 77341 1 507
2 77342 1 507
2 77343 1 507
2 77344 1 507
2 77345 1 507
2 77346 1 507
2 77347 1 507
2 77348 1 507
2 77349 1 507
2 77350 1 507
2 77351 1 507
2 77352 1 507
2 77353 1 507
2 77354 1 507
2 77355 1 507
2 77356 1 507
2 77357 1 507
2 77358 1 507
2 77359 1 507
2 77360 1 507
2 77361 1 507
2 77362 1 507
2 77363 1 507
2 77364 1 507
2 77365 1 507
2 77366 1 507
2 77367 1 507
2 77368 1 507
2 77369 1 507
2 77370 1 507
2 77371 1 507
2 77372 1 507
2 77373 1 507
2 77374 1 507
2 77375 1 507
2 77376 1 507
2 77377 1 507
2 77378 1 507
2 77379 1 507
2 77380 1 507
2 77381 1 507
2 77382 1 507
2 77383 1 507
2 77384 1 507
2 77385 1 507
2 77386 1 507
2 77387 1 507
2 77388 1 508
2 77389 1 508
2 77390 1 508
2 77391 1 508
2 77392 1 508
2 77393 1 508
2 77394 1 508
2 77395 1 508
2 77396 1 508
2 77397 1 508
2 77398 1 508
2 77399 1 508
2 77400 1 508
2 77401 1 508
2 77402 1 508
2 77403 1 508
2 77404 1 508
2 77405 1 508
2 77406 1 508
2 77407 1 508
2 77408 1 508
2 77409 1 508
2 77410 1 508
2 77411 1 508
2 77412 1 508
2 77413 1 508
2 77414 1 508
2 77415 1 508
2 77416 1 508
2 77417 1 508
2 77418 1 508
2 77419 1 508
2 77420 1 508
2 77421 1 508
2 77422 1 508
2 77423 1 508
2 77424 1 508
2 77425 1 508
2 77426 1 508
2 77427 1 508
2 77428 1 508
2 77429 1 508
2 77430 1 508
2 77431 1 508
2 77432 1 508
2 77433 1 508
2 77434 1 508
2 77435 1 508
2 77436 1 508
2 77437 1 508
2 77438 1 508
2 77439 1 508
2 77440 1 508
2 77441 1 508
2 77442 1 508
2 77443 1 508
2 77444 1 508
2 77445 1 508
2 77446 1 508
2 77447 1 508
2 77448 1 508
2 77449 1 508
2 77450 1 508
2 77451 1 508
2 77452 1 508
2 77453 1 508
2 77454 1 508
2 77455 1 508
2 77456 1 508
2 77457 1 508
2 77458 1 508
2 77459 1 508
2 77460 1 508
2 77461 1 508
2 77462 1 508
2 77463 1 508
2 77464 1 508
2 77465 1 508
2 77466 1 508
2 77467 1 508
2 77468 1 508
2 77469 1 508
2 77470 1 508
2 77471 1 508
2 77472 1 508
2 77473 1 508
2 77474 1 508
2 77475 1 508
2 77476 1 508
2 77477 1 508
2 77478 1 508
2 77479 1 508
2 77480 1 508
2 77481 1 508
2 77482 1 508
2 77483 1 508
2 77484 1 508
2 77485 1 508
2 77486 1 508
2 77487 1 508
2 77488 1 508
2 77489 1 508
2 77490 1 508
2 77491 1 508
2 77492 1 508
2 77493 1 510
2 77494 1 510
2 77495 1 511
2 77496 1 511
2 77497 1 511
2 77498 1 511
2 77499 1 511
2 77500 1 511
2 77501 1 511
2 77502 1 511
2 77503 1 511
2 77504 1 511
2 77505 1 512
2 77506 1 512
2 77507 1 515
2 77508 1 515
2 77509 1 515
2 77510 1 515
2 77511 1 516
2 77512 1 516
2 77513 1 518
2 77514 1 518
2 77515 1 518
2 77516 1 518
2 77517 1 520
2 77518 1 520
2 77519 1 520
2 77520 1 520
2 77521 1 520
2 77522 1 520
2 77523 1 520
2 77524 1 520
2 77525 1 520
2 77526 1 520
2 77527 1 520
2 77528 1 520
2 77529 1 520
2 77530 1 520
2 77531 1 529
2 77532 1 529
2 77533 1 529
2 77534 1 529
2 77535 1 529
2 77536 1 529
2 77537 1 529
2 77538 1 529
2 77539 1 529
2 77540 1 529
2 77541 1 529
2 77542 1 529
2 77543 1 529
2 77544 1 529
2 77545 1 529
2 77546 1 529
2 77547 1 529
2 77548 1 530
2 77549 1 530
2 77550 1 530
2 77551 1 530
2 77552 1 530
2 77553 1 530
2 77554 1 530
2 77555 1 530
2 77556 1 531
2 77557 1 531
2 77558 1 531
2 77559 1 531
2 77560 1 531
2 77561 1 531
2 77562 1 532
2 77563 1 532
2 77564 1 532
2 77565 1 532
2 77566 1 532
2 77567 1 532
2 77568 1 532
2 77569 1 532
2 77570 1 532
2 77571 1 532
2 77572 1 532
2 77573 1 533
2 77574 1 533
2 77575 1 533
2 77576 1 535
2 77577 1 535
2 77578 1 535
2 77579 1 536
2 77580 1 536
2 77581 1 539
2 77582 1 539
2 77583 1 539
2 77584 1 540
2 77585 1 540
2 77586 1 540
2 77587 1 540
2 77588 1 540
2 77589 1 540
2 77590 1 540
2 77591 1 544
2 77592 1 544
2 77593 1 547
2 77594 1 547
2 77595 1 547
2 77596 1 547
2 77597 1 547
2 77598 1 547
2 77599 1 547
2 77600 1 547
2 77601 1 547
2 77602 1 547
2 77603 1 548
2 77604 1 548
2 77605 1 548
2 77606 1 548
2 77607 1 548
2 77608 1 548
2 77609 1 548
2 77610 1 548
2 77611 1 548
2 77612 1 548
2 77613 1 548
2 77614 1 548
2 77615 1 548
2 77616 1 548
2 77617 1 550
2 77618 1 550
2 77619 1 551
2 77620 1 551
2 77621 1 552
2 77622 1 552
2 77623 1 559
2 77624 1 559
2 77625 1 559
2 77626 1 560
2 77627 1 560
2 77628 1 560
2 77629 1 560
2 77630 1 560
2 77631 1 560
2 77632 1 560
2 77633 1 563
2 77634 1 563
2 77635 1 563
2 77636 1 563
2 77637 1 563
2 77638 1 563
2 77639 1 563
2 77640 1 563
2 77641 1 564
2 77642 1 564
2 77643 1 564
2 77644 1 564
2 77645 1 566
2 77646 1 566
2 77647 1 567
2 77648 1 567
2 77649 1 567
2 77650 1 567
2 77651 1 567
2 77652 1 567
2 77653 1 567
2 77654 1 567
2 77655 1 567
2 77656 1 567
2 77657 1 567
2 77658 1 567
2 77659 1 567
2 77660 1 567
2 77661 1 567
2 77662 1 567
2 77663 1 567
2 77664 1 567
2 77665 1 567
2 77666 1 567
2 77667 1 567
2 77668 1 567
2 77669 1 567
2 77670 1 567
2 77671 1 567
2 77672 1 567
2 77673 1 567
2 77674 1 567
2 77675 1 567
2 77676 1 567
2 77677 1 567
2 77678 1 567
2 77679 1 567
2 77680 1 567
2 77681 1 567
2 77682 1 567
2 77683 1 567
2 77684 1 567
2 77685 1 568
2 77686 1 568
2 77687 1 568
2 77688 1 568
2 77689 1 568
2 77690 1 568
2 77691 1 568
2 77692 1 568
2 77693 1 568
2 77694 1 569
2 77695 1 569
2 77696 1 569
2 77697 1 569
2 77698 1 569
2 77699 1 569
2 77700 1 569
2 77701 1 569
2 77702 1 569
2 77703 1 570
2 77704 1 570
2 77705 1 570
2 77706 1 570
2 77707 1 578
2 77708 1 578
2 77709 1 578
2 77710 1 578
2 77711 1 578
2 77712 1 578
2 77713 1 578
2 77714 1 578
2 77715 1 578
2 77716 1 578
2 77717 1 578
2 77718 1 579
2 77719 1 579
2 77720 1 579
2 77721 1 579
2 77722 1 579
2 77723 1 579
2 77724 1 579
2 77725 1 579
2 77726 1 579
2 77727 1 579
2 77728 1 579
2 77729 1 579
2 77730 1 579
2 77731 1 579
2 77732 1 579
2 77733 1 579
2 77734 1 579
2 77735 1 579
2 77736 1 580
2 77737 1 580
2 77738 1 580
2 77739 1 581
2 77740 1 581
2 77741 1 583
2 77742 1 583
2 77743 1 583
2 77744 1 583
2 77745 1 583
2 77746 1 583
2 77747 1 583
2 77748 1 583
2 77749 1 583
2 77750 1 583
2 77751 1 583
2 77752 1 583
2 77753 1 583
2 77754 1 583
2 77755 1 583
2 77756 1 583
2 77757 1 583
2 77758 1 583
2 77759 1 584
2 77760 1 584
2 77761 1 584
2 77762 1 599
2 77763 1 599
2 77764 1 599
2 77765 1 600
2 77766 1 600
2 77767 1 600
2 77768 1 600
2 77769 1 600
2 77770 1 600
2 77771 1 600
2 77772 1 600
2 77773 1 600
2 77774 1 600
2 77775 1 600
2 77776 1 600
2 77777 1 600
2 77778 1 600
2 77779 1 600
2 77780 1 600
2 77781 1 600
2 77782 1 601
2 77783 1 601
2 77784 1 601
2 77785 1 601
2 77786 1 601
2 77787 1 602
2 77788 1 602
2 77789 1 603
2 77790 1 603
2 77791 1 603
2 77792 1 603
2 77793 1 603
2 77794 1 603
2 77795 1 604
2 77796 1 604
2 77797 1 604
2 77798 1 604
2 77799 1 604
2 77800 1 604
2 77801 1 604
2 77802 1 604
2 77803 1 604
2 77804 1 604
2 77805 1 604
2 77806 1 604
2 77807 1 604
2 77808 1 604
2 77809 1 604
2 77810 1 604
2 77811 1 606
2 77812 1 606
2 77813 1 606
2 77814 1 606
2 77815 1 606
2 77816 1 618
2 77817 1 618
2 77818 1 618
2 77819 1 618
2 77820 1 618
2 77821 1 618
2 77822 1 618
2 77823 1 618
2 77824 1 618
2 77825 1 618
2 77826 1 618
2 77827 1 618
2 77828 1 618
2 77829 1 618
2 77830 1 618
2 77831 1 618
2 77832 1 618
2 77833 1 618
2 77834 1 618
2 77835 1 618
2 77836 1 618
2 77837 1 619
2 77838 1 619
2 77839 1 619
2 77840 1 619
2 77841 1 619
2 77842 1 619
2 77843 1 620
2 77844 1 620
2 77845 1 621
2 77846 1 621
2 77847 1 624
2 77848 1 624
2 77849 1 624
2 77850 1 624
2 77851 1 624
2 77852 1 624
2 77853 1 625
2 77854 1 625
2 77855 1 625
2 77856 1 626
2 77857 1 626
2 77858 1 626
2 77859 1 626
2 77860 1 626
2 77861 1 626
2 77862 1 626
2 77863 1 626
2 77864 1 626
2 77865 1 626
2 77866 1 626
2 77867 1 626
2 77868 1 626
2 77869 1 626
2 77870 1 626
2 77871 1 626
2 77872 1 626
2 77873 1 626
2 77874 1 626
2 77875 1 626
2 77876 1 626
2 77877 1 626
2 77878 1 626
2 77879 1 627
2 77880 1 627
2 77881 1 627
2 77882 1 628
2 77883 1 628
2 77884 1 628
2 77885 1 628
2 77886 1 628
2 77887 1 628
2 77888 1 632
2 77889 1 632
2 77890 1 640
2 77891 1 640
2 77892 1 640
2 77893 1 640
2 77894 1 640
2 77895 1 640
2 77896 1 640
2 77897 1 640
2 77898 1 640
2 77899 1 640
2 77900 1 640
2 77901 1 640
2 77902 1 640
2 77903 1 640
2 77904 1 640
2 77905 1 640
2 77906 1 640
2 77907 1 640
2 77908 1 640
2 77909 1 640
2 77910 1 640
2 77911 1 640
2 77912 1 640
2 77913 1 640
2 77914 1 640
2 77915 1 641
2 77916 1 641
2 77917 1 641
2 77918 1 641
2 77919 1 641
2 77920 1 641
2 77921 1 641
2 77922 1 641
2 77923 1 642
2 77924 1 642
2 77925 1 642
2 77926 1 643
2 77927 1 643
2 77928 1 643
2 77929 1 643
2 77930 1 645
2 77931 1 645
2 77932 1 645
2 77933 1 645
2 77934 1 646
2 77935 1 646
2 77936 1 646
2 77937 1 646
2 77938 1 646
2 77939 1 646
2 77940 1 646
2 77941 1 647
2 77942 1 647
2 77943 1 647
2 77944 1 647
2 77945 1 651
2 77946 1 651
2 77947 1 651
2 77948 1 651
2 77949 1 651
2 77950 1 651
2 77951 1 651
2 77952 1 651
2 77953 1 651
2 77954 1 652
2 77955 1 652
2 77956 1 653
2 77957 1 653
2 77958 1 653
2 77959 1 653
2 77960 1 653
2 77961 1 653
2 77962 1 653
2 77963 1 653
2 77964 1 653
2 77965 1 653
2 77966 1 653
2 77967 1 655
2 77968 1 655
2 77969 1 655
2 77970 1 663
2 77971 1 663
2 77972 1 663
2 77973 1 663
2 77974 1 663
2 77975 1 663
2 77976 1 663
2 77977 1 663
2 77978 1 663
2 77979 1 663
2 77980 1 665
2 77981 1 665
2 77982 1 666
2 77983 1 666
2 77984 1 666
2 77985 1 666
2 77986 1 666
2 77987 1 666
2 77988 1 666
2 77989 1 666
2 77990 1 666
2 77991 1 666
2 77992 1 666
2 77993 1 666
2 77994 1 666
2 77995 1 666
2 77996 1 666
2 77997 1 666
2 77998 1 666
2 77999 1 667
2 78000 1 667
2 78001 1 667
2 78002 1 667
2 78003 1 667
2 78004 1 671
2 78005 1 671
2 78006 1 671
2 78007 1 671
2 78008 1 673
2 78009 1 673
2 78010 1 673
2 78011 1 673
2 78012 1 673
2 78013 1 673
2 78014 1 673
2 78015 1 673
2 78016 1 673
2 78017 1 673
2 78018 1 673
2 78019 1 673
2 78020 1 673
2 78021 1 673
2 78022 1 673
2 78023 1 674
2 78024 1 674
2 78025 1 674
2 78026 1 674
2 78027 1 675
2 78028 1 675
2 78029 1 675
2 78030 1 675
2 78031 1 675
2 78032 1 675
2 78033 1 675
2 78034 1 676
2 78035 1 676
2 78036 1 676
2 78037 1 678
2 78038 1 678
2 78039 1 684
2 78040 1 684
2 78041 1 684
2 78042 1 685
2 78043 1 685
2 78044 1 685
2 78045 1 687
2 78046 1 687
2 78047 1 687
2 78048 1 687
2 78049 1 689
2 78050 1 689
2 78051 1 694
2 78052 1 694
2 78053 1 694
2 78054 1 694
2 78055 1 694
2 78056 1 695
2 78057 1 695
2 78058 1 696
2 78059 1 696
2 78060 1 696
2 78061 1 696
2 78062 1 696
2 78063 1 697
2 78064 1 697
2 78065 1 698
2 78066 1 698
2 78067 1 720
2 78068 1 720
2 78069 1 720
2 78070 1 720
2 78071 1 720
2 78072 1 720
2 78073 1 720
2 78074 1 720
2 78075 1 720
2 78076 1 720
2 78077 1 720
2 78078 1 720
2 78079 1 720
2 78080 1 720
2 78081 1 720
2 78082 1 720
2 78083 1 720
2 78084 1 720
2 78085 1 720
2 78086 1 721
2 78087 1 721
2 78088 1 721
2 78089 1 721
2 78090 1 721
2 78091 1 721
2 78092 1 721
2 78093 1 721
2 78094 1 721
2 78095 1 721
2 78096 1 721
2 78097 1 721
2 78098 1 721
2 78099 1 721
2 78100 1 721
2 78101 1 721
2 78102 1 722
2 78103 1 722
2 78104 1 722
2 78105 1 722
2 78106 1 722
2 78107 1 723
2 78108 1 723
2 78109 1 723
2 78110 1 723
2 78111 1 723
2 78112 1 723
2 78113 1 723
2 78114 1 723
2 78115 1 723
2 78116 1 723
2 78117 1 724
2 78118 1 724
2 78119 1 724
2 78120 1 728
2 78121 1 728
2 78122 1 728
2 78123 1 728
2 78124 1 728
2 78125 1 728
2 78126 1 728
2 78127 1 728
2 78128 1 728
2 78129 1 728
2 78130 1 728
2 78131 1 728
2 78132 1 728
2 78133 1 728
2 78134 1 728
2 78135 1 728
2 78136 1 729
2 78137 1 729
2 78138 1 729
2 78139 1 729
2 78140 1 729
2 78141 1 729
2 78142 1 730
2 78143 1 730
2 78144 1 730
2 78145 1 730
2 78146 1 730
2 78147 1 730
2 78148 1 730
2 78149 1 730
2 78150 1 730
2 78151 1 730
2 78152 1 732
2 78153 1 732
2 78154 1 732
2 78155 1 732
2 78156 1 732
2 78157 1 732
2 78158 1 732
2 78159 1 732
2 78160 1 732
2 78161 1 732
2 78162 1 732
2 78163 1 732
2 78164 1 732
2 78165 1 732
2 78166 1 732
2 78167 1 732
2 78168 1 732
2 78169 1 732
2 78170 1 732
2 78171 1 732
2 78172 1 732
2 78173 1 732
2 78174 1 732
2 78175 1 732
2 78176 1 732
2 78177 1 732
2 78178 1 732
2 78179 1 732
2 78180 1 732
2 78181 1 732
2 78182 1 732
2 78183 1 732
2 78184 1 732
2 78185 1 732
2 78186 1 732
2 78187 1 732
2 78188 1 732
2 78189 1 733
2 78190 1 733
2 78191 1 733
2 78192 1 733
2 78193 1 733
2 78194 1 733
2 78195 1 733
2 78196 1 733
2 78197 1 733
2 78198 1 733
2 78199 1 733
2 78200 1 733
2 78201 1 733
2 78202 1 733
2 78203 1 733
2 78204 1 733
2 78205 1 733
2 78206 1 733
2 78207 1 733
2 78208 1 733
2 78209 1 733
2 78210 1 733
2 78211 1 733
2 78212 1 733
2 78213 1 733
2 78214 1 733
2 78215 1 733
2 78216 1 733
2 78217 1 733
2 78218 1 733
2 78219 1 733
2 78220 1 733
2 78221 1 733
2 78222 1 733
2 78223 1 733
2 78224 1 733
2 78225 1 733
2 78226 1 733
2 78227 1 733
2 78228 1 733
2 78229 1 733
2 78230 1 733
2 78231 1 733
2 78232 1 733
2 78233 1 733
2 78234 1 733
2 78235 1 733
2 78236 1 733
2 78237 1 733
2 78238 1 733
2 78239 1 733
2 78240 1 733
2 78241 1 733
2 78242 1 733
2 78243 1 733
2 78244 1 733
2 78245 1 733
2 78246 1 733
2 78247 1 733
2 78248 1 733
2 78249 1 733
2 78250 1 733
2 78251 1 733
2 78252 1 733
2 78253 1 733
2 78254 1 733
2 78255 1 733
2 78256 1 733
2 78257 1 733
2 78258 1 733
2 78259 1 733
2 78260 1 733
2 78261 1 733
2 78262 1 733
2 78263 1 733
2 78264 1 733
2 78265 1 733
2 78266 1 733
2 78267 1 733
2 78268 1 733
2 78269 1 733
2 78270 1 733
2 78271 1 733
2 78272 1 733
2 78273 1 733
2 78274 1 733
2 78275 1 733
2 78276 1 733
2 78277 1 733
2 78278 1 733
2 78279 1 733
2 78280 1 734
2 78281 1 734
2 78282 1 735
2 78283 1 735
2 78284 1 739
2 78285 1 739
2 78286 1 739
2 78287 1 739
2 78288 1 739
2 78289 1 739
2 78290 1 739
2 78291 1 739
2 78292 1 741
2 78293 1 741
2 78294 1 741
2 78295 1 741
2 78296 1 741
2 78297 1 741
2 78298 1 742
2 78299 1 742
2 78300 1 742
2 78301 1 742
2 78302 1 743
2 78303 1 743
2 78304 1 745
2 78305 1 745
2 78306 1 745
2 78307 1 745
2 78308 1 745
2 78309 1 745
2 78310 1 745
2 78311 1 745
2 78312 1 745
2 78313 1 745
2 78314 1 745
2 78315 1 745
2 78316 1 745
2 78317 1 745
2 78318 1 745
2 78319 1 745
2 78320 1 745
2 78321 1 745
2 78322 1 745
2 78323 1 745
2 78324 1 745
2 78325 1 745
2 78326 1 745
2 78327 1 746
2 78328 1 746
2 78329 1 746
2 78330 1 746
2 78331 1 746
2 78332 1 747
2 78333 1 747
2 78334 1 747
2 78335 1 747
2 78336 1 747
2 78337 1 748
2 78338 1 748
2 78339 1 748
2 78340 1 748
2 78341 1 748
2 78342 1 748
2 78343 1 748
2 78344 1 748
2 78345 1 748
2 78346 1 748
2 78347 1 748
2 78348 1 748
2 78349 1 748
2 78350 1 748
2 78351 1 748
2 78352 1 748
2 78353 1 748
2 78354 1 749
2 78355 1 749
2 78356 1 749
2 78357 1 749
2 78358 1 750
2 78359 1 750
2 78360 1 750
2 78361 1 750
2 78362 1 750
2 78363 1 750
2 78364 1 750
2 78365 1 750
2 78366 1 750
2 78367 1 750
2 78368 1 750
2 78369 1 759
2 78370 1 759
2 78371 1 759
2 78372 1 759
2 78373 1 759
2 78374 1 759
2 78375 1 759
2 78376 1 759
2 78377 1 759
2 78378 1 759
2 78379 1 759
2 78380 1 759
2 78381 1 759
2 78382 1 759
2 78383 1 759
2 78384 1 759
2 78385 1 759
2 78386 1 759
2 78387 1 759
2 78388 1 760
2 78389 1 760
2 78390 1 760
2 78391 1 761
2 78392 1 761
2 78393 1 761
2 78394 1 761
2 78395 1 761
2 78396 1 761
2 78397 1 761
2 78398 1 764
2 78399 1 764
2 78400 1 764
2 78401 1 764
2 78402 1 764
2 78403 1 764
2 78404 1 764
2 78405 1 764
2 78406 1 764
2 78407 1 764
2 78408 1 764
2 78409 1 764
2 78410 1 764
2 78411 1 764
2 78412 1 764
2 78413 1 764
2 78414 1 764
2 78415 1 764
2 78416 1 764
2 78417 1 764
2 78418 1 764
2 78419 1 764
2 78420 1 764
2 78421 1 765
2 78422 1 765
2 78423 1 765
2 78424 1 766
2 78425 1 766
2 78426 1 766
2 78427 1 766
2 78428 1 766
2 78429 1 766
2 78430 1 766
2 78431 1 766
2 78432 1 766
2 78433 1 766
2 78434 1 766
2 78435 1 766
2 78436 1 766
2 78437 1 766
2 78438 1 766
2 78439 1 766
2 78440 1 766
2 78441 1 766
2 78442 1 767
2 78443 1 767
2 78444 1 767
2 78445 1 767
2 78446 1 767
2 78447 1 767
2 78448 1 767
2 78449 1 767
2 78450 1 767
2 78451 1 768
2 78452 1 768
2 78453 1 768
2 78454 1 769
2 78455 1 769
2 78456 1 769
2 78457 1 769
2 78458 1 769
2 78459 1 769
2 78460 1 769
2 78461 1 769
2 78462 1 769
2 78463 1 769
2 78464 1 770
2 78465 1 770
2 78466 1 771
2 78467 1 771
2 78468 1 772
2 78469 1 772
2 78470 1 772
2 78471 1 772
2 78472 1 772
2 78473 1 772
2 78474 1 772
2 78475 1 772
2 78476 1 772
2 78477 1 772
2 78478 1 772
2 78479 1 772
2 78480 1 772
2 78481 1 772
2 78482 1 772
2 78483 1 772
2 78484 1 772
2 78485 1 772
2 78486 1 772
2 78487 1 772
2 78488 1 772
2 78489 1 772
2 78490 1 772
2 78491 1 772
2 78492 1 772
2 78493 1 772
2 78494 1 773
2 78495 1 773
2 78496 1 773
2 78497 1 773
2 78498 1 773
2 78499 1 774
2 78500 1 774
2 78501 1 774
2 78502 1 775
2 78503 1 775
2 78504 1 777
2 78505 1 777
2 78506 1 777
2 78507 1 777
2 78508 1 777
2 78509 1 777
2 78510 1 777
2 78511 1 777
2 78512 1 777
2 78513 1 777
2 78514 1 777
2 78515 1 777
2 78516 1 777
2 78517 1 777
2 78518 1 777
2 78519 1 777
2 78520 1 777
2 78521 1 777
2 78522 1 777
2 78523 1 777
2 78524 1 778
2 78525 1 778
2 78526 1 784
2 78527 1 784
2 78528 1 784
2 78529 1 784
2 78530 1 789
2 78531 1 789
2 78532 1 792
2 78533 1 792
2 78534 1 792
2 78535 1 792
2 78536 1 792
2 78537 1 792
2 78538 1 792
2 78539 1 792
2 78540 1 792
2 78541 1 792
2 78542 1 792
2 78543 1 792
2 78544 1 793
2 78545 1 793
2 78546 1 793
2 78547 1 793
2 78548 1 793
2 78549 1 793
2 78550 1 793
2 78551 1 793
2 78552 1 793
2 78553 1 793
2 78554 1 793
2 78555 1 793
2 78556 1 793
2 78557 1 793
2 78558 1 793
2 78559 1 794
2 78560 1 794
2 78561 1 796
2 78562 1 796
2 78563 1 796
2 78564 1 796
2 78565 1 796
2 78566 1 796
2 78567 1 796
2 78568 1 796
2 78569 1 796
2 78570 1 796
2 78571 1 796
2 78572 1 796
2 78573 1 796
2 78574 1 796
2 78575 1 796
2 78576 1 796
2 78577 1 796
2 78578 1 796
2 78579 1 796
2 78580 1 796
2 78581 1 796
2 78582 1 796
2 78583 1 796
2 78584 1 796
2 78585 1 796
2 78586 1 797
2 78587 1 797
2 78588 1 797
2 78589 1 797
2 78590 1 797
2 78591 1 797
2 78592 1 797
2 78593 1 797
2 78594 1 797
2 78595 1 797
2 78596 1 797
2 78597 1 797
2 78598 1 797
2 78599 1 797
2 78600 1 798
2 78601 1 798
2 78602 1 798
2 78603 1 805
2 78604 1 805
2 78605 1 815
2 78606 1 815
2 78607 1 815
2 78608 1 815
2 78609 1 815
2 78610 1 815
2 78611 1 815
2 78612 1 815
2 78613 1 815
2 78614 1 815
2 78615 1 815
2 78616 1 815
2 78617 1 815
2 78618 1 815
2 78619 1 815
2 78620 1 815
2 78621 1 815
2 78622 1 815
2 78623 1 815
2 78624 1 815
2 78625 1 815
2 78626 1 815
2 78627 1 815
2 78628 1 815
2 78629 1 815
2 78630 1 815
2 78631 1 815
2 78632 1 815
2 78633 1 815
2 78634 1 815
2 78635 1 815
2 78636 1 815
2 78637 1 815
2 78638 1 815
2 78639 1 815
2 78640 1 815
2 78641 1 815
2 78642 1 815
2 78643 1 815
2 78644 1 815
2 78645 1 815
2 78646 1 815
2 78647 1 815
2 78648 1 815
2 78649 1 815
2 78650 1 815
2 78651 1 815
2 78652 1 815
2 78653 1 815
2 78654 1 815
2 78655 1 815
2 78656 1 815
2 78657 1 815
2 78658 1 815
2 78659 1 815
2 78660 1 815
2 78661 1 815
2 78662 1 815
2 78663 1 815
2 78664 1 815
2 78665 1 815
2 78666 1 815
2 78667 1 815
2 78668 1 815
2 78669 1 815
2 78670 1 815
2 78671 1 816
2 78672 1 816
2 78673 1 816
2 78674 1 816
2 78675 1 816
2 78676 1 816
2 78677 1 816
2 78678 1 816
2 78679 1 816
2 78680 1 816
2 78681 1 816
2 78682 1 816
2 78683 1 816
2 78684 1 816
2 78685 1 816
2 78686 1 816
2 78687 1 816
2 78688 1 816
2 78689 1 816
2 78690 1 816
2 78691 1 816
2 78692 1 816
2 78693 1 816
2 78694 1 816
2 78695 1 816
2 78696 1 816
2 78697 1 816
2 78698 1 816
2 78699 1 816
2 78700 1 816
2 78701 1 816
2 78702 1 816
2 78703 1 816
2 78704 1 816
2 78705 1 816
2 78706 1 816
2 78707 1 816
2 78708 1 816
2 78709 1 816
2 78710 1 816
2 78711 1 816
2 78712 1 816
2 78713 1 816
2 78714 1 819
2 78715 1 819
2 78716 1 824
2 78717 1 824
2 78718 1 824
2 78719 1 824
2 78720 1 824
2 78721 1 824
2 78722 1 824
2 78723 1 824
2 78724 1 824
2 78725 1 824
2 78726 1 824
2 78727 1 824
2 78728 1 824
2 78729 1 824
2 78730 1 824
2 78731 1 824
2 78732 1 832
2 78733 1 832
2 78734 1 833
2 78735 1 833
2 78736 1 833
2 78737 1 833
2 78738 1 833
2 78739 1 833
2 78740 1 833
2 78741 1 833
2 78742 1 833
2 78743 1 833
2 78744 1 833
2 78745 1 833
2 78746 1 833
2 78747 1 833
2 78748 1 833
2 78749 1 833
2 78750 1 833
2 78751 1 834
2 78752 1 834
2 78753 1 834
2 78754 1 834
2 78755 1 835
2 78756 1 835
2 78757 1 835
2 78758 1 836
2 78759 1 836
2 78760 1 836
2 78761 1 836
2 78762 1 836
2 78763 1 836
2 78764 1 836
2 78765 1 837
2 78766 1 837
2 78767 1 838
2 78768 1 838
2 78769 1 838
2 78770 1 845
2 78771 1 845
2 78772 1 848
2 78773 1 848
2 78774 1 848
2 78775 1 848
2 78776 1 848
2 78777 1 850
2 78778 1 850
2 78779 1 852
2 78780 1 852
2 78781 1 858
2 78782 1 858
2 78783 1 858
2 78784 1 858
2 78785 1 858
2 78786 1 858
2 78787 1 859
2 78788 1 859
2 78789 1 859
2 78790 1 859
2 78791 1 861
2 78792 1 861
2 78793 1 861
2 78794 1 861
2 78795 1 861
2 78796 1 861
2 78797 1 861
2 78798 1 861
2 78799 1 861
2 78800 1 861
2 78801 1 861
2 78802 1 861
2 78803 1 861
2 78804 1 861
2 78805 1 861
2 78806 1 861
2 78807 1 861
2 78808 1 861
2 78809 1 861
2 78810 1 861
2 78811 1 863
2 78812 1 863
2 78813 1 864
2 78814 1 864
2 78815 1 879
2 78816 1 879
2 78817 1 879
2 78818 1 879
2 78819 1 879
2 78820 1 879
2 78821 1 879
2 78822 1 879
2 78823 1 880
2 78824 1 880
2 78825 1 880
2 78826 1 880
2 78827 1 880
2 78828 1 880
2 78829 1 881
2 78830 1 881
2 78831 1 881
2 78832 1 881
2 78833 1 881
2 78834 1 881
2 78835 1 881
2 78836 1 881
2 78837 1 881
2 78838 1 882
2 78839 1 882
2 78840 1 884
2 78841 1 884
2 78842 1 885
2 78843 1 885
2 78844 1 885
2 78845 1 885
2 78846 1 885
2 78847 1 885
2 78848 1 897
2 78849 1 897
2 78850 1 897
2 78851 1 897
2 78852 1 897
2 78853 1 897
2 78854 1 897
2 78855 1 897
2 78856 1 897
2 78857 1 897
2 78858 1 897
2 78859 1 897
2 78860 1 897
2 78861 1 897
2 78862 1 897
2 78863 1 897
2 78864 1 897
2 78865 1 897
2 78866 1 897
2 78867 1 897
2 78868 1 897
2 78869 1 897
2 78870 1 897
2 78871 1 897
2 78872 1 897
2 78873 1 897
2 78874 1 897
2 78875 1 897
2 78876 1 897
2 78877 1 897
2 78878 1 897
2 78879 1 897
2 78880 1 897
2 78881 1 897
2 78882 1 897
2 78883 1 897
2 78884 1 897
2 78885 1 897
2 78886 1 897
2 78887 1 897
2 78888 1 897
2 78889 1 897
2 78890 1 899
2 78891 1 899
2 78892 1 899
2 78893 1 899
2 78894 1 899
2 78895 1 899
2 78896 1 899
2 78897 1 899
2 78898 1 899
2 78899 1 899
2 78900 1 901
2 78901 1 901
2 78902 1 901
2 78903 1 901
2 78904 1 901
2 78905 1 901
2 78906 1 901
2 78907 1 901
2 78908 1 902
2 78909 1 902
2 78910 1 904
2 78911 1 904
2 78912 1 904
2 78913 1 904
2 78914 1 904
2 78915 1 904
2 78916 1 905
2 78917 1 905
2 78918 1 907
2 78919 1 907
2 78920 1 907
2 78921 1 907
2 78922 1 907
2 78923 1 907
2 78924 1 907
2 78925 1 907
2 78926 1 909
2 78927 1 909
2 78928 1 909
2 78929 1 909
2 78930 1 909
2 78931 1 910
2 78932 1 910
2 78933 1 910
2 78934 1 910
2 78935 1 910
2 78936 1 910
2 78937 1 910
2 78938 1 910
2 78939 1 910
2 78940 1 912
2 78941 1 912
2 78942 1 913
2 78943 1 913
2 78944 1 915
2 78945 1 915
2 78946 1 921
2 78947 1 921
2 78948 1 921
2 78949 1 921
2 78950 1 921
2 78951 1 921
2 78952 1 921
2 78953 1 921
2 78954 1 921
2 78955 1 921
2 78956 1 921
2 78957 1 922
2 78958 1 922
2 78959 1 922
2 78960 1 922
2 78961 1 923
2 78962 1 923
2 78963 1 924
2 78964 1 924
2 78965 1 928
2 78966 1 928
2 78967 1 932
2 78968 1 932
2 78969 1 934
2 78970 1 934
2 78971 1 934
2 78972 1 935
2 78973 1 935
2 78974 1 951
2 78975 1 951
2 78976 1 951
2 78977 1 951
2 78978 1 951
2 78979 1 951
2 78980 1 951
2 78981 1 951
2 78982 1 951
2 78983 1 951
2 78984 1 951
2 78985 1 951
2 78986 1 951
2 78987 1 951
2 78988 1 951
2 78989 1 951
2 78990 1 951
2 78991 1 951
2 78992 1 951
2 78993 1 951
2 78994 1 951
2 78995 1 951
2 78996 1 951
2 78997 1 951
2 78998 1 951
2 78999 1 951
2 79000 1 951
2 79001 1 951
2 79002 1 951
2 79003 1 952
2 79004 1 952
2 79005 1 952
2 79006 1 952
2 79007 1 953
2 79008 1 953
2 79009 1 953
2 79010 1 953
2 79011 1 953
2 79012 1 954
2 79013 1 954
2 79014 1 954
2 79015 1 954
2 79016 1 955
2 79017 1 955
2 79018 1 959
2 79019 1 959
2 79020 1 959
2 79021 1 959
2 79022 1 959
2 79023 1 959
2 79024 1 959
2 79025 1 959
2 79026 1 959
2 79027 1 959
2 79028 1 959
2 79029 1 959
2 79030 1 959
2 79031 1 959
2 79032 1 959
2 79033 1 959
2 79034 1 959
2 79035 1 959
2 79036 1 959
2 79037 1 959
2 79038 1 959
2 79039 1 960
2 79040 1 960
2 79041 1 961
2 79042 1 961
2 79043 1 961
2 79044 1 961
2 79045 1 961
2 79046 1 962
2 79047 1 962
2 79048 1 962
2 79049 1 962
2 79050 1 962
2 79051 1 962
2 79052 1 962
2 79053 1 962
2 79054 1 962
2 79055 1 962
2 79056 1 962
2 79057 1 962
2 79058 1 970
2 79059 1 970
2 79060 1 970
2 79061 1 970
2 79062 1 970
2 79063 1 970
2 79064 1 970
2 79065 1 970
2 79066 1 970
2 79067 1 970
2 79068 1 970
2 79069 1 970
2 79070 1 970
2 79071 1 970
2 79072 1 970
2 79073 1 970
2 79074 1 971
2 79075 1 971
2 79076 1 974
2 79077 1 974
2 79078 1 974
2 79079 1 975
2 79080 1 975
2 79081 1 975
2 79082 1 975
2 79083 1 975
2 79084 1 975
2 79085 1 975
2 79086 1 975
2 79087 1 975
2 79088 1 975
2 79089 1 975
2 79090 1 975
2 79091 1 975
2 79092 1 975
2 79093 1 975
2 79094 1 975
2 79095 1 987
2 79096 1 987
2 79097 1 989
2 79098 1 989
2 79099 1 989
2 79100 1 989
2 79101 1 989
2 79102 1 989
2 79103 1 989
2 79104 1 989
2 79105 1 989
2 79106 1 989
2 79107 1 989
2 79108 1 989
2 79109 1 989
2 79110 1 989
2 79111 1 989
2 79112 1 989
2 79113 1 989
2 79114 1 989
2 79115 1 989
2 79116 1 989
2 79117 1 989
2 79118 1 990
2 79119 1 990
2 79120 1 990
2 79121 1 990
2 79122 1 990
2 79123 1 990
2 79124 1 990
2 79125 1 990
2 79126 1 998
2 79127 1 998
2 79128 1 998
2 79129 1 998
2 79130 1 998
2 79131 1 998
2 79132 1 998
2 79133 1 998
2 79134 1 998
2 79135 1 998
2 79136 1 998
2 79137 1 998
2 79138 1 998
2 79139 1 998
2 79140 1 998
2 79141 1 998
2 79142 1 998
2 79143 1 998
2 79144 1 998
2 79145 1 998
2 79146 1 998
2 79147 1 998
2 79148 1 998
2 79149 1 998
2 79150 1 998
2 79151 1 998
2 79152 1 998
2 79153 1 998
2 79154 1 998
2 79155 1 998
2 79156 1 998
2 79157 1 998
2 79158 1 999
2 79159 1 999
2 79160 1 999
2 79161 1 999
2 79162 1 1004
2 79163 1 1004
2 79164 1 1004
2 79165 1 1004
2 79166 1 1004
2 79167 1 1004
2 79168 1 1004
2 79169 1 1004
2 79170 1 1004
2 79171 1 1004
2 79172 1 1006
2 79173 1 1006
2 79174 1 1006
2 79175 1 1006
2 79176 1 1006
2 79177 1 1007
2 79178 1 1007
2 79179 1 1007
2 79180 1 1007
2 79181 1 1007
2 79182 1 1008
2 79183 1 1008
2 79184 1 1008
2 79185 1 1008
2 79186 1 1008
2 79187 1 1008
2 79188 1 1009
2 79189 1 1009
2 79190 1 1009
2 79191 1 1009
2 79192 1 1013
2 79193 1 1013
2 79194 1 1013
2 79195 1 1013
2 79196 1 1013
2 79197 1 1013
2 79198 1 1013
2 79199 1 1013
2 79200 1 1013
2 79201 1 1013
2 79202 1 1013
2 79203 1 1014
2 79204 1 1014
2 79205 1 1017
2 79206 1 1017
2 79207 1 1017
2 79208 1 1017
2 79209 1 1017
2 79210 1 1017
2 79211 1 1017
2 79212 1 1017
2 79213 1 1017
2 79214 1 1018
2 79215 1 1018
2 79216 1 1018
2 79217 1 1018
2 79218 1 1019
2 79219 1 1019
2 79220 1 1019
2 79221 1 1019
2 79222 1 1019
2 79223 1 1019
2 79224 1 1019
2 79225 1 1019
2 79226 1 1019
2 79227 1 1019
2 79228 1 1019
2 79229 1 1019
2 79230 1 1019
2 79231 1 1019
2 79232 1 1019
2 79233 1 1019
2 79234 1 1019
2 79235 1 1019
2 79236 1 1020
2 79237 1 1020
2 79238 1 1020
2 79239 1 1022
2 79240 1 1022
2 79241 1 1022
2 79242 1 1022
2 79243 1 1022
2 79244 1 1023
2 79245 1 1023
2 79246 1 1023
2 79247 1 1023
2 79248 1 1023
2 79249 1 1023
2 79250 1 1023
2 79251 1 1023
2 79252 1 1024
2 79253 1 1024
2 79254 1 1024
2 79255 1 1025
2 79256 1 1025
2 79257 1 1025
2 79258 1 1025
2 79259 1 1025
2 79260 1 1025
2 79261 1 1025
2 79262 1 1025
2 79263 1 1025
2 79264 1 1026
2 79265 1 1026
2 79266 1 1035
2 79267 1 1035
2 79268 1 1035
2 79269 1 1035
2 79270 1 1035
2 79271 1 1035
2 79272 1 1035
2 79273 1 1035
2 79274 1 1035
2 79275 1 1035
2 79276 1 1035
2 79277 1 1035
2 79278 1 1035
2 79279 1 1035
2 79280 1 1035
2 79281 1 1035
2 79282 1 1035
2 79283 1 1035
2 79284 1 1035
2 79285 1 1035
2 79286 1 1035
2 79287 1 1035
2 79288 1 1035
2 79289 1 1035
2 79290 1 1035
2 79291 1 1035
2 79292 1 1035
2 79293 1 1036
2 79294 1 1036
2 79295 1 1037
2 79296 1 1037
2 79297 1 1037
2 79298 1 1037
2 79299 1 1037
2 79300 1 1038
2 79301 1 1038
2 79302 1 1038
2 79303 1 1039
2 79304 1 1039
2 79305 1 1039
2 79306 1 1040
2 79307 1 1040
2 79308 1 1040
2 79309 1 1043
2 79310 1 1043
2 79311 1 1043
2 79312 1 1043
2 79313 1 1043
2 79314 1 1043
2 79315 1 1043
2 79316 1 1044
2 79317 1 1044
2 79318 1 1046
2 79319 1 1046
2 79320 1 1054
2 79321 1 1054
2 79322 1 1054
2 79323 1 1054
2 79324 1 1054
2 79325 1 1054
2 79326 1 1054
2 79327 1 1054
2 79328 1 1054
2 79329 1 1054
2 79330 1 1054
2 79331 1 1055
2 79332 1 1055
2 79333 1 1055
2 79334 1 1055
2 79335 1 1057
2 79336 1 1057
2 79337 1 1057
2 79338 1 1057
2 79339 1 1057
2 79340 1 1057
2 79341 1 1058
2 79342 1 1058
2 79343 1 1058
2 79344 1 1058
2 79345 1 1058
2 79346 1 1070
2 79347 1 1070
2 79348 1 1070
2 79349 1 1070
2 79350 1 1070
2 79351 1 1070
2 79352 1 1070
2 79353 1 1070
2 79354 1 1070
2 79355 1 1070
2 79356 1 1070
2 79357 1 1071
2 79358 1 1071
2 79359 1 1071
2 79360 1 1071
2 79361 1 1071
2 79362 1 1071
2 79363 1 1071
2 79364 1 1071
2 79365 1 1071
2 79366 1 1071
2 79367 1 1071
2 79368 1 1071
2 79369 1 1071
2 79370 1 1071
2 79371 1 1071
2 79372 1 1071
2 79373 1 1071
2 79374 1 1071
2 79375 1 1071
2 79376 1 1071
2 79377 1 1071
2 79378 1 1071
2 79379 1 1071
2 79380 1 1071
2 79381 1 1071
2 79382 1 1071
2 79383 1 1071
2 79384 1 1071
2 79385 1 1071
2 79386 1 1072
2 79387 1 1072
2 79388 1 1072
2 79389 1 1072
2 79390 1 1072
2 79391 1 1072
2 79392 1 1072
2 79393 1 1072
2 79394 1 1072
2 79395 1 1073
2 79396 1 1073
2 79397 1 1073
2 79398 1 1073
2 79399 1 1073
2 79400 1 1073
2 79401 1 1073
2 79402 1 1073
2 79403 1 1074
2 79404 1 1074
2 79405 1 1074
2 79406 1 1075
2 79407 1 1075
2 79408 1 1075
2 79409 1 1075
2 79410 1 1075
2 79411 1 1075
2 79412 1 1075
2 79413 1 1075
2 79414 1 1075
2 79415 1 1075
2 79416 1 1075
2 79417 1 1075
2 79418 1 1075
2 79419 1 1076
2 79420 1 1076
2 79421 1 1076
2 79422 1 1076
2 79423 1 1076
2 79424 1 1076
2 79425 1 1076
2 79426 1 1076
2 79427 1 1077
2 79428 1 1077
2 79429 1 1078
2 79430 1 1078
2 79431 1 1078
2 79432 1 1078
2 79433 1 1078
2 79434 1 1078
2 79435 1 1080
2 79436 1 1080
2 79437 1 1087
2 79438 1 1087
2 79439 1 1089
2 79440 1 1089
2 79441 1 1090
2 79442 1 1090
2 79443 1 1100
2 79444 1 1100
2 79445 1 1100
2 79446 1 1100
2 79447 1 1100
2 79448 1 1100
2 79449 1 1100
2 79450 1 1100
2 79451 1 1100
2 79452 1 1100
2 79453 1 1101
2 79454 1 1101
2 79455 1 1101
2 79456 1 1101
2 79457 1 1101
2 79458 1 1103
2 79459 1 1103
2 79460 1 1103
2 79461 1 1103
2 79462 1 1103
2 79463 1 1103
2 79464 1 1103
2 79465 1 1103
2 79466 1 1103
2 79467 1 1103
2 79468 1 1103
2 79469 1 1103
2 79470 1 1103
2 79471 1 1103
2 79472 1 1103
2 79473 1 1103
2 79474 1 1103
2 79475 1 1103
2 79476 1 1103
2 79477 1 1103
2 79478 1 1103
2 79479 1 1103
2 79480 1 1103
2 79481 1 1103
2 79482 1 1103
2 79483 1 1104
2 79484 1 1104
2 79485 1 1105
2 79486 1 1105
2 79487 1 1105
2 79488 1 1105
2 79489 1 1118
2 79490 1 1118
2 79491 1 1119
2 79492 1 1119
2 79493 1 1122
2 79494 1 1122
2 79495 1 1122
2 79496 1 1123
2 79497 1 1123
2 79498 1 1123
2 79499 1 1123
2 79500 1 1123
2 79501 1 1123
2 79502 1 1123
2 79503 1 1123
2 79504 1 1123
2 79505 1 1123
2 79506 1 1123
2 79507 1 1123
2 79508 1 1123
2 79509 1 1123
2 79510 1 1123
2 79511 1 1123
2 79512 1 1123
2 79513 1 1124
2 79514 1 1124
2 79515 1 1124
2 79516 1 1124
2 79517 1 1124
2 79518 1 1124
2 79519 1 1124
2 79520 1 1124
2 79521 1 1124
2 79522 1 1124
2 79523 1 1125
2 79524 1 1125
2 79525 1 1125
2 79526 1 1125
2 79527 1 1137
2 79528 1 1137
2 79529 1 1137
2 79530 1 1138
2 79531 1 1138
2 79532 1 1138
2 79533 1 1148
2 79534 1 1148
2 79535 1 1148
2 79536 1 1149
2 79537 1 1149
2 79538 1 1149
2 79539 1 1149
2 79540 1 1150
2 79541 1 1150
2 79542 1 1151
2 79543 1 1151
2 79544 1 1151
2 79545 1 1151
2 79546 1 1151
2 79547 1 1152
2 79548 1 1152
2 79549 1 1153
2 79550 1 1153
2 79551 1 1154
2 79552 1 1154
2 79553 1 1154
2 79554 1 1154
2 79555 1 1154
2 79556 1 1154
2 79557 1 1154
2 79558 1 1154
2 79559 1 1154
2 79560 1 1154
2 79561 1 1154
2 79562 1 1154
2 79563 1 1155
2 79564 1 1155
2 79565 1 1156
2 79566 1 1156
2 79567 1 1156
2 79568 1 1156
2 79569 1 1156
2 79570 1 1156
2 79571 1 1156
2 79572 1 1156
2 79573 1 1156
2 79574 1 1156
2 79575 1 1156
2 79576 1 1156
2 79577 1 1156
2 79578 1 1156
2 79579 1 1156
2 79580 1 1156
2 79581 1 1156
2 79582 1 1156
2 79583 1 1156
2 79584 1 1158
2 79585 1 1158
2 79586 1 1159
2 79587 1 1159
2 79588 1 1159
2 79589 1 1161
2 79590 1 1161
2 79591 1 1161
2 79592 1 1166
2 79593 1 1166
2 79594 1 1166
2 79595 1 1166
2 79596 1 1166
2 79597 1 1166
2 79598 1 1166
2 79599 1 1167
2 79600 1 1167
2 79601 1 1167
2 79602 1 1167
2 79603 1 1167
2 79604 1 1168
2 79605 1 1168
2 79606 1 1168
2 79607 1 1176
2 79608 1 1176
2 79609 1 1176
2 79610 1 1177
2 79611 1 1177
2 79612 1 1178
2 79613 1 1178
2 79614 1 1178
2 79615 1 1178
2 79616 1 1178
2 79617 1 1178
2 79618 1 1179
2 79619 1 1179
2 79620 1 1179
2 79621 1 1179
2 79622 1 1187
2 79623 1 1187
2 79624 1 1187
2 79625 1 1187
2 79626 1 1187
2 79627 1 1187
2 79628 1 1187
2 79629 1 1187
2 79630 1 1187
2 79631 1 1187
2 79632 1 1187
2 79633 1 1187
2 79634 1 1187
2 79635 1 1187
2 79636 1 1187
2 79637 1 1187
2 79638 1 1187
2 79639 1 1187
2 79640 1 1187
2 79641 1 1187
2 79642 1 1187
2 79643 1 1187
2 79644 1 1187
2 79645 1 1187
2 79646 1 1187
2 79647 1 1187
2 79648 1 1187
2 79649 1 1187
2 79650 1 1187
2 79651 1 1188
2 79652 1 1188
2 79653 1 1188
2 79654 1 1188
2 79655 1 1188
2 79656 1 1188
2 79657 1 1188
2 79658 1 1188
2 79659 1 1188
2 79660 1 1188
2 79661 1 1188
2 79662 1 1188
2 79663 1 1188
2 79664 1 1188
2 79665 1 1188
2 79666 1 1188
2 79667 1 1188
2 79668 1 1189
2 79669 1 1189
2 79670 1 1190
2 79671 1 1190
2 79672 1 1191
2 79673 1 1191
2 79674 1 1191
2 79675 1 1198
2 79676 1 1198
2 79677 1 1198
2 79678 1 1198
2 79679 1 1199
2 79680 1 1199
2 79681 1 1199
2 79682 1 1199
2 79683 1 1199
2 79684 1 1199
2 79685 1 1200
2 79686 1 1200
2 79687 1 1200
2 79688 1 1201
2 79689 1 1201
2 79690 1 1201
2 79691 1 1201
2 79692 1 1201
2 79693 1 1201
2 79694 1 1201
2 79695 1 1202
2 79696 1 1202
2 79697 1 1202
2 79698 1 1203
2 79699 1 1203
2 79700 1 1203
2 79701 1 1203
2 79702 1 1203
2 79703 1 1203
2 79704 1 1203
2 79705 1 1203
2 79706 1 1203
2 79707 1 1204
2 79708 1 1204
2 79709 1 1204
2 79710 1 1212
2 79711 1 1212
2 79712 1 1212
2 79713 1 1212
2 79714 1 1212
2 79715 1 1212
2 79716 1 1212
2 79717 1 1212
2 79718 1 1212
2 79719 1 1212
2 79720 1 1212
2 79721 1 1212
2 79722 1 1212
2 79723 1 1212
2 79724 1 1212
2 79725 1 1212
2 79726 1 1212
2 79727 1 1212
2 79728 1 1212
2 79729 1 1212
2 79730 1 1212
2 79731 1 1212
2 79732 1 1212
2 79733 1 1212
2 79734 1 1212
2 79735 1 1212
2 79736 1 1212
2 79737 1 1212
2 79738 1 1212
2 79739 1 1212
2 79740 1 1212
2 79741 1 1212
2 79742 1 1212
2 79743 1 1212
2 79744 1 1213
2 79745 1 1213
2 79746 1 1214
2 79747 1 1214
2 79748 1 1215
2 79749 1 1215
2 79750 1 1215
2 79751 1 1221
2 79752 1 1221
2 79753 1 1221
2 79754 1 1221
2 79755 1 1221
2 79756 1 1222
2 79757 1 1222
2 79758 1 1222
2 79759 1 1222
2 79760 1 1222
2 79761 1 1222
2 79762 1 1222
2 79763 1 1222
2 79764 1 1222
2 79765 1 1222
2 79766 1 1222
2 79767 1 1222
2 79768 1 1222
2 79769 1 1222
2 79770 1 1222
2 79771 1 1222
2 79772 1 1222
2 79773 1 1222
2 79774 1 1222
2 79775 1 1222
2 79776 1 1222
2 79777 1 1227
2 79778 1 1227
2 79779 1 1228
2 79780 1 1228
2 79781 1 1228
2 79782 1 1228
2 79783 1 1228
2 79784 1 1228
2 79785 1 1228
2 79786 1 1228
2 79787 1 1228
2 79788 1 1230
2 79789 1 1230
2 79790 1 1230
2 79791 1 1230
2 79792 1 1230
2 79793 1 1230
2 79794 1 1230
2 79795 1 1230
2 79796 1 1230
2 79797 1 1243
2 79798 1 1243
2 79799 1 1243
2 79800 1 1243
2 79801 1 1243
2 79802 1 1243
2 79803 1 1243
2 79804 1 1243
2 79805 1 1243
2 79806 1 1243
2 79807 1 1243
2 79808 1 1243
2 79809 1 1243
2 79810 1 1243
2 79811 1 1243
2 79812 1 1243
2 79813 1 1243
2 79814 1 1243
2 79815 1 1243
2 79816 1 1244
2 79817 1 1244
2 79818 1 1244
2 79819 1 1244
2 79820 1 1244
2 79821 1 1244
2 79822 1 1244
2 79823 1 1245
2 79824 1 1245
2 79825 1 1245
2 79826 1 1245
2 79827 1 1245
2 79828 1 1245
2 79829 1 1245
2 79830 1 1245
2 79831 1 1246
2 79832 1 1246
2 79833 1 1246
2 79834 1 1246
2 79835 1 1246
2 79836 1 1246
2 79837 1 1246
2 79838 1 1246
2 79839 1 1246
2 79840 1 1246
2 79841 1 1246
2 79842 1 1246
2 79843 1 1246
2 79844 1 1246
2 79845 1 1246
2 79846 1 1246
2 79847 1 1246
2 79848 1 1246
2 79849 1 1246
2 79850 1 1246
2 79851 1 1246
2 79852 1 1246
2 79853 1 1246
2 79854 1 1246
2 79855 1 1246
2 79856 1 1246
2 79857 1 1246
2 79858 1 1246
2 79859 1 1246
2 79860 1 1247
2 79861 1 1247
2 79862 1 1247
2 79863 1 1247
2 79864 1 1248
2 79865 1 1248
2 79866 1 1250
2 79867 1 1250
2 79868 1 1250
2 79869 1 1259
2 79870 1 1259
2 79871 1 1259
2 79872 1 1260
2 79873 1 1260
2 79874 1 1260
2 79875 1 1261
2 79876 1 1261
2 79877 1 1262
2 79878 1 1262
2 79879 1 1264
2 79880 1 1264
2 79881 1 1264
2 79882 1 1264
2 79883 1 1267
2 79884 1 1267
2 79885 1 1267
2 79886 1 1267
2 79887 1 1268
2 79888 1 1268
2 79889 1 1268
2 79890 1 1268
2 79891 1 1271
2 79892 1 1271
2 79893 1 1271
2 79894 1 1271
2 79895 1 1272
2 79896 1 1272
2 79897 1 1280
2 79898 1 1280
2 79899 1 1280
2 79900 1 1280
2 79901 1 1280
2 79902 1 1280
2 79903 1 1281
2 79904 1 1281
2 79905 1 1281
2 79906 1 1281
2 79907 1 1281
2 79908 1 1281
2 79909 1 1281
2 79910 1 1281
2 79911 1 1281
2 79912 1 1281
2 79913 1 1281
2 79914 1 1282
2 79915 1 1282
2 79916 1 1284
2 79917 1 1284
2 79918 1 1284
2 79919 1 1284
2 79920 1 1288
2 79921 1 1288
2 79922 1 1288
2 79923 1 1288
2 79924 1 1288
2 79925 1 1288
2 79926 1 1288
2 79927 1 1288
2 79928 1 1289
2 79929 1 1289
2 79930 1 1289
2 79931 1 1289
2 79932 1 1290
2 79933 1 1290
2 79934 1 1305
2 79935 1 1305
2 79936 1 1305
2 79937 1 1305
2 79938 1 1305
2 79939 1 1306
2 79940 1 1306
2 79941 1 1306
2 79942 1 1307
2 79943 1 1307
2 79944 1 1307
2 79945 1 1307
2 79946 1 1307
2 79947 1 1307
2 79948 1 1307
2 79949 1 1308
2 79950 1 1308
2 79951 1 1308
2 79952 1 1308
2 79953 1 1308
2 79954 1 1308
2 79955 1 1308
2 79956 1 1308
2 79957 1 1308
2 79958 1 1308
2 79959 1 1308
2 79960 1 1308
2 79961 1 1308
2 79962 1 1308
2 79963 1 1308
2 79964 1 1308
2 79965 1 1308
2 79966 1 1308
2 79967 1 1308
2 79968 1 1308
2 79969 1 1308
2 79970 1 1308
2 79971 1 1308
2 79972 1 1308
2 79973 1 1308
2 79974 1 1316
2 79975 1 1316
2 79976 1 1319
2 79977 1 1319
2 79978 1 1319
2 79979 1 1319
2 79980 1 1319
2 79981 1 1319
2 79982 1 1319
2 79983 1 1319
2 79984 1 1319
2 79985 1 1319
2 79986 1 1328
2 79987 1 1328
2 79988 1 1328
2 79989 1 1328
2 79990 1 1328
2 79991 1 1329
2 79992 1 1329
2 79993 1 1329
2 79994 1 1329
2 79995 1 1329
2 79996 1 1329
2 79997 1 1330
2 79998 1 1330
2 79999 1 1330
2 80000 1 1330
2 80001 1 1330
2 80002 1 1331
2 80003 1 1331
2 80004 1 1334
2 80005 1 1334
2 80006 1 1335
2 80007 1 1335
2 80008 1 1335
2 80009 1 1335
2 80010 1 1335
2 80011 1 1335
2 80012 1 1335
2 80013 1 1335
2 80014 1 1335
2 80015 1 1335
2 80016 1 1335
2 80017 1 1335
2 80018 1 1335
2 80019 1 1335
2 80020 1 1335
2 80021 1 1335
2 80022 1 1335
2 80023 1 1335
2 80024 1 1335
2 80025 1 1335
2 80026 1 1335
2 80027 1 1335
2 80028 1 1335
2 80029 1 1335
2 80030 1 1335
2 80031 1 1335
2 80032 1 1335
2 80033 1 1335
2 80034 1 1335
2 80035 1 1335
2 80036 1 1335
2 80037 1 1335
2 80038 1 1335
2 80039 1 1336
2 80040 1 1336
2 80041 1 1336
2 80042 1 1338
2 80043 1 1338
2 80044 1 1341
2 80045 1 1341
2 80046 1 1341
2 80047 1 1341
2 80048 1 1341
2 80049 1 1342
2 80050 1 1342
2 80051 1 1342
2 80052 1 1343
2 80053 1 1343
2 80054 1 1344
2 80055 1 1344
2 80056 1 1347
2 80057 1 1347
2 80058 1 1350
2 80059 1 1350
2 80060 1 1350
2 80061 1 1350
2 80062 1 1350
2 80063 1 1350
2 80064 1 1350
2 80065 1 1350
2 80066 1 1351
2 80067 1 1351
2 80068 1 1351
2 80069 1 1351
2 80070 1 1351
2 80071 1 1351
2 80072 1 1351
2 80073 1 1351
2 80074 1 1351
2 80075 1 1351
2 80076 1 1351
2 80077 1 1351
2 80078 1 1351
2 80079 1 1351
2 80080 1 1351
2 80081 1 1351
2 80082 1 1351
2 80083 1 1351
2 80084 1 1351
2 80085 1 1351
2 80086 1 1351
2 80087 1 1353
2 80088 1 1353
2 80089 1 1353
2 80090 1 1353
2 80091 1 1353
2 80092 1 1353
2 80093 1 1353
2 80094 1 1354
2 80095 1 1354
2 80096 1 1354
2 80097 1 1354
2 80098 1 1354
2 80099 1 1354
2 80100 1 1354
2 80101 1 1354
2 80102 1 1354
2 80103 1 1354
2 80104 1 1354
2 80105 1 1354
2 80106 1 1355
2 80107 1 1355
2 80108 1 1355
2 80109 1 1355
2 80110 1 1359
2 80111 1 1359
2 80112 1 1359
2 80113 1 1359
2 80114 1 1359
2 80115 1 1359
2 80116 1 1359
2 80117 1 1359
2 80118 1 1359
2 80119 1 1359
2 80120 1 1359
2 80121 1 1359
2 80122 1 1359
2 80123 1 1359
2 80124 1 1359
2 80125 1 1359
2 80126 1 1359
2 80127 1 1359
2 80128 1 1359
2 80129 1 1359
2 80130 1 1359
2 80131 1 1359
2 80132 1 1359
2 80133 1 1360
2 80134 1 1360
2 80135 1 1360
2 80136 1 1360
2 80137 1 1361
2 80138 1 1361
2 80139 1 1361
2 80140 1 1367
2 80141 1 1367
2 80142 1 1367
2 80143 1 1367
2 80144 1 1368
2 80145 1 1368
2 80146 1 1370
2 80147 1 1370
2 80148 1 1380
2 80149 1 1380
2 80150 1 1380
2 80151 1 1380
2 80152 1 1380
2 80153 1 1380
2 80154 1 1380
2 80155 1 1380
2 80156 1 1381
2 80157 1 1381
2 80158 1 1381
2 80159 1 1381
2 80160 1 1381
2 80161 1 1381
2 80162 1 1381
2 80163 1 1381
2 80164 1 1381
2 80165 1 1381
2 80166 1 1381
2 80167 1 1381
2 80168 1 1381
2 80169 1 1381
2 80170 1 1382
2 80171 1 1382
2 80172 1 1382
2 80173 1 1382
2 80174 1 1382
2 80175 1 1382
2 80176 1 1382
2 80177 1 1382
2 80178 1 1382
2 80179 1 1382
2 80180 1 1382
2 80181 1 1382
2 80182 1 1383
2 80183 1 1383
2 80184 1 1386
2 80185 1 1386
2 80186 1 1404
2 80187 1 1404
2 80188 1 1404
2 80189 1 1404
2 80190 1 1404
2 80191 1 1404
2 80192 1 1404
2 80193 1 1404
2 80194 1 1404
2 80195 1 1404
2 80196 1 1405
2 80197 1 1405
2 80198 1 1405
2 80199 1 1405
2 80200 1 1405
2 80201 1 1405
2 80202 1 1405
2 80203 1 1405
2 80204 1 1405
2 80205 1 1405
2 80206 1 1405
2 80207 1 1406
2 80208 1 1406
2 80209 1 1406
2 80210 1 1406
2 80211 1 1406
2 80212 1 1406
2 80213 1 1406
2 80214 1 1406
2 80215 1 1406
2 80216 1 1406
2 80217 1 1407
2 80218 1 1407
2 80219 1 1408
2 80220 1 1408
2 80221 1 1408
2 80222 1 1410
2 80223 1 1410
2 80224 1 1410
2 80225 1 1410
2 80226 1 1410
2 80227 1 1410
2 80228 1 1410
2 80229 1 1410
2 80230 1 1410
2 80231 1 1410
2 80232 1 1410
2 80233 1 1410
2 80234 1 1410
2 80235 1 1410
2 80236 1 1410
2 80237 1 1410
2 80238 1 1410
2 80239 1 1411
2 80240 1 1411
2 80241 1 1411
2 80242 1 1411
2 80243 1 1411
2 80244 1 1411
2 80245 1 1411
2 80246 1 1411
2 80247 1 1411
2 80248 1 1411
2 80249 1 1411
2 80250 1 1411
2 80251 1 1412
2 80252 1 1412
2 80253 1 1412
2 80254 1 1413
2 80255 1 1413
2 80256 1 1413
2 80257 1 1413
2 80258 1 1414
2 80259 1 1414
2 80260 1 1414
2 80261 1 1415
2 80262 1 1415
2 80263 1 1415
2 80264 1 1415
2 80265 1 1415
2 80266 1 1415
2 80267 1 1415
2 80268 1 1415
2 80269 1 1415
2 80270 1 1415
2 80271 1 1415
2 80272 1 1416
2 80273 1 1416
2 80274 1 1416
2 80275 1 1416
2 80276 1 1418
2 80277 1 1418
2 80278 1 1418
2 80279 1 1418
2 80280 1 1418
2 80281 1 1418
2 80282 1 1418
2 80283 1 1425
2 80284 1 1425
2 80285 1 1425
2 80286 1 1425
2 80287 1 1425
2 80288 1 1425
2 80289 1 1425
2 80290 1 1425
2 80291 1 1425
2 80292 1 1425
2 80293 1 1425
2 80294 1 1425
2 80295 1 1425
2 80296 1 1425
2 80297 1 1425
2 80298 1 1425
2 80299 1 1425
2 80300 1 1425
2 80301 1 1425
2 80302 1 1425
2 80303 1 1425
2 80304 1 1425
2 80305 1 1425
2 80306 1 1426
2 80307 1 1426
2 80308 1 1426
2 80309 1 1427
2 80310 1 1427
2 80311 1 1429
2 80312 1 1429
2 80313 1 1429
2 80314 1 1429
2 80315 1 1429
2 80316 1 1429
2 80317 1 1429
2 80318 1 1429
2 80319 1 1429
2 80320 1 1429
2 80321 1 1429
2 80322 1 1431
2 80323 1 1431
2 80324 1 1439
2 80325 1 1439
2 80326 1 1439
2 80327 1 1439
2 80328 1 1439
2 80329 1 1439
2 80330 1 1441
2 80331 1 1441
2 80332 1 1441
2 80333 1 1441
2 80334 1 1441
2 80335 1 1441
2 80336 1 1441
2 80337 1 1441
2 80338 1 1441
2 80339 1 1441
2 80340 1 1441
2 80341 1 1441
2 80342 1 1441
2 80343 1 1441
2 80344 1 1441
2 80345 1 1441
2 80346 1 1441
2 80347 1 1441
2 80348 1 1441
2 80349 1 1441
2 80350 1 1441
2 80351 1 1441
2 80352 1 1441
2 80353 1 1441
2 80354 1 1441
2 80355 1 1441
2 80356 1 1441
2 80357 1 1441
2 80358 1 1441
2 80359 1 1441
2 80360 1 1441
2 80361 1 1441
2 80362 1 1441
2 80363 1 1441
2 80364 1 1441
2 80365 1 1441
2 80366 1 1441
2 80367 1 1441
2 80368 1 1441
2 80369 1 1441
2 80370 1 1441
2 80371 1 1441
2 80372 1 1441
2 80373 1 1441
2 80374 1 1441
2 80375 1 1441
2 80376 1 1441
2 80377 1 1441
2 80378 1 1441
2 80379 1 1441
2 80380 1 1441
2 80381 1 1441
2 80382 1 1441
2 80383 1 1442
2 80384 1 1442
2 80385 1 1442
2 80386 1 1442
2 80387 1 1442
2 80388 1 1442
2 80389 1 1442
2 80390 1 1442
2 80391 1 1442
2 80392 1 1442
2 80393 1 1442
2 80394 1 1442
2 80395 1 1442
2 80396 1 1442
2 80397 1 1442
2 80398 1 1442
2 80399 1 1442
2 80400 1 1442
2 80401 1 1442
2 80402 1 1442
2 80403 1 1442
2 80404 1 1442
2 80405 1 1442
2 80406 1 1442
2 80407 1 1442
2 80408 1 1442
2 80409 1 1442
2 80410 1 1442
2 80411 1 1442
2 80412 1 1442
2 80413 1 1442
2 80414 1 1442
2 80415 1 1442
2 80416 1 1442
2 80417 1 1442
2 80418 1 1442
2 80419 1 1442
2 80420 1 1442
2 80421 1 1442
2 80422 1 1442
2 80423 1 1442
2 80424 1 1442
2 80425 1 1442
2 80426 1 1442
2 80427 1 1442
2 80428 1 1442
2 80429 1 1442
2 80430 1 1442
2 80431 1 1442
2 80432 1 1442
2 80433 1 1442
2 80434 1 1443
2 80435 1 1443
2 80436 1 1443
2 80437 1 1443
2 80438 1 1443
2 80439 1 1444
2 80440 1 1444
2 80441 1 1444
2 80442 1 1444
2 80443 1 1444
2 80444 1 1444
2 80445 1 1444
2 80446 1 1444
2 80447 1 1444
2 80448 1 1445
2 80449 1 1445
2 80450 1 1446
2 80451 1 1446
2 80452 1 1446
2 80453 1 1446
2 80454 1 1446
2 80455 1 1449
2 80456 1 1449
2 80457 1 1449
2 80458 1 1449
2 80459 1 1449
2 80460 1 1451
2 80461 1 1451
2 80462 1 1451
2 80463 1 1451
2 80464 1 1451
2 80465 1 1451
2 80466 1 1451
2 80467 1 1451
2 80468 1 1451
2 80469 1 1451
2 80470 1 1452
2 80471 1 1452
2 80472 1 1452
2 80473 1 1452
2 80474 1 1453
2 80475 1 1453
2 80476 1 1453
2 80477 1 1453
2 80478 1 1453
2 80479 1 1453
2 80480 1 1453
2 80481 1 1453
2 80482 1 1453
2 80483 1 1454
2 80484 1 1454
2 80485 1 1456
2 80486 1 1456
2 80487 1 1456
2 80488 1 1457
2 80489 1 1457
2 80490 1 1457
2 80491 1 1457
2 80492 1 1457
2 80493 1 1458
2 80494 1 1458
2 80495 1 1458
2 80496 1 1458
2 80497 1 1458
2 80498 1 1458
2 80499 1 1458
2 80500 1 1458
2 80501 1 1458
2 80502 1 1459
2 80503 1 1459
2 80504 1 1459
2 80505 1 1459
2 80506 1 1459
2 80507 1 1459
2 80508 1 1459
2 80509 1 1460
2 80510 1 1460
2 80511 1 1460
2 80512 1 1460
2 80513 1 1460
2 80514 1 1460
2 80515 1 1460
2 80516 1 1460
2 80517 1 1460
2 80518 1 1460
2 80519 1 1460
2 80520 1 1460
2 80521 1 1460
2 80522 1 1460
2 80523 1 1460
2 80524 1 1460
2 80525 1 1460
2 80526 1 1460
2 80527 1 1460
2 80528 1 1460
2 80529 1 1460
2 80530 1 1460
2 80531 1 1460
2 80532 1 1461
2 80533 1 1461
2 80534 1 1462
2 80535 1 1462
2 80536 1 1462
2 80537 1 1462
2 80538 1 1462
2 80539 1 1469
2 80540 1 1469
2 80541 1 1469
2 80542 1 1469
2 80543 1 1469
2 80544 1 1469
2 80545 1 1469
2 80546 1 1469
2 80547 1 1469
2 80548 1 1469
2 80549 1 1469
2 80550 1 1471
2 80551 1 1471
2 80552 1 1471
2 80553 1 1471
2 80554 1 1471
2 80555 1 1471
2 80556 1 1471
2 80557 1 1471
2 80558 1 1484
2 80559 1 1484
2 80560 1 1484
2 80561 1 1485
2 80562 1 1485
2 80563 1 1485
2 80564 1 1485
2 80565 1 1485
2 80566 1 1485
2 80567 1 1485
2 80568 1 1485
2 80569 1 1485
2 80570 1 1485
2 80571 1 1485
2 80572 1 1485
2 80573 1 1485
2 80574 1 1485
2 80575 1 1485
2 80576 1 1485
2 80577 1 1485
2 80578 1 1485
2 80579 1 1485
2 80580 1 1485
2 80581 1 1485
2 80582 1 1485
2 80583 1 1485
2 80584 1 1485
2 80585 1 1485
2 80586 1 1485
2 80587 1 1485
2 80588 1 1485
2 80589 1 1485
2 80590 1 1485
2 80591 1 1485
2 80592 1 1485
2 80593 1 1485
2 80594 1 1485
2 80595 1 1485
2 80596 1 1485
2 80597 1 1485
2 80598 1 1485
2 80599 1 1485
2 80600 1 1485
2 80601 1 1485
2 80602 1 1485
2 80603 1 1485
2 80604 1 1485
2 80605 1 1485
2 80606 1 1485
2 80607 1 1485
2 80608 1 1485
2 80609 1 1485
2 80610 1 1485
2 80611 1 1485
2 80612 1 1485
2 80613 1 1485
2 80614 1 1485
2 80615 1 1485
2 80616 1 1485
2 80617 1 1485
2 80618 1 1485
2 80619 1 1485
2 80620 1 1485
2 80621 1 1485
2 80622 1 1485
2 80623 1 1485
2 80624 1 1485
2 80625 1 1485
2 80626 1 1485
2 80627 1 1485
2 80628 1 1485
2 80629 1 1485
2 80630 1 1485
2 80631 1 1485
2 80632 1 1485
2 80633 1 1485
2 80634 1 1485
2 80635 1 1485
2 80636 1 1485
2 80637 1 1485
2 80638 1 1485
2 80639 1 1485
2 80640 1 1485
2 80641 1 1485
2 80642 1 1485
2 80643 1 1485
2 80644 1 1485
2 80645 1 1485
2 80646 1 1485
2 80647 1 1485
2 80648 1 1485
2 80649 1 1485
2 80650 1 1485
2 80651 1 1485
2 80652 1 1485
2 80653 1 1485
2 80654 1 1485
2 80655 1 1485
2 80656 1 1485
2 80657 1 1485
2 80658 1 1485
2 80659 1 1485
2 80660 1 1485
2 80661 1 1485
2 80662 1 1485
2 80663 1 1485
2 80664 1 1485
2 80665 1 1485
2 80666 1 1485
2 80667 1 1485
2 80668 1 1485
2 80669 1 1486
2 80670 1 1486
2 80671 1 1486
2 80672 1 1486
2 80673 1 1486
2 80674 1 1486
2 80675 1 1486
2 80676 1 1486
2 80677 1 1486
2 80678 1 1486
2 80679 1 1486
2 80680 1 1486
2 80681 1 1486
2 80682 1 1486
2 80683 1 1486
2 80684 1 1486
2 80685 1 1486
2 80686 1 1486
2 80687 1 1486
2 80688 1 1486
2 80689 1 1486
2 80690 1 1486
2 80691 1 1486
2 80692 1 1486
2 80693 1 1486
2 80694 1 1486
2 80695 1 1486
2 80696 1 1486
2 80697 1 1486
2 80698 1 1486
2 80699 1 1486
2 80700 1 1486
2 80701 1 1486
2 80702 1 1486
2 80703 1 1486
2 80704 1 1486
2 80705 1 1486
2 80706 1 1486
2 80707 1 1486
2 80708 1 1486
2 80709 1 1486
2 80710 1 1486
2 80711 1 1486
2 80712 1 1486
2 80713 1 1486
2 80714 1 1486
2 80715 1 1486
2 80716 1 1486
2 80717 1 1486
2 80718 1 1486
2 80719 1 1486
2 80720 1 1486
2 80721 1 1486
2 80722 1 1486
2 80723 1 1486
2 80724 1 1486
2 80725 1 1486
2 80726 1 1486
2 80727 1 1486
2 80728 1 1486
2 80729 1 1486
2 80730 1 1486
2 80731 1 1486
2 80732 1 1486
2 80733 1 1486
2 80734 1 1486
2 80735 1 1486
2 80736 1 1486
2 80737 1 1486
2 80738 1 1486
2 80739 1 1486
2 80740 1 1486
2 80741 1 1486
2 80742 1 1486
2 80743 1 1486
2 80744 1 1486
2 80745 1 1486
2 80746 1 1486
2 80747 1 1486
2 80748 1 1486
2 80749 1 1486
2 80750 1 1486
2 80751 1 1486
2 80752 1 1486
2 80753 1 1486
2 80754 1 1486
2 80755 1 1486
2 80756 1 1486
2 80757 1 1486
2 80758 1 1486
2 80759 1 1486
2 80760 1 1486
2 80761 1 1486
2 80762 1 1486
2 80763 1 1486
2 80764 1 1486
2 80765 1 1486
2 80766 1 1486
2 80767 1 1486
2 80768 1 1486
2 80769 1 1486
2 80770 1 1486
2 80771 1 1486
2 80772 1 1486
2 80773 1 1486
2 80774 1 1486
2 80775 1 1486
2 80776 1 1486
2 80777 1 1486
2 80778 1 1486
2 80779 1 1486
2 80780 1 1486
2 80781 1 1486
2 80782 1 1486
2 80783 1 1486
2 80784 1 1486
2 80785 1 1486
2 80786 1 1486
2 80787 1 1486
2 80788 1 1487
2 80789 1 1487
2 80790 1 1487
2 80791 1 1487
2 80792 1 1487
2 80793 1 1489
2 80794 1 1489
2 80795 1 1489
2 80796 1 1489
2 80797 1 1489
2 80798 1 1489
2 80799 1 1490
2 80800 1 1490
2 80801 1 1490
2 80802 1 1490
2 80803 1 1490
2 80804 1 1492
2 80805 1 1492
2 80806 1 1492
2 80807 1 1493
2 80808 1 1493
2 80809 1 1493
2 80810 1 1493
2 80811 1 1493
2 80812 1 1493
2 80813 1 1493
2 80814 1 1493
2 80815 1 1494
2 80816 1 1494
2 80817 1 1496
2 80818 1 1496
2 80819 1 1497
2 80820 1 1497
2 80821 1 1498
2 80822 1 1498
2 80823 1 1498
2 80824 1 1509
2 80825 1 1509
2 80826 1 1509
2 80827 1 1509
2 80828 1 1509
2 80829 1 1509
2 80830 1 1509
2 80831 1 1509
2 80832 1 1509
2 80833 1 1509
2 80834 1 1509
2 80835 1 1509
2 80836 1 1509
2 80837 1 1509
2 80838 1 1509
2 80839 1 1509
2 80840 1 1509
2 80841 1 1509
2 80842 1 1511
2 80843 1 1511
2 80844 1 1512
2 80845 1 1512
2 80846 1 1512
2 80847 1 1512
2 80848 1 1512
2 80849 1 1512
2 80850 1 1512
2 80851 1 1512
2 80852 1 1512
2 80853 1 1512
2 80854 1 1512
2 80855 1 1512
2 80856 1 1512
2 80857 1 1512
2 80858 1 1512
2 80859 1 1513
2 80860 1 1513
2 80861 1 1513
2 80862 1 1513
2 80863 1 1513
2 80864 1 1513
2 80865 1 1513
2 80866 1 1513
2 80867 1 1513
2 80868 1 1513
2 80869 1 1513
2 80870 1 1513
2 80871 1 1513
2 80872 1 1513
2 80873 1 1513
2 80874 1 1513
2 80875 1 1513
2 80876 1 1513
2 80877 1 1513
2 80878 1 1514
2 80879 1 1514
2 80880 1 1514
2 80881 1 1514
2 80882 1 1514
2 80883 1 1514
2 80884 1 1514
2 80885 1 1514
2 80886 1 1515
2 80887 1 1515
2 80888 1 1515
2 80889 1 1517
2 80890 1 1517
2 80891 1 1520
2 80892 1 1520
2 80893 1 1520
2 80894 1 1520
2 80895 1 1520
2 80896 1 1520
2 80897 1 1520
2 80898 1 1520
2 80899 1 1520
2 80900 1 1520
2 80901 1 1520
2 80902 1 1520
2 80903 1 1521
2 80904 1 1521
2 80905 1 1522
2 80906 1 1522
2 80907 1 1522
2 80908 1 1522
2 80909 1 1522
2 80910 1 1522
2 80911 1 1523
2 80912 1 1523
2 80913 1 1533
2 80914 1 1533
2 80915 1 1549
2 80916 1 1549
2 80917 1 1549
2 80918 1 1550
2 80919 1 1550
2 80920 1 1550
2 80921 1 1550
2 80922 1 1550
2 80923 1 1550
2 80924 1 1550
2 80925 1 1550
2 80926 1 1550
2 80927 1 1550
2 80928 1 1550
2 80929 1 1551
2 80930 1 1551
2 80931 1 1552
2 80932 1 1552
2 80933 1 1552
2 80934 1 1552
2 80935 1 1552
2 80936 1 1552
2 80937 1 1552
2 80938 1 1552
2 80939 1 1552
2 80940 1 1552
2 80941 1 1552
2 80942 1 1552
2 80943 1 1552
2 80944 1 1552
2 80945 1 1552
2 80946 1 1552
2 80947 1 1552
2 80948 1 1552
2 80949 1 1552
2 80950 1 1553
2 80951 1 1553
2 80952 1 1553
2 80953 1 1557
2 80954 1 1557
2 80955 1 1557
2 80956 1 1565
2 80957 1 1565
2 80958 1 1565
2 80959 1 1565
2 80960 1 1565
2 80961 1 1566
2 80962 1 1566
2 80963 1 1567
2 80964 1 1567
2 80965 1 1570
2 80966 1 1570
2 80967 1 1570
2 80968 1 1570
2 80969 1 1578
2 80970 1 1578
2 80971 1 1578
2 80972 1 1578
2 80973 1 1578
2 80974 1 1578
2 80975 1 1578
2 80976 1 1578
2 80977 1 1579
2 80978 1 1579
2 80979 1 1583
2 80980 1 1583
2 80981 1 1583
2 80982 1 1583
2 80983 1 1583
2 80984 1 1583
2 80985 1 1583
2 80986 1 1583
2 80987 1 1583
2 80988 1 1583
2 80989 1 1583
2 80990 1 1583
2 80991 1 1583
2 80992 1 1583
2 80993 1 1583
2 80994 1 1583
2 80995 1 1583
2 80996 1 1583
2 80997 1 1584
2 80998 1 1584
2 80999 1 1584
2 81000 1 1584
2 81001 1 1585
2 81002 1 1585
2 81003 1 1585
2 81004 1 1585
2 81005 1 1585
2 81006 1 1585
2 81007 1 1585
2 81008 1 1585
2 81009 1 1585
2 81010 1 1585
2 81011 1 1585
2 81012 1 1585
2 81013 1 1586
2 81014 1 1586
2 81015 1 1586
2 81016 1 1586
2 81017 1 1586
2 81018 1 1586
2 81019 1 1586
2 81020 1 1586
2 81021 1 1586
2 81022 1 1586
2 81023 1 1586
2 81024 1 1586
2 81025 1 1586
2 81026 1 1586
2 81027 1 1586
2 81028 1 1586
2 81029 1 1586
2 81030 1 1586
2 81031 1 1586
2 81032 1 1586
2 81033 1 1586
2 81034 1 1586
2 81035 1 1586
2 81036 1 1586
2 81037 1 1586
2 81038 1 1586
2 81039 1 1586
2 81040 1 1586
2 81041 1 1586
2 81042 1 1586
2 81043 1 1586
2 81044 1 1586
2 81045 1 1586
2 81046 1 1586
2 81047 1 1586
2 81048 1 1586
2 81049 1 1586
2 81050 1 1586
2 81051 1 1586
2 81052 1 1586
2 81053 1 1586
2 81054 1 1586
2 81055 1 1586
2 81056 1 1586
2 81057 1 1586
2 81058 1 1586
2 81059 1 1586
2 81060 1 1586
2 81061 1 1586
2 81062 1 1586
2 81063 1 1586
2 81064 1 1586
2 81065 1 1586
2 81066 1 1586
2 81067 1 1586
2 81068 1 1586
2 81069 1 1586
2 81070 1 1586
2 81071 1 1586
2 81072 1 1586
2 81073 1 1586
2 81074 1 1586
2 81075 1 1586
2 81076 1 1586
2 81077 1 1586
2 81078 1 1586
2 81079 1 1586
2 81080 1 1586
2 81081 1 1586
2 81082 1 1586
2 81083 1 1586
2 81084 1 1586
2 81085 1 1586
2 81086 1 1586
2 81087 1 1587
2 81088 1 1587
2 81089 1 1587
2 81090 1 1587
2 81091 1 1589
2 81092 1 1589
2 81093 1 1589
2 81094 1 1589
2 81095 1 1591
2 81096 1 1591
2 81097 1 1591
2 81098 1 1597
2 81099 1 1597
2 81100 1 1597
2 81101 1 1606
2 81102 1 1606
2 81103 1 1606
2 81104 1 1606
2 81105 1 1606
2 81106 1 1606
2 81107 1 1606
2 81108 1 1606
2 81109 1 1606
2 81110 1 1606
2 81111 1 1606
2 81112 1 1607
2 81113 1 1607
2 81114 1 1607
2 81115 1 1607
2 81116 1 1607
2 81117 1 1608
2 81118 1 1608
2 81119 1 1608
2 81120 1 1617
2 81121 1 1617
2 81122 1 1617
2 81123 1 1617
2 81124 1 1617
2 81125 1 1628
2 81126 1 1628
2 81127 1 1628
2 81128 1 1628
2 81129 1 1628
2 81130 1 1628
2 81131 1 1628
2 81132 1 1628
2 81133 1 1628
2 81134 1 1628
2 81135 1 1628
2 81136 1 1628
2 81137 1 1628
2 81138 1 1628
2 81139 1 1628
2 81140 1 1628
2 81141 1 1628
2 81142 1 1628
2 81143 1 1628
2 81144 1 1628
2 81145 1 1629
2 81146 1 1629
2 81147 1 1630
2 81148 1 1630
2 81149 1 1630
2 81150 1 1630
2 81151 1 1642
2 81152 1 1642
2 81153 1 1642
2 81154 1 1642
2 81155 1 1642
2 81156 1 1642
2 81157 1 1642
2 81158 1 1642
2 81159 1 1642
2 81160 1 1642
2 81161 1 1642
2 81162 1 1642
2 81163 1 1642
2 81164 1 1645
2 81165 1 1645
2 81166 1 1646
2 81167 1 1646
2 81168 1 1647
2 81169 1 1647
2 81170 1 1647
2 81171 1 1649
2 81172 1 1649
2 81173 1 1649
2 81174 1 1649
2 81175 1 1649
2 81176 1 1649
2 81177 1 1649
2 81178 1 1649
2 81179 1 1650
2 81180 1 1650
2 81181 1 1650
2 81182 1 1650
2 81183 1 1650
2 81184 1 1650
2 81185 1 1650
2 81186 1 1651
2 81187 1 1651
2 81188 1 1651
2 81189 1 1651
2 81190 1 1651
2 81191 1 1652
2 81192 1 1652
2 81193 1 1652
2 81194 1 1652
2 81195 1 1652
2 81196 1 1652
2 81197 1 1660
2 81198 1 1660
2 81199 1 1660
2 81200 1 1661
2 81201 1 1661
2 81202 1 1661
2 81203 1 1661
2 81204 1 1661
2 81205 1 1661
2 81206 1 1661
2 81207 1 1661
2 81208 1 1661
2 81209 1 1661
2 81210 1 1661
2 81211 1 1661
2 81212 1 1661
2 81213 1 1661
2 81214 1 1661
2 81215 1 1661
2 81216 1 1661
2 81217 1 1661
2 81218 1 1661
2 81219 1 1662
2 81220 1 1662
2 81221 1 1662
2 81222 1 1662
2 81223 1 1662
2 81224 1 1662
2 81225 1 1662
2 81226 1 1667
2 81227 1 1667
2 81228 1 1667
2 81229 1 1667
2 81230 1 1667
2 81231 1 1667
2 81232 1 1667
2 81233 1 1667
2 81234 1 1667
2 81235 1 1667
2 81236 1 1667
2 81237 1 1667
2 81238 1 1667
2 81239 1 1667
2 81240 1 1667
2 81241 1 1667
2 81242 1 1667
2 81243 1 1667
2 81244 1 1668
2 81245 1 1668
2 81246 1 1668
2 81247 1 1668
2 81248 1 1668
2 81249 1 1668
2 81250 1 1668
2 81251 1 1668
2 81252 1 1668
2 81253 1 1674
2 81254 1 1674
2 81255 1 1676
2 81256 1 1676
2 81257 1 1682
2 81258 1 1682
2 81259 1 1682
2 81260 1 1682
2 81261 1 1682
2 81262 1 1682
2 81263 1 1682
2 81264 1 1682
2 81265 1 1683
2 81266 1 1683
2 81267 1 1683
2 81268 1 1683
2 81269 1 1684
2 81270 1 1684
2 81271 1 1684
2 81272 1 1685
2 81273 1 1685
2 81274 1 1686
2 81275 1 1686
2 81276 1 1687
2 81277 1 1687
2 81278 1 1687
2 81279 1 1687
2 81280 1 1687
2 81281 1 1687
2 81282 1 1687
2 81283 1 1687
2 81284 1 1687
2 81285 1 1687
2 81286 1 1687
2 81287 1 1687
2 81288 1 1687
2 81289 1 1687
2 81290 1 1687
2 81291 1 1687
2 81292 1 1687
2 81293 1 1688
2 81294 1 1688
2 81295 1 1693
2 81296 1 1693
2 81297 1 1696
2 81298 1 1696
2 81299 1 1696
2 81300 1 1696
2 81301 1 1696
2 81302 1 1696
2 81303 1 1696
2 81304 1 1696
2 81305 1 1705
2 81306 1 1705
2 81307 1 1705
2 81308 1 1705
2 81309 1 1705
2 81310 1 1705
2 81311 1 1705
2 81312 1 1705
2 81313 1 1705
2 81314 1 1705
2 81315 1 1706
2 81316 1 1706
2 81317 1 1706
2 81318 1 1706
2 81319 1 1706
2 81320 1 1706
2 81321 1 1706
2 81322 1 1706
2 81323 1 1707
2 81324 1 1707
2 81325 1 1707
2 81326 1 1708
2 81327 1 1708
2 81328 1 1708
2 81329 1 1708
2 81330 1 1708
2 81331 1 1710
2 81332 1 1710
2 81333 1 1710
2 81334 1 1710
2 81335 1 1710
2 81336 1 1712
2 81337 1 1712
2 81338 1 1729
2 81339 1 1729
2 81340 1 1729
2 81341 1 1729
2 81342 1 1729
2 81343 1 1729
2 81344 1 1729
2 81345 1 1729
2 81346 1 1729
2 81347 1 1729
2 81348 1 1729
2 81349 1 1729
2 81350 1 1729
2 81351 1 1729
2 81352 1 1730
2 81353 1 1730
2 81354 1 1730
2 81355 1 1732
2 81356 1 1732
2 81357 1 1732
2 81358 1 1732
2 81359 1 1732
2 81360 1 1732
2 81361 1 1732
2 81362 1 1732
2 81363 1 1732
2 81364 1 1732
2 81365 1 1732
2 81366 1 1733
2 81367 1 1733
2 81368 1 1733
2 81369 1 1733
2 81370 1 1733
2 81371 1 1735
2 81372 1 1735
2 81373 1 1735
2 81374 1 1735
2 81375 1 1735
2 81376 1 1735
2 81377 1 1735
2 81378 1 1736
2 81379 1 1736
2 81380 1 1737
2 81381 1 1737
2 81382 1 1738
2 81383 1 1738
2 81384 1 1743
2 81385 1 1743
2 81386 1 1752
2 81387 1 1752
2 81388 1 1752
2 81389 1 1752
2 81390 1 1752
2 81391 1 1752
2 81392 1 1752
2 81393 1 1752
2 81394 1 1752
2 81395 1 1752
2 81396 1 1752
2 81397 1 1752
2 81398 1 1752
2 81399 1 1752
2 81400 1 1752
2 81401 1 1752
2 81402 1 1752
2 81403 1 1752
2 81404 1 1752
2 81405 1 1752
2 81406 1 1752
2 81407 1 1754
2 81408 1 1754
2 81409 1 1754
2 81410 1 1754
2 81411 1 1754
2 81412 1 1754
2 81413 1 1754
2 81414 1 1754
2 81415 1 1754
2 81416 1 1754
2 81417 1 1754
2 81418 1 1754
2 81419 1 1754
2 81420 1 1754
2 81421 1 1754
2 81422 1 1754
2 81423 1 1754
2 81424 1 1754
2 81425 1 1755
2 81426 1 1755
2 81427 1 1755
2 81428 1 1755
2 81429 1 1755
2 81430 1 1755
2 81431 1 1755
2 81432 1 1755
2 81433 1 1755
2 81434 1 1755
2 81435 1 1755
2 81436 1 1755
2 81437 1 1755
2 81438 1 1755
2 81439 1 1755
2 81440 1 1755
2 81441 1 1755
2 81442 1 1755
2 81443 1 1755
2 81444 1 1755
2 81445 1 1755
2 81446 1 1758
2 81447 1 1758
2 81448 1 1763
2 81449 1 1763
2 81450 1 1764
2 81451 1 1764
2 81452 1 1774
2 81453 1 1774
2 81454 1 1774
2 81455 1 1774
2 81456 1 1774
2 81457 1 1774
2 81458 1 1774
2 81459 1 1774
2 81460 1 1774
2 81461 1 1774
2 81462 1 1774
2 81463 1 1774
2 81464 1 1774
2 81465 1 1774
2 81466 1 1774
2 81467 1 1774
2 81468 1 1774
2 81469 1 1774
2 81470 1 1774
2 81471 1 1774
2 81472 1 1774
2 81473 1 1774
2 81474 1 1774
2 81475 1 1774
2 81476 1 1774
2 81477 1 1774
2 81478 1 1774
2 81479 1 1774
2 81480 1 1774
2 81481 1 1774
2 81482 1 1774
2 81483 1 1774
2 81484 1 1774
2 81485 1 1774
2 81486 1 1774
2 81487 1 1774
2 81488 1 1774
2 81489 1 1774
2 81490 1 1774
2 81491 1 1775
2 81492 1 1775
2 81493 1 1775
2 81494 1 1775
2 81495 1 1775
2 81496 1 1776
2 81497 1 1776
2 81498 1 1776
2 81499 1 1776
2 81500 1 1776
2 81501 1 1776
2 81502 1 1776
2 81503 1 1776
2 81504 1 1776
2 81505 1 1776
2 81506 1 1776
2 81507 1 1776
2 81508 1 1776
2 81509 1 1776
2 81510 1 1776
2 81511 1 1779
2 81512 1 1779
2 81513 1 1787
2 81514 1 1787
2 81515 1 1788
2 81516 1 1788
2 81517 1 1788
2 81518 1 1788
2 81519 1 1788
2 81520 1 1788
2 81521 1 1788
2 81522 1 1788
2 81523 1 1788
2 81524 1 1788
2 81525 1 1788
2 81526 1 1788
2 81527 1 1788
2 81528 1 1788
2 81529 1 1788
2 81530 1 1788
2 81531 1 1788
2 81532 1 1788
2 81533 1 1788
2 81534 1 1788
2 81535 1 1788
2 81536 1 1788
2 81537 1 1788
2 81538 1 1788
2 81539 1 1788
2 81540 1 1788
2 81541 1 1788
2 81542 1 1788
2 81543 1 1789
2 81544 1 1789
2 81545 1 1789
2 81546 1 1798
2 81547 1 1798
2 81548 1 1800
2 81549 1 1800
2 81550 1 1800
2 81551 1 1800
2 81552 1 1800
2 81553 1 1802
2 81554 1 1802
2 81555 1 1802
2 81556 1 1802
2 81557 1 1802
2 81558 1 1802
2 81559 1 1802
2 81560 1 1803
2 81561 1 1803
2 81562 1 1806
2 81563 1 1806
2 81564 1 1806
2 81565 1 1806
2 81566 1 1806
2 81567 1 1816
2 81568 1 1816
2 81569 1 1816
2 81570 1 1816
2 81571 1 1816
2 81572 1 1816
2 81573 1 1816
2 81574 1 1816
2 81575 1 1816
2 81576 1 1816
2 81577 1 1816
2 81578 1 1817
2 81579 1 1817
2 81580 1 1817
2 81581 1 1817
2 81582 1 1817
2 81583 1 1817
2 81584 1 1817
2 81585 1 1817
2 81586 1 1817
2 81587 1 1817
2 81588 1 1817
2 81589 1 1818
2 81590 1 1818
2 81591 1 1818
2 81592 1 1819
2 81593 1 1819
2 81594 1 1819
2 81595 1 1819
2 81596 1 1819
2 81597 1 1819
2 81598 1 1819
2 81599 1 1828
2 81600 1 1828
2 81601 1 1828
2 81602 1 1828
2 81603 1 1828
2 81604 1 1828
2 81605 1 1828
2 81606 1 1841
2 81607 1 1841
2 81608 1 1841
2 81609 1 1841
2 81610 1 1841
2 81611 1 1841
2 81612 1 1841
2 81613 1 1841
2 81614 1 1841
2 81615 1 1841
2 81616 1 1842
2 81617 1 1842
2 81618 1 1842
2 81619 1 1842
2 81620 1 1843
2 81621 1 1843
2 81622 1 1843
2 81623 1 1844
2 81624 1 1844
2 81625 1 1844
2 81626 1 1845
2 81627 1 1845
2 81628 1 1845
2 81629 1 1850
2 81630 1 1850
2 81631 1 1851
2 81632 1 1851
2 81633 1 1851
2 81634 1 1852
2 81635 1 1852
2 81636 1 1867
2 81637 1 1867
2 81638 1 1868
2 81639 1 1868
2 81640 1 1868
2 81641 1 1870
2 81642 1 1870
2 81643 1 1877
2 81644 1 1877
2 81645 1 1877
2 81646 1 1877
2 81647 1 1877
2 81648 1 1877
2 81649 1 1877
2 81650 1 1877
2 81651 1 1878
2 81652 1 1878
2 81653 1 1878
2 81654 1 1880
2 81655 1 1880
2 81656 1 1880
2 81657 1 1880
2 81658 1 1881
2 81659 1 1881
2 81660 1 1881
2 81661 1 1883
2 81662 1 1883
2 81663 1 1898
2 81664 1 1898
2 81665 1 1898
2 81666 1 1898
2 81667 1 1898
2 81668 1 1898
2 81669 1 1899
2 81670 1 1899
2 81671 1 1899
2 81672 1 1922
2 81673 1 1922
2 81674 1 1922
2 81675 1 1922
2 81676 1 1922
2 81677 1 1922
2 81678 1 1922
2 81679 1 1922
2 81680 1 1922
2 81681 1 1922
2 81682 1 1922
2 81683 1 1922
2 81684 1 1922
2 81685 1 1922
2 81686 1 1922
2 81687 1 1922
2 81688 1 1922
2 81689 1 1922
2 81690 1 1922
2 81691 1 1922
2 81692 1 1922
2 81693 1 1922
2 81694 1 1922
2 81695 1 1922
2 81696 1 1922
2 81697 1 1922
2 81698 1 1922
2 81699 1 1922
2 81700 1 1922
2 81701 1 1922
2 81702 1 1922
2 81703 1 1922
2 81704 1 1922
2 81705 1 1922
2 81706 1 1922
2 81707 1 1922
2 81708 1 1922
2 81709 1 1922
2 81710 1 1922
2 81711 1 1922
2 81712 1 1922
2 81713 1 1922
2 81714 1 1922
2 81715 1 1922
2 81716 1 1922
2 81717 1 1922
2 81718 1 1922
2 81719 1 1922
2 81720 1 1922
2 81721 1 1922
2 81722 1 1922
2 81723 1 1922
2 81724 1 1922
2 81725 1 1922
2 81726 1 1922
2 81727 1 1922
2 81728 1 1922
2 81729 1 1922
2 81730 1 1922
2 81731 1 1922
2 81732 1 1922
2 81733 1 1922
2 81734 1 1922
2 81735 1 1922
2 81736 1 1922
2 81737 1 1922
2 81738 1 1922
2 81739 1 1922
2 81740 1 1922
2 81741 1 1922
2 81742 1 1922
2 81743 1 1922
2 81744 1 1922
2 81745 1 1922
2 81746 1 1922
2 81747 1 1922
2 81748 1 1922
2 81749 1 1922
2 81750 1 1922
2 81751 1 1922
2 81752 1 1922
2 81753 1 1922
2 81754 1 1922
2 81755 1 1922
2 81756 1 1922
2 81757 1 1922
2 81758 1 1922
2 81759 1 1922
2 81760 1 1922
2 81761 1 1922
2 81762 1 1922
2 81763 1 1922
2 81764 1 1922
2 81765 1 1922
2 81766 1 1922
2 81767 1 1922
2 81768 1 1922
2 81769 1 1922
2 81770 1 1922
2 81771 1 1922
2 81772 1 1922
2 81773 1 1922
2 81774 1 1922
2 81775 1 1922
2 81776 1 1922
2 81777 1 1922
2 81778 1 1922
2 81779 1 1922
2 81780 1 1922
2 81781 1 1922
2 81782 1 1922
2 81783 1 1922
2 81784 1 1922
2 81785 1 1922
2 81786 1 1922
2 81787 1 1922
2 81788 1 1922
2 81789 1 1922
2 81790 1 1922
2 81791 1 1922
2 81792 1 1922
2 81793 1 1922
2 81794 1 1922
2 81795 1 1922
2 81796 1 1922
2 81797 1 1922
2 81798 1 1922
2 81799 1 1922
2 81800 1 1922
2 81801 1 1922
2 81802 1 1922
2 81803 1 1922
2 81804 1 1922
2 81805 1 1922
2 81806 1 1922
2 81807 1 1922
2 81808 1 1922
2 81809 1 1923
2 81810 1 1923
2 81811 1 1923
2 81812 1 1923
2 81813 1 1923
2 81814 1 1923
2 81815 1 1923
2 81816 1 1923
2 81817 1 1923
2 81818 1 1923
2 81819 1 1923
2 81820 1 1923
2 81821 1 1923
2 81822 1 1923
2 81823 1 1923
2 81824 1 1923
2 81825 1 1923
2 81826 1 1923
2 81827 1 1923
2 81828 1 1923
2 81829 1 1923
2 81830 1 1923
2 81831 1 1923
2 81832 1 1923
2 81833 1 1923
2 81834 1 1923
2 81835 1 1923
2 81836 1 1923
2 81837 1 1923
2 81838 1 1923
2 81839 1 1923
2 81840 1 1923
2 81841 1 1923
2 81842 1 1923
2 81843 1 1923
2 81844 1 1923
2 81845 1 1923
2 81846 1 1923
2 81847 1 1923
2 81848 1 1923
2 81849 1 1923
2 81850 1 1923
2 81851 1 1923
2 81852 1 1923
2 81853 1 1923
2 81854 1 1923
2 81855 1 1923
2 81856 1 1923
2 81857 1 1923
2 81858 1 1923
2 81859 1 1923
2 81860 1 1923
2 81861 1 1923
2 81862 1 1923
2 81863 1 1923
2 81864 1 1923
2 81865 1 1923
2 81866 1 1923
2 81867 1 1923
2 81868 1 1923
2 81869 1 1923
2 81870 1 1923
2 81871 1 1923
2 81872 1 1923
2 81873 1 1923
2 81874 1 1923
2 81875 1 1923
2 81876 1 1923
2 81877 1 1923
2 81878 1 1923
2 81879 1 1923
2 81880 1 1923
2 81881 1 1923
2 81882 1 1923
2 81883 1 1923
2 81884 1 1923
2 81885 1 1923
2 81886 1 1923
2 81887 1 1923
2 81888 1 1923
2 81889 1 1923
2 81890 1 1923
2 81891 1 1923
2 81892 1 1923
2 81893 1 1923
2 81894 1 1923
2 81895 1 1923
2 81896 1 1923
2 81897 1 1923
2 81898 1 1923
2 81899 1 1923
2 81900 1 1923
2 81901 1 1923
2 81902 1 1923
2 81903 1 1923
2 81904 1 1923
2 81905 1 1923
2 81906 1 1923
2 81907 1 1923
2 81908 1 1923
2 81909 1 1923
2 81910 1 1923
2 81911 1 1923
2 81912 1 1923
2 81913 1 1923
2 81914 1 1923
2 81915 1 1923
2 81916 1 1923
2 81917 1 1923
2 81918 1 1923
2 81919 1 1923
2 81920 1 1923
2 81921 1 1923
2 81922 1 1923
2 81923 1 1923
2 81924 1 1923
2 81925 1 1923
2 81926 1 1923
2 81927 1 1923
2 81928 1 1923
2 81929 1 1923
2 81930 1 1923
2 81931 1 1923
2 81932 1 1923
2 81933 1 1923
2 81934 1 1923
2 81935 1 1923
2 81936 1 1923
2 81937 1 1923
2 81938 1 1923
2 81939 1 1923
2 81940 1 1923
2 81941 1 1923
2 81942 1 1923
2 81943 1 1923
2 81944 1 1923
2 81945 1 1923
2 81946 1 1923
2 81947 1 1923
2 81948 1 1923
2 81949 1 1923
2 81950 1 1923
2 81951 1 1923
2 81952 1 1923
2 81953 1 1923
2 81954 1 1924
2 81955 1 1924
2 81956 1 1924
2 81957 1 1924
2 81958 1 1924
2 81959 1 1924
2 81960 1 1924
2 81961 1 1924
2 81962 1 1924
2 81963 1 1924
2 81964 1 1924
2 81965 1 1924
2 81966 1 1924
2 81967 1 1924
2 81968 1 1924
2 81969 1 1924
2 81970 1 1924
2 81971 1 1924
2 81972 1 1924
2 81973 1 1924
2 81974 1 1926
2 81975 1 1926
2 81976 1 1926
2 81977 1 1928
2 81978 1 1928
2 81979 1 1935
2 81980 1 1935
2 81981 1 1936
2 81982 1 1936
2 81983 1 1936
2 81984 1 1936
2 81985 1 1936
2 81986 1 1936
2 81987 1 1936
2 81988 1 1937
2 81989 1 1937
2 81990 1 1937
2 81991 1 1937
2 81992 1 1938
2 81993 1 1938
2 81994 1 1938
2 81995 1 1938
2 81996 1 1943
2 81997 1 1943
2 81998 1 1946
2 81999 1 1946
2 82000 1 1946
2 82001 1 1946
2 82002 1 1946
2 82003 1 1946
2 82004 1 1946
2 82005 1 1946
2 82006 1 1946
2 82007 1 1946
2 82008 1 1946
2 82009 1 1946
2 82010 1 1946
2 82011 1 1946
2 82012 1 1946
2 82013 1 1946
2 82014 1 1946
2 82015 1 1946
2 82016 1 1946
2 82017 1 1947
2 82018 1 1947
2 82019 1 1948
2 82020 1 1948
2 82021 1 1948
2 82022 1 1956
2 82023 1 1956
2 82024 1 1956
2 82025 1 1956
2 82026 1 1956
2 82027 1 1956
2 82028 1 1956
2 82029 1 1956
2 82030 1 1956
2 82031 1 1956
2 82032 1 1956
2 82033 1 1956
2 82034 1 1957
2 82035 1 1957
2 82036 1 1957
2 82037 1 1957
2 82038 1 1957
2 82039 1 1957
2 82040 1 1957
2 82041 1 1957
2 82042 1 1957
2 82043 1 1957
2 82044 1 1957
2 82045 1 1957
2 82046 1 1957
2 82047 1 1957
2 82048 1 1957
2 82049 1 1957
2 82050 1 1958
2 82051 1 1958
2 82052 1 1958
2 82053 1 1958
2 82054 1 1958
2 82055 1 1958
2 82056 1 1958
2 82057 1 1958
2 82058 1 1958
2 82059 1 1958
2 82060 1 1959
2 82061 1 1959
2 82062 1 1959
2 82063 1 1959
2 82064 1 1961
2 82065 1 1961
2 82066 1 1963
2 82067 1 1963
2 82068 1 1971
2 82069 1 1971
2 82070 1 1971
2 82071 1 1972
2 82072 1 1972
2 82073 1 1973
2 82074 1 1973
2 82075 1 1977
2 82076 1 1977
2 82077 1 1977
2 82078 1 1977
2 82079 1 1977
2 82080 1 1977
2 82081 1 1977
2 82082 1 1977
2 82083 1 1977
2 82084 1 1977
2 82085 1 1979
2 82086 1 1979
2 82087 1 1979
2 82088 1 1981
2 82089 1 1981
2 82090 1 1982
2 82091 1 1982
2 82092 1 1989
2 82093 1 1989
2 82094 1 1989
2 82095 1 1989
2 82096 1 1989
2 82097 1 1989
2 82098 1 1989
2 82099 1 1989
2 82100 1 1989
2 82101 1 1989
2 82102 1 1989
2 82103 1 1989
2 82104 1 1989
2 82105 1 1989
2 82106 1 1989
2 82107 1 1989
2 82108 1 1989
2 82109 1 1989
2 82110 1 1989
2 82111 1 1989
2 82112 1 1989
2 82113 1 1989
2 82114 1 1989
2 82115 1 1989
2 82116 1 1989
2 82117 1 1989
2 82118 1 1989
2 82119 1 1989
2 82120 1 1989
2 82121 1 1989
2 82122 1 1989
2 82123 1 1989
2 82124 1 1989
2 82125 1 1989
2 82126 1 1989
2 82127 1 1990
2 82128 1 1990
2 82129 1 1991
2 82130 1 1991
2 82131 1 1991
2 82132 1 1991
2 82133 1 1991
2 82134 1 1991
2 82135 1 1991
2 82136 1 1991
2 82137 1 1991
2 82138 1 1991
2 82139 1 1991
2 82140 1 1991
2 82141 1 1991
2 82142 1 1991
2 82143 1 1991
2 82144 1 1991
2 82145 1 1991
2 82146 1 1991
2 82147 1 1991
2 82148 1 1991
2 82149 1 1991
2 82150 1 1992
2 82151 1 1992
2 82152 1 1992
2 82153 1 1993
2 82154 1 1993
2 82155 1 1996
2 82156 1 1996
2 82157 1 1996
2 82158 1 1996
2 82159 1 1996
2 82160 1 1996
2 82161 1 1998
2 82162 1 1998
2 82163 1 1999
2 82164 1 1999
2 82165 1 1999
2 82166 1 1999
2 82167 1 1999
2 82168 1 1999
2 82169 1 1999
2 82170 1 1999
2 82171 1 1999
2 82172 1 1999
2 82173 1 1999
2 82174 1 1999
2 82175 1 1999
2 82176 1 2000
2 82177 1 2000
2 82178 1 2000
2 82179 1 2000
2 82180 1 2000
2 82181 1 2000
2 82182 1 2000
2 82183 1 2001
2 82184 1 2001
2 82185 1 2001
2 82186 1 2001
2 82187 1 2001
2 82188 1 2001
2 82189 1 2001
2 82190 1 2001
2 82191 1 2001
2 82192 1 2001
2 82193 1 2001
2 82194 1 2001
2 82195 1 2001
2 82196 1 2001
2 82197 1 2001
2 82198 1 2001
2 82199 1 2001
2 82200 1 2001
2 82201 1 2001
2 82202 1 2001
2 82203 1 2001
2 82204 1 2001
2 82205 1 2001
2 82206 1 2003
2 82207 1 2003
2 82208 1 2003
2 82209 1 2016
2 82210 1 2016
2 82211 1 2017
2 82212 1 2017
2 82213 1 2017
2 82214 1 2017
2 82215 1 2017
2 82216 1 2017
2 82217 1 2017
2 82218 1 2017
2 82219 1 2017
2 82220 1 2017
2 82221 1 2031
2 82222 1 2031
2 82223 1 2031
2 82224 1 2031
2 82225 1 2031
2 82226 1 2031
2 82227 1 2031
2 82228 1 2031
2 82229 1 2031
2 82230 1 2032
2 82231 1 2032
2 82232 1 2033
2 82233 1 2033
2 82234 1 2035
2 82235 1 2035
2 82236 1 2035
2 82237 1 2035
2 82238 1 2035
2 82239 1 2035
2 82240 1 2035
2 82241 1 2035
2 82242 1 2035
2 82243 1 2035
2 82244 1 2035
2 82245 1 2035
2 82246 1 2035
2 82247 1 2035
2 82248 1 2035
2 82249 1 2035
2 82250 1 2035
2 82251 1 2035
2 82252 1 2035
2 82253 1 2035
2 82254 1 2037
2 82255 1 2037
2 82256 1 2050
2 82257 1 2050
2 82258 1 2050
2 82259 1 2057
2 82260 1 2057
2 82261 1 2057
2 82262 1 2057
2 82263 1 2059
2 82264 1 2059
2 82265 1 2059
2 82266 1 2060
2 82267 1 2060
2 82268 1 2062
2 82269 1 2062
2 82270 1 2063
2 82271 1 2063
2 82272 1 2063
2 82273 1 2063
2 82274 1 2063
2 82275 1 2063
2 82276 1 2063
2 82277 1 2063
2 82278 1 2063
2 82279 1 2063
2 82280 1 2064
2 82281 1 2064
2 82282 1 2064
2 82283 1 2064
2 82284 1 2064
2 82285 1 2064
2 82286 1 2064
2 82287 1 2073
2 82288 1 2073
2 82289 1 2077
2 82290 1 2077
2 82291 1 2077
2 82292 1 2077
2 82293 1 2078
2 82294 1 2078
2 82295 1 2078
2 82296 1 2078
2 82297 1 2078
2 82298 1 2078
2 82299 1 2078
2 82300 1 2078
2 82301 1 2078
2 82302 1 2078
2 82303 1 2083
2 82304 1 2083
2 82305 1 2083
2 82306 1 2083
2 82307 1 2083
2 82308 1 2083
2 82309 1 2083
2 82310 1 2083
2 82311 1 2083
2 82312 1 2084
2 82313 1 2084
2 82314 1 2084
2 82315 1 2084
2 82316 1 2084
2 82317 1 2084
2 82318 1 2084
2 82319 1 2084
2 82320 1 2084
2 82321 1 2084
2 82322 1 2084
2 82323 1 2084
2 82324 1 2084
2 82325 1 2084
2 82326 1 2084
2 82327 1 2084
2 82328 1 2084
2 82329 1 2084
2 82330 1 2084
2 82331 1 2084
2 82332 1 2084
2 82333 1 2084
2 82334 1 2086
2 82335 1 2086
2 82336 1 2096
2 82337 1 2096
2 82338 1 2096
2 82339 1 2096
2 82340 1 2096
2 82341 1 2096
2 82342 1 2096
2 82343 1 2096
2 82344 1 2096
2 82345 1 2096
2 82346 1 2096
2 82347 1 2096
2 82348 1 2096
2 82349 1 2096
2 82350 1 2096
2 82351 1 2096
2 82352 1 2096
2 82353 1 2096
2 82354 1 2096
2 82355 1 2096
2 82356 1 2096
2 82357 1 2096
2 82358 1 2096
2 82359 1 2096
2 82360 1 2096
2 82361 1 2097
2 82362 1 2097
2 82363 1 2097
2 82364 1 2097
2 82365 1 2097
2 82366 1 2097
2 82367 1 2097
2 82368 1 2097
2 82369 1 2097
2 82370 1 2097
2 82371 1 2097
2 82372 1 2097
2 82373 1 2097
2 82374 1 2097
2 82375 1 2098
2 82376 1 2098
2 82377 1 2098
2 82378 1 2098
2 82379 1 2098
2 82380 1 2098
2 82381 1 2098
2 82382 1 2098
2 82383 1 2098
2 82384 1 2098
2 82385 1 2098
2 82386 1 2098
2 82387 1 2098
2 82388 1 2098
2 82389 1 2098
2 82390 1 2098
2 82391 1 2098
2 82392 1 2098
2 82393 1 2098
2 82394 1 2099
2 82395 1 2099
2 82396 1 2099
2 82397 1 2100
2 82398 1 2100
2 82399 1 2100
2 82400 1 2102
2 82401 1 2102
2 82402 1 2102
2 82403 1 2102
2 82404 1 2102
2 82405 1 2102
2 82406 1 2104
2 82407 1 2104
2 82408 1 2112
2 82409 1 2112
2 82410 1 2112
2 82411 1 2112
2 82412 1 2112
2 82413 1 2112
2 82414 1 2112
2 82415 1 2112
2 82416 1 2112
2 82417 1 2112
2 82418 1 2113
2 82419 1 2113
2 82420 1 2114
2 82421 1 2114
2 82422 1 2117
2 82423 1 2117
2 82424 1 2117
2 82425 1 2117
2 82426 1 2117
2 82427 1 2117
2 82428 1 2117
2 82429 1 2117
2 82430 1 2117
2 82431 1 2117
2 82432 1 2117
2 82433 1 2117
2 82434 1 2117
2 82435 1 2117
2 82436 1 2117
2 82437 1 2117
2 82438 1 2117
2 82439 1 2117
2 82440 1 2117
2 82441 1 2117
2 82442 1 2117
2 82443 1 2117
2 82444 1 2117
2 82445 1 2117
2 82446 1 2117
2 82447 1 2117
2 82448 1 2117
2 82449 1 2117
2 82450 1 2117
2 82451 1 2117
2 82452 1 2117
2 82453 1 2117
2 82454 1 2117
2 82455 1 2117
2 82456 1 2117
2 82457 1 2117
2 82458 1 2117
2 82459 1 2117
2 82460 1 2117
2 82461 1 2117
2 82462 1 2117
2 82463 1 2117
2 82464 1 2117
2 82465 1 2117
2 82466 1 2117
2 82467 1 2117
2 82468 1 2117
2 82469 1 2117
2 82470 1 2117
2 82471 1 2117
2 82472 1 2117
2 82473 1 2117
2 82474 1 2117
2 82475 1 2117
2 82476 1 2117
2 82477 1 2117
2 82478 1 2117
2 82479 1 2117
2 82480 1 2117
2 82481 1 2117
2 82482 1 2117
2 82483 1 2118
2 82484 1 2118
2 82485 1 2118
2 82486 1 2118
2 82487 1 2118
2 82488 1 2118
2 82489 1 2118
2 82490 1 2118
2 82491 1 2118
2 82492 1 2118
2 82493 1 2118
2 82494 1 2118
2 82495 1 2118
2 82496 1 2118
2 82497 1 2118
2 82498 1 2118
2 82499 1 2118
2 82500 1 2118
2 82501 1 2118
2 82502 1 2118
2 82503 1 2118
2 82504 1 2118
2 82505 1 2118
2 82506 1 2118
2 82507 1 2118
2 82508 1 2118
2 82509 1 2118
2 82510 1 2118
2 82511 1 2118
2 82512 1 2118
2 82513 1 2118
2 82514 1 2118
2 82515 1 2118
2 82516 1 2119
2 82517 1 2119
2 82518 1 2120
2 82519 1 2120
2 82520 1 2120
2 82521 1 2120
2 82522 1 2123
2 82523 1 2123
2 82524 1 2123
2 82525 1 2123
2 82526 1 2123
2 82527 1 2123
2 82528 1 2123
2 82529 1 2123
2 82530 1 2123
2 82531 1 2123
2 82532 1 2123
2 82533 1 2125
2 82534 1 2125
2 82535 1 2125
2 82536 1 2125
2 82537 1 2125
2 82538 1 2125
2 82539 1 2125
2 82540 1 2138
2 82541 1 2138
2 82542 1 2138
2 82543 1 2138
2 82544 1 2138
2 82545 1 2138
2 82546 1 2138
2 82547 1 2138
2 82548 1 2138
2 82549 1 2138
2 82550 1 2138
2 82551 1 2138
2 82552 1 2138
2 82553 1 2138
2 82554 1 2138
2 82555 1 2139
2 82556 1 2139
2 82557 1 2139
2 82558 1 2140
2 82559 1 2140
2 82560 1 2140
2 82561 1 2140
2 82562 1 2140
2 82563 1 2140
2 82564 1 2140
2 82565 1 2140
2 82566 1 2140
2 82567 1 2140
2 82568 1 2140
2 82569 1 2142
2 82570 1 2142
2 82571 1 2142
2 82572 1 2143
2 82573 1 2143
2 82574 1 2143
2 82575 1 2144
2 82576 1 2144
2 82577 1 2144
2 82578 1 2144
2 82579 1 2144
2 82580 1 2144
2 82581 1 2144
2 82582 1 2144
2 82583 1 2144
2 82584 1 2146
2 82585 1 2146
2 82586 1 2146
2 82587 1 2146
2 82588 1 2146
2 82589 1 2146
2 82590 1 2146
2 82591 1 2146
2 82592 1 2146
2 82593 1 2146
2 82594 1 2146
2 82595 1 2146
2 82596 1 2146
2 82597 1 2146
2 82598 1 2146
2 82599 1 2146
2 82600 1 2146
2 82601 1 2146
2 82602 1 2146
2 82603 1 2146
2 82604 1 2146
2 82605 1 2146
2 82606 1 2146
2 82607 1 2146
2 82608 1 2146
2 82609 1 2146
2 82610 1 2146
2 82611 1 2146
2 82612 1 2146
2 82613 1 2147
2 82614 1 2147
2 82615 1 2147
2 82616 1 2147
2 82617 1 2147
2 82618 1 2147
2 82619 1 2147
2 82620 1 2147
2 82621 1 2147
2 82622 1 2147
2 82623 1 2147
2 82624 1 2147
2 82625 1 2147
2 82626 1 2147
2 82627 1 2147
2 82628 1 2148
2 82629 1 2148
2 82630 1 2148
2 82631 1 2148
2 82632 1 2148
2 82633 1 2148
2 82634 1 2148
2 82635 1 2148
2 82636 1 2148
2 82637 1 2148
2 82638 1 2148
2 82639 1 2148
2 82640 1 2148
2 82641 1 2148
2 82642 1 2149
2 82643 1 2149
2 82644 1 2149
2 82645 1 2149
2 82646 1 2149
2 82647 1 2149
2 82648 1 2149
2 82649 1 2149
2 82650 1 2149
2 82651 1 2149
2 82652 1 2149
2 82653 1 2149
2 82654 1 2149
2 82655 1 2149
2 82656 1 2149
2 82657 1 2149
2 82658 1 2150
2 82659 1 2150
2 82660 1 2150
2 82661 1 2151
2 82662 1 2151
2 82663 1 2158
2 82664 1 2158
2 82665 1 2158
2 82666 1 2158
2 82667 1 2158
2 82668 1 2158
2 82669 1 2158
2 82670 1 2158
2 82671 1 2158
2 82672 1 2158
2 82673 1 2158
2 82674 1 2159
2 82675 1 2159
2 82676 1 2161
2 82677 1 2161
2 82678 1 2161
2 82679 1 2161
2 82680 1 2161
2 82681 1 2161
2 82682 1 2161
2 82683 1 2161
2 82684 1 2161
2 82685 1 2162
2 82686 1 2162
2 82687 1 2165
2 82688 1 2165
2 82689 1 2165
2 82690 1 2168
2 82691 1 2168
2 82692 1 2168
2 82693 1 2168
2 82694 1 2168
2 82695 1 2168
2 82696 1 2168
2 82697 1 2168
2 82698 1 2168
2 82699 1 2168
2 82700 1 2168
2 82701 1 2169
2 82702 1 2169
2 82703 1 2169
2 82704 1 2169
2 82705 1 2169
2 82706 1 2169
2 82707 1 2170
2 82708 1 2170
2 82709 1 2170
2 82710 1 2170
2 82711 1 2177
2 82712 1 2177
2 82713 1 2177
2 82714 1 2178
2 82715 1 2178
2 82716 1 2179
2 82717 1 2179
2 82718 1 2180
2 82719 1 2180
2 82720 1 2192
2 82721 1 2192
2 82722 1 2192
2 82723 1 2192
2 82724 1 2192
2 82725 1 2192
2 82726 1 2192
2 82727 1 2192
2 82728 1 2192
2 82729 1 2193
2 82730 1 2193
2 82731 1 2193
2 82732 1 2193
2 82733 1 2193
2 82734 1 2193
2 82735 1 2193
2 82736 1 2193
2 82737 1 2193
2 82738 1 2193
2 82739 1 2193
2 82740 1 2193
2 82741 1 2193
2 82742 1 2193
2 82743 1 2193
2 82744 1 2193
2 82745 1 2193
2 82746 1 2194
2 82747 1 2194
2 82748 1 2195
2 82749 1 2195
2 82750 1 2196
2 82751 1 2196
2 82752 1 2207
2 82753 1 2207
2 82754 1 2207
2 82755 1 2207
2 82756 1 2207
2 82757 1 2207
2 82758 1 2207
2 82759 1 2207
2 82760 1 2207
2 82761 1 2207
2 82762 1 2207
2 82763 1 2207
2 82764 1 2207
2 82765 1 2207
2 82766 1 2207
2 82767 1 2208
2 82768 1 2208
2 82769 1 2208
2 82770 1 2208
2 82771 1 2208
2 82772 1 2216
2 82773 1 2216
2 82774 1 2216
2 82775 1 2216
2 82776 1 2216
2 82777 1 2216
2 82778 1 2216
2 82779 1 2216
2 82780 1 2216
2 82781 1 2217
2 82782 1 2217
2 82783 1 2217
2 82784 1 2220
2 82785 1 2220
2 82786 1 2220
2 82787 1 2220
2 82788 1 2220
2 82789 1 2220
2 82790 1 2220
2 82791 1 2220
2 82792 1 2220
2 82793 1 2220
2 82794 1 2221
2 82795 1 2221
2 82796 1 2221
2 82797 1 2221
2 82798 1 2221
2 82799 1 2222
2 82800 1 2222
2 82801 1 2222
2 82802 1 2222
2 82803 1 2223
2 82804 1 2223
2 82805 1 2224
2 82806 1 2224
2 82807 1 2232
2 82808 1 2232
2 82809 1 2232
2 82810 1 2232
2 82811 1 2232
2 82812 1 2232
2 82813 1 2232
2 82814 1 2232
2 82815 1 2232
2 82816 1 2232
2 82817 1 2232
2 82818 1 2232
2 82819 1 2232
2 82820 1 2232
2 82821 1 2232
2 82822 1 2232
2 82823 1 2232
2 82824 1 2232
2 82825 1 2232
2 82826 1 2232
2 82827 1 2232
2 82828 1 2232
2 82829 1 2232
2 82830 1 2232
2 82831 1 2232
2 82832 1 2233
2 82833 1 2233
2 82834 1 2233
2 82835 1 2233
2 82836 1 2233
2 82837 1 2234
2 82838 1 2234
2 82839 1 2234
2 82840 1 2234
2 82841 1 2234
2 82842 1 2234
2 82843 1 2234
2 82844 1 2234
2 82845 1 2236
2 82846 1 2236
2 82847 1 2236
2 82848 1 2237
2 82849 1 2237
2 82850 1 2237
2 82851 1 2237
2 82852 1 2237
2 82853 1 2237
2 82854 1 2237
2 82855 1 2237
2 82856 1 2237
2 82857 1 2238
2 82858 1 2238
2 82859 1 2239
2 82860 1 2239
2 82861 1 2239
2 82862 1 2239
2 82863 1 2240
2 82864 1 2240
2 82865 1 2241
2 82866 1 2241
2 82867 1 2242
2 82868 1 2242
2 82869 1 2242
2 82870 1 2242
2 82871 1 2242
2 82872 1 2242
2 82873 1 2242
2 82874 1 2242
2 82875 1 2242
2 82876 1 2242
2 82877 1 2242
2 82878 1 2242
2 82879 1 2242
2 82880 1 2244
2 82881 1 2244
2 82882 1 2244
2 82883 1 2244
2 82884 1 2244
2 82885 1 2244
2 82886 1 2244
2 82887 1 2244
2 82888 1 2244
2 82889 1 2244
2 82890 1 2244
2 82891 1 2244
2 82892 1 2244
2 82893 1 2244
2 82894 1 2244
2 82895 1 2244
2 82896 1 2244
2 82897 1 2244
2 82898 1 2244
2 82899 1 2244
2 82900 1 2244
2 82901 1 2244
2 82902 1 2244
2 82903 1 2244
2 82904 1 2244
2 82905 1 2244
2 82906 1 2244
2 82907 1 2244
2 82908 1 2244
2 82909 1 2244
2 82910 1 2244
2 82911 1 2244
2 82912 1 2244
2 82913 1 2244
2 82914 1 2244
2 82915 1 2244
2 82916 1 2244
2 82917 1 2244
2 82918 1 2244
2 82919 1 2244
2 82920 1 2244
2 82921 1 2244
2 82922 1 2244
2 82923 1 2244
2 82924 1 2244
2 82925 1 2244
2 82926 1 2244
2 82927 1 2244
2 82928 1 2244
2 82929 1 2244
2 82930 1 2244
2 82931 1 2244
2 82932 1 2244
2 82933 1 2244
2 82934 1 2244
2 82935 1 2244
2 82936 1 2244
2 82937 1 2244
2 82938 1 2244
2 82939 1 2244
2 82940 1 2244
2 82941 1 2244
2 82942 1 2245
2 82943 1 2245
2 82944 1 2245
2 82945 1 2245
2 82946 1 2245
2 82947 1 2245
2 82948 1 2245
2 82949 1 2245
2 82950 1 2245
2 82951 1 2245
2 82952 1 2245
2 82953 1 2245
2 82954 1 2245
2 82955 1 2245
2 82956 1 2245
2 82957 1 2245
2 82958 1 2245
2 82959 1 2245
2 82960 1 2245
2 82961 1 2245
2 82962 1 2245
2 82963 1 2245
2 82964 1 2245
2 82965 1 2245
2 82966 1 2245
2 82967 1 2245
2 82968 1 2245
2 82969 1 2245
2 82970 1 2245
2 82971 1 2245
2 82972 1 2245
2 82973 1 2245
2 82974 1 2245
2 82975 1 2245
2 82976 1 2245
2 82977 1 2245
2 82978 1 2245
2 82979 1 2245
2 82980 1 2245
2 82981 1 2245
2 82982 1 2245
2 82983 1 2245
2 82984 1 2245
2 82985 1 2245
2 82986 1 2245
2 82987 1 2245
2 82988 1 2245
2 82989 1 2245
2 82990 1 2245
2 82991 1 2245
2 82992 1 2245
2 82993 1 2245
2 82994 1 2245
2 82995 1 2245
2 82996 1 2245
2 82997 1 2245
2 82998 1 2245
2 82999 1 2245
2 83000 1 2246
2 83001 1 2246
2 83002 1 2246
2 83003 1 2246
2 83004 1 2246
2 83005 1 2246
2 83006 1 2246
2 83007 1 2246
2 83008 1 2246
2 83009 1 2247
2 83010 1 2247
2 83011 1 2247
2 83012 1 2247
2 83013 1 2247
2 83014 1 2262
2 83015 1 2262
2 83016 1 2262
2 83017 1 2262
2 83018 1 2265
2 83019 1 2265
2 83020 1 2265
2 83021 1 2272
2 83022 1 2272
2 83023 1 2274
2 83024 1 2274
2 83025 1 2274
2 83026 1 2274
2 83027 1 2274
2 83028 1 2274
2 83029 1 2274
2 83030 1 2274
2 83031 1 2274
2 83032 1 2276
2 83033 1 2276
2 83034 1 2291
2 83035 1 2291
2 83036 1 2291
2 83037 1 2291
2 83038 1 2291
2 83039 1 2291
2 83040 1 2291
2 83041 1 2291
2 83042 1 2291
2 83043 1 2291
2 83044 1 2291
2 83045 1 2291
2 83046 1 2291
2 83047 1 2291
2 83048 1 2291
2 83049 1 2291
2 83050 1 2291
2 83051 1 2291
2 83052 1 2292
2 83053 1 2292
2 83054 1 2292
2 83055 1 2292
2 83056 1 2292
2 83057 1 2292
2 83058 1 2295
2 83059 1 2295
2 83060 1 2295
2 83061 1 2295
2 83062 1 2295
2 83063 1 2295
2 83064 1 2295
2 83065 1 2295
2 83066 1 2295
2 83067 1 2295
2 83068 1 2295
2 83069 1 2295
2 83070 1 2295
2 83071 1 2295
2 83072 1 2295
2 83073 1 2295
2 83074 1 2295
2 83075 1 2296
2 83076 1 2296
2 83077 1 2296
2 83078 1 2296
2 83079 1 2296
2 83080 1 2296
2 83081 1 2301
2 83082 1 2301
2 83083 1 2304
2 83084 1 2304
2 83085 1 2304
2 83086 1 2304
2 83087 1 2304
2 83088 1 2304
2 83089 1 2305
2 83090 1 2305
2 83091 1 2305
2 83092 1 2305
2 83093 1 2305
2 83094 1 2305
2 83095 1 2306
2 83096 1 2306
2 83097 1 2306
2 83098 1 2307
2 83099 1 2307
2 83100 1 2307
2 83101 1 2307
2 83102 1 2307
2 83103 1 2320
2 83104 1 2320
2 83105 1 2320
2 83106 1 2320
2 83107 1 2320
2 83108 1 2321
2 83109 1 2321
2 83110 1 2321
2 83111 1 2321
2 83112 1 2321
2 83113 1 2321
2 83114 1 2321
2 83115 1 2321
2 83116 1 2322
2 83117 1 2322
2 83118 1 2322
2 83119 1 2322
2 83120 1 2322
2 83121 1 2322
2 83122 1 2322
2 83123 1 2322
2 83124 1 2323
2 83125 1 2323
2 83126 1 2326
2 83127 1 2326
2 83128 1 2331
2 83129 1 2331
2 83130 1 2331
2 83131 1 2331
2 83132 1 2333
2 83133 1 2333
2 83134 1 2333
2 83135 1 2333
2 83136 1 2333
2 83137 1 2333
2 83138 1 2333
2 83139 1 2333
2 83140 1 2333
2 83141 1 2333
2 83142 1 2333
2 83143 1 2334
2 83144 1 2334
2 83145 1 2334
2 83146 1 2355
2 83147 1 2355
2 83148 1 2355
2 83149 1 2355
2 83150 1 2355
2 83151 1 2355
2 83152 1 2355
2 83153 1 2355
2 83154 1 2355
2 83155 1 2356
2 83156 1 2356
2 83157 1 2356
2 83158 1 2356
2 83159 1 2356
2 83160 1 2356
2 83161 1 2357
2 83162 1 2357
2 83163 1 2358
2 83164 1 2358
2 83165 1 2358
2 83166 1 2358
2 83167 1 2358
2 83168 1 2363
2 83169 1 2363
2 83170 1 2363
2 83171 1 2363
2 83172 1 2363
2 83173 1 2363
2 83174 1 2363
2 83175 1 2364
2 83176 1 2364
2 83177 1 2370
2 83178 1 2370
2 83179 1 2370
2 83180 1 2370
2 83181 1 2370
2 83182 1 2370
2 83183 1 2370
2 83184 1 2370
2 83185 1 2370
2 83186 1 2370
2 83187 1 2370
2 83188 1 2370
2 83189 1 2370
2 83190 1 2370
2 83191 1 2370
2 83192 1 2370
2 83193 1 2370
2 83194 1 2372
2 83195 1 2372
2 83196 1 2372
2 83197 1 2372
2 83198 1 2372
2 83199 1 2372
2 83200 1 2372
2 83201 1 2372
2 83202 1 2372
2 83203 1 2372
2 83204 1 2372
2 83205 1 2372
2 83206 1 2372
2 83207 1 2372
2 83208 1 2382
2 83209 1 2382
2 83210 1 2382
2 83211 1 2383
2 83212 1 2383
2 83213 1 2383
2 83214 1 2383
2 83215 1 2383
2 83216 1 2383
2 83217 1 2383
2 83218 1 2383
2 83219 1 2383
2 83220 1 2383
2 83221 1 2383
2 83222 1 2383
2 83223 1 2383
2 83224 1 2383
2 83225 1 2383
2 83226 1 2385
2 83227 1 2385
2 83228 1 2393
2 83229 1 2393
2 83230 1 2393
2 83231 1 2393
2 83232 1 2394
2 83233 1 2394
2 83234 1 2394
2 83235 1 2396
2 83236 1 2396
2 83237 1 2399
2 83238 1 2399
2 83239 1 2399
2 83240 1 2399
2 83241 1 2399
2 83242 1 2399
2 83243 1 2399
2 83244 1 2399
2 83245 1 2399
2 83246 1 2399
2 83247 1 2399
2 83248 1 2399
2 83249 1 2400
2 83250 1 2400
2 83251 1 2400
2 83252 1 2402
2 83253 1 2402
2 83254 1 2402
2 83255 1 2402
2 83256 1 2402
2 83257 1 2402
2 83258 1 2402
2 83259 1 2402
2 83260 1 2402
2 83261 1 2402
2 83262 1 2402
2 83263 1 2402
2 83264 1 2403
2 83265 1 2403
2 83266 1 2403
2 83267 1 2403
2 83268 1 2411
2 83269 1 2411
2 83270 1 2411
2 83271 1 2411
2 83272 1 2411
2 83273 1 2411
2 83274 1 2412
2 83275 1 2412
2 83276 1 2413
2 83277 1 2413
2 83278 1 2413
2 83279 1 2413
2 83280 1 2421
2 83281 1 2421
2 83282 1 2421
2 83283 1 2421
2 83284 1 2421
2 83285 1 2421
2 83286 1 2422
2 83287 1 2422
2 83288 1 2434
2 83289 1 2434
2 83290 1 2434
2 83291 1 2434
2 83292 1 2434
2 83293 1 2434
2 83294 1 2434
2 83295 1 2434
2 83296 1 2434
2 83297 1 2434
2 83298 1 2434
2 83299 1 2434
2 83300 1 2434
2 83301 1 2434
2 83302 1 2434
2 83303 1 2436
2 83304 1 2436
2 83305 1 2436
2 83306 1 2437
2 83307 1 2437
2 83308 1 2437
2 83309 1 2438
2 83310 1 2438
2 83311 1 2438
2 83312 1 2438
2 83313 1 2438
2 83314 1 2439
2 83315 1 2439
2 83316 1 2439
2 83317 1 2439
2 83318 1 2439
2 83319 1 2439
2 83320 1 2439
2 83321 1 2439
2 83322 1 2439
2 83323 1 2439
2 83324 1 2439
2 83325 1 2439
2 83326 1 2439
2 83327 1 2439
2 83328 1 2439
2 83329 1 2439
2 83330 1 2439
2 83331 1 2439
2 83332 1 2439
2 83333 1 2439
2 83334 1 2439
2 83335 1 2439
2 83336 1 2439
2 83337 1 2439
2 83338 1 2439
2 83339 1 2439
2 83340 1 2441
2 83341 1 2441
2 83342 1 2441
2 83343 1 2441
2 83344 1 2441
2 83345 1 2441
2 83346 1 2441
2 83347 1 2441
2 83348 1 2441
2 83349 1 2441
2 83350 1 2441
2 83351 1 2441
2 83352 1 2441
2 83353 1 2444
2 83354 1 2444
2 83355 1 2444
2 83356 1 2449
2 83357 1 2449
2 83358 1 2450
2 83359 1 2450
2 83360 1 2450
2 83361 1 2450
2 83362 1 2450
2 83363 1 2450
2 83364 1 2451
2 83365 1 2451
2 83366 1 2451
2 83367 1 2452
2 83368 1 2452
2 83369 1 2452
2 83370 1 2452
2 83371 1 2452
2 83372 1 2452
2 83373 1 2452
2 83374 1 2452
2 83375 1 2452
2 83376 1 2452
2 83377 1 2452
2 83378 1 2452
2 83379 1 2453
2 83380 1 2453
2 83381 1 2453
2 83382 1 2453
2 83383 1 2453
2 83384 1 2455
2 83385 1 2455
2 83386 1 2455
2 83387 1 2467
2 83388 1 2467
2 83389 1 2471
2 83390 1 2471
2 83391 1 2471
2 83392 1 2471
2 83393 1 2471
2 83394 1 2471
2 83395 1 2471
2 83396 1 2471
2 83397 1 2471
2 83398 1 2471
2 83399 1 2471
2 83400 1 2471
2 83401 1 2472
2 83402 1 2472
2 83403 1 2472
2 83404 1 2472
2 83405 1 2481
2 83406 1 2481
2 83407 1 2481
2 83408 1 2481
2 83409 1 2481
2 83410 1 2481
2 83411 1 2481
2 83412 1 2481
2 83413 1 2481
2 83414 1 2490
2 83415 1 2490
2 83416 1 2490
2 83417 1 2490
2 83418 1 2490
2 83419 1 2490
2 83420 1 2490
2 83421 1 2490
2 83422 1 2490
2 83423 1 2490
2 83424 1 2490
2 83425 1 2490
2 83426 1 2490
2 83427 1 2491
2 83428 1 2491
2 83429 1 2493
2 83430 1 2493
2 83431 1 2493
2 83432 1 2493
2 83433 1 2494
2 83434 1 2494
2 83435 1 2494
2 83436 1 2494
2 83437 1 2494
2 83438 1 2494
2 83439 1 2494
2 83440 1 2494
2 83441 1 2494
2 83442 1 2495
2 83443 1 2495
2 83444 1 2495
2 83445 1 2495
2 83446 1 2496
2 83447 1 2496
2 83448 1 2496
2 83449 1 2496
2 83450 1 2496
2 83451 1 2496
2 83452 1 2497
2 83453 1 2497
2 83454 1 2497
2 83455 1 2497
2 83456 1 2497
2 83457 1 2497
2 83458 1 2497
2 83459 1 2497
2 83460 1 2498
2 83461 1 2498
2 83462 1 2499
2 83463 1 2499
2 83464 1 2499
2 83465 1 2499
2 83466 1 2499
2 83467 1 2504
2 83468 1 2504
2 83469 1 2510
2 83470 1 2510
2 83471 1 2510
2 83472 1 2510
2 83473 1 2510
2 83474 1 2510
2 83475 1 2511
2 83476 1 2511
2 83477 1 2511
2 83478 1 2511
2 83479 1 2511
2 83480 1 2511
2 83481 1 2511
2 83482 1 2512
2 83483 1 2512
2 83484 1 2512
2 83485 1 2513
2 83486 1 2513
2 83487 1 2513
2 83488 1 2513
2 83489 1 2513
2 83490 1 2513
2 83491 1 2516
2 83492 1 2516
2 83493 1 2527
2 83494 1 2527
2 83495 1 2527
2 83496 1 2527
2 83497 1 2527
2 83498 1 2527
2 83499 1 2527
2 83500 1 2527
2 83501 1 2527
2 83502 1 2527
2 83503 1 2527
2 83504 1 2527
2 83505 1 2527
2 83506 1 2527
2 83507 1 2527
2 83508 1 2528
2 83509 1 2528
2 83510 1 2529
2 83511 1 2529
2 83512 1 2529
2 83513 1 2529
2 83514 1 2530
2 83515 1 2530
2 83516 1 2530
2 83517 1 2531
2 83518 1 2531
2 83519 1 2532
2 83520 1 2532
2 83521 1 2532
2 83522 1 2532
2 83523 1 2532
2 83524 1 2533
2 83525 1 2533
2 83526 1 2533
2 83527 1 2533
2 83528 1 2533
2 83529 1 2533
2 83530 1 2533
2 83531 1 2533
2 83532 1 2533
2 83533 1 2533
2 83534 1 2533
2 83535 1 2533
2 83536 1 2534
2 83537 1 2534
2 83538 1 2535
2 83539 1 2535
2 83540 1 2535
2 83541 1 2535
2 83542 1 2535
2 83543 1 2535
2 83544 1 2535
2 83545 1 2535
2 83546 1 2535
2 83547 1 2535
2 83548 1 2535
2 83549 1 2535
2 83550 1 2535
2 83551 1 2535
2 83552 1 2535
2 83553 1 2537
2 83554 1 2537
2 83555 1 2537
2 83556 1 2537
2 83557 1 2538
2 83558 1 2538
2 83559 1 2538
2 83560 1 2538
2 83561 1 2538
2 83562 1 2538
2 83563 1 2538
2 83564 1 2538
2 83565 1 2538
2 83566 1 2538
2 83567 1 2538
2 83568 1 2539
2 83569 1 2539
2 83570 1 2539
2 83571 1 2540
2 83572 1 2540
2 83573 1 2540
2 83574 1 2541
2 83575 1 2541
2 83576 1 2541
2 83577 1 2541
2 83578 1 2553
2 83579 1 2553
2 83580 1 2553
2 83581 1 2553
2 83582 1 2553
2 83583 1 2553
2 83584 1 2553
2 83585 1 2553
2 83586 1 2553
2 83587 1 2554
2 83588 1 2554
2 83589 1 2555
2 83590 1 2555
2 83591 1 2555
2 83592 1 2557
2 83593 1 2557
2 83594 1 2564
2 83595 1 2564
2 83596 1 2564
2 83597 1 2564
2 83598 1 2564
2 83599 1 2564
2 83600 1 2564
2 83601 1 2564
2 83602 1 2564
2 83603 1 2564
2 83604 1 2564
2 83605 1 2564
2 83606 1 2564
2 83607 1 2565
2 83608 1 2565
2 83609 1 2565
2 83610 1 2566
2 83611 1 2566
2 83612 1 2566
2 83613 1 2566
2 83614 1 2572
2 83615 1 2572
2 83616 1 2572
2 83617 1 2572
2 83618 1 2572
2 83619 1 2572
2 83620 1 2572
2 83621 1 2572
2 83622 1 2572
2 83623 1 2572
2 83624 1 2572
2 83625 1 2572
2 83626 1 2583
2 83627 1 2583
2 83628 1 2583
2 83629 1 2597
2 83630 1 2597
2 83631 1 2597
2 83632 1 2597
2 83633 1 2597
2 83634 1 2597
2 83635 1 2597
2 83636 1 2597
2 83637 1 2598
2 83638 1 2598
2 83639 1 2599
2 83640 1 2599
2 83641 1 2602
2 83642 1 2602
2 83643 1 2602
2 83644 1 2603
2 83645 1 2603
2 83646 1 2608
2 83647 1 2608
2 83648 1 2608
2 83649 1 2608
2 83650 1 2609
2 83651 1 2609
2 83652 1 2609
2 83653 1 2609
2 83654 1 2610
2 83655 1 2610
2 83656 1 2611
2 83657 1 2611
2 83658 1 2621
2 83659 1 2621
2 83660 1 2629
2 83661 1 2629
2 83662 1 2629
2 83663 1 2629
2 83664 1 2629
2 83665 1 2629
2 83666 1 2629
2 83667 1 2629
2 83668 1 2629
2 83669 1 2629
2 83670 1 2629
2 83671 1 2629
2 83672 1 2630
2 83673 1 2630
2 83674 1 2630
2 83675 1 2632
2 83676 1 2632
2 83677 1 2633
2 83678 1 2633
2 83679 1 2633
2 83680 1 2633
2 83681 1 2633
2 83682 1 2633
2 83683 1 2634
2 83684 1 2634
2 83685 1 2634
2 83686 1 2634
2 83687 1 2636
2 83688 1 2636
2 83689 1 2643
2 83690 1 2643
2 83691 1 2643
2 83692 1 2643
2 83693 1 2643
2 83694 1 2644
2 83695 1 2644
2 83696 1 2644
2 83697 1 2644
2 83698 1 2644
2 83699 1 2644
2 83700 1 2644
2 83701 1 2644
2 83702 1 2644
2 83703 1 2644
2 83704 1 2644
2 83705 1 2644
2 83706 1 2644
2 83707 1 2644
2 83708 1 2644
2 83709 1 2645
2 83710 1 2645
2 83711 1 2645
2 83712 1 2645
2 83713 1 2654
2 83714 1 2654
2 83715 1 2655
2 83716 1 2655
2 83717 1 2664
2 83718 1 2664
2 83719 1 2664
2 83720 1 2664
2 83721 1 2664
2 83722 1 2664
2 83723 1 2664
2 83724 1 2664
2 83725 1 2664
2 83726 1 2664
2 83727 1 2664
2 83728 1 2664
2 83729 1 2664
2 83730 1 2664
2 83731 1 2664
2 83732 1 2664
2 83733 1 2664
2 83734 1 2664
2 83735 1 2664
2 83736 1 2665
2 83737 1 2665
2 83738 1 2665
2 83739 1 2665
2 83740 1 2666
2 83741 1 2666
2 83742 1 2666
2 83743 1 2666
2 83744 1 2666
2 83745 1 2666
2 83746 1 2666
2 83747 1 2666
2 83748 1 2666
2 83749 1 2666
2 83750 1 2666
2 83751 1 2666
2 83752 1 2666
2 83753 1 2666
2 83754 1 2666
2 83755 1 2666
2 83756 1 2666
2 83757 1 2666
2 83758 1 2666
2 83759 1 2666
2 83760 1 2666
2 83761 1 2666
2 83762 1 2666
2 83763 1 2666
2 83764 1 2666
2 83765 1 2666
2 83766 1 2668
2 83767 1 2668
2 83768 1 2669
2 83769 1 2669
2 83770 1 2670
2 83771 1 2670
2 83772 1 2674
2 83773 1 2674
2 83774 1 2674
2 83775 1 2674
2 83776 1 2674
2 83777 1 2675
2 83778 1 2675
2 83779 1 2675
2 83780 1 2675
2 83781 1 2675
2 83782 1 2675
2 83783 1 2676
2 83784 1 2676
2 83785 1 2676
2 83786 1 2676
2 83787 1 2676
2 83788 1 2676
2 83789 1 2676
2 83790 1 2676
2 83791 1 2676
2 83792 1 2676
2 83793 1 2676
2 83794 1 2676
2 83795 1 2678
2 83796 1 2678
2 83797 1 2679
2 83798 1 2679
2 83799 1 2696
2 83800 1 2696
2 83801 1 2708
2 83802 1 2708
2 83803 1 2708
2 83804 1 2708
2 83805 1 2708
2 83806 1 2709
2 83807 1 2709
2 83808 1 2709
2 83809 1 2709
2 83810 1 2709
2 83811 1 2709
2 83812 1 2709
2 83813 1 2709
2 83814 1 2709
2 83815 1 2709
2 83816 1 2709
2 83817 1 2709
2 83818 1 2710
2 83819 1 2710
2 83820 1 2712
2 83821 1 2712
2 83822 1 2712
2 83823 1 2712
2 83824 1 2712
2 83825 1 2713
2 83826 1 2713
2 83827 1 2713
2 83828 1 2713
2 83829 1 2713
2 83830 1 2715
2 83831 1 2715
2 83832 1 2716
2 83833 1 2716
2 83834 1 2717
2 83835 1 2717
2 83836 1 2726
2 83837 1 2726
2 83838 1 2734
2 83839 1 2734
2 83840 1 2736
2 83841 1 2736
2 83842 1 2737
2 83843 1 2737
2 83844 1 2737
2 83845 1 2737
2 83846 1 2737
2 83847 1 2737
2 83848 1 2737
2 83849 1 2737
2 83850 1 2737
2 83851 1 2738
2 83852 1 2738
2 83853 1 2738
2 83854 1 2738
2 83855 1 2739
2 83856 1 2739
2 83857 1 2739
2 83858 1 2739
2 83859 1 2739
2 83860 1 2740
2 83861 1 2740
2 83862 1 2742
2 83863 1 2742
2 83864 1 2746
2 83865 1 2746
2 83866 1 2746
2 83867 1 2746
2 83868 1 2749
2 83869 1 2749
2 83870 1 2755
2 83871 1 2755
2 83872 1 2762
2 83873 1 2762
2 83874 1 2775
2 83875 1 2775
2 83876 1 2775
2 83877 1 2775
2 83878 1 2776
2 83879 1 2776
2 83880 1 2776
2 83881 1 2776
2 83882 1 2776
2 83883 1 2776
2 83884 1 2776
2 83885 1 2776
2 83886 1 2776
2 83887 1 2777
2 83888 1 2777
2 83889 1 2777
2 83890 1 2777
2 83891 1 2777
2 83892 1 2777
2 83893 1 2777
2 83894 1 2777
2 83895 1 2777
2 83896 1 2777
2 83897 1 2777
2 83898 1 2777
2 83899 1 2777
2 83900 1 2777
2 83901 1 2777
2 83902 1 2777
2 83903 1 2777
2 83904 1 2777
2 83905 1 2777
2 83906 1 2777
2 83907 1 2777
2 83908 1 2777
2 83909 1 2777
2 83910 1 2777
2 83911 1 2777
2 83912 1 2777
2 83913 1 2777
2 83914 1 2777
2 83915 1 2777
2 83916 1 2777
2 83917 1 2778
2 83918 1 2778
2 83919 1 2778
2 83920 1 2779
2 83921 1 2779
2 83922 1 2789
2 83923 1 2789
2 83924 1 2792
2 83925 1 2792
2 83926 1 2799
2 83927 1 2799
2 83928 1 2801
2 83929 1 2801
2 83930 1 2801
2 83931 1 2801
2 83932 1 2801
2 83933 1 2802
2 83934 1 2802
2 83935 1 2810
2 83936 1 2810
2 83937 1 2810
2 83938 1 2810
2 83939 1 2810
2 83940 1 2810
2 83941 1 2810
2 83942 1 2810
2 83943 1 2810
2 83944 1 2810
2 83945 1 2811
2 83946 1 2811
2 83947 1 2811
2 83948 1 2811
2 83949 1 2811
2 83950 1 2812
2 83951 1 2812
2 83952 1 2812
2 83953 1 2812
2 83954 1 2812
2 83955 1 2812
2 83956 1 2812
2 83957 1 2812
2 83958 1 2814
2 83959 1 2814
2 83960 1 2828
2 83961 1 2828
2 83962 1 2828
2 83963 1 2828
2 83964 1 2828
2 83965 1 2828
2 83966 1 2828
2 83967 1 2828
2 83968 1 2828
2 83969 1 2828
2 83970 1 2828
2 83971 1 2828
2 83972 1 2828
2 83973 1 2828
2 83974 1 2828
2 83975 1 2828
2 83976 1 2828
2 83977 1 2828
2 83978 1 2828
2 83979 1 2828
2 83980 1 2829
2 83981 1 2829
2 83982 1 2831
2 83983 1 2831
2 83984 1 2832
2 83985 1 2832
2 83986 1 2832
2 83987 1 2832
2 83988 1 2832
2 83989 1 2832
2 83990 1 2832
2 83991 1 2832
2 83992 1 2832
2 83993 1 2832
2 83994 1 2832
2 83995 1 2832
2 83996 1 2832
2 83997 1 2832
2 83998 1 2832
2 83999 1 2832
2 84000 1 2832
2 84001 1 2832
2 84002 1 2832
2 84003 1 2832
2 84004 1 2833
2 84005 1 2833
2 84006 1 2834
2 84007 1 2834
2 84008 1 2836
2 84009 1 2836
2 84010 1 2839
2 84011 1 2839
2 84012 1 2839
2 84013 1 2847
2 84014 1 2847
2 84015 1 2847
2 84016 1 2847
2 84017 1 2847
2 84018 1 2847
2 84019 1 2847
2 84020 1 2847
2 84021 1 2848
2 84022 1 2848
2 84023 1 2848
2 84024 1 2849
2 84025 1 2849
2 84026 1 2850
2 84027 1 2850
2 84028 1 2870
2 84029 1 2870
2 84030 1 2870
2 84031 1 2882
2 84032 1 2882
2 84033 1 2885
2 84034 1 2885
2 84035 1 2885
2 84036 1 2885
2 84037 1 2885
2 84038 1 2885
2 84039 1 2885
2 84040 1 2885
2 84041 1 2887
2 84042 1 2887
2 84043 1 2893
2 84044 1 2893
2 84045 1 2893
2 84046 1 2893
2 84047 1 2894
2 84048 1 2894
2 84049 1 2895
2 84050 1 2895
2 84051 1 2902
2 84052 1 2902
2 84053 1 2902
2 84054 1 2902
2 84055 1 2902
2 84056 1 2902
2 84057 1 2902
2 84058 1 2902
2 84059 1 2902
2 84060 1 2903
2 84061 1 2903
2 84062 1 2903
2 84063 1 2903
2 84064 1 2903
2 84065 1 2903
2 84066 1 2903
2 84067 1 2903
2 84068 1 2903
2 84069 1 2903
2 84070 1 2903
2 84071 1 2903
2 84072 1 2903
2 84073 1 2903
2 84074 1 2903
2 84075 1 2903
2 84076 1 2903
2 84077 1 2911
2 84078 1 2911
2 84079 1 2911
2 84080 1 2911
2 84081 1 2911
2 84082 1 2911
2 84083 1 2911
2 84084 1 2911
2 84085 1 2911
2 84086 1 2911
2 84087 1 2912
2 84088 1 2912
2 84089 1 2912
2 84090 1 2912
2 84091 1 2913
2 84092 1 2913
2 84093 1 2914
2 84094 1 2914
2 84095 1 2914
2 84096 1 2917
2 84097 1 2917
2 84098 1 2917
2 84099 1 2917
2 84100 1 2917
2 84101 1 2917
2 84102 1 2917
2 84103 1 2917
2 84104 1 2917
2 84105 1 2917
2 84106 1 2917
2 84107 1 2917
2 84108 1 2918
2 84109 1 2918
2 84110 1 2919
2 84111 1 2919
2 84112 1 2919
2 84113 1 2919
2 84114 1 2920
2 84115 1 2920
2 84116 1 2920
2 84117 1 2920
2 84118 1 2920
2 84119 1 2922
2 84120 1 2922
2 84121 1 2922
2 84122 1 2922
2 84123 1 2922
2 84124 1 2927
2 84125 1 2927
2 84126 1 2927
2 84127 1 2927
2 84128 1 2927
2 84129 1 2927
2 84130 1 2927
2 84131 1 2927
2 84132 1 2927
2 84133 1 2927
2 84134 1 2927
2 84135 1 2927
2 84136 1 2927
2 84137 1 2927
2 84138 1 2927
2 84139 1 2927
2 84140 1 2929
2 84141 1 2929
2 84142 1 2929
2 84143 1 2929
2 84144 1 2929
2 84145 1 2930
2 84146 1 2930
2 84147 1 2930
2 84148 1 2930
2 84149 1 2930
2 84150 1 2939
2 84151 1 2939
2 84152 1 2939
2 84153 1 2939
2 84154 1 2939
2 84155 1 2939
2 84156 1 2940
2 84157 1 2940
2 84158 1 2940
2 84159 1 2940
2 84160 1 2940
2 84161 1 2940
2 84162 1 2940
2 84163 1 2940
2 84164 1 2940
2 84165 1 2940
2 84166 1 2940
2 84167 1 2941
2 84168 1 2941
2 84169 1 2942
2 84170 1 2942
2 84171 1 2943
2 84172 1 2943
2 84173 1 2943
2 84174 1 2943
2 84175 1 2943
2 84176 1 2943
2 84177 1 2943
2 84178 1 2943
2 84179 1 2944
2 84180 1 2944
2 84181 1 2944
2 84182 1 2944
2 84183 1 2944
2 84184 1 2944
2 84185 1 2944
2 84186 1 2944
2 84187 1 2944
2 84188 1 2944
2 84189 1 2944
2 84190 1 2946
2 84191 1 2946
2 84192 1 2948
2 84193 1 2948
2 84194 1 2948
2 84195 1 2948
2 84196 1 2948
2 84197 1 2962
2 84198 1 2962
2 84199 1 2963
2 84200 1 2963
2 84201 1 2963
2 84202 1 2963
2 84203 1 2964
2 84204 1 2964
2 84205 1 2964
2 84206 1 2964
2 84207 1 2964
2 84208 1 2964
2 84209 1 2964
2 84210 1 2964
2 84211 1 2964
2 84212 1 2967
2 84213 1 2967
2 84214 1 2967
2 84215 1 2967
2 84216 1 2967
2 84217 1 2967
2 84218 1 2967
2 84219 1 2974
2 84220 1 2974
2 84221 1 2974
2 84222 1 2979
2 84223 1 2979
2 84224 1 2980
2 84225 1 2980
2 84226 1 2981
2 84227 1 2981
2 84228 1 2981
2 84229 1 2981
2 84230 1 2982
2 84231 1 2982
2 84232 1 2982
2 84233 1 2982
2 84234 1 2982
2 84235 1 2982
2 84236 1 2982
2 84237 1 2982
2 84238 1 2983
2 84239 1 2983
2 84240 1 2990
2 84241 1 2990
2 84242 1 2990
2 84243 1 2990
2 84244 1 2990
2 84245 1 2990
2 84246 1 2990
2 84247 1 2991
2 84248 1 2991
2 84249 1 2991
2 84250 1 2991
2 84251 1 2991
2 84252 1 2991
2 84253 1 2991
2 84254 1 2991
2 84255 1 2991
2 84256 1 2991
2 84257 1 2991
2 84258 1 2991
2 84259 1 2991
2 84260 1 2991
2 84261 1 2991
2 84262 1 2991
2 84263 1 2992
2 84264 1 2992
2 84265 1 2992
2 84266 1 2992
2 84267 1 2994
2 84268 1 2994
2 84269 1 2994
2 84270 1 2995
2 84271 1 2995
2 84272 1 2995
2 84273 1 2995
2 84274 1 2996
2 84275 1 2996
2 84276 1 2996
2 84277 1 3005
2 84278 1 3005
2 84279 1 3005
2 84280 1 3005
2 84281 1 3005
2 84282 1 3005
2 84283 1 3005
2 84284 1 3005
2 84285 1 3005
2 84286 1 3005
2 84287 1 3005
2 84288 1 3005
2 84289 1 3005
2 84290 1 3005
2 84291 1 3005
2 84292 1 3005
2 84293 1 3005
2 84294 1 3005
2 84295 1 3005
2 84296 1 3005
2 84297 1 3005
2 84298 1 3005
2 84299 1 3005
2 84300 1 3005
2 84301 1 3005
2 84302 1 3005
2 84303 1 3005
2 84304 1 3005
2 84305 1 3005
2 84306 1 3005
2 84307 1 3005
2 84308 1 3006
2 84309 1 3006
2 84310 1 3007
2 84311 1 3007
2 84312 1 3008
2 84313 1 3008
2 84314 1 3009
2 84315 1 3009
2 84316 1 3009
2 84317 1 3009
2 84318 1 3009
2 84319 1 3009
2 84320 1 3009
2 84321 1 3009
2 84322 1 3009
2 84323 1 3009
2 84324 1 3009
2 84325 1 3009
2 84326 1 3009
2 84327 1 3009
2 84328 1 3009
2 84329 1 3009
2 84330 1 3009
2 84331 1 3009
2 84332 1 3009
2 84333 1 3010
2 84334 1 3010
2 84335 1 3014
2 84336 1 3014
2 84337 1 3014
2 84338 1 3014
2 84339 1 3014
2 84340 1 3014
2 84341 1 3014
2 84342 1 3014
2 84343 1 3014
2 84344 1 3014
2 84345 1 3016
2 84346 1 3016
2 84347 1 3016
2 84348 1 3018
2 84349 1 3018
2 84350 1 3018
2 84351 1 3018
2 84352 1 3018
2 84353 1 3018
2 84354 1 3018
2 84355 1 3018
2 84356 1 3018
2 84357 1 3018
2 84358 1 3018
2 84359 1 3018
2 84360 1 3018
2 84361 1 3018
2 84362 1 3019
2 84363 1 3019
2 84364 1 3019
2 84365 1 3019
2 84366 1 3019
2 84367 1 3021
2 84368 1 3021
2 84369 1 3021
2 84370 1 3021
2 84371 1 3021
2 84372 1 3021
2 84373 1 3021
2 84374 1 3022
2 84375 1 3022
2 84376 1 3022
2 84377 1 3022
2 84378 1 3022
2 84379 1 3022
2 84380 1 3022
2 84381 1 3022
2 84382 1 3022
2 84383 1 3022
2 84384 1 3022
2 84385 1 3023
2 84386 1 3023
2 84387 1 3031
2 84388 1 3031
2 84389 1 3031
2 84390 1 3031
2 84391 1 3032
2 84392 1 3032
2 84393 1 3033
2 84394 1 3033
2 84395 1 3033
2 84396 1 3035
2 84397 1 3035
2 84398 1 3036
2 84399 1 3036
2 84400 1 3036
2 84401 1 3036
2 84402 1 3037
2 84403 1 3037
2 84404 1 3037
2 84405 1 3037
2 84406 1 3037
2 84407 1 3037
2 84408 1 3037
2 84409 1 3037
2 84410 1 3037
2 84411 1 3037
2 84412 1 3037
2 84413 1 3040
2 84414 1 3040
2 84415 1 3043
2 84416 1 3043
2 84417 1 3045
2 84418 1 3045
2 84419 1 3045
2 84420 1 3045
2 84421 1 3045
2 84422 1 3045
2 84423 1 3045
2 84424 1 3045
2 84425 1 3045
2 84426 1 3046
2 84427 1 3046
2 84428 1 3046
2 84429 1 3046
2 84430 1 3046
2 84431 1 3056
2 84432 1 3056
2 84433 1 3056
2 84434 1 3059
2 84435 1 3059
2 84436 1 3059
2 84437 1 3059
2 84438 1 3059
2 84439 1 3060
2 84440 1 3060
2 84441 1 3060
2 84442 1 3060
2 84443 1 3060
2 84444 1 3060
2 84445 1 3060
2 84446 1 3061
2 84447 1 3061
2 84448 1 3061
2 84449 1 3061
2 84450 1 3072
2 84451 1 3072
2 84452 1 3072
2 84453 1 3072
2 84454 1 3072
2 84455 1 3072
2 84456 1 3072
2 84457 1 3072
2 84458 1 3072
2 84459 1 3072
2 84460 1 3072
2 84461 1 3072
2 84462 1 3072
2 84463 1 3072
2 84464 1 3072
2 84465 1 3072
2 84466 1 3074
2 84467 1 3074
2 84468 1 3075
2 84469 1 3075
2 84470 1 3076
2 84471 1 3076
2 84472 1 3076
2 84473 1 3076
2 84474 1 3076
2 84475 1 3080
2 84476 1 3080
2 84477 1 3081
2 84478 1 3081
2 84479 1 3081
2 84480 1 3081
2 84481 1 3081
2 84482 1 3081
2 84483 1 3081
2 84484 1 3081
2 84485 1 3081
2 84486 1 3081
2 84487 1 3081
2 84488 1 3081
2 84489 1 3081
2 84490 1 3081
2 84491 1 3081
2 84492 1 3081
2 84493 1 3081
2 84494 1 3081
2 84495 1 3082
2 84496 1 3082
2 84497 1 3083
2 84498 1 3083
2 84499 1 3083
2 84500 1 3083
2 84501 1 3083
2 84502 1 3083
2 84503 1 3085
2 84504 1 3085
2 84505 1 3085
2 84506 1 3094
2 84507 1 3094
2 84508 1 3094
2 84509 1 3094
2 84510 1 3094
2 84511 1 3094
2 84512 1 3094
2 84513 1 3097
2 84514 1 3097
2 84515 1 3097
2 84516 1 3097
2 84517 1 3097
2 84518 1 3097
2 84519 1 3098
2 84520 1 3098
2 84521 1 3098
2 84522 1 3099
2 84523 1 3099
2 84524 1 3099
2 84525 1 3099
2 84526 1 3099
2 84527 1 3099
2 84528 1 3099
2 84529 1 3099
2 84530 1 3099
2 84531 1 3099
2 84532 1 3099
2 84533 1 3099
2 84534 1 3100
2 84535 1 3100
2 84536 1 3100
2 84537 1 3114
2 84538 1 3114
2 84539 1 3114
2 84540 1 3114
2 84541 1 3114
2 84542 1 3114
2 84543 1 3114
2 84544 1 3114
2 84545 1 3114
2 84546 1 3114
2 84547 1 3114
2 84548 1 3114
2 84549 1 3114
2 84550 1 3114
2 84551 1 3114
2 84552 1 3114
2 84553 1 3114
2 84554 1 3114
2 84555 1 3114
2 84556 1 3114
2 84557 1 3114
2 84558 1 3114
2 84559 1 3114
2 84560 1 3114
2 84561 1 3115
2 84562 1 3115
2 84563 1 3115
2 84564 1 3115
2 84565 1 3115
2 84566 1 3119
2 84567 1 3119
2 84568 1 3119
2 84569 1 3119
2 84570 1 3119
2 84571 1 3119
2 84572 1 3119
2 84573 1 3119
2 84574 1 3119
2 84575 1 3119
2 84576 1 3119
2 84577 1 3119
2 84578 1 3119
2 84579 1 3120
2 84580 1 3120
2 84581 1 3120
2 84582 1 3121
2 84583 1 3121
2 84584 1 3121
2 84585 1 3121
2 84586 1 3121
2 84587 1 3121
2 84588 1 3121
2 84589 1 3121
2 84590 1 3121
2 84591 1 3122
2 84592 1 3122
2 84593 1 3122
2 84594 1 3122
2 84595 1 3122
2 84596 1 3122
2 84597 1 3122
2 84598 1 3122
2 84599 1 3122
2 84600 1 3122
2 84601 1 3122
2 84602 1 3122
2 84603 1 3122
2 84604 1 3131
2 84605 1 3131
2 84606 1 3132
2 84607 1 3132
2 84608 1 3132
2 84609 1 3132
2 84610 1 3132
2 84611 1 3132
2 84612 1 3132
2 84613 1 3133
2 84614 1 3133
2 84615 1 3134
2 84616 1 3134
2 84617 1 3134
2 84618 1 3134
2 84619 1 3134
2 84620 1 3134
2 84621 1 3134
2 84622 1 3134
2 84623 1 3134
2 84624 1 3134
2 84625 1 3142
2 84626 1 3142
2 84627 1 3142
2 84628 1 3142
2 84629 1 3142
2 84630 1 3143
2 84631 1 3143
2 84632 1 3145
2 84633 1 3145
2 84634 1 3149
2 84635 1 3149
2 84636 1 3149
2 84637 1 3150
2 84638 1 3150
2 84639 1 3150
2 84640 1 3150
2 84641 1 3150
2 84642 1 3150
2 84643 1 3150
2 84644 1 3150
2 84645 1 3150
2 84646 1 3150
2 84647 1 3150
2 84648 1 3150
2 84649 1 3150
2 84650 1 3150
2 84651 1 3150
2 84652 1 3159
2 84653 1 3159
2 84654 1 3160
2 84655 1 3160
2 84656 1 3160
2 84657 1 3160
2 84658 1 3160
2 84659 1 3160
2 84660 1 3160
2 84661 1 3160
2 84662 1 3160
2 84663 1 3160
2 84664 1 3160
2 84665 1 3160
2 84666 1 3160
2 84667 1 3160
2 84668 1 3160
2 84669 1 3160
2 84670 1 3160
2 84671 1 3160
2 84672 1 3160
2 84673 1 3160
2 84674 1 3160
2 84675 1 3160
2 84676 1 3160
2 84677 1 3160
2 84678 1 3160
2 84679 1 3160
2 84680 1 3160
2 84681 1 3160
2 84682 1 3160
2 84683 1 3160
2 84684 1 3160
2 84685 1 3160
2 84686 1 3160
2 84687 1 3160
2 84688 1 3160
2 84689 1 3160
2 84690 1 3160
2 84691 1 3160
2 84692 1 3161
2 84693 1 3161
2 84694 1 3161
2 84695 1 3161
2 84696 1 3162
2 84697 1 3162
2 84698 1 3162
2 84699 1 3162
2 84700 1 3163
2 84701 1 3163
2 84702 1 3163
2 84703 1 3163
2 84704 1 3163
2 84705 1 3163
2 84706 1 3163
2 84707 1 3163
2 84708 1 3163
2 84709 1 3163
2 84710 1 3163
2 84711 1 3163
2 84712 1 3163
2 84713 1 3163
2 84714 1 3163
2 84715 1 3163
2 84716 1 3163
2 84717 1 3164
2 84718 1 3164
2 84719 1 3174
2 84720 1 3174
2 84721 1 3174
2 84722 1 3175
2 84723 1 3175
2 84724 1 3176
2 84725 1 3176
2 84726 1 3176
2 84727 1 3176
2 84728 1 3178
2 84729 1 3178
2 84730 1 3178
2 84731 1 3181
2 84732 1 3181
2 84733 1 3181
2 84734 1 3182
2 84735 1 3182
2 84736 1 3182
2 84737 1 3182
2 84738 1 3182
2 84739 1 3182
2 84740 1 3182
2 84741 1 3182
2 84742 1 3182
2 84743 1 3182
2 84744 1 3182
2 84745 1 3182
2 84746 1 3182
2 84747 1 3182
2 84748 1 3182
2 84749 1 3183
2 84750 1 3183
2 84751 1 3183
2 84752 1 3183
2 84753 1 3183
2 84754 1 3185
2 84755 1 3185
2 84756 1 3185
2 84757 1 3185
2 84758 1 3185
2 84759 1 3185
2 84760 1 3186
2 84761 1 3186
2 84762 1 3186
2 84763 1 3186
2 84764 1 3188
2 84765 1 3188
2 84766 1 3188
2 84767 1 3188
2 84768 1 3188
2 84769 1 3189
2 84770 1 3189
2 84771 1 3189
2 84772 1 3189
2 84773 1 3191
2 84774 1 3191
2 84775 1 3191
2 84776 1 3191
2 84777 1 3191
2 84778 1 3191
2 84779 1 3191
2 84780 1 3192
2 84781 1 3192
2 84782 1 3192
2 84783 1 3193
2 84784 1 3193
2 84785 1 3193
2 84786 1 3201
2 84787 1 3201
2 84788 1 3201
2 84789 1 3201
2 84790 1 3201
2 84791 1 3201
2 84792 1 3201
2 84793 1 3201
2 84794 1 3201
2 84795 1 3202
2 84796 1 3202
2 84797 1 3202
2 84798 1 3202
2 84799 1 3203
2 84800 1 3203
2 84801 1 3203
2 84802 1 3203
2 84803 1 3203
2 84804 1 3203
2 84805 1 3204
2 84806 1 3204
2 84807 1 3204
2 84808 1 3204
2 84809 1 3204
2 84810 1 3204
2 84811 1 3204
2 84812 1 3204
2 84813 1 3204
2 84814 1 3204
2 84815 1 3204
2 84816 1 3204
2 84817 1 3204
2 84818 1 3204
2 84819 1 3204
2 84820 1 3204
2 84821 1 3204
2 84822 1 3204
2 84823 1 3204
2 84824 1 3204
2 84825 1 3204
2 84826 1 3204
2 84827 1 3204
2 84828 1 3204
2 84829 1 3204
2 84830 1 3204
2 84831 1 3204
2 84832 1 3204
2 84833 1 3204
2 84834 1 3204
2 84835 1 3204
2 84836 1 3204
2 84837 1 3204
2 84838 1 3204
2 84839 1 3204
2 84840 1 3204
2 84841 1 3204
2 84842 1 3204
2 84843 1 3204
2 84844 1 3204
2 84845 1 3204
2 84846 1 3204
2 84847 1 3204
2 84848 1 3204
2 84849 1 3204
2 84850 1 3204
2 84851 1 3204
2 84852 1 3204
2 84853 1 3204
2 84854 1 3204
2 84855 1 3204
2 84856 1 3204
2 84857 1 3204
2 84858 1 3204
2 84859 1 3204
2 84860 1 3204
2 84861 1 3204
2 84862 1 3204
2 84863 1 3204
2 84864 1 3204
2 84865 1 3204
2 84866 1 3204
2 84867 1 3204
2 84868 1 3204
2 84869 1 3204
2 84870 1 3204
2 84871 1 3204
2 84872 1 3204
2 84873 1 3204
2 84874 1 3204
2 84875 1 3204
2 84876 1 3204
2 84877 1 3204
2 84878 1 3204
2 84879 1 3204
2 84880 1 3204
2 84881 1 3204
2 84882 1 3204
2 84883 1 3204
2 84884 1 3204
2 84885 1 3204
2 84886 1 3204
2 84887 1 3204
2 84888 1 3204
2 84889 1 3204
2 84890 1 3204
2 84891 1 3204
2 84892 1 3204
2 84893 1 3204
2 84894 1 3204
2 84895 1 3205
2 84896 1 3205
2 84897 1 3205
2 84898 1 3205
2 84899 1 3205
2 84900 1 3205
2 84901 1 3205
2 84902 1 3205
2 84903 1 3205
2 84904 1 3205
2 84905 1 3205
2 84906 1 3205
2 84907 1 3205
2 84908 1 3205
2 84909 1 3205
2 84910 1 3205
2 84911 1 3205
2 84912 1 3205
2 84913 1 3205
2 84914 1 3205
2 84915 1 3205
2 84916 1 3205
2 84917 1 3205
2 84918 1 3205
2 84919 1 3205
2 84920 1 3205
2 84921 1 3205
2 84922 1 3206
2 84923 1 3206
2 84924 1 3206
2 84925 1 3206
2 84926 1 3207
2 84927 1 3207
2 84928 1 3209
2 84929 1 3209
2 84930 1 3209
2 84931 1 3209
2 84932 1 3209
2 84933 1 3209
2 84934 1 3209
2 84935 1 3209
2 84936 1 3209
2 84937 1 3209
2 84938 1 3209
2 84939 1 3209
2 84940 1 3209
2 84941 1 3209
2 84942 1 3209
2 84943 1 3209
2 84944 1 3209
2 84945 1 3209
2 84946 1 3210
2 84947 1 3210
2 84948 1 3214
2 84949 1 3214
2 84950 1 3217
2 84951 1 3217
2 84952 1 3217
2 84953 1 3217
2 84954 1 3217
2 84955 1 3217
2 84956 1 3219
2 84957 1 3219
2 84958 1 3220
2 84959 1 3220
2 84960 1 3220
2 84961 1 3220
2 84962 1 3220
2 84963 1 3220
2 84964 1 3220
2 84965 1 3220
2 84966 1 3220
2 84967 1 3220
2 84968 1 3220
2 84969 1 3221
2 84970 1 3221
2 84971 1 3221
2 84972 1 3221
2 84973 1 3221
2 84974 1 3221
2 84975 1 3221
2 84976 1 3221
2 84977 1 3221
2 84978 1 3221
2 84979 1 3221
2 84980 1 3221
2 84981 1 3222
2 84982 1 3222
2 84983 1 3223
2 84984 1 3223
2 84985 1 3223
2 84986 1 3223
2 84987 1 3235
2 84988 1 3235
2 84989 1 3235
2 84990 1 3235
2 84991 1 3235
2 84992 1 3235
2 84993 1 3235
2 84994 1 3235
2 84995 1 3235
2 84996 1 3235
2 84997 1 3235
2 84998 1 3235
2 84999 1 3235
2 85000 1 3235
2 85001 1 3235
2 85002 1 3235
2 85003 1 3235
2 85004 1 3235
2 85005 1 3235
2 85006 1 3235
2 85007 1 3235
2 85008 1 3235
2 85009 1 3235
2 85010 1 3235
2 85011 1 3235
2 85012 1 3235
2 85013 1 3235
2 85014 1 3235
2 85015 1 3235
2 85016 1 3235
2 85017 1 3235
2 85018 1 3235
2 85019 1 3235
2 85020 1 3235
2 85021 1 3235
2 85022 1 3235
2 85023 1 3235
2 85024 1 3235
2 85025 1 3235
2 85026 1 3235
2 85027 1 3235
2 85028 1 3235
2 85029 1 3235
2 85030 1 3235
2 85031 1 3235
2 85032 1 3235
2 85033 1 3235
2 85034 1 3235
2 85035 1 3235
2 85036 1 3235
2 85037 1 3235
2 85038 1 3235
2 85039 1 3235
2 85040 1 3235
2 85041 1 3235
2 85042 1 3237
2 85043 1 3237
2 85044 1 3237
2 85045 1 3237
2 85046 1 3237
2 85047 1 3238
2 85048 1 3238
2 85049 1 3238
2 85050 1 3238
2 85051 1 3238
2 85052 1 3238
2 85053 1 3238
2 85054 1 3239
2 85055 1 3239
2 85056 1 3239
2 85057 1 3239
2 85058 1 3240
2 85059 1 3240
2 85060 1 3242
2 85061 1 3242
2 85062 1 3242
2 85063 1 3242
2 85064 1 3242
2 85065 1 3246
2 85066 1 3246
2 85067 1 3246
2 85068 1 3246
2 85069 1 3246
2 85070 1 3246
2 85071 1 3248
2 85072 1 3248
2 85073 1 3251
2 85074 1 3251
2 85075 1 3251
2 85076 1 3251
2 85077 1 3251
2 85078 1 3251
2 85079 1 3251
2 85080 1 3251
2 85081 1 3251
2 85082 1 3251
2 85083 1 3251
2 85084 1 3251
2 85085 1 3251
2 85086 1 3251
2 85087 1 3251
2 85088 1 3251
2 85089 1 3251
2 85090 1 3252
2 85091 1 3252
2 85092 1 3252
2 85093 1 3252
2 85094 1 3252
2 85095 1 3254
2 85096 1 3254
2 85097 1 3257
2 85098 1 3257
2 85099 1 3257
2 85100 1 3257
2 85101 1 3257
2 85102 1 3257
2 85103 1 3257
2 85104 1 3257
2 85105 1 3257
2 85106 1 3257
2 85107 1 3257
2 85108 1 3257
2 85109 1 3257
2 85110 1 3257
2 85111 1 3258
2 85112 1 3258
2 85113 1 3258
2 85114 1 3258
2 85115 1 3258
2 85116 1 3258
2 85117 1 3258
2 85118 1 3258
2 85119 1 3258
2 85120 1 3258
2 85121 1 3258
2 85122 1 3258
2 85123 1 3258
2 85124 1 3258
2 85125 1 3258
2 85126 1 3258
2 85127 1 3258
2 85128 1 3258
2 85129 1 3258
2 85130 1 3258
2 85131 1 3258
2 85132 1 3258
2 85133 1 3258
2 85134 1 3258
2 85135 1 3258
2 85136 1 3258
2 85137 1 3258
2 85138 1 3258
2 85139 1 3258
2 85140 1 3258
2 85141 1 3258
2 85142 1 3258
2 85143 1 3258
2 85144 1 3258
2 85145 1 3258
2 85146 1 3258
2 85147 1 3258
2 85148 1 3258
2 85149 1 3258
2 85150 1 3258
2 85151 1 3258
2 85152 1 3258
2 85153 1 3258
2 85154 1 3258
2 85155 1 3258
2 85156 1 3258
2 85157 1 3258
2 85158 1 3258
2 85159 1 3258
2 85160 1 3258
2 85161 1 3258
2 85162 1 3258
2 85163 1 3258
2 85164 1 3258
2 85165 1 3258
2 85166 1 3258
2 85167 1 3258
2 85168 1 3258
2 85169 1 3258
2 85170 1 3258
2 85171 1 3258
2 85172 1 3258
2 85173 1 3258
2 85174 1 3258
2 85175 1 3258
2 85176 1 3258
2 85177 1 3258
2 85178 1 3258
2 85179 1 3258
2 85180 1 3258
2 85181 1 3259
2 85182 1 3259
2 85183 1 3259
2 85184 1 3260
2 85185 1 3260
2 85186 1 3261
2 85187 1 3261
2 85188 1 3261
2 85189 1 3265
2 85190 1 3265
2 85191 1 3265
2 85192 1 3265
2 85193 1 3273
2 85194 1 3273
2 85195 1 3273
2 85196 1 3273
2 85197 1 3273
2 85198 1 3273
2 85199 1 3273
2 85200 1 3273
2 85201 1 3273
2 85202 1 3273
2 85203 1 3273
2 85204 1 3273
2 85205 1 3273
2 85206 1 3273
2 85207 1 3273
2 85208 1 3273
2 85209 1 3273
2 85210 1 3273
2 85211 1 3273
2 85212 1 3273
2 85213 1 3273
2 85214 1 3273
2 85215 1 3273
2 85216 1 3273
2 85217 1 3273
2 85218 1 3273
2 85219 1 3273
2 85220 1 3273
2 85221 1 3273
2 85222 1 3273
2 85223 1 3273
2 85224 1 3273
2 85225 1 3273
2 85226 1 3273
2 85227 1 3273
2 85228 1 3273
2 85229 1 3273
2 85230 1 3273
2 85231 1 3273
2 85232 1 3273
2 85233 1 3273
2 85234 1 3273
2 85235 1 3273
2 85236 1 3273
2 85237 1 3273
2 85238 1 3273
2 85239 1 3273
2 85240 1 3273
2 85241 1 3273
2 85242 1 3273
2 85243 1 3273
2 85244 1 3273
2 85245 1 3273
2 85246 1 3273
2 85247 1 3273
2 85248 1 3273
2 85249 1 3273
2 85250 1 3273
2 85251 1 3273
2 85252 1 3273
2 85253 1 3273
2 85254 1 3273
2 85255 1 3273
2 85256 1 3273
2 85257 1 3273
2 85258 1 3273
2 85259 1 3273
2 85260 1 3273
2 85261 1 3273
2 85262 1 3273
2 85263 1 3273
2 85264 1 3273
2 85265 1 3273
2 85266 1 3273
2 85267 1 3273
2 85268 1 3273
2 85269 1 3273
2 85270 1 3273
2 85271 1 3273
2 85272 1 3273
2 85273 1 3273
2 85274 1 3273
2 85275 1 3273
2 85276 1 3273
2 85277 1 3273
2 85278 1 3273
2 85279 1 3273
2 85280 1 3273
2 85281 1 3273
2 85282 1 3273
2 85283 1 3273
2 85284 1 3273
2 85285 1 3273
2 85286 1 3273
2 85287 1 3273
2 85288 1 3273
2 85289 1 3273
2 85290 1 3273
2 85291 1 3273
2 85292 1 3273
2 85293 1 3273
2 85294 1 3273
2 85295 1 3273
2 85296 1 3273
2 85297 1 3273
2 85298 1 3273
2 85299 1 3273
2 85300 1 3273
2 85301 1 3273
2 85302 1 3273
2 85303 1 3273
2 85304 1 3273
2 85305 1 3273
2 85306 1 3273
2 85307 1 3273
2 85308 1 3273
2 85309 1 3273
2 85310 1 3273
2 85311 1 3273
2 85312 1 3273
2 85313 1 3273
2 85314 1 3273
2 85315 1 3273
2 85316 1 3273
2 85317 1 3273
2 85318 1 3273
2 85319 1 3273
2 85320 1 3273
2 85321 1 3273
2 85322 1 3273
2 85323 1 3273
2 85324 1 3273
2 85325 1 3273
2 85326 1 3273
2 85327 1 3273
2 85328 1 3273
2 85329 1 3273
2 85330 1 3273
2 85331 1 3273
2 85332 1 3273
2 85333 1 3273
2 85334 1 3273
2 85335 1 3273
2 85336 1 3273
2 85337 1 3273
2 85338 1 3273
2 85339 1 3273
2 85340 1 3273
2 85341 1 3273
2 85342 1 3273
2 85343 1 3273
2 85344 1 3273
2 85345 1 3273
2 85346 1 3273
2 85347 1 3273
2 85348 1 3273
2 85349 1 3273
2 85350 1 3273
2 85351 1 3273
2 85352 1 3273
2 85353 1 3274
2 85354 1 3274
2 85355 1 3274
2 85356 1 3274
2 85357 1 3274
2 85358 1 3274
2 85359 1 3274
2 85360 1 3274
2 85361 1 3274
2 85362 1 3274
2 85363 1 3274
2 85364 1 3274
2 85365 1 3274
2 85366 1 3276
2 85367 1 3276
2 85368 1 3276
2 85369 1 3276
2 85370 1 3276
2 85371 1 3284
2 85372 1 3284
2 85373 1 3284
2 85374 1 3284
2 85375 1 3285
2 85376 1 3285
2 85377 1 3285
2 85378 1 3285
2 85379 1 3285
2 85380 1 3286
2 85381 1 3286
2 85382 1 3286
2 85383 1 3286
2 85384 1 3287
2 85385 1 3287
2 85386 1 3290
2 85387 1 3290
2 85388 1 3290
2 85389 1 3290
2 85390 1 3292
2 85391 1 3292
2 85392 1 3292
2 85393 1 3293
2 85394 1 3293
2 85395 1 3301
2 85396 1 3301
2 85397 1 3301
2 85398 1 3303
2 85399 1 3303
2 85400 1 3316
2 85401 1 3316
2 85402 1 3316
2 85403 1 3316
2 85404 1 3316
2 85405 1 3316
2 85406 1 3316
2 85407 1 3317
2 85408 1 3317
2 85409 1 3323
2 85410 1 3323
2 85411 1 3323
2 85412 1 3323
2 85413 1 3323
2 85414 1 3332
2 85415 1 3332
2 85416 1 3332
2 85417 1 3332
2 85418 1 3332
2 85419 1 3332
2 85420 1 3332
2 85421 1 3332
2 85422 1 3333
2 85423 1 3333
2 85424 1 3333
2 85425 1 3334
2 85426 1 3334
2 85427 1 3334
2 85428 1 3334
2 85429 1 3334
2 85430 1 3355
2 85431 1 3355
2 85432 1 3355
2 85433 1 3355
2 85434 1 3355
2 85435 1 3355
2 85436 1 3355
2 85437 1 3355
2 85438 1 3355
2 85439 1 3355
2 85440 1 3355
2 85441 1 3355
2 85442 1 3355
2 85443 1 3355
2 85444 1 3355
2 85445 1 3355
2 85446 1 3357
2 85447 1 3357
2 85448 1 3357
2 85449 1 3357
2 85450 1 3357
2 85451 1 3357
2 85452 1 3357
2 85453 1 3357
2 85454 1 3357
2 85455 1 3357
2 85456 1 3357
2 85457 1 3357
2 85458 1 3357
2 85459 1 3357
2 85460 1 3357
2 85461 1 3357
2 85462 1 3357
2 85463 1 3357
2 85464 1 3357
2 85465 1 3357
2 85466 1 3357
2 85467 1 3357
2 85468 1 3357
2 85469 1 3357
2 85470 1 3357
2 85471 1 3357
2 85472 1 3357
2 85473 1 3357
2 85474 1 3359
2 85475 1 3359
2 85476 1 3359
2 85477 1 3359
2 85478 1 3359
2 85479 1 3359
2 85480 1 3360
2 85481 1 3360
2 85482 1 3360
2 85483 1 3360
2 85484 1 3360
2 85485 1 3360
2 85486 1 3360
2 85487 1 3360
2 85488 1 3360
2 85489 1 3360
2 85490 1 3360
2 85491 1 3360
2 85492 1 3360
2 85493 1 3360
2 85494 1 3360
2 85495 1 3360
2 85496 1 3360
2 85497 1 3360
2 85498 1 3360
2 85499 1 3360
2 85500 1 3360
2 85501 1 3360
2 85502 1 3360
2 85503 1 3360
2 85504 1 3360
2 85505 1 3360
2 85506 1 3360
2 85507 1 3360
2 85508 1 3360
2 85509 1 3360
2 85510 1 3360
2 85511 1 3360
2 85512 1 3360
2 85513 1 3360
2 85514 1 3360
2 85515 1 3360
2 85516 1 3360
2 85517 1 3360
2 85518 1 3360
2 85519 1 3360
2 85520 1 3360
2 85521 1 3360
2 85522 1 3360
2 85523 1 3360
2 85524 1 3360
2 85525 1 3360
2 85526 1 3360
2 85527 1 3360
2 85528 1 3360
2 85529 1 3360
2 85530 1 3360
2 85531 1 3360
2 85532 1 3360
2 85533 1 3360
2 85534 1 3360
2 85535 1 3360
2 85536 1 3360
2 85537 1 3360
2 85538 1 3360
2 85539 1 3360
2 85540 1 3360
2 85541 1 3360
2 85542 1 3360
2 85543 1 3360
2 85544 1 3360
2 85545 1 3360
2 85546 1 3360
2 85547 1 3360
2 85548 1 3360
2 85549 1 3360
2 85550 1 3360
2 85551 1 3360
2 85552 1 3360
2 85553 1 3360
2 85554 1 3360
2 85555 1 3360
2 85556 1 3360
2 85557 1 3360
2 85558 1 3360
2 85559 1 3360
2 85560 1 3360
2 85561 1 3360
2 85562 1 3360
2 85563 1 3360
2 85564 1 3360
2 85565 1 3360
2 85566 1 3360
2 85567 1 3361
2 85568 1 3361
2 85569 1 3361
2 85570 1 3361
2 85571 1 3361
2 85572 1 3361
2 85573 1 3361
2 85574 1 3361
2 85575 1 3361
2 85576 1 3363
2 85577 1 3363
2 85578 1 3363
2 85579 1 3363
2 85580 1 3363
2 85581 1 3363
2 85582 1 3363
2 85583 1 3363
2 85584 1 3363
2 85585 1 3363
2 85586 1 3364
2 85587 1 3364
2 85588 1 3364
2 85589 1 3365
2 85590 1 3365
2 85591 1 3372
2 85592 1 3372
2 85593 1 3372
2 85594 1 3372
2 85595 1 3373
2 85596 1 3373
2 85597 1 3373
2 85598 1 3373
2 85599 1 3373
2 85600 1 3376
2 85601 1 3376
2 85602 1 3377
2 85603 1 3377
2 85604 1 3378
2 85605 1 3378
2 85606 1 3381
2 85607 1 3381
2 85608 1 3389
2 85609 1 3389
2 85610 1 3389
2 85611 1 3389
2 85612 1 3389
2 85613 1 3389
2 85614 1 3389
2 85615 1 3389
2 85616 1 3389
2 85617 1 3389
2 85618 1 3389
2 85619 1 3390
2 85620 1 3390
2 85621 1 3390
2 85622 1 3390
2 85623 1 3390
2 85624 1 3390
2 85625 1 3390
2 85626 1 3390
2 85627 1 3390
2 85628 1 3390
2 85629 1 3390
2 85630 1 3390
2 85631 1 3390
2 85632 1 3390
2 85633 1 3390
2 85634 1 3390
2 85635 1 3390
2 85636 1 3390
2 85637 1 3390
2 85638 1 3390
2 85639 1 3390
2 85640 1 3390
2 85641 1 3390
2 85642 1 3390
2 85643 1 3390
2 85644 1 3390
2 85645 1 3391
2 85646 1 3391
2 85647 1 3391
2 85648 1 3391
2 85649 1 3391
2 85650 1 3391
2 85651 1 3391
2 85652 1 3391
2 85653 1 3391
2 85654 1 3391
2 85655 1 3391
2 85656 1 3391
2 85657 1 3391
2 85658 1 3391
2 85659 1 3392
2 85660 1 3392
2 85661 1 3392
2 85662 1 3392
2 85663 1 3392
2 85664 1 3392
2 85665 1 3392
2 85666 1 3392
2 85667 1 3392
2 85668 1 3392
2 85669 1 3392
2 85670 1 3392
2 85671 1 3392
2 85672 1 3392
2 85673 1 3392
2 85674 1 3392
2 85675 1 3392
2 85676 1 3392
2 85677 1 3392
2 85678 1 3392
2 85679 1 3392
2 85680 1 3392
2 85681 1 3392
2 85682 1 3392
2 85683 1 3392
2 85684 1 3392
2 85685 1 3392
2 85686 1 3392
2 85687 1 3392
2 85688 1 3392
2 85689 1 3392
2 85690 1 3392
2 85691 1 3392
2 85692 1 3392
2 85693 1 3392
2 85694 1 3392
2 85695 1 3392
2 85696 1 3392
2 85697 1 3392
2 85698 1 3392
2 85699 1 3392
2 85700 1 3392
2 85701 1 3392
2 85702 1 3392
2 85703 1 3392
2 85704 1 3392
2 85705 1 3392
2 85706 1 3392
2 85707 1 3392
2 85708 1 3392
2 85709 1 3392
2 85710 1 3392
2 85711 1 3392
2 85712 1 3392
2 85713 1 3392
2 85714 1 3392
2 85715 1 3392
2 85716 1 3392
2 85717 1 3392
2 85718 1 3392
2 85719 1 3393
2 85720 1 3393
2 85721 1 3393
2 85722 1 3393
2 85723 1 3394
2 85724 1 3394
2 85725 1 3395
2 85726 1 3395
2 85727 1 3396
2 85728 1 3396
2 85729 1 3399
2 85730 1 3399
2 85731 1 3403
2 85732 1 3403
2 85733 1 3403
2 85734 1 3403
2 85735 1 3403
2 85736 1 3403
2 85737 1 3403
2 85738 1 3403
2 85739 1 3403
2 85740 1 3403
2 85741 1 3403
2 85742 1 3403
2 85743 1 3403
2 85744 1 3403
2 85745 1 3403
2 85746 1 3403
2 85747 1 3403
2 85748 1 3403
2 85749 1 3403
2 85750 1 3403
2 85751 1 3403
2 85752 1 3403
2 85753 1 3404
2 85754 1 3404
2 85755 1 3404
2 85756 1 3404
2 85757 1 3404
2 85758 1 3406
2 85759 1 3406
2 85760 1 3406
2 85761 1 3406
2 85762 1 3407
2 85763 1 3407
2 85764 1 3407
2 85765 1 3407
2 85766 1 3407
2 85767 1 3407
2 85768 1 3407
2 85769 1 3408
2 85770 1 3408
2 85771 1 3408
2 85772 1 3409
2 85773 1 3409
2 85774 1 3409
2 85775 1 3414
2 85776 1 3414
2 85777 1 3414
2 85778 1 3417
2 85779 1 3417
2 85780 1 3417
2 85781 1 3419
2 85782 1 3419
2 85783 1 3421
2 85784 1 3421
2 85785 1 3424
2 85786 1 3424
2 85787 1 3424
2 85788 1 3424
2 85789 1 3424
2 85790 1 3424
2 85791 1 3425
2 85792 1 3425
2 85793 1 3425
2 85794 1 3426
2 85795 1 3426
2 85796 1 3427
2 85797 1 3427
2 85798 1 3432
2 85799 1 3432
2 85800 1 3432
2 85801 1 3433
2 85802 1 3433
2 85803 1 3436
2 85804 1 3436
2 85805 1 3446
2 85806 1 3446
2 85807 1 3446
2 85808 1 3446
2 85809 1 3446
2 85810 1 3447
2 85811 1 3447
2 85812 1 3447
2 85813 1 3447
2 85814 1 3449
2 85815 1 3449
2 85816 1 3455
2 85817 1 3455
2 85818 1 3467
2 85819 1 3467
2 85820 1 3467
2 85821 1 3467
2 85822 1 3467
2 85823 1 3467
2 85824 1 3467
2 85825 1 3470
2 85826 1 3470
2 85827 1 3470
2 85828 1 3470
2 85829 1 3470
2 85830 1 3470
2 85831 1 3470
2 85832 1 3477
2 85833 1 3477
2 85834 1 3477
2 85835 1 3477
2 85836 1 3489
2 85837 1 3489
2 85838 1 3489
2 85839 1 3495
2 85840 1 3495
2 85841 1 3505
2 85842 1 3505
2 85843 1 3505
2 85844 1 3505
2 85845 1 3505
2 85846 1 3505
2 85847 1 3505
2 85848 1 3505
2 85849 1 3508
2 85850 1 3508
2 85851 1 3508
2 85852 1 3508
2 85853 1 3508
2 85854 1 3508
2 85855 1 3508
2 85856 1 3508
2 85857 1 3508
2 85858 1 3508
2 85859 1 3508
2 85860 1 3508
2 85861 1 3508
2 85862 1 3508
2 85863 1 3508
2 85864 1 3508
2 85865 1 3508
2 85866 1 3508
2 85867 1 3508
2 85868 1 3508
2 85869 1 3508
2 85870 1 3508
2 85871 1 3508
2 85872 1 3508
2 85873 1 3508
2 85874 1 3508
2 85875 1 3508
2 85876 1 3508
2 85877 1 3508
2 85878 1 3508
2 85879 1 3508
2 85880 1 3508
2 85881 1 3508
2 85882 1 3508
2 85883 1 3508
2 85884 1 3508
2 85885 1 3508
2 85886 1 3508
2 85887 1 3508
2 85888 1 3508
2 85889 1 3508
2 85890 1 3508
2 85891 1 3508
2 85892 1 3508
2 85893 1 3508
2 85894 1 3508
2 85895 1 3508
2 85896 1 3508
2 85897 1 3508
2 85898 1 3508
2 85899 1 3508
2 85900 1 3508
2 85901 1 3508
2 85902 1 3508
2 85903 1 3508
2 85904 1 3508
2 85905 1 3508
2 85906 1 3508
2 85907 1 3508
2 85908 1 3508
2 85909 1 3508
2 85910 1 3508
2 85911 1 3508
2 85912 1 3508
2 85913 1 3508
2 85914 1 3508
2 85915 1 3508
2 85916 1 3508
2 85917 1 3508
2 85918 1 3508
2 85919 1 3508
2 85920 1 3508
2 85921 1 3508
2 85922 1 3508
2 85923 1 3508
2 85924 1 3508
2 85925 1 3508
2 85926 1 3508
2 85927 1 3508
2 85928 1 3508
2 85929 1 3508
2 85930 1 3508
2 85931 1 3508
2 85932 1 3508
2 85933 1 3508
2 85934 1 3508
2 85935 1 3508
2 85936 1 3508
2 85937 1 3508
2 85938 1 3508
2 85939 1 3508
2 85940 1 3508
2 85941 1 3508
2 85942 1 3508
2 85943 1 3508
2 85944 1 3508
2 85945 1 3508
2 85946 1 3508
2 85947 1 3508
2 85948 1 3508
2 85949 1 3508
2 85950 1 3508
2 85951 1 3508
2 85952 1 3508
2 85953 1 3508
2 85954 1 3508
2 85955 1 3508
2 85956 1 3508
2 85957 1 3508
2 85958 1 3508
2 85959 1 3508
2 85960 1 3508
2 85961 1 3508
2 85962 1 3508
2 85963 1 3508
2 85964 1 3508
2 85965 1 3508
2 85966 1 3508
2 85967 1 3508
2 85968 1 3508
2 85969 1 3508
2 85970 1 3523
2 85971 1 3523
2 85972 1 3523
2 85973 1 3533
2 85974 1 3533
2 85975 1 3549
2 85976 1 3549
2 85977 1 3549
2 85978 1 3549
2 85979 1 3549
2 85980 1 3549
2 85981 1 3549
2 85982 1 3549
2 85983 1 3551
2 85984 1 3551
2 85985 1 3551
2 85986 1 3551
2 85987 1 3551
2 85988 1 3551
2 85989 1 3551
2 85990 1 3551
2 85991 1 3552
2 85992 1 3552
2 85993 1 3558
2 85994 1 3558
2 85995 1 3558
2 85996 1 3559
2 85997 1 3559
2 85998 1 3560
2 85999 1 3560
2 86000 1 3560
2 86001 1 3560
2 86002 1 3560
2 86003 1 3560
2 86004 1 3560
2 86005 1 3560
2 86006 1 3560
2 86007 1 3560
2 86008 1 3562
2 86009 1 3562
2 86010 1 3562
2 86011 1 3562
2 86012 1 3580
2 86013 1 3580
2 86014 1 3587
2 86015 1 3587
2 86016 1 3588
2 86017 1 3588
2 86018 1 3598
2 86019 1 3598
2 86020 1 3599
2 86021 1 3599
2 86022 1 3599
2 86023 1 3599
2 86024 1 3599
2 86025 1 3599
2 86026 1 3599
2 86027 1 3599
2 86028 1 3599
2 86029 1 3600
2 86030 1 3600
2 86031 1 3600
2 86032 1 3600
2 86033 1 3600
2 86034 1 3600
2 86035 1 3600
2 86036 1 3600
2 86037 1 3600
2 86038 1 3601
2 86039 1 3601
2 86040 1 3601
2 86041 1 3601
2 86042 1 3601
2 86043 1 3601
2 86044 1 3601
2 86045 1 3601
2 86046 1 3601
2 86047 1 3601
2 86048 1 3601
2 86049 1 3601
2 86050 1 3601
2 86051 1 3601
2 86052 1 3601
2 86053 1 3601
2 86054 1 3601
2 86055 1 3601
2 86056 1 3601
2 86057 1 3601
2 86058 1 3601
2 86059 1 3601
2 86060 1 3601
2 86061 1 3601
2 86062 1 3601
2 86063 1 3601
2 86064 1 3601
2 86065 1 3601
2 86066 1 3601
2 86067 1 3601
2 86068 1 3601
2 86069 1 3601
2 86070 1 3601
2 86071 1 3601
2 86072 1 3601
2 86073 1 3601
2 86074 1 3601
2 86075 1 3601
2 86076 1 3601
2 86077 1 3601
2 86078 1 3601
2 86079 1 3601
2 86080 1 3602
2 86081 1 3602
2 86082 1 3602
2 86083 1 3610
2 86084 1 3610
2 86085 1 3610
2 86086 1 3611
2 86087 1 3611
2 86088 1 3611
2 86089 1 3611
2 86090 1 3611
2 86091 1 3611
2 86092 1 3611
2 86093 1 3613
2 86094 1 3613
2 86095 1 3613
2 86096 1 3613
2 86097 1 3613
2 86098 1 3614
2 86099 1 3614
2 86100 1 3614
2 86101 1 3614
2 86102 1 3614
2 86103 1 3615
2 86104 1 3615
2 86105 1 3615
2 86106 1 3615
2 86107 1 3615
2 86108 1 3623
2 86109 1 3623
2 86110 1 3623
2 86111 1 3623
2 86112 1 3624
2 86113 1 3624
2 86114 1 3624
2 86115 1 3625
2 86116 1 3625
2 86117 1 3625
2 86118 1 3625
2 86119 1 3625
2 86120 1 3626
2 86121 1 3626
2 86122 1 3627
2 86123 1 3627
2 86124 1 3628
2 86125 1 3628
2 86126 1 3628
2 86127 1 3636
2 86128 1 3636
2 86129 1 3643
2 86130 1 3643
2 86131 1 3643
2 86132 1 3643
2 86133 1 3643
2 86134 1 3643
2 86135 1 3643
2 86136 1 3643
2 86137 1 3643
2 86138 1 3643
2 86139 1 3643
2 86140 1 3643
2 86141 1 3643
2 86142 1 3643
2 86143 1 3644
2 86144 1 3644
2 86145 1 3644
2 86146 1 3645
2 86147 1 3645
2 86148 1 3645
2 86149 1 3645
2 86150 1 3646
2 86151 1 3646
2 86152 1 3647
2 86153 1 3647
2 86154 1 3648
2 86155 1 3648
2 86156 1 3648
2 86157 1 3650
2 86158 1 3650
2 86159 1 3651
2 86160 1 3651
2 86161 1 3651
2 86162 1 3651
2 86163 1 3654
2 86164 1 3654
2 86165 1 3658
2 86166 1 3658
2 86167 1 3659
2 86168 1 3659
2 86169 1 3659
2 86170 1 3659
2 86171 1 3661
2 86172 1 3661
2 86173 1 3661
2 86174 1 3661
2 86175 1 3662
2 86176 1 3662
2 86177 1 3662
2 86178 1 3662
2 86179 1 3665
2 86180 1 3665
2 86181 1 3666
2 86182 1 3666
2 86183 1 3671
2 86184 1 3671
2 86185 1 3671
2 86186 1 3672
2 86187 1 3672
2 86188 1 3673
2 86189 1 3673
2 86190 1 3673
2 86191 1 3674
2 86192 1 3674
2 86193 1 3674
2 86194 1 3687
2 86195 1 3687
2 86196 1 3687
2 86197 1 3687
2 86198 1 3687
2 86199 1 3687
2 86200 1 3687
2 86201 1 3687
2 86202 1 3697
2 86203 1 3697
2 86204 1 3697
2 86205 1 3698
2 86206 1 3698
2 86207 1 3698
2 86208 1 3698
2 86209 1 3698
2 86210 1 3698
2 86211 1 3698
2 86212 1 3698
2 86213 1 3698
2 86214 1 3698
2 86215 1 3698
2 86216 1 3698
2 86217 1 3698
2 86218 1 3698
2 86219 1 3698
2 86220 1 3698
2 86221 1 3698
2 86222 1 3698
2 86223 1 3698
2 86224 1 3698
2 86225 1 3698
2 86226 1 3699
2 86227 1 3699
2 86228 1 3699
2 86229 1 3699
2 86230 1 3699
2 86231 1 3699
2 86232 1 3700
2 86233 1 3700
2 86234 1 3701
2 86235 1 3701
2 86236 1 3702
2 86237 1 3702
2 86238 1 3702
2 86239 1 3702
2 86240 1 3712
2 86241 1 3712
2 86242 1 3720
2 86243 1 3720
2 86244 1 3720
2 86245 1 3720
2 86246 1 3720
2 86247 1 3728
2 86248 1 3728
2 86249 1 3728
2 86250 1 3728
2 86251 1 3728
2 86252 1 3728
2 86253 1 3728
2 86254 1 3728
2 86255 1 3728
2 86256 1 3728
2 86257 1 3728
2 86258 1 3728
2 86259 1 3729
2 86260 1 3729
2 86261 1 3729
2 86262 1 3729
2 86263 1 3729
2 86264 1 3729
2 86265 1 3729
2 86266 1 3729
2 86267 1 3729
2 86268 1 3729
2 86269 1 3729
2 86270 1 3729
2 86271 1 3729
2 86272 1 3729
2 86273 1 3729
2 86274 1 3729
2 86275 1 3729
2 86276 1 3729
2 86277 1 3729
2 86278 1 3729
2 86279 1 3729
2 86280 1 3731
2 86281 1 3731
2 86282 1 3736
2 86283 1 3736
2 86284 1 3737
2 86285 1 3737
2 86286 1 3737
2 86287 1 3739
2 86288 1 3739
2 86289 1 3741
2 86290 1 3741
2 86291 1 3744
2 86292 1 3744
2 86293 1 3744
2 86294 1 3744
2 86295 1 3746
2 86296 1 3746
2 86297 1 3746
2 86298 1 3747
2 86299 1 3747
2 86300 1 3747
2 86301 1 3747
2 86302 1 3747
2 86303 1 3747
2 86304 1 3747
2 86305 1 3747
2 86306 1 3748
2 86307 1 3748
2 86308 1 3748
2 86309 1 3748
2 86310 1 3749
2 86311 1 3749
2 86312 1 3753
2 86313 1 3753
2 86314 1 3754
2 86315 1 3754
2 86316 1 3755
2 86317 1 3755
2 86318 1 3760
2 86319 1 3760
2 86320 1 3760
2 86321 1 3760
2 86322 1 3760
2 86323 1 3760
2 86324 1 3761
2 86325 1 3761
2 86326 1 3761
2 86327 1 3761
2 86328 1 3761
2 86329 1 3761
2 86330 1 3762
2 86331 1 3762
2 86332 1 3763
2 86333 1 3763
2 86334 1 3763
2 86335 1 3763
2 86336 1 3763
2 86337 1 3763
2 86338 1 3763
2 86339 1 3763
2 86340 1 3763
2 86341 1 3763
2 86342 1 3763
2 86343 1 3763
2 86344 1 3763
2 86345 1 3763
2 86346 1 3763
2 86347 1 3763
2 86348 1 3763
2 86349 1 3763
2 86350 1 3763
2 86351 1 3763
2 86352 1 3763
2 86353 1 3763
2 86354 1 3763
2 86355 1 3763
2 86356 1 3763
2 86357 1 3764
2 86358 1 3764
2 86359 1 3764
2 86360 1 3764
2 86361 1 3764
2 86362 1 3764
2 86363 1 3764
2 86364 1 3764
2 86365 1 3764
2 86366 1 3764
2 86367 1 3764
2 86368 1 3764
2 86369 1 3764
2 86370 1 3764
2 86371 1 3764
2 86372 1 3764
2 86373 1 3765
2 86374 1 3765
2 86375 1 3765
2 86376 1 3771
2 86377 1 3771
2 86378 1 3771
2 86379 1 3771
2 86380 1 3771
2 86381 1 3771
2 86382 1 3772
2 86383 1 3772
2 86384 1 3772
2 86385 1 3782
2 86386 1 3782
2 86387 1 3783
2 86388 1 3783
2 86389 1 3783
2 86390 1 3783
2 86391 1 3783
2 86392 1 3792
2 86393 1 3792
2 86394 1 3792
2 86395 1 3792
2 86396 1 3792
2 86397 1 3792
2 86398 1 3792
2 86399 1 3792
2 86400 1 3792
2 86401 1 3792
2 86402 1 3792
2 86403 1 3792
2 86404 1 3792
2 86405 1 3792
2 86406 1 3792
2 86407 1 3792
2 86408 1 3792
2 86409 1 3792
2 86410 1 3792
2 86411 1 3792
2 86412 1 3793
2 86413 1 3793
2 86414 1 3793
2 86415 1 3793
2 86416 1 3793
2 86417 1 3793
2 86418 1 3793
2 86419 1 3793
2 86420 1 3793
2 86421 1 3793
2 86422 1 3794
2 86423 1 3794
2 86424 1 3794
2 86425 1 3794
2 86426 1 3794
2 86427 1 3794
2 86428 1 3795
2 86429 1 3795
2 86430 1 3795
2 86431 1 3795
2 86432 1 3795
2 86433 1 3796
2 86434 1 3796
2 86435 1 3804
2 86436 1 3804
2 86437 1 3804
2 86438 1 3805
2 86439 1 3805
2 86440 1 3806
2 86441 1 3806
2 86442 1 3807
2 86443 1 3807
2 86444 1 3807
2 86445 1 3807
2 86446 1 3807
2 86447 1 3808
2 86448 1 3808
2 86449 1 3808
2 86450 1 3808
2 86451 1 3808
2 86452 1 3810
2 86453 1 3810
2 86454 1 3812
2 86455 1 3812
2 86456 1 3813
2 86457 1 3813
2 86458 1 3813
2 86459 1 3813
2 86460 1 3813
2 86461 1 3814
2 86462 1 3814
2 86463 1 3814
2 86464 1 3815
2 86465 1 3815
2 86466 1 3815
2 86467 1 3816
2 86468 1 3816
2 86469 1 3818
2 86470 1 3818
2 86471 1 3820
2 86472 1 3820
2 86473 1 3821
2 86474 1 3821
2 86475 1 3821
2 86476 1 3821
2 86477 1 3821
2 86478 1 3821
2 86479 1 3821
2 86480 1 3823
2 86481 1 3823
2 86482 1 3826
2 86483 1 3826
2 86484 1 3828
2 86485 1 3828
2 86486 1 3835
2 86487 1 3835
2 86488 1 3835
2 86489 1 3835
2 86490 1 3835
2 86491 1 3835
2 86492 1 3835
2 86493 1 3835
2 86494 1 3836
2 86495 1 3836
2 86496 1 3837
2 86497 1 3837
2 86498 1 3837
2 86499 1 3837
2 86500 1 3837
2 86501 1 3837
2 86502 1 3837
2 86503 1 3837
2 86504 1 3837
2 86505 1 3837
2 86506 1 3837
2 86507 1 3837
2 86508 1 3837
2 86509 1 3837
2 86510 1 3837
2 86511 1 3846
2 86512 1 3846
2 86513 1 3847
2 86514 1 3847
2 86515 1 3847
2 86516 1 3848
2 86517 1 3848
2 86518 1 3857
2 86519 1 3857
2 86520 1 3857
2 86521 1 3858
2 86522 1 3858
2 86523 1 3858
2 86524 1 3858
2 86525 1 3859
2 86526 1 3859
2 86527 1 3859
2 86528 1 3859
2 86529 1 3859
2 86530 1 3859
2 86531 1 3859
2 86532 1 3859
2 86533 1 3859
2 86534 1 3859
2 86535 1 3870
2 86536 1 3870
2 86537 1 3870
2 86538 1 3870
2 86539 1 3870
2 86540 1 3870
2 86541 1 3870
2 86542 1 3870
2 86543 1 3870
2 86544 1 3870
2 86545 1 3870
2 86546 1 3870
2 86547 1 3870
2 86548 1 3870
2 86549 1 3870
2 86550 1 3871
2 86551 1 3871
2 86552 1 3872
2 86553 1 3872
2 86554 1 3880
2 86555 1 3880
2 86556 1 3880
2 86557 1 3880
2 86558 1 3880
2 86559 1 3880
2 86560 1 3881
2 86561 1 3881
2 86562 1 3890
2 86563 1 3890
2 86564 1 3890
2 86565 1 3890
2 86566 1 3890
2 86567 1 3890
2 86568 1 3890
2 86569 1 3890
2 86570 1 3890
2 86571 1 3890
2 86572 1 3890
2 86573 1 3891
2 86574 1 3891
2 86575 1 3891
2 86576 1 3892
2 86577 1 3892
2 86578 1 3897
2 86579 1 3897
2 86580 1 3897
2 86581 1 3914
2 86582 1 3914
2 86583 1 3914
2 86584 1 3915
2 86585 1 3915
2 86586 1 3916
2 86587 1 3916
2 86588 1 3916
2 86589 1 3916
2 86590 1 3919
2 86591 1 3919
2 86592 1 3919
2 86593 1 3927
2 86594 1 3927
2 86595 1 3927
2 86596 1 3927
2 86597 1 3928
2 86598 1 3928
2 86599 1 3928
2 86600 1 3928
2 86601 1 3928
2 86602 1 3928
2 86603 1 3941
2 86604 1 3941
2 86605 1 3941
2 86606 1 3941
2 86607 1 3941
2 86608 1 3941
2 86609 1 3941
2 86610 1 3941
2 86611 1 3941
2 86612 1 3941
2 86613 1 3941
2 86614 1 3941
2 86615 1 3941
2 86616 1 3941
2 86617 1 3942
2 86618 1 3942
2 86619 1 3943
2 86620 1 3943
2 86621 1 3944
2 86622 1 3944
2 86623 1 3944
2 86624 1 3945
2 86625 1 3945
2 86626 1 3949
2 86627 1 3949
2 86628 1 3962
2 86629 1 3962
2 86630 1 3963
2 86631 1 3963
2 86632 1 3964
2 86633 1 3964
2 86634 1 3964
2 86635 1 3964
2 86636 1 3965
2 86637 1 3965
2 86638 1 3966
2 86639 1 3966
2 86640 1 3966
2 86641 1 3966
2 86642 1 3967
2 86643 1 3967
2 86644 1 3982
2 86645 1 3982
2 86646 1 3983
2 86647 1 3983
2 86648 1 3984
2 86649 1 3984
2 86650 1 3984
2 86651 1 3984
2 86652 1 3984
2 86653 1 3984
2 86654 1 3984
2 86655 1 3984
2 86656 1 3984
2 86657 1 3988
2 86658 1 3988
2 86659 1 3990
2 86660 1 3990
2 86661 1 3991
2 86662 1 3991
2 86663 1 3991
2 86664 1 3998
2 86665 1 3998
2 86666 1 3998
2 86667 1 3998
2 86668 1 3998
2 86669 1 3998
2 86670 1 3998
2 86671 1 3998
2 86672 1 3998
2 86673 1 3998
2 86674 1 3998
2 86675 1 3998
2 86676 1 3998
2 86677 1 3998
2 86678 1 3998
2 86679 1 3998
2 86680 1 3998
2 86681 1 3998
2 86682 1 3998
2 86683 1 3998
2 86684 1 3998
2 86685 1 3999
2 86686 1 3999
2 86687 1 3999
2 86688 1 3999
2 86689 1 4001
2 86690 1 4001
2 86691 1 4001
2 86692 1 4002
2 86693 1 4002
2 86694 1 4002
2 86695 1 4002
2 86696 1 4002
2 86697 1 4002
2 86698 1 4002
2 86699 1 4002
2 86700 1 4002
2 86701 1 4002
2 86702 1 4002
2 86703 1 4018
2 86704 1 4018
2 86705 1 4018
2 86706 1 4024
2 86707 1 4024
2 86708 1 4024
2 86709 1 4024
2 86710 1 4024
2 86711 1 4026
2 86712 1 4026
2 86713 1 4027
2 86714 1 4027
2 86715 1 4027
2 86716 1 4027
2 86717 1 4028
2 86718 1 4028
2 86719 1 4036
2 86720 1 4036
2 86721 1 4036
2 86722 1 4036
2 86723 1 4046
2 86724 1 4046
2 86725 1 4046
2 86726 1 4046
2 86727 1 4046
2 86728 1 4047
2 86729 1 4047
2 86730 1 4047
2 86731 1 4047
2 86732 1 4047
2 86733 1 4047
2 86734 1 4049
2 86735 1 4049
2 86736 1 4056
2 86737 1 4056
2 86738 1 4057
2 86739 1 4057
2 86740 1 4057
2 86741 1 4057
2 86742 1 4058
2 86743 1 4058
2 86744 1 4070
2 86745 1 4070
2 86746 1 4070
2 86747 1 4072
2 86748 1 4072
2 86749 1 4072
2 86750 1 4072
2 86751 1 4072
2 86752 1 4072
2 86753 1 4073
2 86754 1 4073
2 86755 1 4073
2 86756 1 4076
2 86757 1 4076
2 86758 1 4076
2 86759 1 4077
2 86760 1 4077
2 86761 1 4100
2 86762 1 4100
2 86763 1 4100
2 86764 1 4100
2 86765 1 4100
2 86766 1 4100
2 86767 1 4100
2 86768 1 4100
2 86769 1 4100
2 86770 1 4100
2 86771 1 4100
2 86772 1 4101
2 86773 1 4101
2 86774 1 4101
2 86775 1 4101
2 86776 1 4101
2 86777 1 4101
2 86778 1 4101
2 86779 1 4101
2 86780 1 4101
2 86781 1 4101
2 86782 1 4102
2 86783 1 4102
2 86784 1 4102
2 86785 1 4102
2 86786 1 4102
2 86787 1 4103
2 86788 1 4103
2 86789 1 4103
2 86790 1 4103
2 86791 1 4103
2 86792 1 4103
2 86793 1 4103
2 86794 1 4103
2 86795 1 4105
2 86796 1 4105
2 86797 1 4105
2 86798 1 4105
2 86799 1 4106
2 86800 1 4106
2 86801 1 4109
2 86802 1 4109
2 86803 1 4112
2 86804 1 4112
2 86805 1 4112
2 86806 1 4112
2 86807 1 4112
2 86808 1 4113
2 86809 1 4113
2 86810 1 4113
2 86811 1 4113
2 86812 1 4113
2 86813 1 4113
2 86814 1 4115
2 86815 1 4115
2 86816 1 4115
2 86817 1 4116
2 86818 1 4116
2 86819 1 4117
2 86820 1 4117
2 86821 1 4120
2 86822 1 4120
2 86823 1 4120
2 86824 1 4120
2 86825 1 4121
2 86826 1 4121
2 86827 1 4121
2 86828 1 4121
2 86829 1 4121
2 86830 1 4121
2 86831 1 4131
2 86832 1 4131
2 86833 1 4131
2 86834 1 4131
2 86835 1 4131
2 86836 1 4131
2 86837 1 4131
2 86838 1 4131
2 86839 1 4132
2 86840 1 4132
2 86841 1 4132
2 86842 1 4132
2 86843 1 4132
2 86844 1 4132
2 86845 1 4132
2 86846 1 4133
2 86847 1 4133
2 86848 1 4133
2 86849 1 4133
2 86850 1 4133
2 86851 1 4134
2 86852 1 4134
2 86853 1 4136
2 86854 1 4136
2 86855 1 4145
2 86856 1 4145
2 86857 1 4145
2 86858 1 4145
2 86859 1 4145
2 86860 1 4146
2 86861 1 4146
2 86862 1 4149
2 86863 1 4149
2 86864 1 4150
2 86865 1 4150
2 86866 1 4150
2 86867 1 4150
2 86868 1 4150
2 86869 1 4150
2 86870 1 4160
2 86871 1 4160
2 86872 1 4160
2 86873 1 4161
2 86874 1 4161
2 86875 1 4161
2 86876 1 4163
2 86877 1 4163
2 86878 1 4167
2 86879 1 4167
2 86880 1 4173
2 86881 1 4173
2 86882 1 4177
2 86883 1 4177
2 86884 1 4177
2 86885 1 4177
2 86886 1 4178
2 86887 1 4178
2 86888 1 4179
2 86889 1 4179
2 86890 1 4180
2 86891 1 4180
2 86892 1 4180
2 86893 1 4181
2 86894 1 4181
2 86895 1 4181
2 86896 1 4181
2 86897 1 4181
2 86898 1 4181
2 86899 1 4181
2 86900 1 4181
2 86901 1 4181
2 86902 1 4181
2 86903 1 4182
2 86904 1 4182
2 86905 1 4183
2 86906 1 4183
2 86907 1 4183
2 86908 1 4184
2 86909 1 4184
2 86910 1 4184
2 86911 1 4189
2 86912 1 4189
2 86913 1 4196
2 86914 1 4196
2 86915 1 4196
2 86916 1 4197
2 86917 1 4197
2 86918 1 4206
2 86919 1 4206
2 86920 1 4206
2 86921 1 4206
2 86922 1 4207
2 86923 1 4207
2 86924 1 4208
2 86925 1 4208
2 86926 1 4208
2 86927 1 4209
2 86928 1 4209
2 86929 1 4209
2 86930 1 4211
2 86931 1 4211
2 86932 1 4211
2 86933 1 4212
2 86934 1 4212
2 86935 1 4212
2 86936 1 4212
2 86937 1 4212
2 86938 1 4213
2 86939 1 4213
2 86940 1 4214
2 86941 1 4214
2 86942 1 4214
2 86943 1 4214
2 86944 1 4214
2 86945 1 4214
2 86946 1 4214
2 86947 1 4216
2 86948 1 4216
2 86949 1 4216
2 86950 1 4216
2 86951 1 4216
2 86952 1 4217
2 86953 1 4217
2 86954 1 4217
2 86955 1 4219
2 86956 1 4219
2 86957 1 4222
2 86958 1 4222
2 86959 1 4222
2 86960 1 4223
2 86961 1 4223
2 86962 1 4226
2 86963 1 4226
2 86964 1 4230
2 86965 1 4230
2 86966 1 4233
2 86967 1 4233
2 86968 1 4233
2 86969 1 4234
2 86970 1 4234
2 86971 1 4234
2 86972 1 4234
2 86973 1 4234
2 86974 1 4234
2 86975 1 4234
2 86976 1 4235
2 86977 1 4235
2 86978 1 4235
2 86979 1 4235
2 86980 1 4235
2 86981 1 4235
2 86982 1 4235
2 86983 1 4235
2 86984 1 4235
2 86985 1 4235
2 86986 1 4235
2 86987 1 4235
2 86988 1 4235
2 86989 1 4237
2 86990 1 4237
2 86991 1 4237
2 86992 1 4237
2 86993 1 4237
2 86994 1 4238
2 86995 1 4238
2 86996 1 4238
2 86997 1 4238
2 86998 1 4238
2 86999 1 4239
2 87000 1 4239
2 87001 1 4240
2 87002 1 4240
2 87003 1 4249
2 87004 1 4249
2 87005 1 4249
2 87006 1 4257
2 87007 1 4257
2 87008 1 4257
2 87009 1 4257
2 87010 1 4257
2 87011 1 4257
2 87012 1 4257
2 87013 1 4257
2 87014 1 4257
2 87015 1 4257
2 87016 1 4257
2 87017 1 4257
2 87018 1 4257
2 87019 1 4258
2 87020 1 4258
2 87021 1 4258
2 87022 1 4259
2 87023 1 4259
2 87024 1 4276
2 87025 1 4276
2 87026 1 4276
2 87027 1 4276
2 87028 1 4276
2 87029 1 4277
2 87030 1 4277
2 87031 1 4277
2 87032 1 4277
2 87033 1 4277
2 87034 1 4277
2 87035 1 4277
2 87036 1 4277
2 87037 1 4277
2 87038 1 4277
2 87039 1 4277
2 87040 1 4277
2 87041 1 4277
2 87042 1 4277
2 87043 1 4280
2 87044 1 4280
2 87045 1 4291
2 87046 1 4291
2 87047 1 4291
2 87048 1 4291
2 87049 1 4291
2 87050 1 4291
2 87051 1 4291
2 87052 1 4291
2 87053 1 4291
2 87054 1 4291
2 87055 1 4292
2 87056 1 4292
2 87057 1 4292
2 87058 1 4294
2 87059 1 4294
2 87060 1 4294
2 87061 1 4294
2 87062 1 4294
2 87063 1 4294
2 87064 1 4296
2 87065 1 4296
2 87066 1 4297
2 87067 1 4297
2 87068 1 4297
2 87069 1 4297
2 87070 1 4297
2 87071 1 4297
2 87072 1 4297
2 87073 1 4297
2 87074 1 4298
2 87075 1 4298
2 87076 1 4298
2 87077 1 4300
2 87078 1 4300
2 87079 1 4302
2 87080 1 4302
2 87081 1 4305
2 87082 1 4305
2 87083 1 4305
2 87084 1 4305
2 87085 1 4305
2 87086 1 4305
2 87087 1 4305
2 87088 1 4306
2 87089 1 4306
2 87090 1 4307
2 87091 1 4307
2 87092 1 4314
2 87093 1 4314
2 87094 1 4314
2 87095 1 4315
2 87096 1 4315
2 87097 1 4315
2 87098 1 4315
2 87099 1 4336
2 87100 1 4336
2 87101 1 4336
2 87102 1 4336
2 87103 1 4336
2 87104 1 4336
2 87105 1 4336
2 87106 1 4336
2 87107 1 4336
2 87108 1 4336
2 87109 1 4337
2 87110 1 4337
2 87111 1 4337
2 87112 1 4337
2 87113 1 4341
2 87114 1 4341
2 87115 1 4342
2 87116 1 4342
2 87117 1 4351
2 87118 1 4351
2 87119 1 4352
2 87120 1 4352
2 87121 1 4352
2 87122 1 4352
2 87123 1 4352
2 87124 1 4352
2 87125 1 4352
2 87126 1 4352
2 87127 1 4352
2 87128 1 4352
2 87129 1 4352
2 87130 1 4352
2 87131 1 4352
2 87132 1 4352
2 87133 1 4352
2 87134 1 4352
2 87135 1 4352
2 87136 1 4353
2 87137 1 4353
2 87138 1 4353
2 87139 1 4365
2 87140 1 4365
2 87141 1 4366
2 87142 1 4366
2 87143 1 4366
2 87144 1 4377
2 87145 1 4377
2 87146 1 4378
2 87147 1 4378
2 87148 1 4378
2 87149 1 4379
2 87150 1 4379
2 87151 1 4379
2 87152 1 4379
2 87153 1 4386
2 87154 1 4386
2 87155 1 4386
2 87156 1 4387
2 87157 1 4387
2 87158 1 4387
2 87159 1 4387
2 87160 1 4396
2 87161 1 4396
2 87162 1 4396
2 87163 1 4404
2 87164 1 4404
2 87165 1 4404
2 87166 1 4404
2 87167 1 4404
2 87168 1 4404
2 87169 1 4404
2 87170 1 4406
2 87171 1 4406
2 87172 1 4406
2 87173 1 4407
2 87174 1 4407
2 87175 1 4407
2 87176 1 4441
2 87177 1 4441
2 87178 1 4441
2 87179 1 4441
2 87180 1 4445
2 87181 1 4445
2 87182 1 4445
2 87183 1 4445
2 87184 1 4445
2 87185 1 4445
2 87186 1 4445
2 87187 1 4445
2 87188 1 4445
2 87189 1 4445
2 87190 1 4445
2 87191 1 4445
2 87192 1 4445
2 87193 1 4445
2 87194 1 4445
2 87195 1 4445
2 87196 1 4447
2 87197 1 4447
2 87198 1 4457
2 87199 1 4457
2 87200 1 4457
2 87201 1 4457
2 87202 1 4457
2 87203 1 4457
2 87204 1 4457
2 87205 1 4457
2 87206 1 4457
2 87207 1 4457
2 87208 1 4457
2 87209 1 4457
2 87210 1 4458
2 87211 1 4458
2 87212 1 4458
2 87213 1 4459
2 87214 1 4459
2 87215 1 4459
2 87216 1 4459
2 87217 1 4459
2 87218 1 4460
2 87219 1 4460
2 87220 1 4466
2 87221 1 4466
2 87222 1 4466
2 87223 1 4467
2 87224 1 4467
2 87225 1 4467
2 87226 1 4467
2 87227 1 4467
2 87228 1 4467
2 87229 1 4467
2 87230 1 4467
2 87231 1 4467
2 87232 1 4467
2 87233 1 4467
2 87234 1 4467
2 87235 1 4467
2 87236 1 4467
2 87237 1 4467
2 87238 1 4467
2 87239 1 4468
2 87240 1 4468
2 87241 1 4468
2 87242 1 4468
2 87243 1 4468
2 87244 1 4468
2 87245 1 4468
2 87246 1 4468
2 87247 1 4468
2 87248 1 4468
2 87249 1 4468
2 87250 1 4468
2 87251 1 4468
2 87252 1 4468
2 87253 1 4475
2 87254 1 4475
2 87255 1 4475
2 87256 1 4475
2 87257 1 4475
2 87258 1 4475
2 87259 1 4475
2 87260 1 4475
2 87261 1 4477
2 87262 1 4477
2 87263 1 4478
2 87264 1 4478
2 87265 1 4492
2 87266 1 4492
2 87267 1 4492
2 87268 1 4492
2 87269 1 4492
2 87270 1 4495
2 87271 1 4495
2 87272 1 4495
2 87273 1 4495
2 87274 1 4496
2 87275 1 4496
2 87276 1 4496
2 87277 1 4503
2 87278 1 4503
2 87279 1 4503
2 87280 1 4503
2 87281 1 4503
2 87282 1 4504
2 87283 1 4504
2 87284 1 4504
2 87285 1 4504
2 87286 1 4504
2 87287 1 4504
2 87288 1 4504
2 87289 1 4504
2 87290 1 4504
2 87291 1 4504
2 87292 1 4504
2 87293 1 4504
2 87294 1 4504
2 87295 1 4505
2 87296 1 4505
2 87297 1 4505
2 87298 1 4513
2 87299 1 4513
2 87300 1 4516
2 87301 1 4516
2 87302 1 4516
2 87303 1 4516
2 87304 1 4517
2 87305 1 4517
2 87306 1 4518
2 87307 1 4518
2 87308 1 4518
2 87309 1 4520
2 87310 1 4520
2 87311 1 4520
2 87312 1 4520
2 87313 1 4520
2 87314 1 4520
2 87315 1 4532
2 87316 1 4532
2 87317 1 4532
2 87318 1 4532
2 87319 1 4532
2 87320 1 4532
2 87321 1 4534
2 87322 1 4534
2 87323 1 4537
2 87324 1 4537
2 87325 1 4540
2 87326 1 4540
2 87327 1 4546
2 87328 1 4546
2 87329 1 4546
2 87330 1 4546
2 87331 1 4546
2 87332 1 4546
2 87333 1 4546
2 87334 1 4546
2 87335 1 4546
2 87336 1 4546
2 87337 1 4546
2 87338 1 4546
2 87339 1 4546
2 87340 1 4546
2 87341 1 4546
2 87342 1 4546
2 87343 1 4546
2 87344 1 4547
2 87345 1 4547
2 87346 1 4548
2 87347 1 4548
2 87348 1 4548
2 87349 1 4548
2 87350 1 4549
2 87351 1 4549
2 87352 1 4549
2 87353 1 4549
2 87354 1 4549
2 87355 1 4551
2 87356 1 4551
2 87357 1 4551
2 87358 1 4551
2 87359 1 4551
2 87360 1 4551
2 87361 1 4551
2 87362 1 4551
2 87363 1 4551
2 87364 1 4551
2 87365 1 4551
2 87366 1 4555
2 87367 1 4555
2 87368 1 4558
2 87369 1 4558
2 87370 1 4559
2 87371 1 4559
2 87372 1 4560
2 87373 1 4560
2 87374 1 4560
2 87375 1 4560
2 87376 1 4560
2 87377 1 4560
2 87378 1 4560
2 87379 1 4560
2 87380 1 4560
2 87381 1 4560
2 87382 1 4560
2 87383 1 4560
2 87384 1 4560
2 87385 1 4560
2 87386 1 4560
2 87387 1 4561
2 87388 1 4561
2 87389 1 4564
2 87390 1 4564
2 87391 1 4564
2 87392 1 4564
2 87393 1 4565
2 87394 1 4565
2 87395 1 4579
2 87396 1 4579
2 87397 1 4579
2 87398 1 4579
2 87399 1 4579
2 87400 1 4579
2 87401 1 4579
2 87402 1 4579
2 87403 1 4579
2 87404 1 4579
2 87405 1 4579
2 87406 1 4579
2 87407 1 4579
2 87408 1 4579
2 87409 1 4579
2 87410 1 4579
2 87411 1 4579
2 87412 1 4579
2 87413 1 4579
2 87414 1 4579
2 87415 1 4579
2 87416 1 4579
2 87417 1 4579
2 87418 1 4579
2 87419 1 4579
2 87420 1 4579
2 87421 1 4579
2 87422 1 4579
2 87423 1 4579
2 87424 1 4579
2 87425 1 4580
2 87426 1 4580
2 87427 1 4580
2 87428 1 4580
2 87429 1 4580
2 87430 1 4580
2 87431 1 4581
2 87432 1 4581
2 87433 1 4590
2 87434 1 4590
2 87435 1 4590
2 87436 1 4590
2 87437 1 4590
2 87438 1 4590
2 87439 1 4590
2 87440 1 4590
2 87441 1 4590
2 87442 1 4590
2 87443 1 4591
2 87444 1 4591
2 87445 1 4599
2 87446 1 4599
2 87447 1 4600
2 87448 1 4600
2 87449 1 4600
2 87450 1 4600
2 87451 1 4600
2 87452 1 4600
2 87453 1 4600
2 87454 1 4600
2 87455 1 4600
2 87456 1 4600
2 87457 1 4600
2 87458 1 4600
2 87459 1 4600
2 87460 1 4600
2 87461 1 4600
2 87462 1 4600
2 87463 1 4601
2 87464 1 4601
2 87465 1 4602
2 87466 1 4602
2 87467 1 4603
2 87468 1 4603
2 87469 1 4603
2 87470 1 4603
2 87471 1 4603
2 87472 1 4603
2 87473 1 4603
2 87474 1 4603
2 87475 1 4603
2 87476 1 4603
2 87477 1 4603
2 87478 1 4603
2 87479 1 4603
2 87480 1 4604
2 87481 1 4604
2 87482 1 4604
2 87483 1 4604
2 87484 1 4604
2 87485 1 4604
2 87486 1 4607
2 87487 1 4607
2 87488 1 4607
2 87489 1 4607
2 87490 1 4607
2 87491 1 4620
2 87492 1 4620
2 87493 1 4620
2 87494 1 4620
2 87495 1 4620
2 87496 1 4630
2 87497 1 4630
2 87498 1 4633
2 87499 1 4633
2 87500 1 4634
2 87501 1 4634
2 87502 1 4634
2 87503 1 4634
2 87504 1 4634
2 87505 1 4634
2 87506 1 4634
2 87507 1 4634
2 87508 1 4634
2 87509 1 4634
2 87510 1 4634
2 87511 1 4634
2 87512 1 4634
2 87513 1 4634
2 87514 1 4634
2 87515 1 4634
2 87516 1 4634
2 87517 1 4636
2 87518 1 4636
2 87519 1 4643
2 87520 1 4643
2 87521 1 4643
2 87522 1 4650
2 87523 1 4650
2 87524 1 4651
2 87525 1 4651
2 87526 1 4651
2 87527 1 4651
2 87528 1 4651
2 87529 1 4662
2 87530 1 4662
2 87531 1 4663
2 87532 1 4663
2 87533 1 4667
2 87534 1 4667
2 87535 1 4668
2 87536 1 4668
2 87537 1 4668
2 87538 1 4675
2 87539 1 4675
2 87540 1 4675
2 87541 1 4675
2 87542 1 4676
2 87543 1 4676
2 87544 1 4678
2 87545 1 4678
2 87546 1 4678
2 87547 1 4678
2 87548 1 4678
2 87549 1 4678
2 87550 1 4678
2 87551 1 4678
2 87552 1 4678
2 87553 1 4679
2 87554 1 4679
2 87555 1 4681
2 87556 1 4681
2 87557 1 4686
2 87558 1 4686
2 87559 1 4701
2 87560 1 4701
2 87561 1 4702
2 87562 1 4702
2 87563 1 4702
2 87564 1 4703
2 87565 1 4703
2 87566 1 4703
2 87567 1 4703
2 87568 1 4703
2 87569 1 4704
2 87570 1 4704
2 87571 1 4704
2 87572 1 4704
2 87573 1 4704
2 87574 1 4704
2 87575 1 4705
2 87576 1 4705
2 87577 1 4708
2 87578 1 4708
2 87579 1 4709
2 87580 1 4709
2 87581 1 4709
2 87582 1 4709
2 87583 1 4709
2 87584 1 4717
2 87585 1 4717
2 87586 1 4718
2 87587 1 4718
2 87588 1 4718
2 87589 1 4718
2 87590 1 4719
2 87591 1 4719
2 87592 1 4728
2 87593 1 4728
2 87594 1 4739
2 87595 1 4739
2 87596 1 4739
2 87597 1 4739
2 87598 1 4739
2 87599 1 4739
2 87600 1 4740
2 87601 1 4740
2 87602 1 4740
2 87603 1 4744
2 87604 1 4744
2 87605 1 4744
2 87606 1 4744
2 87607 1 4745
2 87608 1 4745
2 87609 1 4745
2 87610 1 4746
2 87611 1 4746
2 87612 1 4746
2 87613 1 4746
2 87614 1 4754
2 87615 1 4754
2 87616 1 4754
2 87617 1 4754
2 87618 1 4755
2 87619 1 4755
2 87620 1 4757
2 87621 1 4757
2 87622 1 4757
2 87623 1 4765
2 87624 1 4765
2 87625 1 4765
2 87626 1 4765
2 87627 1 4765
2 87628 1 4765
2 87629 1 4765
2 87630 1 4765
2 87631 1 4765
2 87632 1 4766
2 87633 1 4766
2 87634 1 4766
2 87635 1 4766
2 87636 1 4766
2 87637 1 4766
2 87638 1 4766
2 87639 1 4766
2 87640 1 4766
2 87641 1 4766
2 87642 1 4766
2 87643 1 4766
2 87644 1 4767
2 87645 1 4767
2 87646 1 4767
2 87647 1 4767
2 87648 1 4767
2 87649 1 4767
2 87650 1 4767
2 87651 1 4767
2 87652 1 4767
2 87653 1 4767
2 87654 1 4767
2 87655 1 4768
2 87656 1 4768
2 87657 1 4768
2 87658 1 4768
2 87659 1 4769
2 87660 1 4769
2 87661 1 4769
2 87662 1 4771
2 87663 1 4771
2 87664 1 4771
2 87665 1 4771
2 87666 1 4771
2 87667 1 4771
2 87668 1 4771
2 87669 1 4771
2 87670 1 4771
2 87671 1 4771
2 87672 1 4771
2 87673 1 4771
2 87674 1 4786
2 87675 1 4786
2 87676 1 4787
2 87677 1 4787
2 87678 1 4799
2 87679 1 4799
2 87680 1 4801
2 87681 1 4801
2 87682 1 4807
2 87683 1 4807
2 87684 1 4807
2 87685 1 4811
2 87686 1 4811
2 87687 1 4815
2 87688 1 4815
2 87689 1 4815
2 87690 1 4816
2 87691 1 4816
2 87692 1 4816
2 87693 1 4816
2 87694 1 4816
2 87695 1 4816
2 87696 1 4816
2 87697 1 4816
2 87698 1 4816
2 87699 1 4816
2 87700 1 4816
2 87701 1 4816
2 87702 1 4816
2 87703 1 4816
2 87704 1 4816
2 87705 1 4816
2 87706 1 4816
2 87707 1 4816
2 87708 1 4816
2 87709 1 4816
2 87710 1 4816
2 87711 1 4816
2 87712 1 4816
2 87713 1 4817
2 87714 1 4817
2 87715 1 4820
2 87716 1 4820
2 87717 1 4832
2 87718 1 4832
2 87719 1 4833
2 87720 1 4833
2 87721 1 4833
2 87722 1 4833
2 87723 1 4833
2 87724 1 4833
2 87725 1 4833
2 87726 1 4833
2 87727 1 4833
2 87728 1 4833
2 87729 1 4833
2 87730 1 4833
2 87731 1 4833
2 87732 1 4833
2 87733 1 4833
2 87734 1 4833
2 87735 1 4833
2 87736 1 4833
2 87737 1 4833
2 87738 1 4833
2 87739 1 4833
2 87740 1 4833
2 87741 1 4833
2 87742 1 4833
2 87743 1 4833
2 87744 1 4833
2 87745 1 4833
2 87746 1 4833
2 87747 1 4833
2 87748 1 4833
2 87749 1 4833
2 87750 1 4833
2 87751 1 4833
2 87752 1 4833
2 87753 1 4833
2 87754 1 4833
2 87755 1 4833
2 87756 1 4833
2 87757 1 4833
2 87758 1 4833
2 87759 1 4834
2 87760 1 4834
2 87761 1 4834
2 87762 1 4834
2 87763 1 4834
2 87764 1 4835
2 87765 1 4835
2 87766 1 4835
2 87767 1 4838
2 87768 1 4838
2 87769 1 4838
2 87770 1 4839
2 87771 1 4839
2 87772 1 4839
2 87773 1 4841
2 87774 1 4841
2 87775 1 4841
2 87776 1 4841
2 87777 1 4842
2 87778 1 4842
2 87779 1 4842
2 87780 1 4842
2 87781 1 4843
2 87782 1 4843
2 87783 1 4843
2 87784 1 4843
2 87785 1 4843
2 87786 1 4843
2 87787 1 4843
2 87788 1 4843
2 87789 1 4843
2 87790 1 4843
2 87791 1 4843
2 87792 1 4843
2 87793 1 4843
2 87794 1 4843
2 87795 1 4843
2 87796 1 4843
2 87797 1 4843
2 87798 1 4843
2 87799 1 4843
2 87800 1 4843
2 87801 1 4843
2 87802 1 4843
2 87803 1 4843
2 87804 1 4843
2 87805 1 4843
2 87806 1 4843
2 87807 1 4843
2 87808 1 4843
2 87809 1 4843
2 87810 1 4843
2 87811 1 4843
2 87812 1 4843
2 87813 1 4843
2 87814 1 4844
2 87815 1 4844
2 87816 1 4844
2 87817 1 4844
2 87818 1 4846
2 87819 1 4846
2 87820 1 4851
2 87821 1 4851
2 87822 1 4851
2 87823 1 4852
2 87824 1 4852
2 87825 1 4852
2 87826 1 4857
2 87827 1 4857
2 87828 1 4857
2 87829 1 4861
2 87830 1 4861
2 87831 1 4861
2 87832 1 4861
2 87833 1 4861
2 87834 1 4861
2 87835 1 4862
2 87836 1 4862
2 87837 1 4862
2 87838 1 4871
2 87839 1 4871
2 87840 1 4873
2 87841 1 4873
2 87842 1 4873
2 87843 1 4873
2 87844 1 4873
2 87845 1 4874
2 87846 1 4874
2 87847 1 4878
2 87848 1 4878
2 87849 1 4881
2 87850 1 4881
2 87851 1 4882
2 87852 1 4882
2 87853 1 4885
2 87854 1 4885
2 87855 1 4886
2 87856 1 4886
2 87857 1 4894
2 87858 1 4894
2 87859 1 4894
2 87860 1 4896
2 87861 1 4896
2 87862 1 4896
2 87863 1 4906
2 87864 1 4906
2 87865 1 4906
2 87866 1 4906
2 87867 1 4906
2 87868 1 4906
2 87869 1 4906
2 87870 1 4906
2 87871 1 4907
2 87872 1 4907
2 87873 1 4907
2 87874 1 4915
2 87875 1 4915
2 87876 1 4918
2 87877 1 4918
2 87878 1 4921
2 87879 1 4921
2 87880 1 4921
2 87881 1 4921
2 87882 1 4921
2 87883 1 4921
2 87884 1 4921
2 87885 1 4921
2 87886 1 4921
2 87887 1 4921
2 87888 1 4921
2 87889 1 4922
2 87890 1 4922
2 87891 1 4925
2 87892 1 4925
2 87893 1 4939
2 87894 1 4939
2 87895 1 4939
2 87896 1 4939
2 87897 1 4939
2 87898 1 4941
2 87899 1 4941
2 87900 1 4941
2 87901 1 4941
2 87902 1 4943
2 87903 1 4943
2 87904 1 4946
2 87905 1 4946
2 87906 1 4947
2 87907 1 4947
2 87908 1 4947
2 87909 1 4947
2 87910 1 4947
2 87911 1 4947
2 87912 1 4947
2 87913 1 4947
2 87914 1 4947
2 87915 1 4948
2 87916 1 4948
2 87917 1 4948
2 87918 1 4948
2 87919 1 4948
2 87920 1 4948
2 87921 1 4948
2 87922 1 4948
2 87923 1 4948
2 87924 1 4948
2 87925 1 4948
2 87926 1 4948
2 87927 1 4948
2 87928 1 4948
2 87929 1 4948
2 87930 1 4948
2 87931 1 4948
2 87932 1 4949
2 87933 1 4949
2 87934 1 4949
2 87935 1 4961
2 87936 1 4961
2 87937 1 4962
2 87938 1 4962
2 87939 1 4965
2 87940 1 4965
2 87941 1 4967
2 87942 1 4967
2 87943 1 4968
2 87944 1 4968
2 87945 1 4968
2 87946 1 4969
2 87947 1 4969
2 87948 1 4972
2 87949 1 4972
2 87950 1 4973
2 87951 1 4973
2 87952 1 4973
2 87953 1 4973
2 87954 1 4973
2 87955 1 4973
2 87956 1 4973
2 87957 1 4973
2 87958 1 4973
2 87959 1 4973
2 87960 1 4973
2 87961 1 4973
2 87962 1 4973
2 87963 1 4973
2 87964 1 4973
2 87965 1 4973
2 87966 1 4973
2 87967 1 4974
2 87968 1 4974
2 87969 1 4998
2 87970 1 4998
2 87971 1 4999
2 87972 1 4999
2 87973 1 4999
2 87974 1 4999
2 87975 1 5000
2 87976 1 5000
2 87977 1 5000
2 87978 1 5000
2 87979 1 5001
2 87980 1 5001
2 87981 1 5006
2 87982 1 5006
2 87983 1 5022
2 87984 1 5022
2 87985 1 5022
2 87986 1 5022
2 87987 1 5022
2 87988 1 5022
2 87989 1 5022
2 87990 1 5023
2 87991 1 5023
2 87992 1 5023
2 87993 1 5026
2 87994 1 5026
2 87995 1 5026
2 87996 1 5026
2 87997 1 5026
2 87998 1 5026
2 87999 1 5026
2 88000 1 5026
2 88001 1 5026
2 88002 1 5026
2 88003 1 5026
2 88004 1 5026
2 88005 1 5026
2 88006 1 5027
2 88007 1 5027
2 88008 1 5032
2 88009 1 5032
2 88010 1 5032
2 88011 1 5042
2 88012 1 5042
2 88013 1 5042
2 88014 1 5042
2 88015 1 5042
2 88016 1 5042
2 88017 1 5042
2 88018 1 5042
2 88019 1 5042
2 88020 1 5042
2 88021 1 5042
2 88022 1 5042
2 88023 1 5042
2 88024 1 5042
2 88025 1 5042
2 88026 1 5042
2 88027 1 5042
2 88028 1 5042
2 88029 1 5042
2 88030 1 5042
2 88031 1 5042
2 88032 1 5042
2 88033 1 5042
2 88034 1 5042
2 88035 1 5042
2 88036 1 5042
2 88037 1 5042
2 88038 1 5043
2 88039 1 5043
2 88040 1 5043
2 88041 1 5043
2 88042 1 5043
2 88043 1 5043
2 88044 1 5043
2 88045 1 5043
2 88046 1 5044
2 88047 1 5044
2 88048 1 5044
2 88049 1 5044
2 88050 1 5044
2 88051 1 5044
2 88052 1 5044
2 88053 1 5044
2 88054 1 5044
2 88055 1 5044
2 88056 1 5045
2 88057 1 5045
2 88058 1 5045
2 88059 1 5045
2 88060 1 5045
2 88061 1 5045
2 88062 1 5045
2 88063 1 5045
2 88064 1 5045
2 88065 1 5045
2 88066 1 5045
2 88067 1 5045
2 88068 1 5045
2 88069 1 5045
2 88070 1 5045
2 88071 1 5045
2 88072 1 5045
2 88073 1 5045
2 88074 1 5045
2 88075 1 5045
2 88076 1 5045
2 88077 1 5045
2 88078 1 5045
2 88079 1 5045
2 88080 1 5045
2 88081 1 5045
2 88082 1 5045
2 88083 1 5045
2 88084 1 5045
2 88085 1 5045
2 88086 1 5045
2 88087 1 5045
2 88088 1 5046
2 88089 1 5046
2 88090 1 5046
2 88091 1 5046
2 88092 1 5046
2 88093 1 5046
2 88094 1 5046
2 88095 1 5046
2 88096 1 5046
2 88097 1 5046
2 88098 1 5046
2 88099 1 5046
2 88100 1 5046
2 88101 1 5046
2 88102 1 5046
2 88103 1 5046
2 88104 1 5046
2 88105 1 5046
2 88106 1 5046
2 88107 1 5046
2 88108 1 5046
2 88109 1 5046
2 88110 1 5046
2 88111 1 5046
2 88112 1 5046
2 88113 1 5046
2 88114 1 5046
2 88115 1 5046
2 88116 1 5046
2 88117 1 5046
2 88118 1 5046
2 88119 1 5046
2 88120 1 5046
2 88121 1 5046
2 88122 1 5046
2 88123 1 5046
2 88124 1 5046
2 88125 1 5046
2 88126 1 5046
2 88127 1 5046
2 88128 1 5046
2 88129 1 5046
2 88130 1 5046
2 88131 1 5046
2 88132 1 5046
2 88133 1 5046
2 88134 1 5046
2 88135 1 5046
2 88136 1 5046
2 88137 1 5046
2 88138 1 5046
2 88139 1 5046
2 88140 1 5046
2 88141 1 5046
2 88142 1 5046
2 88143 1 5046
2 88144 1 5046
2 88145 1 5046
2 88146 1 5046
2 88147 1 5046
2 88148 1 5046
2 88149 1 5046
2 88150 1 5046
2 88151 1 5046
2 88152 1 5046
2 88153 1 5046
2 88154 1 5046
2 88155 1 5046
2 88156 1 5046
2 88157 1 5046
2 88158 1 5046
2 88159 1 5046
2 88160 1 5046
2 88161 1 5046
2 88162 1 5046
2 88163 1 5046
2 88164 1 5046
2 88165 1 5046
2 88166 1 5046
2 88167 1 5046
2 88168 1 5046
2 88169 1 5046
2 88170 1 5046
2 88171 1 5046
2 88172 1 5046
2 88173 1 5046
2 88174 1 5046
2 88175 1 5046
2 88176 1 5046
2 88177 1 5046
2 88178 1 5046
2 88179 1 5046
2 88180 1 5046
2 88181 1 5046
2 88182 1 5046
2 88183 1 5046
2 88184 1 5046
2 88185 1 5046
2 88186 1 5046
2 88187 1 5046
2 88188 1 5046
2 88189 1 5046
2 88190 1 5046
2 88191 1 5046
2 88192 1 5046
2 88193 1 5046
2 88194 1 5046
2 88195 1 5046
2 88196 1 5046
2 88197 1 5046
2 88198 1 5046
2 88199 1 5046
2 88200 1 5046
2 88201 1 5046
2 88202 1 5046
2 88203 1 5046
2 88204 1 5046
2 88205 1 5046
2 88206 1 5046
2 88207 1 5046
2 88208 1 5046
2 88209 1 5046
2 88210 1 5046
2 88211 1 5046
2 88212 1 5046
2 88213 1 5046
2 88214 1 5046
2 88215 1 5046
2 88216 1 5046
2 88217 1 5046
2 88218 1 5046
2 88219 1 5046
2 88220 1 5046
2 88221 1 5046
2 88222 1 5046
2 88223 1 5046
2 88224 1 5046
2 88225 1 5046
2 88226 1 5046
2 88227 1 5046
2 88228 1 5046
2 88229 1 5046
2 88230 1 5046
2 88231 1 5046
2 88232 1 5046
2 88233 1 5046
2 88234 1 5046
2 88235 1 5046
2 88236 1 5046
2 88237 1 5046
2 88238 1 5046
2 88239 1 5046
2 88240 1 5046
2 88241 1 5046
2 88242 1 5046
2 88243 1 5046
2 88244 1 5046
2 88245 1 5046
2 88246 1 5046
2 88247 1 5046
2 88248 1 5046
2 88249 1 5046
2 88250 1 5046
2 88251 1 5046
2 88252 1 5046
2 88253 1 5046
2 88254 1 5046
2 88255 1 5046
2 88256 1 5046
2 88257 1 5046
2 88258 1 5046
2 88259 1 5046
2 88260 1 5046
2 88261 1 5046
2 88262 1 5046
2 88263 1 5046
2 88264 1 5046
2 88265 1 5046
2 88266 1 5046
2 88267 1 5046
2 88268 1 5046
2 88269 1 5046
2 88270 1 5046
2 88271 1 5046
2 88272 1 5046
2 88273 1 5046
2 88274 1 5046
2 88275 1 5046
2 88276 1 5046
2 88277 1 5046
2 88278 1 5046
2 88279 1 5046
2 88280 1 5046
2 88281 1 5046
2 88282 1 5046
2 88283 1 5047
2 88284 1 5047
2 88285 1 5047
2 88286 1 5047
2 88287 1 5047
2 88288 1 5047
2 88289 1 5047
2 88290 1 5047
2 88291 1 5047
2 88292 1 5047
2 88293 1 5047
2 88294 1 5047
2 88295 1 5049
2 88296 1 5049
2 88297 1 5050
2 88298 1 5050
2 88299 1 5050
2 88300 1 5050
2 88301 1 5051
2 88302 1 5051
2 88303 1 5051
2 88304 1 5058
2 88305 1 5058
2 88306 1 5058
2 88307 1 5058
2 88308 1 5058
2 88309 1 5058
2 88310 1 5058
2 88311 1 5059
2 88312 1 5059
2 88313 1 5059
2 88314 1 5067
2 88315 1 5067
2 88316 1 5067
2 88317 1 5069
2 88318 1 5069
2 88319 1 5076
2 88320 1 5076
2 88321 1 5076
2 88322 1 5076
2 88323 1 5076
2 88324 1 5076
2 88325 1 5089
2 88326 1 5089
2 88327 1 5092
2 88328 1 5092
2 88329 1 5092
2 88330 1 5092
2 88331 1 5092
2 88332 1 5099
2 88333 1 5099
2 88334 1 5099
2 88335 1 5099
2 88336 1 5099
2 88337 1 5099
2 88338 1 5100
2 88339 1 5100
2 88340 1 5101
2 88341 1 5101
2 88342 1 5101
2 88343 1 5101
2 88344 1 5101
2 88345 1 5103
2 88346 1 5103
2 88347 1 5103
2 88348 1 5103
2 88349 1 5103
2 88350 1 5103
2 88351 1 5103
2 88352 1 5103
2 88353 1 5103
2 88354 1 5103
2 88355 1 5103
2 88356 1 5103
2 88357 1 5103
2 88358 1 5104
2 88359 1 5104
2 88360 1 5105
2 88361 1 5105
2 88362 1 5105
2 88363 1 5128
2 88364 1 5128
2 88365 1 5128
2 88366 1 5128
2 88367 1 5128
2 88368 1 5128
2 88369 1 5128
2 88370 1 5128
2 88371 1 5128
2 88372 1 5128
2 88373 1 5128
2 88374 1 5129
2 88375 1 5129
2 88376 1 5129
2 88377 1 5129
2 88378 1 5129
2 88379 1 5129
2 88380 1 5129
2 88381 1 5129
2 88382 1 5130
2 88383 1 5130
2 88384 1 5130
2 88385 1 5130
2 88386 1 5130
2 88387 1 5131
2 88388 1 5131
2 88389 1 5131
2 88390 1 5131
2 88391 1 5131
2 88392 1 5131
2 88393 1 5131
2 88394 1 5131
2 88395 1 5131
2 88396 1 5131
2 88397 1 5131
2 88398 1 5131
2 88399 1 5131
2 88400 1 5131
2 88401 1 5131
2 88402 1 5131
2 88403 1 5131
2 88404 1 5131
2 88405 1 5131
2 88406 1 5131
2 88407 1 5131
2 88408 1 5131
2 88409 1 5131
2 88410 1 5131
2 88411 1 5131
2 88412 1 5132
2 88413 1 5132
2 88414 1 5132
2 88415 1 5134
2 88416 1 5134
2 88417 1 5135
2 88418 1 5135
2 88419 1 5135
2 88420 1 5135
2 88421 1 5136
2 88422 1 5136
2 88423 1 5139
2 88424 1 5139
2 88425 1 5145
2 88426 1 5145
2 88427 1 5146
2 88428 1 5146
2 88429 1 5146
2 88430 1 5146
2 88431 1 5146
2 88432 1 5153
2 88433 1 5153
2 88434 1 5153
2 88435 1 5153
2 88436 1 5154
2 88437 1 5154
2 88438 1 5156
2 88439 1 5156
2 88440 1 5173
2 88441 1 5173
2 88442 1 5174
2 88443 1 5174
2 88444 1 5174
2 88445 1 5174
2 88446 1 5175
2 88447 1 5175
2 88448 1 5175
2 88449 1 5176
2 88450 1 5176
2 88451 1 5176
2 88452 1 5176
2 88453 1 5176
2 88454 1 5182
2 88455 1 5182
2 88456 1 5182
2 88457 1 5182
2 88458 1 5182
2 88459 1 5182
2 88460 1 5182
2 88461 1 5182
2 88462 1 5182
2 88463 1 5183
2 88464 1 5183
2 88465 1 5200
2 88466 1 5200
2 88467 1 5200
2 88468 1 5200
2 88469 1 5205
2 88470 1 5205
2 88471 1 5205
2 88472 1 5205
2 88473 1 5205
2 88474 1 5205
2 88475 1 5208
2 88476 1 5208
2 88477 1 5209
2 88478 1 5209
2 88479 1 5230
2 88480 1 5230
2 88481 1 5230
2 88482 1 5230
2 88483 1 5230
2 88484 1 5230
2 88485 1 5230
2 88486 1 5230
2 88487 1 5230
2 88488 1 5230
2 88489 1 5230
2 88490 1 5230
2 88491 1 5230
2 88492 1 5230
2 88493 1 5230
2 88494 1 5230
2 88495 1 5230
2 88496 1 5230
2 88497 1 5230
2 88498 1 5230
2 88499 1 5230
2 88500 1 5230
2 88501 1 5230
2 88502 1 5230
2 88503 1 5230
2 88504 1 5230
2 88505 1 5230
2 88506 1 5230
2 88507 1 5230
2 88508 1 5230
2 88509 1 5230
2 88510 1 5230
2 88511 1 5230
2 88512 1 5230
2 88513 1 5230
2 88514 1 5230
2 88515 1 5230
2 88516 1 5230
2 88517 1 5230
2 88518 1 5230
2 88519 1 5230
2 88520 1 5230
2 88521 1 5230
2 88522 1 5230
2 88523 1 5230
2 88524 1 5230
2 88525 1 5230
2 88526 1 5230
2 88527 1 5230
2 88528 1 5230
2 88529 1 5230
2 88530 1 5230
2 88531 1 5230
2 88532 1 5230
2 88533 1 5230
2 88534 1 5230
2 88535 1 5230
2 88536 1 5230
2 88537 1 5230
2 88538 1 5230
2 88539 1 5230
2 88540 1 5230
2 88541 1 5230
2 88542 1 5230
2 88543 1 5230
2 88544 1 5230
2 88545 1 5230
2 88546 1 5230
2 88547 1 5230
2 88548 1 5230
2 88549 1 5230
2 88550 1 5230
2 88551 1 5230
2 88552 1 5230
2 88553 1 5230
2 88554 1 5230
2 88555 1 5230
2 88556 1 5230
2 88557 1 5230
2 88558 1 5230
2 88559 1 5230
2 88560 1 5230
2 88561 1 5230
2 88562 1 5230
2 88563 1 5230
2 88564 1 5230
2 88565 1 5230
2 88566 1 5230
2 88567 1 5230
2 88568 1 5230
2 88569 1 5230
2 88570 1 5230
2 88571 1 5230
2 88572 1 5230
2 88573 1 5230
2 88574 1 5230
2 88575 1 5230
2 88576 1 5230
2 88577 1 5230
2 88578 1 5230
2 88579 1 5230
2 88580 1 5230
2 88581 1 5230
2 88582 1 5230
2 88583 1 5230
2 88584 1 5230
2 88585 1 5230
2 88586 1 5230
2 88587 1 5230
2 88588 1 5230
2 88589 1 5230
2 88590 1 5230
2 88591 1 5230
2 88592 1 5230
2 88593 1 5230
2 88594 1 5230
2 88595 1 5230
2 88596 1 5230
2 88597 1 5230
2 88598 1 5230
2 88599 1 5230
2 88600 1 5230
2 88601 1 5230
2 88602 1 5230
2 88603 1 5230
2 88604 1 5230
2 88605 1 5230
2 88606 1 5230
2 88607 1 5230
2 88608 1 5230
2 88609 1 5230
2 88610 1 5230
2 88611 1 5230
2 88612 1 5230
2 88613 1 5230
2 88614 1 5230
2 88615 1 5230
2 88616 1 5230
2 88617 1 5230
2 88618 1 5230
2 88619 1 5230
2 88620 1 5230
2 88621 1 5230
2 88622 1 5230
2 88623 1 5230
2 88624 1 5230
2 88625 1 5230
2 88626 1 5230
2 88627 1 5230
2 88628 1 5230
2 88629 1 5230
2 88630 1 5230
2 88631 1 5230
2 88632 1 5230
2 88633 1 5230
2 88634 1 5230
2 88635 1 5230
2 88636 1 5230
2 88637 1 5230
2 88638 1 5230
2 88639 1 5232
2 88640 1 5232
2 88641 1 5232
2 88642 1 5232
2 88643 1 5234
2 88644 1 5234
2 88645 1 5234
2 88646 1 5234
2 88647 1 5234
2 88648 1 5235
2 88649 1 5235
2 88650 1 5237
2 88651 1 5237
2 88652 1 5237
2 88653 1 5237
2 88654 1 5237
2 88655 1 5238
2 88656 1 5238
2 88657 1 5239
2 88658 1 5239
2 88659 1 5241
2 88660 1 5241
2 88661 1 5241
2 88662 1 5244
2 88663 1 5244
2 88664 1 5245
2 88665 1 5245
2 88666 1 5252
2 88667 1 5252
2 88668 1 5253
2 88669 1 5253
2 88670 1 5255
2 88671 1 5255
2 88672 1 5262
2 88673 1 5262
2 88674 1 5264
2 88675 1 5264
2 88676 1 5264
2 88677 1 5264
2 88678 1 5264
2 88679 1 5264
2 88680 1 5264
2 88681 1 5264
2 88682 1 5264
2 88683 1 5264
2 88684 1 5264
2 88685 1 5265
2 88686 1 5265
2 88687 1 5265
2 88688 1 5265
2 88689 1 5265
2 88690 1 5265
2 88691 1 5265
2 88692 1 5265
2 88693 1 5265
2 88694 1 5265
2 88695 1 5265
2 88696 1 5265
2 88697 1 5266
2 88698 1 5266
2 88699 1 5266
2 88700 1 5277
2 88701 1 5277
2 88702 1 5277
2 88703 1 5277
2 88704 1 5277
2 88705 1 5277
2 88706 1 5277
2 88707 1 5277
2 88708 1 5277
2 88709 1 5277
2 88710 1 5277
2 88711 1 5277
2 88712 1 5278
2 88713 1 5278
2 88714 1 5279
2 88715 1 5279
2 88716 1 5286
2 88717 1 5286
2 88718 1 5286
2 88719 1 5293
2 88720 1 5293
2 88721 1 5293
2 88722 1 5293
2 88723 1 5293
2 88724 1 5294
2 88725 1 5294
2 88726 1 5295
2 88727 1 5295
2 88728 1 5295
2 88729 1 5295
2 88730 1 5295
2 88731 1 5295
2 88732 1 5301
2 88733 1 5301
2 88734 1 5312
2 88735 1 5312
2 88736 1 5312
2 88737 1 5313
2 88738 1 5313
2 88739 1 5315
2 88740 1 5315
2 88741 1 5316
2 88742 1 5316
2 88743 1 5322
2 88744 1 5322
2 88745 1 5323
2 88746 1 5323
2 88747 1 5323
2 88748 1 5334
2 88749 1 5334
2 88750 1 5334
2 88751 1 5334
2 88752 1 5334
2 88753 1 5335
2 88754 1 5335
2 88755 1 5347
2 88756 1 5347
2 88757 1 5347
2 88758 1 5347
2 88759 1 5347
2 88760 1 5347
2 88761 1 5347
2 88762 1 5347
2 88763 1 5347
2 88764 1 5347
2 88765 1 5347
2 88766 1 5347
2 88767 1 5347
2 88768 1 5348
2 88769 1 5348
2 88770 1 5348
2 88771 1 5348
2 88772 1 5348
2 88773 1 5348
2 88774 1 5351
2 88775 1 5351
2 88776 1 5352
2 88777 1 5352
2 88778 1 5352
2 88779 1 5374
2 88780 1 5374
2 88781 1 5375
2 88782 1 5375
2 88783 1 5397
2 88784 1 5397
2 88785 1 5400
2 88786 1 5400
2 88787 1 5400
2 88788 1 5401
2 88789 1 5401
2 88790 1 5401
2 88791 1 5401
2 88792 1 5402
2 88793 1 5402
2 88794 1 5417
2 88795 1 5417
2 88796 1 5418
2 88797 1 5418
2 88798 1 5418
2 88799 1 5418
2 88800 1 5424
2 88801 1 5424
2 88802 1 5425
2 88803 1 5425
2 88804 1 5452
2 88805 1 5452
2 88806 1 5473
2 88807 1 5473
2 88808 1 5474
2 88809 1 5474
2 88810 1 5474
2 88811 1 5479
2 88812 1 5479
2 88813 1 5479
2 88814 1 5479
2 88815 1 5479
2 88816 1 5481
2 88817 1 5481
2 88818 1 5481
2 88819 1 5508
2 88820 1 5508
2 88821 1 5508
2 88822 1 5508
2 88823 1 5508
2 88824 1 5508
2 88825 1 5508
2 88826 1 5508
2 88827 1 5508
2 88828 1 5508
2 88829 1 5509
2 88830 1 5509
2 88831 1 5509
2 88832 1 5509
2 88833 1 5510
2 88834 1 5510
2 88835 1 5511
2 88836 1 5511
2 88837 1 5511
2 88838 1 5514
2 88839 1 5514
2 88840 1 5515
2 88841 1 5515
2 88842 1 5522
2 88843 1 5522
2 88844 1 5523
2 88845 1 5523
2 88846 1 5523
2 88847 1 5547
2 88848 1 5547
2 88849 1 5547
2 88850 1 5547
2 88851 1 5547
2 88852 1 5548
2 88853 1 5548
2 88854 1 5550
2 88855 1 5550
2 88856 1 5563
2 88857 1 5563
2 88858 1 5564
2 88859 1 5564
2 88860 1 5564
2 88861 1 5566
2 88862 1 5566
2 88863 1 5569
2 88864 1 5569
2 88865 1 5569
2 88866 1 5569
2 88867 1 5569
2 88868 1 5569
2 88869 1 5569
2 88870 1 5569
2 88871 1 5569
2 88872 1 5583
2 88873 1 5583
2 88874 1 5586
2 88875 1 5586
2 88876 1 5601
2 88877 1 5601
2 88878 1 5601
2 88879 1 5601
2 88880 1 5601
2 88881 1 5601
2 88882 1 5613
2 88883 1 5613
2 88884 1 5613
2 88885 1 5613
2 88886 1 5613
2 88887 1 5613
2 88888 1 5631
2 88889 1 5631
2 88890 1 5631
2 88891 1 5631
2 88892 1 5631
2 88893 1 5631
2 88894 1 5631
2 88895 1 5631
2 88896 1 5631
2 88897 1 5631
2 88898 1 5631
2 88899 1 5631
2 88900 1 5631
2 88901 1 5631
2 88902 1 5632
2 88903 1 5632
2 88904 1 5632
2 88905 1 5632
2 88906 1 5632
2 88907 1 5633
2 88908 1 5633
2 88909 1 5633
2 88910 1 5633
2 88911 1 5633
2 88912 1 5633
2 88913 1 5633
2 88914 1 5633
2 88915 1 5633
2 88916 1 5633
2 88917 1 5633
2 88918 1 5633
2 88919 1 5633
2 88920 1 5633
2 88921 1 5633
2 88922 1 5633
2 88923 1 5633
2 88924 1 5633
2 88925 1 5633
2 88926 1 5633
2 88927 1 5633
2 88928 1 5633
2 88929 1 5633
2 88930 1 5633
2 88931 1 5633
2 88932 1 5633
2 88933 1 5634
2 88934 1 5634
2 88935 1 5634
2 88936 1 5635
2 88937 1 5635
2 88938 1 5635
2 88939 1 5635
2 88940 1 5635
2 88941 1 5635
2 88942 1 5635
2 88943 1 5635
2 88944 1 5635
2 88945 1 5635
2 88946 1 5635
2 88947 1 5635
2 88948 1 5635
2 88949 1 5635
2 88950 1 5635
2 88951 1 5635
2 88952 1 5635
2 88953 1 5635
2 88954 1 5635
2 88955 1 5635
2 88956 1 5635
2 88957 1 5635
2 88958 1 5635
2 88959 1 5635
2 88960 1 5635
2 88961 1 5635
2 88962 1 5635
2 88963 1 5635
2 88964 1 5635
2 88965 1 5635
2 88966 1 5635
2 88967 1 5635
2 88968 1 5635
2 88969 1 5635
2 88970 1 5635
2 88971 1 5635
2 88972 1 5635
2 88973 1 5635
2 88974 1 5635
2 88975 1 5635
2 88976 1 5635
2 88977 1 5635
2 88978 1 5635
2 88979 1 5635
2 88980 1 5635
2 88981 1 5635
2 88982 1 5635
2 88983 1 5635
2 88984 1 5635
2 88985 1 5635
2 88986 1 5635
2 88987 1 5635
2 88988 1 5635
2 88989 1 5635
2 88990 1 5635
2 88991 1 5635
2 88992 1 5635
2 88993 1 5635
2 88994 1 5635
2 88995 1 5635
2 88996 1 5635
2 88997 1 5635
2 88998 1 5635
2 88999 1 5635
2 89000 1 5635
2 89001 1 5635
2 89002 1 5635
2 89003 1 5635
2 89004 1 5635
2 89005 1 5635
2 89006 1 5635
2 89007 1 5635
2 89008 1 5635
2 89009 1 5636
2 89010 1 5636
2 89011 1 5636
2 89012 1 5636
2 89013 1 5636
2 89014 1 5636
2 89015 1 5636
2 89016 1 5637
2 89017 1 5637
2 89018 1 5640
2 89019 1 5640
2 89020 1 5640
2 89021 1 5642
2 89022 1 5642
2 89023 1 5642
2 89024 1 5642
2 89025 1 5642
2 89026 1 5643
2 89027 1 5643
2 89028 1 5643
2 89029 1 5643
2 89030 1 5645
2 89031 1 5645
2 89032 1 5646
2 89033 1 5646
2 89034 1 5648
2 89035 1 5648
2 89036 1 5648
2 89037 1 5648
2 89038 1 5651
2 89039 1 5651
2 89040 1 5651
2 89041 1 5652
2 89042 1 5652
2 89043 1 5652
2 89044 1 5652
2 89045 1 5652
2 89046 1 5652
2 89047 1 5652
2 89048 1 5652
2 89049 1 5652
2 89050 1 5652
2 89051 1 5652
2 89052 1 5655
2 89053 1 5655
2 89054 1 5665
2 89055 1 5665
2 89056 1 5665
2 89057 1 5665
2 89058 1 5665
2 89059 1 5666
2 89060 1 5666
2 89061 1 5668
2 89062 1 5668
2 89063 1 5668
2 89064 1 5671
2 89065 1 5671
2 89066 1 5671
2 89067 1 5672
2 89068 1 5672
2 89069 1 5679
2 89070 1 5679
2 89071 1 5679
2 89072 1 5680
2 89073 1 5680
2 89074 1 5681
2 89075 1 5681
2 89076 1 5681
2 89077 1 5697
2 89078 1 5697
2 89079 1 5697
2 89080 1 5697
2 89081 1 5697
2 89082 1 5697
2 89083 1 5697
2 89084 1 5697
2 89085 1 5697
2 89086 1 5697
2 89087 1 5697
2 89088 1 5697
2 89089 1 5697
2 89090 1 5697
2 89091 1 5697
2 89092 1 5697
2 89093 1 5698
2 89094 1 5698
2 89095 1 5700
2 89096 1 5700
2 89097 1 5702
2 89098 1 5702
2 89099 1 5708
2 89100 1 5708
2 89101 1 5708
2 89102 1 5708
2 89103 1 5709
2 89104 1 5709
2 89105 1 5710
2 89106 1 5710
2 89107 1 5710
2 89108 1 5710
2 89109 1 5710
2 89110 1 5710
2 89111 1 5724
2 89112 1 5724
2 89113 1 5724
2 89114 1 5724
2 89115 1 5725
2 89116 1 5725
2 89117 1 5725
2 89118 1 5725
2 89119 1 5725
2 89120 1 5725
2 89121 1 5725
2 89122 1 5725
2 89123 1 5725
2 89124 1 5725
2 89125 1 5725
2 89126 1 5725
2 89127 1 5725
2 89128 1 5725
2 89129 1 5725
2 89130 1 5725
2 89131 1 5725
2 89132 1 5725
2 89133 1 5725
2 89134 1 5727
2 89135 1 5727
2 89136 1 5728
2 89137 1 5728
2 89138 1 5728
2 89139 1 5728
2 89140 1 5728
2 89141 1 5728
2 89142 1 5728
2 89143 1 5728
2 89144 1 5728
2 89145 1 5743
2 89146 1 5743
2 89147 1 5748
2 89148 1 5748
2 89149 1 5748
2 89150 1 5748
2 89151 1 5748
2 89152 1 5748
2 89153 1 5748
2 89154 1 5748
2 89155 1 5748
2 89156 1 5748
2 89157 1 5748
2 89158 1 5749
2 89159 1 5749
2 89160 1 5750
2 89161 1 5750
2 89162 1 5762
2 89163 1 5762
2 89164 1 5762
2 89165 1 5762
2 89166 1 5762
2 89167 1 5762
2 89168 1 5762
2 89169 1 5762
2 89170 1 5762
2 89171 1 5762
2 89172 1 5762
2 89173 1 5763
2 89174 1 5763
2 89175 1 5763
2 89176 1 5764
2 89177 1 5764
2 89178 1 5764
2 89179 1 5764
2 89180 1 5764
2 89181 1 5764
2 89182 1 5783
2 89183 1 5783
2 89184 1 5783
2 89185 1 5783
2 89186 1 5783
2 89187 1 5783
2 89188 1 5783
2 89189 1 5783
2 89190 1 5783
2 89191 1 5783
2 89192 1 5784
2 89193 1 5784
2 89194 1 5786
2 89195 1 5786
2 89196 1 5793
2 89197 1 5793
2 89198 1 5809
2 89199 1 5809
2 89200 1 5810
2 89201 1 5810
2 89202 1 5810
2 89203 1 5810
2 89204 1 5810
2 89205 1 5811
2 89206 1 5811
2 89207 1 5811
2 89208 1 5812
2 89209 1 5812
2 89210 1 5812
2 89211 1 5812
2 89212 1 5812
2 89213 1 5812
2 89214 1 5812
2 89215 1 5813
2 89216 1 5813
2 89217 1 5813
2 89218 1 5820
2 89219 1 5820
2 89220 1 5820
2 89221 1 5820
2 89222 1 5827
2 89223 1 5827
2 89224 1 5827
2 89225 1 5836
2 89226 1 5836
2 89227 1 5844
2 89228 1 5844
2 89229 1 5850
2 89230 1 5850
2 89231 1 5850
2 89232 1 5850
2 89233 1 5850
2 89234 1 5850
2 89235 1 5850
2 89236 1 5850
2 89237 1 5859
2 89238 1 5859
2 89239 1 5859
2 89240 1 5860
2 89241 1 5860
2 89242 1 5860
2 89243 1 5860
2 89244 1 5861
2 89245 1 5861
2 89246 1 5861
2 89247 1 5861
2 89248 1 5861
2 89249 1 5861
2 89250 1 5868
2 89251 1 5868
2 89252 1 5868
2 89253 1 5870
2 89254 1 5870
2 89255 1 5870
2 89256 1 5870
2 89257 1 5870
2 89258 1 5870
2 89259 1 5870
2 89260 1 5873
2 89261 1 5873
2 89262 1 5886
2 89263 1 5886
2 89264 1 5886
2 89265 1 5886
2 89266 1 5887
2 89267 1 5887
2 89268 1 5887
2 89269 1 5888
2 89270 1 5888
2 89271 1 5889
2 89272 1 5889
2 89273 1 5889
2 89274 1 5889
2 89275 1 5889
2 89276 1 5889
2 89277 1 5889
2 89278 1 5890
2 89279 1 5890
2 89280 1 5890
2 89281 1 5890
2 89282 1 5895
2 89283 1 5895
2 89284 1 5896
2 89285 1 5896
2 89286 1 5905
2 89287 1 5905
2 89288 1 5905
2 89289 1 5905
2 89290 1 5905
2 89291 1 5905
2 89292 1 5905
2 89293 1 5905
2 89294 1 5905
2 89295 1 5905
2 89296 1 5905
2 89297 1 5905
2 89298 1 5909
2 89299 1 5909
2 89300 1 5909
2 89301 1 5909
2 89302 1 5909
2 89303 1 5909
2 89304 1 5909
2 89305 1 5909
2 89306 1 5909
2 89307 1 5909
2 89308 1 5909
2 89309 1 5909
2 89310 1 5909
2 89311 1 5909
2 89312 1 5909
2 89313 1 5909
2 89314 1 5909
2 89315 1 5909
2 89316 1 5909
2 89317 1 5909
2 89318 1 5910
2 89319 1 5910
2 89320 1 5910
2 89321 1 5910
2 89322 1 5910
2 89323 1 5910
2 89324 1 5910
2 89325 1 5910
2 89326 1 5914
2 89327 1 5914
2 89328 1 5914
2 89329 1 5917
2 89330 1 5917
2 89331 1 5917
2 89332 1 5917
2 89333 1 5917
2 89334 1 5917
2 89335 1 5917
2 89336 1 5917
2 89337 1 5924
2 89338 1 5924
2 89339 1 5931
2 89340 1 5931
2 89341 1 5931
2 89342 1 5931
2 89343 1 5939
2 89344 1 5939
2 89345 1 5939
2 89346 1 5939
2 89347 1 5939
2 89348 1 5939
2 89349 1 5939
2 89350 1 5939
2 89351 1 5939
2 89352 1 5939
2 89353 1 5939
2 89354 1 5939
2 89355 1 5939
2 89356 1 5939
2 89357 1 5939
2 89358 1 5939
2 89359 1 5939
2 89360 1 5940
2 89361 1 5940
2 89362 1 5940
2 89363 1 5940
2 89364 1 5940
2 89365 1 5940
2 89366 1 5940
2 89367 1 5941
2 89368 1 5941
2 89369 1 5950
2 89370 1 5950
2 89371 1 5950
2 89372 1 5950
2 89373 1 5951
2 89374 1 5951
2 89375 1 5952
2 89376 1 5952
2 89377 1 5953
2 89378 1 5953
2 89379 1 5965
2 89380 1 5965
2 89381 1 5965
2 89382 1 5965
2 89383 1 5965
2 89384 1 5965
2 89385 1 5965
2 89386 1 5966
2 89387 1 5966
2 89388 1 5966
2 89389 1 5966
2 89390 1 5966
2 89391 1 5966
2 89392 1 5966
2 89393 1 5966
2 89394 1 5966
2 89395 1 5966
2 89396 1 5966
2 89397 1 5966
2 89398 1 5966
2 89399 1 5966
2 89400 1 5967
2 89401 1 5967
2 89402 1 5967
2 89403 1 5970
2 89404 1 5970
2 89405 1 5970
2 89406 1 5970
2 89407 1 5970
2 89408 1 5970
2 89409 1 5970
2 89410 1 5970
2 89411 1 5970
2 89412 1 5978
2 89413 1 5978
2 89414 1 5978
2 89415 1 5978
2 89416 1 5978
2 89417 1 5978
2 89418 1 5978
2 89419 1 5980
2 89420 1 5980
2 89421 1 5980
2 89422 1 5981
2 89423 1 5981
2 89424 1 5981
2 89425 1 5981
2 89426 1 5998
2 89427 1 5998
2 89428 1 5998
2 89429 1 5998
2 89430 1 5998
2 89431 1 5998
2 89432 1 5999
2 89433 1 5999
2 89434 1 5999
2 89435 1 5999
2 89436 1 6004
2 89437 1 6004
2 89438 1 6004
2 89439 1 6004
2 89440 1 6004
2 89441 1 6004
2 89442 1 6014
2 89443 1 6014
2 89444 1 6015
2 89445 1 6015
2 89446 1 6037
2 89447 1 6037
2 89448 1 6040
2 89449 1 6040
2 89450 1 6041
2 89451 1 6041
2 89452 1 6041
2 89453 1 6042
2 89454 1 6042
2 89455 1 6050
2 89456 1 6050
2 89457 1 6050
2 89458 1 6050
2 89459 1 6050
2 89460 1 6050
2 89461 1 6061
2 89462 1 6061
2 89463 1 6061
2 89464 1 6061
2 89465 1 6061
2 89466 1 6061
2 89467 1 6061
2 89468 1 6061
2 89469 1 6061
2 89470 1 6061
2 89471 1 6061
2 89472 1 6061
2 89473 1 6061
2 89474 1 6061
2 89475 1 6071
2 89476 1 6071
2 89477 1 6073
2 89478 1 6073
2 89479 1 6073
2 89480 1 6073
2 89481 1 6073
2 89482 1 6073
2 89483 1 6078
2 89484 1 6078
2 89485 1 6087
2 89486 1 6087
2 89487 1 6087
2 89488 1 6088
2 89489 1 6088
2 89490 1 6091
2 89491 1 6091
2 89492 1 6091
2 89493 1 6109
2 89494 1 6109
2 89495 1 6109
2 89496 1 6109
2 89497 1 6109
2 89498 1 6109
2 89499 1 6109
2 89500 1 6109
2 89501 1 6111
2 89502 1 6111
2 89503 1 6111
2 89504 1 6111
2 89505 1 6111
2 89506 1 6111
2 89507 1 6111
2 89508 1 6111
2 89509 1 6111
2 89510 1 6111
2 89511 1 6111
2 89512 1 6111
2 89513 1 6111
2 89514 1 6111
2 89515 1 6111
2 89516 1 6111
2 89517 1 6111
2 89518 1 6111
2 89519 1 6111
2 89520 1 6111
2 89521 1 6111
2 89522 1 6111
2 89523 1 6111
2 89524 1 6111
2 89525 1 6111
2 89526 1 6111
2 89527 1 6111
2 89528 1 6112
2 89529 1 6112
2 89530 1 6112
2 89531 1 6114
2 89532 1 6114
2 89533 1 6114
2 89534 1 6114
2 89535 1 6114
2 89536 1 6114
2 89537 1 6114
2 89538 1 6114
2 89539 1 6114
2 89540 1 6114
2 89541 1 6114
2 89542 1 6114
2 89543 1 6114
2 89544 1 6114
2 89545 1 6114
2 89546 1 6114
2 89547 1 6114
2 89548 1 6114
2 89549 1 6114
2 89550 1 6114
2 89551 1 6114
2 89552 1 6114
2 89553 1 6115
2 89554 1 6115
2 89555 1 6115
2 89556 1 6115
2 89557 1 6115
2 89558 1 6116
2 89559 1 6116
2 89560 1 6119
2 89561 1 6119
2 89562 1 6119
2 89563 1 6119
2 89564 1 6119
2 89565 1 6119
2 89566 1 6119
2 89567 1 6119
2 89568 1 6119
2 89569 1 6119
2 89570 1 6119
2 89571 1 6119
2 89572 1 6119
2 89573 1 6119
2 89574 1 6119
2 89575 1 6119
2 89576 1 6119
2 89577 1 6119
2 89578 1 6119
2 89579 1 6119
2 89580 1 6119
2 89581 1 6119
2 89582 1 6119
2 89583 1 6119
2 89584 1 6119
2 89585 1 6119
2 89586 1 6119
2 89587 1 6119
2 89588 1 6119
2 89589 1 6119
2 89590 1 6119
2 89591 1 6119
2 89592 1 6120
2 89593 1 6120
2 89594 1 6120
2 89595 1 6124
2 89596 1 6124
2 89597 1 6124
2 89598 1 6140
2 89599 1 6140
2 89600 1 6143
2 89601 1 6143
2 89602 1 6146
2 89603 1 6146
2 89604 1 6146
2 89605 1 6146
2 89606 1 6146
2 89607 1 6146
2 89608 1 6146
2 89609 1 6147
2 89610 1 6147
2 89611 1 6159
2 89612 1 6159
2 89613 1 6159
2 89614 1 6160
2 89615 1 6160
2 89616 1 6168
2 89617 1 6168
2 89618 1 6168
2 89619 1 6169
2 89620 1 6169
2 89621 1 6170
2 89622 1 6170
2 89623 1 6170
2 89624 1 6171
2 89625 1 6171
2 89626 1 6172
2 89627 1 6172
2 89628 1 6172
2 89629 1 6172
2 89630 1 6172
2 89631 1 6172
2 89632 1 6172
2 89633 1 6172
2 89634 1 6172
2 89635 1 6172
2 89636 1 6173
2 89637 1 6173
2 89638 1 6173
2 89639 1 6173
2 89640 1 6173
2 89641 1 6173
2 89642 1 6173
2 89643 1 6173
2 89644 1 6177
2 89645 1 6177
2 89646 1 6177
2 89647 1 6177
2 89648 1 6178
2 89649 1 6178
2 89650 1 6183
2 89651 1 6183
2 89652 1 6187
2 89653 1 6187
2 89654 1 6190
2 89655 1 6190
2 89656 1 6190
2 89657 1 6198
2 89658 1 6198
2 89659 1 6202
2 89660 1 6202
2 89661 1 6211
2 89662 1 6211
2 89663 1 6211
2 89664 1 6212
2 89665 1 6212
2 89666 1 6213
2 89667 1 6213
2 89668 1 6222
2 89669 1 6222
2 89670 1 6222
2 89671 1 6222
2 89672 1 6222
2 89673 1 6222
2 89674 1 6222
2 89675 1 6222
2 89676 1 6222
2 89677 1 6222
2 89678 1 6222
2 89679 1 6223
2 89680 1 6223
2 89681 1 6223
2 89682 1 6223
2 89683 1 6223
2 89684 1 6223
2 89685 1 6232
2 89686 1 6232
2 89687 1 6232
2 89688 1 6232
2 89689 1 6232
2 89690 1 6232
2 89691 1 6232
2 89692 1 6232
2 89693 1 6232
2 89694 1 6232
2 89695 1 6232
2 89696 1 6238
2 89697 1 6238
2 89698 1 6239
2 89699 1 6239
2 89700 1 6239
2 89701 1 6239
2 89702 1 6239
2 89703 1 6239
2 89704 1 6241
2 89705 1 6241
2 89706 1 6241
2 89707 1 6241
2 89708 1 6241
2 89709 1 6242
2 89710 1 6242
2 89711 1 6242
2 89712 1 6251
2 89713 1 6251
2 89714 1 6253
2 89715 1 6253
2 89716 1 6253
2 89717 1 6253
2 89718 1 6253
2 89719 1 6253
2 89720 1 6259
2 89721 1 6259
2 89722 1 6260
2 89723 1 6260
2 89724 1 6260
2 89725 1 6260
2 89726 1 6260
2 89727 1 6260
2 89728 1 6260
2 89729 1 6261
2 89730 1 6261
2 89731 1 6261
2 89732 1 6261
2 89733 1 6261
2 89734 1 6262
2 89735 1 6262
2 89736 1 6263
2 89737 1 6263
2 89738 1 6263
2 89739 1 6264
2 89740 1 6264
2 89741 1 6264
2 89742 1 6264
2 89743 1 6264
2 89744 1 6266
2 89745 1 6266
2 89746 1 6287
2 89747 1 6287
2 89748 1 6287
2 89749 1 6287
2 89750 1 6288
2 89751 1 6288
2 89752 1 6289
2 89753 1 6289
2 89754 1 6289
2 89755 1 6289
2 89756 1 6289
2 89757 1 6289
2 89758 1 6289
2 89759 1 6290
2 89760 1 6290
2 89761 1 6290
2 89762 1 6290
2 89763 1 6290
2 89764 1 6291
2 89765 1 6291
2 89766 1 6291
2 89767 1 6294
2 89768 1 6294
2 89769 1 6294
2 89770 1 6294
2 89771 1 6294
2 89772 1 6303
2 89773 1 6303
2 89774 1 6303
2 89775 1 6303
2 89776 1 6303
2 89777 1 6303
2 89778 1 6303
2 89779 1 6307
2 89780 1 6307
2 89781 1 6319
2 89782 1 6319
2 89783 1 6319
2 89784 1 6326
2 89785 1 6326
2 89786 1 6339
2 89787 1 6339
2 89788 1 6339
2 89789 1 6339
2 89790 1 6339
2 89791 1 6342
2 89792 1 6342
2 89793 1 6342
2 89794 1 6342
2 89795 1 6343
2 89796 1 6343
2 89797 1 6343
2 89798 1 6348
2 89799 1 6348
2 89800 1 6361
2 89801 1 6361
2 89802 1 6361
2 89803 1 6361
2 89804 1 6363
2 89805 1 6363
2 89806 1 6372
2 89807 1 6372
2 89808 1 6372
2 89809 1 6372
2 89810 1 6372
2 89811 1 6382
2 89812 1 6382
2 89813 1 6382
2 89814 1 6382
2 89815 1 6382
2 89816 1 6382
2 89817 1 6382
2 89818 1 6382
2 89819 1 6383
2 89820 1 6383
2 89821 1 6384
2 89822 1 6384
2 89823 1 6385
2 89824 1 6385
2 89825 1 6385
2 89826 1 6385
2 89827 1 6385
2 89828 1 6386
2 89829 1 6386
2 89830 1 6386
2 89831 1 6388
2 89832 1 6388
2 89833 1 6389
2 89834 1 6389
2 89835 1 6391
2 89836 1 6391
2 89837 1 6419
2 89838 1 6419
2 89839 1 6419
2 89840 1 6432
2 89841 1 6432
2 89842 1 6432
2 89843 1 6432
2 89844 1 6432
2 89845 1 6432
2 89846 1 6433
2 89847 1 6433
2 89848 1 6433
2 89849 1 6433
2 89850 1 6435
2 89851 1 6435
2 89852 1 6450
2 89853 1 6450
2 89854 1 6451
2 89855 1 6451
2 89856 1 6451
2 89857 1 6462
2 89858 1 6462
2 89859 1 6462
2 89860 1 6471
2 89861 1 6471
2 89862 1 6471
2 89863 1 6471
2 89864 1 6471
2 89865 1 6471
2 89866 1 6471
2 89867 1 6471
2 89868 1 6471
2 89869 1 6471
2 89870 1 6471
2 89871 1 6471
2 89872 1 6471
2 89873 1 6471
2 89874 1 6472
2 89875 1 6472
2 89876 1 6472
2 89877 1 6472
2 89878 1 6472
2 89879 1 6472
2 89880 1 6472
2 89881 1 6474
2 89882 1 6474
2 89883 1 6474
2 89884 1 6474
2 89885 1 6474
2 89886 1 6475
2 89887 1 6475
2 89888 1 6486
2 89889 1 6486
2 89890 1 6493
2 89891 1 6493
2 89892 1 6493
2 89893 1 6493
2 89894 1 6493
2 89895 1 6493
2 89896 1 6493
2 89897 1 6493
2 89898 1 6493
2 89899 1 6493
2 89900 1 6493
2 89901 1 6493
2 89902 1 6493
2 89903 1 6494
2 89904 1 6494
2 89905 1 6494
2 89906 1 6494
2 89907 1 6494
2 89908 1 6494
2 89909 1 6494
2 89910 1 6502
2 89911 1 6502
2 89912 1 6502
2 89913 1 6502
2 89914 1 6502
2 89915 1 6502
2 89916 1 6502
2 89917 1 6502
2 89918 1 6502
2 89919 1 6522
2 89920 1 6522
2 89921 1 6522
2 89922 1 6523
2 89923 1 6523
2 89924 1 6523
2 89925 1 6523
2 89926 1 6523
2 89927 1 6523
2 89928 1 6523
2 89929 1 6523
2 89930 1 6523
2 89931 1 6523
2 89932 1 6523
2 89933 1 6525
2 89934 1 6525
2 89935 1 6531
2 89936 1 6531
2 89937 1 6539
2 89938 1 6539
2 89939 1 6539
2 89940 1 6539
2 89941 1 6540
2 89942 1 6540
2 89943 1 6551
2 89944 1 6551
2 89945 1 6551
2 89946 1 6552
2 89947 1 6552
2 89948 1 6552
2 89949 1 6554
2 89950 1 6554
2 89951 1 6578
2 89952 1 6578
2 89953 1 6578
2 89954 1 6578
2 89955 1 6578
2 89956 1 6578
2 89957 1 6582
2 89958 1 6582
2 89959 1 6600
2 89960 1 6600
2 89961 1 6600
2 89962 1 6601
2 89963 1 6601
2 89964 1 6610
2 89965 1 6610
2 89966 1 6616
2 89967 1 6616
2 89968 1 6616
2 89969 1 6619
2 89970 1 6619
2 89971 1 6626
2 89972 1 6626
2 89973 1 6626
2 89974 1 6628
2 89975 1 6628
2 89976 1 6647
2 89977 1 6647
2 89978 1 6650
2 89979 1 6650
2 89980 1 6650
2 89981 1 6650
2 89982 1 6650
2 89983 1 6650
2 89984 1 6650
2 89985 1 6650
2 89986 1 6650
2 89987 1 6650
2 89988 1 6650
2 89989 1 6650
2 89990 1 6650
2 89991 1 6651
2 89992 1 6651
2 89993 1 6651
2 89994 1 6651
2 89995 1 6651
2 89996 1 6658
2 89997 1 6658
2 89998 1 6658
2 89999 1 6668
2 90000 1 6668
2 90001 1 6678
2 90002 1 6678
2 90003 1 6679
2 90004 1 6679
2 90005 1 6679
2 90006 1 6679
2 90007 1 6680
2 90008 1 6680
2 90009 1 6680
2 90010 1 6680
2 90011 1 6688
2 90012 1 6688
2 90013 1 6693
2 90014 1 6693
2 90015 1 6693
2 90016 1 6693
2 90017 1 6694
2 90018 1 6694
2 90019 1 6694
2 90020 1 6696
2 90021 1 6696
2 90022 1 6713
2 90023 1 6713
2 90024 1 6718
2 90025 1 6718
2 90026 1 6718
2 90027 1 6718
2 90028 1 6718
2 90029 1 6718
2 90030 1 6718
2 90031 1 6718
2 90032 1 6718
2 90033 1 6718
2 90034 1 6726
2 90035 1 6726
2 90036 1 6726
2 90037 1 6726
2 90038 1 6727
2 90039 1 6727
2 90040 1 6727
2 90041 1 6727
2 90042 1 6727
2 90043 1 6727
2 90044 1 6727
2 90045 1 6727
2 90046 1 6727
2 90047 1 6727
2 90048 1 6727
2 90049 1 6727
2 90050 1 6728
2 90051 1 6728
2 90052 1 6728
2 90053 1 6728
2 90054 1 6728
2 90055 1 6729
2 90056 1 6729
2 90057 1 6729
2 90058 1 6737
2 90059 1 6737
2 90060 1 6737
2 90061 1 6746
2 90062 1 6746
2 90063 1 6746
2 90064 1 6746
2 90065 1 6746
2 90066 1 6746
2 90067 1 6746
2 90068 1 6746
2 90069 1 6746
2 90070 1 6746
2 90071 1 6746
2 90072 1 6746
2 90073 1 6746
2 90074 1 6746
2 90075 1 6746
2 90076 1 6746
2 90077 1 6746
2 90078 1 6746
2 90079 1 6746
2 90080 1 6746
2 90081 1 6746
2 90082 1 6746
2 90083 1 6746
2 90084 1 6746
2 90085 1 6746
2 90086 1 6746
2 90087 1 6746
2 90088 1 6747
2 90089 1 6747
2 90090 1 6747
2 90091 1 6747
2 90092 1 6747
2 90093 1 6748
2 90094 1 6748
2 90095 1 6751
2 90096 1 6751
2 90097 1 6751
2 90098 1 6751
2 90099 1 6751
2 90100 1 6752
2 90101 1 6752
2 90102 1 6753
2 90103 1 6753
2 90104 1 6753
2 90105 1 6753
2 90106 1 6753
2 90107 1 6753
2 90108 1 6754
2 90109 1 6754
2 90110 1 6754
2 90111 1 6754
2 90112 1 6754
2 90113 1 6754
2 90114 1 6754
2 90115 1 6754
2 90116 1 6754
2 90117 1 6756
2 90118 1 6756
2 90119 1 6756
2 90120 1 6756
2 90121 1 6757
2 90122 1 6757
2 90123 1 6757
2 90124 1 6757
2 90125 1 6768
2 90126 1 6768
2 90127 1 6768
2 90128 1 6768
2 90129 1 6768
2 90130 1 6768
2 90131 1 6779
2 90132 1 6779
2 90133 1 6780
2 90134 1 6780
2 90135 1 6802
2 90136 1 6802
2 90137 1 6810
2 90138 1 6810
2 90139 1 6810
2 90140 1 6814
2 90141 1 6814
2 90142 1 6814
2 90143 1 6814
2 90144 1 6837
2 90145 1 6837
2 90146 1 6837
2 90147 1 6837
2 90148 1 6837
2 90149 1 6838
2 90150 1 6838
2 90151 1 6838
2 90152 1 6847
2 90153 1 6847
2 90154 1 6850
2 90155 1 6850
2 90156 1 6851
2 90157 1 6851
2 90158 1 6872
2 90159 1 6872
2 90160 1 6873
2 90161 1 6873
2 90162 1 6875
2 90163 1 6875
2 90164 1 6889
2 90165 1 6889
2 90166 1 6889
2 90167 1 6900
2 90168 1 6900
2 90169 1 6900
2 90170 1 6900
2 90171 1 6900
2 90172 1 6900
2 90173 1 6900
2 90174 1 6900
2 90175 1 6900
2 90176 1 6900
2 90177 1 6901
2 90178 1 6901
2 90179 1 6901
2 90180 1 6903
2 90181 1 6903
2 90182 1 6903
2 90183 1 6903
2 90184 1 6904
2 90185 1 6904
2 90186 1 6904
2 90187 1 6904
2 90188 1 6904
2 90189 1 6904
2 90190 1 6904
2 90191 1 6904
2 90192 1 6904
2 90193 1 6904
2 90194 1 6904
2 90195 1 6906
2 90196 1 6906
2 90197 1 6906
2 90198 1 6907
2 90199 1 6907
2 90200 1 6908
2 90201 1 6908
2 90202 1 6909
2 90203 1 6909
2 90204 1 6909
2 90205 1 6918
2 90206 1 6918
2 90207 1 6934
2 90208 1 6934
2 90209 1 6934
2 90210 1 6934
2 90211 1 6934
2 90212 1 6934
2 90213 1 6934
2 90214 1 6934
2 90215 1 6935
2 90216 1 6935
2 90217 1 6935
2 90218 1 6935
2 90219 1 6935
2 90220 1 6935
2 90221 1 6936
2 90222 1 6936
2 90223 1 6937
2 90224 1 6937
2 90225 1 6943
2 90226 1 6943
2 90227 1 6943
2 90228 1 6960
2 90229 1 6960
2 90230 1 6960
2 90231 1 6960
2 90232 1 6960
2 90233 1 6960
2 90234 1 6960
2 90235 1 6980
2 90236 1 6980
2 90237 1 6980
2 90238 1 6989
2 90239 1 6989
2 90240 1 6990
2 90241 1 6990
2 90242 1 6991
2 90243 1 6991
2 90244 1 6991
2 90245 1 7000
2 90246 1 7000
2 90247 1 7010
2 90248 1 7010
2 90249 1 7010
2 90250 1 7010
2 90251 1 7010
2 90252 1 7010
2 90253 1 7010
2 90254 1 7010
2 90255 1 7011
2 90256 1 7011
2 90257 1 7019
2 90258 1 7019
2 90259 1 7019
2 90260 1 7020
2 90261 1 7020
2 90262 1 7020
2 90263 1 7020
2 90264 1 7028
2 90265 1 7028
2 90266 1 7028
2 90267 1 7028
2 90268 1 7028
2 90269 1 7028
2 90270 1 7028
2 90271 1 7028
2 90272 1 7028
2 90273 1 7029
2 90274 1 7029
2 90275 1 7036
2 90276 1 7036
2 90277 1 7043
2 90278 1 7043
2 90279 1 7047
2 90280 1 7047
2 90281 1 7048
2 90282 1 7048
2 90283 1 7048
2 90284 1 7048
2 90285 1 7048
2 90286 1 7048
2 90287 1 7048
2 90288 1 7048
2 90289 1 7048
2 90290 1 7048
2 90291 1 7048
2 90292 1 7048
2 90293 1 7049
2 90294 1 7049
2 90295 1 7049
2 90296 1 7049
2 90297 1 7050
2 90298 1 7050
2 90299 1 7059
2 90300 1 7059
2 90301 1 7060
2 90302 1 7060
2 90303 1 7060
2 90304 1 7060
2 90305 1 7060
2 90306 1 7067
2 90307 1 7067
2 90308 1 7067
2 90309 1 7067
2 90310 1 7069
2 90311 1 7069
2 90312 1 7069
2 90313 1 7069
2 90314 1 7069
2 90315 1 7069
2 90316 1 7069
2 90317 1 7069
2 90318 1 7069
2 90319 1 7069
2 90320 1 7069
2 90321 1 7069
2 90322 1 7069
2 90323 1 7069
2 90324 1 7070
2 90325 1 7070
2 90326 1 7070
2 90327 1 7070
2 90328 1 7070
2 90329 1 7070
2 90330 1 7070
2 90331 1 7075
2 90332 1 7075
2 90333 1 7075
2 90334 1 7075
2 90335 1 7075
2 90336 1 7075
2 90337 1 7075
2 90338 1 7075
2 90339 1 7075
2 90340 1 7075
2 90341 1 7075
2 90342 1 7075
2 90343 1 7076
2 90344 1 7076
2 90345 1 7076
2 90346 1 7076
2 90347 1 7076
2 90348 1 7076
2 90349 1 7076
2 90350 1 7076
2 90351 1 7076
2 90352 1 7076
2 90353 1 7076
2 90354 1 7076
2 90355 1 7076
2 90356 1 7085
2 90357 1 7085
2 90358 1 7085
2 90359 1 7086
2 90360 1 7086
2 90361 1 7086
2 90362 1 7087
2 90363 1 7087
2 90364 1 7087
2 90365 1 7087
2 90366 1 7087
2 90367 1 7087
2 90368 1 7087
2 90369 1 7088
2 90370 1 7088
2 90371 1 7088
2 90372 1 7088
2 90373 1 7088
2 90374 1 7088
2 90375 1 7088
2 90376 1 7089
2 90377 1 7089
2 90378 1 7089
2 90379 1 7090
2 90380 1 7090
2 90381 1 7090
2 90382 1 7090
2 90383 1 7090
2 90384 1 7090
2 90385 1 7092
2 90386 1 7092
2 90387 1 7095
2 90388 1 7095
2 90389 1 7095
2 90390 1 7095
2 90391 1 7095
2 90392 1 7095
2 90393 1 7095
2 90394 1 7095
2 90395 1 7095
2 90396 1 7095
2 90397 1 7095
2 90398 1 7095
2 90399 1 7095
2 90400 1 7096
2 90401 1 7096
2 90402 1 7097
2 90403 1 7097
2 90404 1 7097
2 90405 1 7097
2 90406 1 7097
2 90407 1 7097
2 90408 1 7097
2 90409 1 7097
2 90410 1 7098
2 90411 1 7098
2 90412 1 7100
2 90413 1 7100
2 90414 1 7104
2 90415 1 7104
2 90416 1 7104
2 90417 1 7104
2 90418 1 7104
2 90419 1 7104
2 90420 1 7104
2 90421 1 7104
2 90422 1 7105
2 90423 1 7105
2 90424 1 7105
2 90425 1 7105
2 90426 1 7105
2 90427 1 7105
2 90428 1 7105
2 90429 1 7106
2 90430 1 7106
2 90431 1 7106
2 90432 1 7107
2 90433 1 7107
2 90434 1 7107
2 90435 1 7107
2 90436 1 7109
2 90437 1 7109
2 90438 1 7109
2 90439 1 7109
2 90440 1 7110
2 90441 1 7110
2 90442 1 7111
2 90443 1 7111
2 90444 1 7111
2 90445 1 7111
2 90446 1 7111
2 90447 1 7111
2 90448 1 7111
2 90449 1 7111
2 90450 1 7112
2 90451 1 7112
2 90452 1 7124
2 90453 1 7124
2 90454 1 7124
2 90455 1 7126
2 90456 1 7126
2 90457 1 7126
2 90458 1 7126
2 90459 1 7134
2 90460 1 7134
2 90461 1 7142
2 90462 1 7142
2 90463 1 7142
2 90464 1 7142
2 90465 1 7142
2 90466 1 7142
2 90467 1 7143
2 90468 1 7143
2 90469 1 7143
2 90470 1 7143
2 90471 1 7143
2 90472 1 7143
2 90473 1 7143
2 90474 1 7143
2 90475 1 7143
2 90476 1 7143
2 90477 1 7143
2 90478 1 7143
2 90479 1 7143
2 90480 1 7143
2 90481 1 7143
2 90482 1 7143
2 90483 1 7143
2 90484 1 7143
2 90485 1 7146
2 90486 1 7146
2 90487 1 7146
2 90488 1 7146
2 90489 1 7146
2 90490 1 7146
2 90491 1 7146
2 90492 1 7146
2 90493 1 7146
2 90494 1 7146
2 90495 1 7146
2 90496 1 7158
2 90497 1 7158
2 90498 1 7162
2 90499 1 7162
2 90500 1 7162
2 90501 1 7163
2 90502 1 7163
2 90503 1 7163
2 90504 1 7163
2 90505 1 7178
2 90506 1 7178
2 90507 1 7178
2 90508 1 7179
2 90509 1 7179
2 90510 1 7180
2 90511 1 7180
2 90512 1 7180
2 90513 1 7180
2 90514 1 7180
2 90515 1 7180
2 90516 1 7180
2 90517 1 7180
2 90518 1 7180
2 90519 1 7181
2 90520 1 7181
2 90521 1 7181
2 90522 1 7181
2 90523 1 7181
2 90524 1 7181
2 90525 1 7181
2 90526 1 7181
2 90527 1 7182
2 90528 1 7182
2 90529 1 7182
2 90530 1 7182
2 90531 1 7182
2 90532 1 7182
2 90533 1 7182
2 90534 1 7182
2 90535 1 7182
2 90536 1 7182
2 90537 1 7190
2 90538 1 7190
2 90539 1 7190
2 90540 1 7190
2 90541 1 7190
2 90542 1 7193
2 90543 1 7193
2 90544 1 7193
2 90545 1 7193
2 90546 1 7193
2 90547 1 7202
2 90548 1 7202
2 90549 1 7202
2 90550 1 7202
2 90551 1 7202
2 90552 1 7202
2 90553 1 7202
2 90554 1 7202
2 90555 1 7204
2 90556 1 7204
2 90557 1 7215
2 90558 1 7215
2 90559 1 7217
2 90560 1 7217
2 90561 1 7217
2 90562 1 7222
2 90563 1 7222
2 90564 1 7223
2 90565 1 7223
2 90566 1 7231
2 90567 1 7231
2 90568 1 7231
2 90569 1 7231
2 90570 1 7235
2 90571 1 7235
2 90572 1 7235
2 90573 1 7235
2 90574 1 7235
2 90575 1 7235
2 90576 1 7235
2 90577 1 7235
2 90578 1 7235
2 90579 1 7235
2 90580 1 7235
2 90581 1 7235
2 90582 1 7235
2 90583 1 7235
2 90584 1 7235
2 90585 1 7235
2 90586 1 7235
2 90587 1 7235
2 90588 1 7235
2 90589 1 7235
2 90590 1 7235
2 90591 1 7235
2 90592 1 7235
2 90593 1 7235
2 90594 1 7235
2 90595 1 7236
2 90596 1 7236
2 90597 1 7236
2 90598 1 7236
2 90599 1 7236
2 90600 1 7236
2 90601 1 7237
2 90602 1 7237
2 90603 1 7238
2 90604 1 7238
2 90605 1 7238
2 90606 1 7238
2 90607 1 7238
2 90608 1 7238
2 90609 1 7239
2 90610 1 7239
2 90611 1 7247
2 90612 1 7247
2 90613 1 7256
2 90614 1 7256
2 90615 1 7256
2 90616 1 7256
2 90617 1 7257
2 90618 1 7257
2 90619 1 7262
2 90620 1 7262
2 90621 1 7270
2 90622 1 7270
2 90623 1 7270
2 90624 1 7270
2 90625 1 7270
2 90626 1 7271
2 90627 1 7271
2 90628 1 7271
2 90629 1 7271
2 90630 1 7271
2 90631 1 7272
2 90632 1 7272
2 90633 1 7273
2 90634 1 7273
2 90635 1 7273
2 90636 1 7274
2 90637 1 7274
2 90638 1 7274
2 90639 1 7274
2 90640 1 7274
2 90641 1 7274
2 90642 1 7286
2 90643 1 7286
2 90644 1 7287
2 90645 1 7287
2 90646 1 7287
2 90647 1 7287
2 90648 1 7287
2 90649 1 7287
2 90650 1 7287
2 90651 1 7287
2 90652 1 7288
2 90653 1 7288
2 90654 1 7288
2 90655 1 7288
2 90656 1 7296
2 90657 1 7296
2 90658 1 7296
2 90659 1 7296
2 90660 1 7297
2 90661 1 7297
2 90662 1 7297
2 90663 1 7297
2 90664 1 7297
2 90665 1 7297
2 90666 1 7306
2 90667 1 7306
2 90668 1 7309
2 90669 1 7309
2 90670 1 7309
2 90671 1 7309
2 90672 1 7310
2 90673 1 7310
2 90674 1 7310
2 90675 1 7311
2 90676 1 7311
2 90677 1 7311
2 90678 1 7311
2 90679 1 7320
2 90680 1 7320
2 90681 1 7321
2 90682 1 7321
2 90683 1 7321
2 90684 1 7321
2 90685 1 7339
2 90686 1 7339
2 90687 1 7340
2 90688 1 7340
2 90689 1 7340
2 90690 1 7340
2 90691 1 7340
2 90692 1 7340
2 90693 1 7340
2 90694 1 7340
2 90695 1 7340
2 90696 1 7340
2 90697 1 7341
2 90698 1 7341
2 90699 1 7341
2 90700 1 7341
2 90701 1 7341
2 90702 1 7341
2 90703 1 7341
2 90704 1 7341
2 90705 1 7346
2 90706 1 7346
2 90707 1 7346
2 90708 1 7346
2 90709 1 7346
2 90710 1 7346
2 90711 1 7346
2 90712 1 7347
2 90713 1 7347
2 90714 1 7347
2 90715 1 7347
2 90716 1 7347
2 90717 1 7347
2 90718 1 7347
2 90719 1 7347
2 90720 1 7347
2 90721 1 7347
2 90722 1 7347
2 90723 1 7347
2 90724 1 7363
2 90725 1 7363
2 90726 1 7364
2 90727 1 7364
2 90728 1 7365
2 90729 1 7365
2 90730 1 7365
2 90731 1 7365
2 90732 1 7365
2 90733 1 7369
2 90734 1 7369
2 90735 1 7369
2 90736 1 7369
2 90737 1 7370
2 90738 1 7370
2 90739 1 7370
2 90740 1 7370
2 90741 1 7383
2 90742 1 7383
2 90743 1 7383
2 90744 1 7383
2 90745 1 7383
2 90746 1 7383
2 90747 1 7383
2 90748 1 7383
2 90749 1 7384
2 90750 1 7384
2 90751 1 7384
2 90752 1 7384
2 90753 1 7384
2 90754 1 7384
2 90755 1 7384
2 90756 1 7384
2 90757 1 7385
2 90758 1 7385
2 90759 1 7385
2 90760 1 7385
2 90761 1 7397
2 90762 1 7397
2 90763 1 7397
2 90764 1 7397
2 90765 1 7397
2 90766 1 7397
2 90767 1 7398
2 90768 1 7398
2 90769 1 7398
2 90770 1 7398
2 90771 1 7398
2 90772 1 7398
2 90773 1 7398
2 90774 1 7398
2 90775 1 7398
2 90776 1 7402
2 90777 1 7402
2 90778 1 7402
2 90779 1 7409
2 90780 1 7409
2 90781 1 7420
2 90782 1 7420
2 90783 1 7428
2 90784 1 7428
2 90785 1 7428
2 90786 1 7428
2 90787 1 7428
2 90788 1 7428
2 90789 1 7428
2 90790 1 7428
2 90791 1 7428
2 90792 1 7428
2 90793 1 7429
2 90794 1 7429
2 90795 1 7436
2 90796 1 7436
2 90797 1 7437
2 90798 1 7437
2 90799 1 7437
2 90800 1 7438
2 90801 1 7438
2 90802 1 7453
2 90803 1 7453
2 90804 1 7457
2 90805 1 7457
2 90806 1 7457
2 90807 1 7457
2 90808 1 7457
2 90809 1 7457
2 90810 1 7457
2 90811 1 7457
2 90812 1 7457
2 90813 1 7457
2 90814 1 7457
2 90815 1 7457
2 90816 1 7457
2 90817 1 7457
2 90818 1 7457
2 90819 1 7457
2 90820 1 7457
2 90821 1 7457
2 90822 1 7458
2 90823 1 7458
2 90824 1 7458
2 90825 1 7458
2 90826 1 7458
2 90827 1 7458
2 90828 1 7458
2 90829 1 7473
2 90830 1 7473
2 90831 1 7473
2 90832 1 7473
2 90833 1 7474
2 90834 1 7474
2 90835 1 7475
2 90836 1 7475
2 90837 1 7475
2 90838 1 7476
2 90839 1 7476
2 90840 1 7483
2 90841 1 7483
2 90842 1 7483
2 90843 1 7495
2 90844 1 7495
2 90845 1 7495
2 90846 1 7495
2 90847 1 7497
2 90848 1 7497
2 90849 1 7497
2 90850 1 7497
2 90851 1 7497
2 90852 1 7517
2 90853 1 7517
2 90854 1 7518
2 90855 1 7518
2 90856 1 7519
2 90857 1 7519
2 90858 1 7523
2 90859 1 7523
2 90860 1 7523
2 90861 1 7523
2 90862 1 7523
2 90863 1 7523
2 90864 1 7523
2 90865 1 7523
2 90866 1 7523
2 90867 1 7523
2 90868 1 7523
2 90869 1 7523
2 90870 1 7526
2 90871 1 7526
2 90872 1 7536
2 90873 1 7536
2 90874 1 7536
2 90875 1 7536
2 90876 1 7536
2 90877 1 7536
2 90878 1 7537
2 90879 1 7537
2 90880 1 7537
2 90881 1 7537
2 90882 1 7537
2 90883 1 7538
2 90884 1 7538
2 90885 1 7543
2 90886 1 7543
2 90887 1 7543
2 90888 1 7544
2 90889 1 7544
2 90890 1 7544
2 90891 1 7544
2 90892 1 7544
2 90893 1 7544
2 90894 1 7544
2 90895 1 7544
2 90896 1 7544
2 90897 1 7544
2 90898 1 7544
2 90899 1 7544
2 90900 1 7546
2 90901 1 7546
2 90902 1 7561
2 90903 1 7561
2 90904 1 7561
2 90905 1 7561
2 90906 1 7561
2 90907 1 7561
2 90908 1 7561
2 90909 1 7561
2 90910 1 7561
2 90911 1 7561
2 90912 1 7561
2 90913 1 7561
2 90914 1 7561
2 90915 1 7562
2 90916 1 7562
2 90917 1 7563
2 90918 1 7563
2 90919 1 7563
2 90920 1 7564
2 90921 1 7564
2 90922 1 7564
2 90923 1 7564
2 90924 1 7564
2 90925 1 7564
2 90926 1 7564
2 90927 1 7567
2 90928 1 7567
2 90929 1 7570
2 90930 1 7570
2 90931 1 7570
2 90932 1 7570
2 90933 1 7570
2 90934 1 7570
2 90935 1 7570
2 90936 1 7571
2 90937 1 7571
2 90938 1 7571
2 90939 1 7571
2 90940 1 7571
2 90941 1 7572
2 90942 1 7572
2 90943 1 7572
2 90944 1 7573
2 90945 1 7573
2 90946 1 7595
2 90947 1 7595
2 90948 1 7597
2 90949 1 7597
2 90950 1 7597
2 90951 1 7597
2 90952 1 7597
2 90953 1 7597
2 90954 1 7598
2 90955 1 7598
2 90956 1 7598
2 90957 1 7598
2 90958 1 7605
2 90959 1 7605
2 90960 1 7605
2 90961 1 7606
2 90962 1 7606
2 90963 1 7606
2 90964 1 7606
2 90965 1 7606
2 90966 1 7606
2 90967 1 7607
2 90968 1 7607
2 90969 1 7630
2 90970 1 7630
2 90971 1 7654
2 90972 1 7654
2 90973 1 7669
2 90974 1 7669
2 90975 1 7669
2 90976 1 7671
2 90977 1 7671
2 90978 1 7672
2 90979 1 7672
2 90980 1 7672
2 90981 1 7672
2 90982 1 7672
2 90983 1 7672
2 90984 1 7679
2 90985 1 7679
2 90986 1 7691
2 90987 1 7691
2 90988 1 7691
2 90989 1 7691
2 90990 1 7691
2 90991 1 7691
2 90992 1 7691
2 90993 1 7711
2 90994 1 7711
2 90995 1 7711
2 90996 1 7711
2 90997 1 7711
2 90998 1 7711
2 90999 1 7711
2 91000 1 7711
2 91001 1 7711
2 91002 1 7711
2 91003 1 7711
2 91004 1 7711
2 91005 1 7711
2 91006 1 7711
2 91007 1 7711
2 91008 1 7711
2 91009 1 7711
2 91010 1 7711
2 91011 1 7711
2 91012 1 7711
2 91013 1 7711
2 91014 1 7711
2 91015 1 7711
2 91016 1 7711
2 91017 1 7711
2 91018 1 7711
2 91019 1 7711
2 91020 1 7711
2 91021 1 7711
2 91022 1 7711
2 91023 1 7711
2 91024 1 7711
2 91025 1 7711
2 91026 1 7712
2 91027 1 7712
2 91028 1 7712
2 91029 1 7712
2 91030 1 7712
2 91031 1 7712
2 91032 1 7713
2 91033 1 7713
2 91034 1 7713
2 91035 1 7713
2 91036 1 7713
2 91037 1 7713
2 91038 1 7713
2 91039 1 7713
2 91040 1 7713
2 91041 1 7713
2 91042 1 7714
2 91043 1 7714
2 91044 1 7720
2 91045 1 7720
2 91046 1 7720
2 91047 1 7720
2 91048 1 7720
2 91049 1 7734
2 91050 1 7734
2 91051 1 7734
2 91052 1 7734
2 91053 1 7734
2 91054 1 7744
2 91055 1 7744
2 91056 1 7753
2 91057 1 7753
2 91058 1 7755
2 91059 1 7755
2 91060 1 7755
2 91061 1 7755
2 91062 1 7763
2 91063 1 7763
2 91064 1 7763
2 91065 1 7763
2 91066 1 7763
2 91067 1 7763
2 91068 1 7763
2 91069 1 7763
2 91070 1 7763
2 91071 1 7763
2 91072 1 7763
2 91073 1 7763
2 91074 1 7763
2 91075 1 7763
2 91076 1 7763
2 91077 1 7763
2 91078 1 7764
2 91079 1 7764
2 91080 1 7767
2 91081 1 7767
2 91082 1 7767
2 91083 1 7768
2 91084 1 7768
2 91085 1 7768
2 91086 1 7779
2 91087 1 7779
2 91088 1 7779
2 91089 1 7781
2 91090 1 7781
2 91091 1 7790
2 91092 1 7790
2 91093 1 7790
2 91094 1 7792
2 91095 1 7792
2 91096 1 7796
2 91097 1 7796
2 91098 1 7810
2 91099 1 7810
2 91100 1 7810
2 91101 1 7813
2 91102 1 7813
2 91103 1 7813
2 91104 1 7813
2 91105 1 7813
2 91106 1 7813
2 91107 1 7813
2 91108 1 7813
2 91109 1 7813
2 91110 1 7813
2 91111 1 7823
2 91112 1 7823
2 91113 1 7832
2 91114 1 7832
2 91115 1 7833
2 91116 1 7833
2 91117 1 7833
2 91118 1 7834
2 91119 1 7834
2 91120 1 7835
2 91121 1 7835
2 91122 1 7851
2 91123 1 7851
2 91124 1 7851
2 91125 1 7851
2 91126 1 7851
2 91127 1 7851
2 91128 1 7851
2 91129 1 7851
2 91130 1 7851
2 91131 1 7851
2 91132 1 7851
2 91133 1 7851
2 91134 1 7851
2 91135 1 7851
2 91136 1 7851
2 91137 1 7851
2 91138 1 7851
2 91139 1 7851
2 91140 1 7851
2 91141 1 7851
2 91142 1 7852
2 91143 1 7852
2 91144 1 7852
2 91145 1 7860
2 91146 1 7860
2 91147 1 7860
2 91148 1 7860
2 91149 1 7860
2 91150 1 7860
2 91151 1 7860
2 91152 1 7860
2 91153 1 7860
2 91154 1 7860
2 91155 1 7860
2 91156 1 7860
2 91157 1 7887
2 91158 1 7887
2 91159 1 7887
2 91160 1 7887
2 91161 1 7887
2 91162 1 7887
2 91163 1 7887
2 91164 1 7887
2 91165 1 7887
2 91166 1 7887
2 91167 1 7887
2 91168 1 7887
2 91169 1 7887
2 91170 1 7887
2 91171 1 7887
2 91172 1 7887
2 91173 1 7887
2 91174 1 7887
2 91175 1 7887
2 91176 1 7887
2 91177 1 7887
2 91178 1 7887
2 91179 1 7887
2 91180 1 7887
2 91181 1 7888
2 91182 1 7888
2 91183 1 7888
2 91184 1 7889
2 91185 1 7889
2 91186 1 7889
2 91187 1 7890
2 91188 1 7890
2 91189 1 7890
2 91190 1 7890
2 91191 1 7892
2 91192 1 7892
2 91193 1 7894
2 91194 1 7894
2 91195 1 7894
2 91196 1 7894
2 91197 1 7894
2 91198 1 7894
2 91199 1 7894
2 91200 1 7894
2 91201 1 7895
2 91202 1 7895
2 91203 1 7905
2 91204 1 7905
2 91205 1 7905
2 91206 1 7905
2 91207 1 7906
2 91208 1 7906
2 91209 1 7906
2 91210 1 7906
2 91211 1 7906
2 91212 1 7907
2 91213 1 7907
2 91214 1 7908
2 91215 1 7908
2 91216 1 7908
2 91217 1 7908
2 91218 1 7908
2 91219 1 7908
2 91220 1 7908
2 91221 1 7908
2 91222 1 7908
2 91223 1 7910
2 91224 1 7910
2 91225 1 7913
2 91226 1 7913
2 91227 1 7913
2 91228 1 7916
2 91229 1 7916
2 91230 1 7916
2 91231 1 7918
2 91232 1 7918
2 91233 1 7918
2 91234 1 7918
2 91235 1 7934
2 91236 1 7934
2 91237 1 7934
2 91238 1 7934
2 91239 1 7934
2 91240 1 7934
2 91241 1 7934
2 91242 1 7934
2 91243 1 7934
2 91244 1 7934
2 91245 1 7934
2 91246 1 7934
2 91247 1 7934
2 91248 1 7935
2 91249 1 7935
2 91250 1 7936
2 91251 1 7936
2 91252 1 7936
2 91253 1 7936
2 91254 1 7936
2 91255 1 7936
2 91256 1 7936
2 91257 1 7936
2 91258 1 7937
2 91259 1 7937
2 91260 1 7937
2 91261 1 7937
2 91262 1 7937
2 91263 1 7941
2 91264 1 7941
2 91265 1 7941
2 91266 1 7941
2 91267 1 7941
2 91268 1 7942
2 91269 1 7942
2 91270 1 7942
2 91271 1 7942
2 91272 1 7942
2 91273 1 7942
2 91274 1 7942
2 91275 1 7944
2 91276 1 7944
2 91277 1 7945
2 91278 1 7945
2 91279 1 7946
2 91280 1 7946
2 91281 1 7946
2 91282 1 7946
2 91283 1 7946
2 91284 1 7946
2 91285 1 7946
2 91286 1 7946
2 91287 1 7946
2 91288 1 7946
2 91289 1 7955
2 91290 1 7955
2 91291 1 7955
2 91292 1 7969
2 91293 1 7969
2 91294 1 7969
2 91295 1 7969
2 91296 1 7972
2 91297 1 7972
2 91298 1 7978
2 91299 1 7978
2 91300 1 7978
2 91301 1 7989
2 91302 1 7989
2 91303 1 7993
2 91304 1 7993
2 91305 1 7993
2 91306 1 7994
2 91307 1 7994
2 91308 1 7994
2 91309 1 7994
2 91310 1 7994
2 91311 1 7994
2 91312 1 7996
2 91313 1 7996
2 91314 1 7996
2 91315 1 7996
2 91316 1 7996
2 91317 1 8000
2 91318 1 8000
2 91319 1 8000
2 91320 1 8002
2 91321 1 8002
2 91322 1 8002
2 91323 1 8012
2 91324 1 8012
2 91325 1 8012
2 91326 1 8012
2 91327 1 8012
2 91328 1 8013
2 91329 1 8013
2 91330 1 8034
2 91331 1 8034
2 91332 1 8034
2 91333 1 8034
2 91334 1 8034
2 91335 1 8035
2 91336 1 8035
2 91337 1 8036
2 91338 1 8036
2 91339 1 8037
2 91340 1 8037
2 91341 1 8037
2 91342 1 8037
2 91343 1 8037
2 91344 1 8037
2 91345 1 8041
2 91346 1 8041
2 91347 1 8041
2 91348 1 8041
2 91349 1 8041
2 91350 1 8041
2 91351 1 8041
2 91352 1 8041
2 91353 1 8041
2 91354 1 8042
2 91355 1 8042
2 91356 1 8042
2 91357 1 8042
2 91358 1 8043
2 91359 1 8043
2 91360 1 8044
2 91361 1 8044
2 91362 1 8044
2 91363 1 8044
2 91364 1 8044
2 91365 1 8044
2 91366 1 8046
2 91367 1 8046
2 91368 1 8046
2 91369 1 8046
2 91370 1 8046
2 91371 1 8046
2 91372 1 8046
2 91373 1 8046
2 91374 1 8046
2 91375 1 8046
2 91376 1 8046
2 91377 1 8046
2 91378 1 8046
2 91379 1 8046
2 91380 1 8046
2 91381 1 8046
2 91382 1 8050
2 91383 1 8050
2 91384 1 8050
2 91385 1 8053
2 91386 1 8053
2 91387 1 8053
2 91388 1 8053
2 91389 1 8053
2 91390 1 8053
2 91391 1 8055
2 91392 1 8055
2 91393 1 8055
2 91394 1 8056
2 91395 1 8056
2 91396 1 8064
2 91397 1 8064
2 91398 1 8064
2 91399 1 8064
2 91400 1 8075
2 91401 1 8075
2 91402 1 8079
2 91403 1 8079
2 91404 1 8079
2 91405 1 8079
2 91406 1 8079
2 91407 1 8080
2 91408 1 8080
2 91409 1 8080
2 91410 1 8080
2 91411 1 8081
2 91412 1 8081
2 91413 1 8081
2 91414 1 8081
2 91415 1 8081
2 91416 1 8081
2 91417 1 8091
2 91418 1 8091
2 91419 1 8091
2 91420 1 8092
2 91421 1 8092
2 91422 1 8092
2 91423 1 8092
2 91424 1 8093
2 91425 1 8093
2 91426 1 8093
2 91427 1 8093
2 91428 1 8102
2 91429 1 8102
2 91430 1 8102
2 91431 1 8102
2 91432 1 8102
2 91433 1 8102
2 91434 1 8102
2 91435 1 8102
2 91436 1 8102
2 91437 1 8102
2 91438 1 8105
2 91439 1 8105
2 91440 1 8108
2 91441 1 8108
2 91442 1 8108
2 91443 1 8108
2 91444 1 8108
2 91445 1 8108
2 91446 1 8108
2 91447 1 8108
2 91448 1 8108
2 91449 1 8108
2 91450 1 8108
2 91451 1 8108
2 91452 1 8108
2 91453 1 8108
2 91454 1 8108
2 91455 1 8110
2 91456 1 8110
2 91457 1 8110
2 91458 1 8110
2 91459 1 8118
2 91460 1 8118
2 91461 1 8118
2 91462 1 8118
2 91463 1 8124
2 91464 1 8124
2 91465 1 8125
2 91466 1 8125
2 91467 1 8125
2 91468 1 8125
2 91469 1 8125
2 91470 1 8125
2 91471 1 8152
2 91472 1 8152
2 91473 1 8152
2 91474 1 8152
2 91475 1 8152
2 91476 1 8152
2 91477 1 8155
2 91478 1 8155
2 91479 1 8155
2 91480 1 8157
2 91481 1 8157
2 91482 1 8157
2 91483 1 8157
2 91484 1 8157
2 91485 1 8157
2 91486 1 8157
2 91487 1 8157
2 91488 1 8157
2 91489 1 8157
2 91490 1 8157
2 91491 1 8158
2 91492 1 8158
2 91493 1 8168
2 91494 1 8168
2 91495 1 8177
2 91496 1 8177
2 91497 1 8177
2 91498 1 8177
2 91499 1 8177
2 91500 1 8177
2 91501 1 8177
2 91502 1 8177
2 91503 1 8177
2 91504 1 8177
2 91505 1 8177
2 91506 1 8177
2 91507 1 8178
2 91508 1 8178
2 91509 1 8178
2 91510 1 8190
2 91511 1 8190
2 91512 1 8190
2 91513 1 8191
2 91514 1 8191
2 91515 1 8191
2 91516 1 8191
2 91517 1 8192
2 91518 1 8192
2 91519 1 8192
2 91520 1 8192
2 91521 1 8193
2 91522 1 8193
2 91523 1 8194
2 91524 1 8194
2 91525 1 8199
2 91526 1 8199
2 91527 1 8200
2 91528 1 8200
2 91529 1 8225
2 91530 1 8225
2 91531 1 8225
2 91532 1 8225
2 91533 1 8225
2 91534 1 8225
2 91535 1 8225
2 91536 1 8225
2 91537 1 8225
2 91538 1 8225
2 91539 1 8225
2 91540 1 8225
2 91541 1 8225
2 91542 1 8225
2 91543 1 8225
2 91544 1 8225
2 91545 1 8225
2 91546 1 8226
2 91547 1 8226
2 91548 1 8227
2 91549 1 8227
2 91550 1 8227
2 91551 1 8230
2 91552 1 8230
2 91553 1 8230
2 91554 1 8230
2 91555 1 8230
2 91556 1 8230
2 91557 1 8230
2 91558 1 8230
2 91559 1 8230
2 91560 1 8230
2 91561 1 8230
2 91562 1 8230
2 91563 1 8230
2 91564 1 8230
2 91565 1 8231
2 91566 1 8231
2 91567 1 8231
2 91568 1 8231
2 91569 1 8231
2 91570 1 8231
2 91571 1 8231
2 91572 1 8231
2 91573 1 8231
2 91574 1 8231
2 91575 1 8231
2 91576 1 8241
2 91577 1 8241
2 91578 1 8242
2 91579 1 8242
2 91580 1 8242
2 91581 1 8242
2 91582 1 8250
2 91583 1 8250
2 91584 1 8253
2 91585 1 8253
2 91586 1 8254
2 91587 1 8254
2 91588 1 8254
2 91589 1 8254
2 91590 1 8254
2 91591 1 8257
2 91592 1 8257
2 91593 1 8264
2 91594 1 8264
2 91595 1 8264
2 91596 1 8264
2 91597 1 8265
2 91598 1 8265
2 91599 1 8265
2 91600 1 8265
2 91601 1 8265
2 91602 1 8265
2 91603 1 8265
2 91604 1 8267
2 91605 1 8267
2 91606 1 8267
2 91607 1 8268
2 91608 1 8268
2 91609 1 8268
2 91610 1 8268
2 91611 1 8268
2 91612 1 8268
2 91613 1 8281
2 91614 1 8281
2 91615 1 8283
2 91616 1 8283
2 91617 1 8283
2 91618 1 8286
2 91619 1 8286
2 91620 1 8286
2 91621 1 8287
2 91622 1 8287
2 91623 1 8287
2 91624 1 8287
2 91625 1 8297
2 91626 1 8297
2 91627 1 8297
2 91628 1 8297
2 91629 1 8299
2 91630 1 8299
2 91631 1 8307
2 91632 1 8307
2 91633 1 8307
2 91634 1 8307
2 91635 1 8307
2 91636 1 8307
2 91637 1 8308
2 91638 1 8308
2 91639 1 8308
2 91640 1 8308
2 91641 1 8308
2 91642 1 8309
2 91643 1 8309
2 91644 1 8309
2 91645 1 8309
2 91646 1 8309
2 91647 1 8309
2 91648 1 8310
2 91649 1 8310
2 91650 1 8310
2 91651 1 8310
2 91652 1 8310
2 91653 1 8311
2 91654 1 8311
2 91655 1 8311
2 91656 1 8320
2 91657 1 8320
2 91658 1 8322
2 91659 1 8322
2 91660 1 8322
2 91661 1 8322
2 91662 1 8323
2 91663 1 8323
2 91664 1 8323
2 91665 1 8344
2 91666 1 8344
2 91667 1 8344
2 91668 1 8344
2 91669 1 8344
2 91670 1 8344
2 91671 1 8345
2 91672 1 8345
2 91673 1 8346
2 91674 1 8346
2 91675 1 8346
2 91676 1 8346
2 91677 1 8346
2 91678 1 8346
2 91679 1 8347
2 91680 1 8347
2 91681 1 8347
2 91682 1 8348
2 91683 1 8348
2 91684 1 8351
2 91685 1 8351
2 91686 1 8351
2 91687 1 8351
2 91688 1 8358
2 91689 1 8358
2 91690 1 8358
2 91691 1 8358
2 91692 1 8358
2 91693 1 8358
2 91694 1 8358
2 91695 1 8358
2 91696 1 8358
2 91697 1 8358
2 91698 1 8358
2 91699 1 8358
2 91700 1 8358
2 91701 1 8360
2 91702 1 8360
2 91703 1 8360
2 91704 1 8360
2 91705 1 8360
2 91706 1 8360
2 91707 1 8360
2 91708 1 8360
2 91709 1 8361
2 91710 1 8361
2 91711 1 8361
2 91712 1 8361
2 91713 1 8361
2 91714 1 8361
2 91715 1 8370
2 91716 1 8370
2 91717 1 8370
2 91718 1 8370
2 91719 1 8371
2 91720 1 8371
2 91721 1 8371
2 91722 1 8371
2 91723 1 8372
2 91724 1 8372
2 91725 1 8373
2 91726 1 8373
2 91727 1 8389
2 91728 1 8389
2 91729 1 8389
2 91730 1 8393
2 91731 1 8393
2 91732 1 8421
2 91733 1 8421
2 91734 1 8421
2 91735 1 8421
2 91736 1 8422
2 91737 1 8422
2 91738 1 8422
2 91739 1 8422
2 91740 1 8422
2 91741 1 8429
2 91742 1 8429
2 91743 1 8429
2 91744 1 8429
2 91745 1 8429
2 91746 1 8429
2 91747 1 8430
2 91748 1 8430
2 91749 1 8430
2 91750 1 8430
2 91751 1 8431
2 91752 1 8431
2 91753 1 8432
2 91754 1 8432
2 91755 1 8432
2 91756 1 8434
2 91757 1 8434
2 91758 1 8442
2 91759 1 8442
2 91760 1 8442
2 91761 1 8442
2 91762 1 8447
2 91763 1 8447
2 91764 1 8448
2 91765 1 8448
2 91766 1 8448
2 91767 1 8448
2 91768 1 8448
2 91769 1 8449
2 91770 1 8449
2 91771 1 8449
2 91772 1 8460
2 91773 1 8460
2 91774 1 8460
2 91775 1 8460
2 91776 1 8460
2 91777 1 8460
2 91778 1 8460
2 91779 1 8461
2 91780 1 8461
2 91781 1 8468
2 91782 1 8468
2 91783 1 8468
2 91784 1 8469
2 91785 1 8469
2 91786 1 8469
2 91787 1 8469
2 91788 1 8472
2 91789 1 8472
2 91790 1 8472
2 91791 1 8473
2 91792 1 8473
2 91793 1 8473
2 91794 1 8473
2 91795 1 8494
2 91796 1 8494
2 91797 1 8509
2 91798 1 8509
2 91799 1 8510
2 91800 1 8510
2 91801 1 8510
2 91802 1 8526
2 91803 1 8526
2 91804 1 8526
2 91805 1 8526
2 91806 1 8527
2 91807 1 8527
2 91808 1 8527
2 91809 1 8534
2 91810 1 8534
2 91811 1 8543
2 91812 1 8543
2 91813 1 8543
2 91814 1 8544
2 91815 1 8544
2 91816 1 8545
2 91817 1 8545
2 91818 1 8546
2 91819 1 8546
2 91820 1 8546
2 91821 1 8546
2 91822 1 8547
2 91823 1 8547
2 91824 1 8547
2 91825 1 8547
2 91826 1 8547
2 91827 1 8567
2 91828 1 8567
2 91829 1 8567
2 91830 1 8567
2 91831 1 8567
2 91832 1 8567
2 91833 1 8567
2 91834 1 8568
2 91835 1 8568
2 91836 1 8568
2 91837 1 8569
2 91838 1 8569
2 91839 1 8579
2 91840 1 8579
2 91841 1 8579
2 91842 1 8579
2 91843 1 8579
2 91844 1 8580
2 91845 1 8580
2 91846 1 8580
2 91847 1 8580
2 91848 1 8593
2 91849 1 8593
2 91850 1 8593
2 91851 1 8593
2 91852 1 8593
2 91853 1 8593
2 91854 1 8594
2 91855 1 8594
2 91856 1 8594
2 91857 1 8596
2 91858 1 8596
2 91859 1 8598
2 91860 1 8598
2 91861 1 8616
2 91862 1 8616
2 91863 1 8639
2 91864 1 8639
2 91865 1 8639
2 91866 1 8639
2 91867 1 8639
2 91868 1 8640
2 91869 1 8640
2 91870 1 8640
2 91871 1 8640
2 91872 1 8640
2 91873 1 8640
2 91874 1 8664
2 91875 1 8664
2 91876 1 8664
2 91877 1 8664
2 91878 1 8664
2 91879 1 8664
2 91880 1 8664
2 91881 1 8664
2 91882 1 8664
2 91883 1 8664
2 91884 1 8664
2 91885 1 8664
2 91886 1 8665
2 91887 1 8665
2 91888 1 8665
2 91889 1 8666
2 91890 1 8666
2 91891 1 8679
2 91892 1 8679
2 91893 1 8679
2 91894 1 8679
2 91895 1 8679
2 91896 1 8679
2 91897 1 8679
2 91898 1 8679
2 91899 1 8679
2 91900 1 8679
2 91901 1 8680
2 91902 1 8680
2 91903 1 8681
2 91904 1 8681
2 91905 1 8681
2 91906 1 8681
2 91907 1 8681
2 91908 1 8681
2 91909 1 8681
2 91910 1 8681
2 91911 1 8681
2 91912 1 8681
2 91913 1 8689
2 91914 1 8689
2 91915 1 8689
2 91916 1 8690
2 91917 1 8690
2 91918 1 8702
2 91919 1 8702
2 91920 1 8717
2 91921 1 8717
2 91922 1 8717
2 91923 1 8735
2 91924 1 8735
2 91925 1 8738
2 91926 1 8738
2 91927 1 8738
2 91928 1 8744
2 91929 1 8744
2 91930 1 8744
2 91931 1 8744
2 91932 1 8752
2 91933 1 8752
2 91934 1 8752
2 91935 1 8752
2 91936 1 8753
2 91937 1 8753
2 91938 1 8753
2 91939 1 8754
2 91940 1 8754
2 91941 1 8756
2 91942 1 8756
2 91943 1 8757
2 91944 1 8757
2 91945 1 8766
2 91946 1 8766
2 91947 1 8766
2 91948 1 8766
2 91949 1 8766
2 91950 1 8766
2 91951 1 8766
2 91952 1 8768
2 91953 1 8768
2 91954 1 8768
2 91955 1 8768
2 91956 1 8786
2 91957 1 8786
2 91958 1 8801
2 91959 1 8801
2 91960 1 8801
2 91961 1 8802
2 91962 1 8802
2 91963 1 8802
2 91964 1 8803
2 91965 1 8803
2 91966 1 8803
2 91967 1 8804
2 91968 1 8804
2 91969 1 8805
2 91970 1 8805
2 91971 1 8805
2 91972 1 8813
2 91973 1 8813
2 91974 1 8820
2 91975 1 8820
2 91976 1 8820
2 91977 1 8821
2 91978 1 8821
2 91979 1 8822
2 91980 1 8822
2 91981 1 8836
2 91982 1 8836
2 91983 1 8836
2 91984 1 8836
2 91985 1 8836
2 91986 1 8837
2 91987 1 8837
2 91988 1 8841
2 91989 1 8841
2 91990 1 8841
2 91991 1 8841
2 91992 1 8844
2 91993 1 8844
2 91994 1 8846
2 91995 1 8846
2 91996 1 8849
2 91997 1 8849
2 91998 1 8849
2 91999 1 8849
2 92000 1 8849
2 92001 1 8849
2 92002 1 8849
2 92003 1 8849
2 92004 1 8849
2 92005 1 8849
2 92006 1 8850
2 92007 1 8850
2 92008 1 8851
2 92009 1 8851
2 92010 1 8851
2 92011 1 8851
2 92012 1 8860
2 92013 1 8860
2 92014 1 8869
2 92015 1 8869
2 92016 1 8880
2 92017 1 8880
2 92018 1 8881
2 92019 1 8881
2 92020 1 8892
2 92021 1 8892
2 92022 1 8892
2 92023 1 8894
2 92024 1 8894
2 92025 1 8917
2 92026 1 8917
2 92027 1 8917
2 92028 1 8918
2 92029 1 8918
2 92030 1 8918
2 92031 1 8918
2 92032 1 8918
2 92033 1 8925
2 92034 1 8925
2 92035 1 8925
2 92036 1 8925
2 92037 1 8926
2 92038 1 8926
2 92039 1 8926
2 92040 1 8929
2 92041 1 8929
2 92042 1 8930
2 92043 1 8930
2 92044 1 8937
2 92045 1 8937
2 92046 1 8945
2 92047 1 8945
2 92048 1 8945
2 92049 1 8949
2 92050 1 8949
2 92051 1 8956
2 92052 1 8956
2 92053 1 8956
2 92054 1 8960
2 92055 1 8960
2 92056 1 8961
2 92057 1 8961
2 92058 1 8961
2 92059 1 8961
2 92060 1 8961
2 92061 1 8961
2 92062 1 8961
2 92063 1 8961
2 92064 1 8961
2 92065 1 8961
2 92066 1 8961
2 92067 1 8961
2 92068 1 8961
2 92069 1 8971
2 92070 1 8971
2 92071 1 8971
2 92072 1 8972
2 92073 1 8972
2 92074 1 8972
2 92075 1 8972
2 92076 1 8972
2 92077 1 8972
2 92078 1 8972
2 92079 1 8982
2 92080 1 8982
2 92081 1 8982
2 92082 1 8983
2 92083 1 8983
2 92084 1 8993
2 92085 1 8993
2 92086 1 8993
2 92087 1 8994
2 92088 1 8994
2 92089 1 8994
2 92090 1 8994
2 92091 1 8997
2 92092 1 8997
2 92093 1 9002
2 92094 1 9002
2 92095 1 9022
2 92096 1 9022
2 92097 1 9037
2 92098 1 9037
2 92099 1 9045
2 92100 1 9045
2 92101 1 9068
2 92102 1 9068
2 92103 1 9070
2 92104 1 9070
2 92105 1 9076
2 92106 1 9076
2 92107 1 9088
2 92108 1 9088
2 92109 1 9088
2 92110 1 9088
2 92111 1 9088
2 92112 1 9088
2 92113 1 9088
2 92114 1 9112
2 92115 1 9112
2 92116 1 9123
2 92117 1 9123
2 92118 1 9123
2 92119 1 9123
2 92120 1 9123
2 92121 1 9123
2 92122 1 9123
2 92123 1 9123
2 92124 1 9123
2 92125 1 9123
2 92126 1 9123
2 92127 1 9123
2 92128 1 9123
2 92129 1 9123
2 92130 1 9123
2 92131 1 9123
2 92132 1 9123
2 92133 1 9123
2 92134 1 9123
2 92135 1 9123
2 92136 1 9123
2 92137 1 9123
2 92138 1 9123
2 92139 1 9123
2 92140 1 9123
2 92141 1 9123
2 92142 1 9123
2 92143 1 9123
2 92144 1 9123
2 92145 1 9124
2 92146 1 9124
2 92147 1 9124
2 92148 1 9124
2 92149 1 9124
2 92150 1 9124
2 92151 1 9125
2 92152 1 9125
2 92153 1 9125
2 92154 1 9127
2 92155 1 9127
2 92156 1 9127
2 92157 1 9150
2 92158 1 9150
2 92159 1 9150
2 92160 1 9150
2 92161 1 9150
2 92162 1 9157
2 92163 1 9157
2 92164 1 9157
2 92165 1 9157
2 92166 1 9157
2 92167 1 9158
2 92168 1 9158
2 92169 1 9158
2 92170 1 9158
2 92171 1 9158
2 92172 1 9159
2 92173 1 9159
2 92174 1 9159
2 92175 1 9160
2 92176 1 9160
2 92177 1 9162
2 92178 1 9162
2 92179 1 9163
2 92180 1 9163
2 92181 1 9163
2 92182 1 9163
2 92183 1 9170
2 92184 1 9170
2 92185 1 9171
2 92186 1 9171
2 92187 1 9181
2 92188 1 9181
2 92189 1 9181
2 92190 1 9181
2 92191 1 9181
2 92192 1 9181
2 92193 1 9181
2 92194 1 9181
2 92195 1 9182
2 92196 1 9182
2 92197 1 9182
2 92198 1 9184
2 92199 1 9184
2 92200 1 9184
2 92201 1 9184
2 92202 1 9185
2 92203 1 9185
2 92204 1 9185
2 92205 1 9185
2 92206 1 9197
2 92207 1 9197
2 92208 1 9201
2 92209 1 9201
2 92210 1 9201
2 92211 1 9212
2 92212 1 9212
2 92213 1 9212
2 92214 1 9232
2 92215 1 9232
2 92216 1 9232
2 92217 1 9243
2 92218 1 9243
2 92219 1 9251
2 92220 1 9251
2 92221 1 9251
2 92222 1 9251
2 92223 1 9251
2 92224 1 9251
2 92225 1 9251
2 92226 1 9257
2 92227 1 9257
2 92228 1 9257
2 92229 1 9257
2 92230 1 9257
2 92231 1 9257
2 92232 1 9257
2 92233 1 9258
2 92234 1 9258
2 92235 1 9258
2 92236 1 9258
2 92237 1 9258
2 92238 1 9258
2 92239 1 9258
2 92240 1 9258
2 92241 1 9258
2 92242 1 9260
2 92243 1 9260
2 92244 1 9260
2 92245 1 9260
2 92246 1 9273
2 92247 1 9273
2 92248 1 9273
2 92249 1 9283
2 92250 1 9283
2 92251 1 9283
2 92252 1 9284
2 92253 1 9284
2 92254 1 9284
2 92255 1 9284
2 92256 1 9284
2 92257 1 9284
2 92258 1 9284
2 92259 1 9284
2 92260 1 9284
2 92261 1 9287
2 92262 1 9287
2 92263 1 9300
2 92264 1 9300
2 92265 1 9300
2 92266 1 9300
2 92267 1 9300
2 92268 1 9300
2 92269 1 9307
2 92270 1 9307
2 92271 1 9309
2 92272 1 9309
2 92273 1 9319
2 92274 1 9319
2 92275 1 9319
2 92276 1 9319
2 92277 1 9319
2 92278 1 9319
2 92279 1 9319
2 92280 1 9319
2 92281 1 9319
2 92282 1 9320
2 92283 1 9320
2 92284 1 9321
2 92285 1 9321
2 92286 1 9321
2 92287 1 9321
2 92288 1 9331
2 92289 1 9331
2 92290 1 9332
2 92291 1 9332
2 92292 1 9332
2 92293 1 9334
2 92294 1 9334
2 92295 1 9335
2 92296 1 9335
2 92297 1 9336
2 92298 1 9336
2 92299 1 9336
2 92300 1 9339
2 92301 1 9339
2 92302 1 9339
2 92303 1 9339
2 92304 1 9339
2 92305 1 9339
2 92306 1 9339
2 92307 1 9339
2 92308 1 9339
2 92309 1 9339
2 92310 1 9339
2 92311 1 9340
2 92312 1 9340
2 92313 1 9340
2 92314 1 9340
2 92315 1 9340
2 92316 1 9340
2 92317 1 9340
2 92318 1 9342
2 92319 1 9342
2 92320 1 9350
2 92321 1 9350
2 92322 1 9351
2 92323 1 9351
2 92324 1 9354
2 92325 1 9354
2 92326 1 9356
2 92327 1 9356
2 92328 1 9364
2 92329 1 9364
2 92330 1 9365
2 92331 1 9365
2 92332 1 9367
2 92333 1 9367
2 92334 1 9367
2 92335 1 9370
2 92336 1 9370
2 92337 1 9370
2 92338 1 9370
2 92339 1 9370
2 92340 1 9370
2 92341 1 9370
2 92342 1 9370
2 92343 1 9370
2 92344 1 9382
2 92345 1 9382
2 92346 1 9382
2 92347 1 9382
2 92348 1 9382
2 92349 1 9382
2 92350 1 9382
2 92351 1 9382
2 92352 1 9382
2 92353 1 9382
2 92354 1 9382
2 92355 1 9382
2 92356 1 9382
2 92357 1 9382
2 92358 1 9383
2 92359 1 9383
2 92360 1 9383
2 92361 1 9383
2 92362 1 9384
2 92363 1 9384
2 92364 1 9384
2 92365 1 9384
2 92366 1 9384
2 92367 1 9384
2 92368 1 9384
2 92369 1 9395
2 92370 1 9395
2 92371 1 9396
2 92372 1 9396
2 92373 1 9396
2 92374 1 9397
2 92375 1 9397
2 92376 1 9397
2 92377 1 9400
2 92378 1 9400
2 92379 1 9400
2 92380 1 9400
2 92381 1 9400
2 92382 1 9400
2 92383 1 9400
2 92384 1 9400
2 92385 1 9400
2 92386 1 9400
2 92387 1 9418
2 92388 1 9418
2 92389 1 9418
2 92390 1 9420
2 92391 1 9420
2 92392 1 9420
2 92393 1 9421
2 92394 1 9421
2 92395 1 9425
2 92396 1 9425
2 92397 1 9436
2 92398 1 9436
2 92399 1 9437
2 92400 1 9437
2 92401 1 9437
2 92402 1 9437
2 92403 1 9437
2 92404 1 9437
2 92405 1 9437
2 92406 1 9439
2 92407 1 9439
2 92408 1 9439
2 92409 1 9439
2 92410 1 9439
2 92411 1 9439
2 92412 1 9439
2 92413 1 9439
2 92414 1 9439
2 92415 1 9439
2 92416 1 9448
2 92417 1 9448
2 92418 1 9448
2 92419 1 9448
2 92420 1 9448
2 92421 1 9448
2 92422 1 9448
2 92423 1 9448
2 92424 1 9457
2 92425 1 9457
2 92426 1 9458
2 92427 1 9458
2 92428 1 9459
2 92429 1 9459
2 92430 1 9459
2 92431 1 9461
2 92432 1 9461
2 92433 1 9464
2 92434 1 9464
2 92435 1 9464
2 92436 1 9464
2 92437 1 9465
2 92438 1 9465
2 92439 1 9465
2 92440 1 9465
2 92441 1 9465
2 92442 1 9465
2 92443 1 9465
2 92444 1 9465
2 92445 1 9465
2 92446 1 9465
2 92447 1 9479
2 92448 1 9479
2 92449 1 9479
2 92450 1 9479
2 92451 1 9479
2 92452 1 9479
2 92453 1 9479
2 92454 1 9479
2 92455 1 9480
2 92456 1 9480
2 92457 1 9480
2 92458 1 9481
2 92459 1 9481
2 92460 1 9482
2 92461 1 9482
2 92462 1 9483
2 92463 1 9483
2 92464 1 9483
2 92465 1 9483
2 92466 1 9483
2 92467 1 9496
2 92468 1 9496
2 92469 1 9496
2 92470 1 9497
2 92471 1 9497
2 92472 1 9497
2 92473 1 9497
2 92474 1 9498
2 92475 1 9498
2 92476 1 9499
2 92477 1 9499
2 92478 1 9499
2 92479 1 9499
2 92480 1 9499
2 92481 1 9500
2 92482 1 9500
2 92483 1 9501
2 92484 1 9501
2 92485 1 9501
2 92486 1 9509
2 92487 1 9509
2 92488 1 9509
2 92489 1 9517
2 92490 1 9517
2 92491 1 9518
2 92492 1 9518
2 92493 1 9518
2 92494 1 9518
2 92495 1 9518
2 92496 1 9519
2 92497 1 9519
2 92498 1 9527
2 92499 1 9527
2 92500 1 9527
2 92501 1 9527
2 92502 1 9536
2 92503 1 9536
2 92504 1 9537
2 92505 1 9537
2 92506 1 9542
2 92507 1 9542
2 92508 1 9542
2 92509 1 9542
2 92510 1 9542
2 92511 1 9542
2 92512 1 9542
2 92513 1 9543
2 92514 1 9543
2 92515 1 9552
2 92516 1 9552
2 92517 1 9552
2 92518 1 9553
2 92519 1 9553
2 92520 1 9553
2 92521 1 9562
2 92522 1 9562
2 92523 1 9562
2 92524 1 9562
2 92525 1 9562
2 92526 1 9562
2 92527 1 9563
2 92528 1 9563
2 92529 1 9564
2 92530 1 9564
2 92531 1 9564
2 92532 1 9570
2 92533 1 9570
2 92534 1 9572
2 92535 1 9572
2 92536 1 9573
2 92537 1 9573
2 92538 1 9573
2 92539 1 9573
2 92540 1 9573
2 92541 1 9583
2 92542 1 9583
2 92543 1 9593
2 92544 1 9593
2 92545 1 9593
2 92546 1 9593
2 92547 1 9593
2 92548 1 9593
2 92549 1 9593
2 92550 1 9593
2 92551 1 9594
2 92552 1 9594
2 92553 1 9594
2 92554 1 9594
2 92555 1 9600
2 92556 1 9600
2 92557 1 9600
2 92558 1 9600
2 92559 1 9601
2 92560 1 9601
2 92561 1 9601
2 92562 1 9601
2 92563 1 9602
2 92564 1 9602
2 92565 1 9602
2 92566 1 9602
2 92567 1 9603
2 92568 1 9603
2 92569 1 9603
2 92570 1 9603
2 92571 1 9603
2 92572 1 9613
2 92573 1 9613
2 92574 1 9623
2 92575 1 9623
2 92576 1 9623
2 92577 1 9623
2 92578 1 9623
2 92579 1 9623
2 92580 1 9623
2 92581 1 9623
2 92582 1 9623
2 92583 1 9623
2 92584 1 9623
2 92585 1 9624
2 92586 1 9624
2 92587 1 9625
2 92588 1 9625
2 92589 1 9628
2 92590 1 9628
2 92591 1 9629
2 92592 1 9629
2 92593 1 9629
2 92594 1 9630
2 92595 1 9630
2 92596 1 9630
2 92597 1 9639
2 92598 1 9639
2 92599 1 9639
2 92600 1 9639
2 92601 1 9639
2 92602 1 9642
2 92603 1 9642
2 92604 1 9643
2 92605 1 9643
2 92606 1 9644
2 92607 1 9644
2 92608 1 9644
2 92609 1 9644
2 92610 1 9655
2 92611 1 9655
2 92612 1 9655
2 92613 1 9655
2 92614 1 9655
2 92615 1 9655
2 92616 1 9655
2 92617 1 9655
2 92618 1 9655
2 92619 1 9655
2 92620 1 9658
2 92621 1 9658
2 92622 1 9658
2 92623 1 9658
2 92624 1 9658
2 92625 1 9658
2 92626 1 9663
2 92627 1 9663
2 92628 1 9663
2 92629 1 9663
2 92630 1 9663
2 92631 1 9663
2 92632 1 9663
2 92633 1 9663
2 92634 1 9663
2 92635 1 9664
2 92636 1 9664
2 92637 1 9664
2 92638 1 9665
2 92639 1 9665
2 92640 1 9665
2 92641 1 9667
2 92642 1 9667
2 92643 1 9667
2 92644 1 9672
2 92645 1 9672
2 92646 1 9672
2 92647 1 9672
2 92648 1 9672
2 92649 1 9672
2 92650 1 9672
2 92651 1 9683
2 92652 1 9683
2 92653 1 9695
2 92654 1 9695
2 92655 1 9695
2 92656 1 9695
2 92657 1 9708
2 92658 1 9708
2 92659 1 9716
2 92660 1 9716
2 92661 1 9717
2 92662 1 9717
2 92663 1 9718
2 92664 1 9718
2 92665 1 9718
2 92666 1 9718
2 92667 1 9718
2 92668 1 9718
2 92669 1 9718
2 92670 1 9718
2 92671 1 9718
2 92672 1 9718
2 92673 1 9718
2 92674 1 9718
2 92675 1 9718
2 92676 1 9718
2 92677 1 9718
2 92678 1 9718
2 92679 1 9724
2 92680 1 9724
2 92681 1 9731
2 92682 1 9731
2 92683 1 9740
2 92684 1 9740
2 92685 1 9740
2 92686 1 9746
2 92687 1 9746
2 92688 1 9746
2 92689 1 9746
2 92690 1 9746
2 92691 1 9746
2 92692 1 9746
2 92693 1 9746
2 92694 1 9746
2 92695 1 9746
2 92696 1 9757
2 92697 1 9757
2 92698 1 9757
2 92699 1 9757
2 92700 1 9757
2 92701 1 9757
2 92702 1 9757
2 92703 1 9761
2 92704 1 9761
2 92705 1 9762
2 92706 1 9762
2 92707 1 9771
2 92708 1 9771
2 92709 1 9775
2 92710 1 9775
2 92711 1 9809
2 92712 1 9809
2 92713 1 9809
2 92714 1 9811
2 92715 1 9811
2 92716 1 9811
2 92717 1 9869
2 92718 1 9869
2 92719 1 9869
2 92720 1 9869
2 92721 1 9869
2 92722 1 9870
2 92723 1 9870
2 92724 1 9872
2 92725 1 9872
2 92726 1 9873
2 92727 1 9873
2 92728 1 9874
2 92729 1 9874
2 92730 1 9876
2 92731 1 9876
2 92732 1 9891
2 92733 1 9891
2 92734 1 9892
2 92735 1 9892
2 92736 1 9893
2 92737 1 9893
2 92738 1 9894
2 92739 1 9894
2 92740 1 9894
2 92741 1 9894
2 92742 1 9895
2 92743 1 9895
2 92744 1 9899
2 92745 1 9899
2 92746 1 9899
2 92747 1 9900
2 92748 1 9900
2 92749 1 9905
2 92750 1 9905
2 92751 1 9908
2 92752 1 9908
2 92753 1 9908
2 92754 1 9908
2 92755 1 9908
2 92756 1 9908
2 92757 1 9908
2 92758 1 9908
2 92759 1 9908
2 92760 1 9908
2 92761 1 9925
2 92762 1 9925
2 92763 1 9925
2 92764 1 9925
2 92765 1 9925
2 92766 1 9925
2 92767 1 9925
2 92768 1 9925
2 92769 1 9925
2 92770 1 9925
2 92771 1 9925
2 92772 1 9925
2 92773 1 9925
2 92774 1 9925
2 92775 1 9925
2 92776 1 9925
2 92777 1 9926
2 92778 1 9926
2 92779 1 9926
2 92780 1 9926
2 92781 1 9926
2 92782 1 9926
2 92783 1 9929
2 92784 1 9929
2 92785 1 9938
2 92786 1 9938
2 92787 1 9938
2 92788 1 9938
2 92789 1 9939
2 92790 1 9939
2 92791 1 9956
2 92792 1 9956
2 92793 1 9960
2 92794 1 9960
2 92795 1 9960
2 92796 1 9960
2 92797 1 9960
2 92798 1 9960
2 92799 1 9969
2 92800 1 9969
2 92801 1 9970
2 92802 1 9970
2 92803 1 9970
2 92804 1 9984
2 92805 1 9984
2 92806 1 9984
2 92807 1 9984
2 92808 1 9984
2 92809 1 9984
2 92810 1 9984
2 92811 1 9985
2 92812 1 9985
2 92813 1 9986
2 92814 1 9986
2 92815 1 9986
2 92816 1 9986
2 92817 1 9989
2 92818 1 9989
2 92819 1 9990
2 92820 1 9990
2 92821 1 9990
2 92822 1 9990
2 92823 1 9990
2 92824 1 9990
2 92825 1 9990
2 92826 1 9990
2 92827 1 9990
2 92828 1 9990
2 92829 1 9990
2 92830 1 9990
2 92831 1 9990
2 92832 1 9992
2 92833 1 9992
2 92834 1 9999
2 92835 1 9999
2 92836 1 10000
2 92837 1 10000
2 92838 1 10000
2 92839 1 10000
2 92840 1 10000
2 92841 1 10000
2 92842 1 10000
2 92843 1 10000
2 92844 1 10000
2 92845 1 10000
2 92846 1 10000
2 92847 1 10001
2 92848 1 10001
2 92849 1 10001
2 92850 1 10002
2 92851 1 10002
2 92852 1 10002
2 92853 1 10002
2 92854 1 10002
2 92855 1 10002
2 92856 1 10002
2 92857 1 10011
2 92858 1 10011
2 92859 1 10011
2 92860 1 10011
2 92861 1 10011
2 92862 1 10011
2 92863 1 10011
2 92864 1 10011
2 92865 1 10019
2 92866 1 10019
2 92867 1 10019
2 92868 1 10019
2 92869 1 10019
2 92870 1 10019
2 92871 1 10019
2 92872 1 10020
2 92873 1 10020
2 92874 1 10033
2 92875 1 10033
2 92876 1 10034
2 92877 1 10034
2 92878 1 10035
2 92879 1 10035
2 92880 1 10035
2 92881 1 10036
2 92882 1 10036
2 92883 1 10037
2 92884 1 10037
2 92885 1 10055
2 92886 1 10055
2 92887 1 10055
2 92888 1 10055
2 92889 1 10067
2 92890 1 10067
2 92891 1 10067
2 92892 1 10073
2 92893 1 10073
2 92894 1 10073
2 92895 1 10073
2 92896 1 10073
2 92897 1 10073
2 92898 1 10073
2 92899 1 10073
2 92900 1 10073
2 92901 1 10074
2 92902 1 10074
2 92903 1 10087
2 92904 1 10087
2 92905 1 10108
2 92906 1 10108
2 92907 1 10108
2 92908 1 10108
2 92909 1 10108
2 92910 1 10108
2 92911 1 10108
2 92912 1 10108
2 92913 1 10108
2 92914 1 10109
2 92915 1 10109
2 92916 1 10110
2 92917 1 10110
2 92918 1 10115
2 92919 1 10115
2 92920 1 10115
2 92921 1 10137
2 92922 1 10137
2 92923 1 10137
2 92924 1 10137
2 92925 1 10137
2 92926 1 10137
2 92927 1 10137
2 92928 1 10137
2 92929 1 10137
2 92930 1 10138
2 92931 1 10138
2 92932 1 10138
2 92933 1 10138
2 92934 1 10140
2 92935 1 10140
2 92936 1 10152
2 92937 1 10152
2 92938 1 10152
2 92939 1 10152
2 92940 1 10152
2 92941 1 10154
2 92942 1 10154
2 92943 1 10154
2 92944 1 10155
2 92945 1 10155
2 92946 1 10155
2 92947 1 10155
2 92948 1 10158
2 92949 1 10158
2 92950 1 10172
2 92951 1 10172
2 92952 1 10172
2 92953 1 10186
2 92954 1 10186
2 92955 1 10186
2 92956 1 10186
2 92957 1 10186
2 92958 1 10187
2 92959 1 10187
2 92960 1 10195
2 92961 1 10195
2 92962 1 10195
2 92963 1 10220
2 92964 1 10220
2 92965 1 10220
2 92966 1 10220
2 92967 1 10220
2 92968 1 10220
2 92969 1 10220
2 92970 1 10220
2 92971 1 10220
2 92972 1 10222
2 92973 1 10222
2 92974 1 10222
2 92975 1 10224
2 92976 1 10224
2 92977 1 10224
2 92978 1 10227
2 92979 1 10227
2 92980 1 10227
2 92981 1 10227
2 92982 1 10227
2 92983 1 10228
2 92984 1 10228
2 92985 1 10228
2 92986 1 10235
2 92987 1 10235
2 92988 1 10235
2 92989 1 10235
2 92990 1 10235
2 92991 1 10236
2 92992 1 10236
2 92993 1 10249
2 92994 1 10249
2 92995 1 10249
2 92996 1 10249
2 92997 1 10251
2 92998 1 10251
2 92999 1 10273
2 93000 1 10273
2 93001 1 10273
2 93002 1 10273
2 93003 1 10273
2 93004 1 10273
2 93005 1 10273
2 93006 1 10273
2 93007 1 10273
2 93008 1 10273
2 93009 1 10273
2 93010 1 10273
2 93011 1 10273
2 93012 1 10273
2 93013 1 10273
2 93014 1 10273
2 93015 1 10273
2 93016 1 10273
2 93017 1 10273
2 93018 1 10273
2 93019 1 10273
2 93020 1 10273
2 93021 1 10273
2 93022 1 10273
2 93023 1 10273
2 93024 1 10273
2 93025 1 10273
2 93026 1 10273
2 93027 1 10274
2 93028 1 10274
2 93029 1 10275
2 93030 1 10275
2 93031 1 10278
2 93032 1 10278
2 93033 1 10278
2 93034 1 10295
2 93035 1 10295
2 93036 1 10299
2 93037 1 10299
2 93038 1 10299
2 93039 1 10299
2 93040 1 10299
2 93041 1 10299
2 93042 1 10299
2 93043 1 10299
2 93044 1 10299
2 93045 1 10299
2 93046 1 10299
2 93047 1 10299
2 93048 1 10300
2 93049 1 10300
2 93050 1 10308
2 93051 1 10308
2 93052 1 10308
2 93053 1 10308
2 93054 1 10308
2 93055 1 10308
2 93056 1 10308
2 93057 1 10308
2 93058 1 10308
2 93059 1 10308
2 93060 1 10308
2 93061 1 10308
2 93062 1 10308
2 93063 1 10308
2 93064 1 10308
2 93065 1 10309
2 93066 1 10309
2 93067 1 10317
2 93068 1 10317
2 93069 1 10317
2 93070 1 10317
2 93071 1 10317
2 93072 1 10320
2 93073 1 10320
2 93074 1 10320
2 93075 1 10333
2 93076 1 10333
2 93077 1 10333
2 93078 1 10333
2 93079 1 10334
2 93080 1 10334
2 93081 1 10334
2 93082 1 10334
2 93083 1 10334
2 93084 1 10337
2 93085 1 10337
2 93086 1 10337
2 93087 1 10337
2 93088 1 10337
2 93089 1 10337
2 93090 1 10337
2 93091 1 10337
2 93092 1 10337
2 93093 1 10337
2 93094 1 10337
2 93095 1 10337
2 93096 1 10338
2 93097 1 10338
2 93098 1 10343
2 93099 1 10343
2 93100 1 10346
2 93101 1 10346
2 93102 1 10346
2 93103 1 10346
2 93104 1 10346
2 93105 1 10346
2 93106 1 10346
2 93107 1 10346
2 93108 1 10346
2 93109 1 10346
2 93110 1 10347
2 93111 1 10347
2 93112 1 10347
2 93113 1 10347
2 93114 1 10347
2 93115 1 10347
2 93116 1 10355
2 93117 1 10355
2 93118 1 10355
2 93119 1 10355
2 93120 1 10355
2 93121 1 10355
2 93122 1 10355
2 93123 1 10356
2 93124 1 10356
2 93125 1 10357
2 93126 1 10357
2 93127 1 10357
2 93128 1 10357
2 93129 1 10357
2 93130 1 10359
2 93131 1 10359
2 93132 1 10361
2 93133 1 10361
2 93134 1 10369
2 93135 1 10369
2 93136 1 10370
2 93137 1 10370
2 93138 1 10370
2 93139 1 10370
2 93140 1 10370
2 93141 1 10370
2 93142 1 10370
2 93143 1 10370
2 93144 1 10370
2 93145 1 10378
2 93146 1 10378
2 93147 1 10378
2 93148 1 10378
2 93149 1 10380
2 93150 1 10380
2 93151 1 10390
2 93152 1 10390
2 93153 1 10390
2 93154 1 10390
2 93155 1 10390
2 93156 1 10390
2 93157 1 10390
2 93158 1 10390
2 93159 1 10390
2 93160 1 10393
2 93161 1 10393
2 93162 1 10393
2 93163 1 10393
2 93164 1 10393
2 93165 1 10394
2 93166 1 10394
2 93167 1 10394
2 93168 1 10401
2 93169 1 10401
2 93170 1 10408
2 93171 1 10408
2 93172 1 10416
2 93173 1 10416
2 93174 1 10416
2 93175 1 10416
2 93176 1 10416
2 93177 1 10424
2 93178 1 10424
2 93179 1 10424
2 93180 1 10435
2 93181 1 10435
2 93182 1 10435
2 93183 1 10435
2 93184 1 10437
2 93185 1 10437
2 93186 1 10437
2 93187 1 10444
2 93188 1 10444
2 93189 1 10444
2 93190 1 10444
2 93191 1 10444
2 93192 1 10444
2 93193 1 10445
2 93194 1 10445
2 93195 1 10445
2 93196 1 10445
2 93197 1 10453
2 93198 1 10453
2 93199 1 10456
2 93200 1 10456
2 93201 1 10456
2 93202 1 10457
2 93203 1 10457
2 93204 1 10470
2 93205 1 10470
2 93206 1 10486
2 93207 1 10486
2 93208 1 10489
2 93209 1 10489
2 93210 1 10489
2 93211 1 10489
2 93212 1 10489
2 93213 1 10489
2 93214 1 10489
2 93215 1 10489
2 93216 1 10489
2 93217 1 10489
2 93218 1 10489
2 93219 1 10489
2 93220 1 10489
2 93221 1 10489
2 93222 1 10489
2 93223 1 10489
2 93224 1 10505
2 93225 1 10505
2 93226 1 10505
2 93227 1 10506
2 93228 1 10506
2 93229 1 10506
2 93230 1 10506
2 93231 1 10507
2 93232 1 10507
2 93233 1 10509
2 93234 1 10509
2 93235 1 10509
2 93236 1 10511
2 93237 1 10511
2 93238 1 10511
2 93239 1 10511
2 93240 1 10511
2 93241 1 10511
2 93242 1 10511
2 93243 1 10511
2 93244 1 10511
2 93245 1 10518
2 93246 1 10518
2 93247 1 10518
2 93248 1 10518
2 93249 1 10518
2 93250 1 10518
2 93251 1 10518
2 93252 1 10518
2 93253 1 10518
2 93254 1 10518
2 93255 1 10518
2 93256 1 10518
2 93257 1 10518
2 93258 1 10518
2 93259 1 10518
2 93260 1 10518
2 93261 1 10518
2 93262 1 10518
2 93263 1 10518
2 93264 1 10518
2 93265 1 10518
2 93266 1 10518
2 93267 1 10520
2 93268 1 10520
2 93269 1 10520
2 93270 1 10548
2 93271 1 10548
2 93272 1 10553
2 93273 1 10553
2 93274 1 10567
2 93275 1 10567
2 93276 1 10568
2 93277 1 10568
2 93278 1 10576
2 93279 1 10576
2 93280 1 10576
2 93281 1 10584
2 93282 1 10584
2 93283 1 10584
2 93284 1 10586
2 93285 1 10586
2 93286 1 10586
2 93287 1 10587
2 93288 1 10587
2 93289 1 10587
2 93290 1 10588
2 93291 1 10588
2 93292 1 10589
2 93293 1 10589
2 93294 1 10593
2 93295 1 10593
2 93296 1 10593
2 93297 1 10593
2 93298 1 10604
2 93299 1 10604
2 93300 1 10607
2 93301 1 10607
2 93302 1 10607
2 93303 1 10651
2 93304 1 10651
2 93305 1 10691
2 93306 1 10691
2 93307 1 10691
2 93308 1 10691
2 93309 1 10691
2 93310 1 10691
2 93311 1 10691
2 93312 1 10691
2 93313 1 10692
2 93314 1 10692
2 93315 1 10692
2 93316 1 10692
2 93317 1 10693
2 93318 1 10693
2 93319 1 10693
2 93320 1 10693
2 93321 1 10693
2 93322 1 10694
2 93323 1 10694
2 93324 1 10694
2 93325 1 10694
2 93326 1 10694
2 93327 1 10694
2 93328 1 10694
2 93329 1 10694
2 93330 1 10705
2 93331 1 10705
2 93332 1 10705
2 93333 1 10721
2 93334 1 10721
2 93335 1 10722
2 93336 1 10722
2 93337 1 10751
2 93338 1 10751
2 93339 1 10751
2 93340 1 10760
2 93341 1 10760
2 93342 1 10760
2 93343 1 10760
2 93344 1 10760
2 93345 1 10760
2 93346 1 10765
2 93347 1 10765
2 93348 1 10765
2 93349 1 10765
2 93350 1 10765
2 93351 1 10765
2 93352 1 10765
2 93353 1 10765
2 93354 1 10765
2 93355 1 10767
2 93356 1 10767
2 93357 1 10767
2 93358 1 10767
2 93359 1 10767
2 93360 1 10776
2 93361 1 10776
2 93362 1 10776
2 93363 1 10776
2 93364 1 10777
2 93365 1 10777
2 93366 1 10778
2 93367 1 10778
2 93368 1 10778
2 93369 1 10824
2 93370 1 10824
2 93371 1 10824
2 93372 1 10844
2 93373 1 10844
2 93374 1 10846
2 93375 1 10846
2 93376 1 10846
2 93377 1 10846
2 93378 1 10846
2 93379 1 10846
2 93380 1 10848
2 93381 1 10848
2 93382 1 10866
2 93383 1 10866
2 93384 1 10866
2 93385 1 10871
2 93386 1 10871
2 93387 1 10871
2 93388 1 10876
2 93389 1 10876
2 93390 1 10876
2 93391 1 10877
2 93392 1 10877
2 93393 1 10877
2 93394 1 10877
2 93395 1 10877
2 93396 1 10877
2 93397 1 10877
2 93398 1 10894
2 93399 1 10894
2 93400 1 10894
2 93401 1 10894
2 93402 1 10894
2 93403 1 10895
2 93404 1 10895
2 93405 1 10896
2 93406 1 10896
2 93407 1 10900
2 93408 1 10900
2 93409 1 10901
2 93410 1 10901
2 93411 1 10901
2 93412 1 10901
2 93413 1 10901
2 93414 1 10915
2 93415 1 10915
2 93416 1 10915
2 93417 1 10915
2 93418 1 10915
2 93419 1 10915
2 93420 1 10920
2 93421 1 10920
2 93422 1 10936
2 93423 1 10936
2 93424 1 10936
2 93425 1 10936
2 93426 1 10936
2 93427 1 10936
2 93428 1 10937
2 93429 1 10937
2 93430 1 10946
2 93431 1 10946
2 93432 1 10947
2 93433 1 10947
2 93434 1 10947
2 93435 1 10947
2 93436 1 10948
2 93437 1 10948
2 93438 1 10948
2 93439 1 10948
2 93440 1 10949
2 93441 1 10949
2 93442 1 10949
2 93443 1 10949
2 93444 1 10954
2 93445 1 10954
2 93446 1 10954
2 93447 1 10954
2 93448 1 10954
2 93449 1 10954
2 93450 1 10954
2 93451 1 10967
2 93452 1 10967
2 93453 1 10967
2 93454 1 10967
2 93455 1 10967
2 93456 1 10967
2 93457 1 10967
2 93458 1 10967
2 93459 1 10967
2 93460 1 10967
2 93461 1 10984
2 93462 1 10984
2 93463 1 10997
2 93464 1 10997
2 93465 1 11013
2 93466 1 11013
2 93467 1 11013
2 93468 1 11013
2 93469 1 11014
2 93470 1 11014
2 93471 1 11028
2 93472 1 11028
2 93473 1 11028
2 93474 1 11028
2 93475 1 11028
2 93476 1 11028
2 93477 1 11028
2 93478 1 11029
2 93479 1 11029
2 93480 1 11029
2 93481 1 11029
2 93482 1 11030
2 93483 1 11030
2 93484 1 11045
2 93485 1 11045
2 93486 1 11062
2 93487 1 11062
2 93488 1 11062
2 93489 1 11062
2 93490 1 11068
2 93491 1 11068
2 93492 1 11076
2 93493 1 11076
2 93494 1 11079
2 93495 1 11079
2 93496 1 11079
2 93497 1 11079
2 93498 1 11079
2 93499 1 11080
2 93500 1 11080
2 93501 1 11096
2 93502 1 11096
2 93503 1 11096
2 93504 1 11096
2 93505 1 11101
2 93506 1 11101
2 93507 1 11118
2 93508 1 11118
2 93509 1 11118
2 93510 1 11119
2 93511 1 11119
2 93512 1 11128
2 93513 1 11128
2 93514 1 11128
2 93515 1 11130
2 93516 1 11130
2 93517 1 11130
2 93518 1 11130
2 93519 1 11130
2 93520 1 11131
2 93521 1 11131
2 93522 1 11131
2 93523 1 11134
2 93524 1 11134
2 93525 1 11134
2 93526 1 11134
2 93527 1 11134
2 93528 1 11134
2 93529 1 11134
2 93530 1 11134
2 93531 1 11134
2 93532 1 11134
2 93533 1 11134
2 93534 1 11135
2 93535 1 11135
2 93536 1 11135
2 93537 1 11135
2 93538 1 11150
2 93539 1 11150
2 93540 1 11151
2 93541 1 11151
2 93542 1 11151
2 93543 1 11165
2 93544 1 11165
2 93545 1 11183
2 93546 1 11183
2 93547 1 11183
2 93548 1 11184
2 93549 1 11184
2 93550 1 11185
2 93551 1 11185
2 93552 1 11193
2 93553 1 11193
2 93554 1 11205
2 93555 1 11205
2 93556 1 11208
2 93557 1 11208
2 93558 1 11208
2 93559 1 11208
2 93560 1 11208
2 93561 1 11208
2 93562 1 11208
2 93563 1 11209
2 93564 1 11209
2 93565 1 11212
2 93566 1 11212
2 93567 1 11220
2 93568 1 11220
2 93569 1 11220
2 93570 1 11220
2 93571 1 11220
2 93572 1 11221
2 93573 1 11221
2 93574 1 11221
2 93575 1 11221
2 93576 1 11221
2 93577 1 11221
2 93578 1 11252
2 93579 1 11252
2 93580 1 11253
2 93581 1 11253
2 93582 1 11253
2 93583 1 11253
2 93584 1 11253
2 93585 1 11253
2 93586 1 11253
2 93587 1 11253
2 93588 1 11253
2 93589 1 11253
2 93590 1 11253
2 93591 1 11254
2 93592 1 11254
2 93593 1 11254
2 93594 1 11254
2 93595 1 11254
2 93596 1 11254
2 93597 1 11254
2 93598 1 11254
2 93599 1 11255
2 93600 1 11255
2 93601 1 11255
2 93602 1 11265
2 93603 1 11265
2 93604 1 11265
2 93605 1 11265
2 93606 1 11265
2 93607 1 11265
2 93608 1 11265
2 93609 1 11265
2 93610 1 11265
2 93611 1 11265
2 93612 1 11265
2 93613 1 11265
2 93614 1 11266
2 93615 1 11266
2 93616 1 11266
2 93617 1 11266
2 93618 1 11266
2 93619 1 11266
2 93620 1 11266
2 93621 1 11266
2 93622 1 11266
2 93623 1 11267
2 93624 1 11267
2 93625 1 11267
2 93626 1 11267
2 93627 1 11267
2 93628 1 11267
2 93629 1 11268
2 93630 1 11268
2 93631 1 11268
2 93632 1 11268
2 93633 1 11286
2 93634 1 11286
2 93635 1 11286
2 93636 1 11297
2 93637 1 11297
2 93638 1 11297
2 93639 1 11297
2 93640 1 11297
2 93641 1 11298
2 93642 1 11298
2 93643 1 11298
2 93644 1 11298
2 93645 1 11298
2 93646 1 11301
2 93647 1 11301
2 93648 1 11301
2 93649 1 11301
2 93650 1 11301
2 93651 1 11301
2 93652 1 11301
2 93653 1 11303
2 93654 1 11303
2 93655 1 11304
2 93656 1 11304
2 93657 1 11304
2 93658 1 11304
2 93659 1 11304
2 93660 1 11304
2 93661 1 11304
2 93662 1 11304
2 93663 1 11304
2 93664 1 11304
2 93665 1 11314
2 93666 1 11314
2 93667 1 11314
2 93668 1 11314
2 93669 1 11314
2 93670 1 11314
2 93671 1 11314
2 93672 1 11314
2 93673 1 11315
2 93674 1 11315
2 93675 1 11316
2 93676 1 11316
2 93677 1 11319
2 93678 1 11319
2 93679 1 11319
2 93680 1 11329
2 93681 1 11329
2 93682 1 11330
2 93683 1 11330
2 93684 1 11330
2 93685 1 11330
2 93686 1 11330
2 93687 1 11330
2 93688 1 11332
2 93689 1 11332
2 93690 1 11332
2 93691 1 11333
2 93692 1 11333
2 93693 1 11333
2 93694 1 11333
2 93695 1 11345
2 93696 1 11345
2 93697 1 11345
2 93698 1 11345
2 93699 1 11345
2 93700 1 11345
2 93701 1 11345
2 93702 1 11345
2 93703 1 11345
2 93704 1 11345
2 93705 1 11345
2 93706 1 11345
2 93707 1 11345
2 93708 1 11345
2 93709 1 11345
2 93710 1 11345
2 93711 1 11345
2 93712 1 11345
2 93713 1 11345
2 93714 1 11345
2 93715 1 11345
2 93716 1 11345
2 93717 1 11345
2 93718 1 11356
2 93719 1 11356
2 93720 1 11356
2 93721 1 11356
2 93722 1 11356
2 93723 1 11356
2 93724 1 11362
2 93725 1 11362
2 93726 1 11362
2 93727 1 11362
2 93728 1 11362
2 93729 1 11362
2 93730 1 11362
2 93731 1 11362
2 93732 1 11362
2 93733 1 11362
2 93734 1 11362
2 93735 1 11362
2 93736 1 11362
2 93737 1 11362
2 93738 1 11362
2 93739 1 11362
2 93740 1 11362
2 93741 1 11362
2 93742 1 11362
2 93743 1 11362
2 93744 1 11363
2 93745 1 11363
2 93746 1 11372
2 93747 1 11372
2 93748 1 11372
2 93749 1 11372
2 93750 1 11372
2 93751 1 11372
2 93752 1 11372
2 93753 1 11372
2 93754 1 11373
2 93755 1 11373
2 93756 1 11373
2 93757 1 11373
2 93758 1 11373
2 93759 1 11373
2 93760 1 11375
2 93761 1 11375
2 93762 1 11376
2 93763 1 11376
2 93764 1 11376
2 93765 1 11376
2 93766 1 11376
2 93767 1 11376
2 93768 1 11376
2 93769 1 11376
2 93770 1 11377
2 93771 1 11377
2 93772 1 11399
2 93773 1 11399
2 93774 1 11399
2 93775 1 11401
2 93776 1 11401
2 93777 1 11402
2 93778 1 11402
2 93779 1 11402
2 93780 1 11403
2 93781 1 11403
2 93782 1 11404
2 93783 1 11404
2 93784 1 11405
2 93785 1 11405
2 93786 1 11406
2 93787 1 11406
2 93788 1 11406
2 93789 1 11408
2 93790 1 11408
2 93791 1 11411
2 93792 1 11411
2 93793 1 11413
2 93794 1 11413
2 93795 1 11413
2 93796 1 11414
2 93797 1 11414
2 93798 1 11414
2 93799 1 11414
2 93800 1 11414
2 93801 1 11421
2 93802 1 11421
2 93803 1 11421
2 93804 1 11421
2 93805 1 11421
2 93806 1 11421
2 93807 1 11422
2 93808 1 11422
2 93809 1 11422
2 93810 1 11422
2 93811 1 11422
2 93812 1 11422
2 93813 1 11422
2 93814 1 11422
2 93815 1 11422
2 93816 1 11422
2 93817 1 11424
2 93818 1 11424
2 93819 1 11424
2 93820 1 11424
2 93821 1 11424
2 93822 1 11425
2 93823 1 11425
2 93824 1 11427
2 93825 1 11427
2 93826 1 11427
2 93827 1 11427
2 93828 1 11427
2 93829 1 11428
2 93830 1 11428
2 93831 1 11428
2 93832 1 11428
2 93833 1 11432
2 93834 1 11432
2 93835 1 11433
2 93836 1 11433
2 93837 1 11433
2 93838 1 11434
2 93839 1 11434
2 93840 1 11434
2 93841 1 11447
2 93842 1 11447
2 93843 1 11447
2 93844 1 11447
2 93845 1 11447
2 93846 1 11447
2 93847 1 11447
2 93848 1 11447
2 93849 1 11447
2 93850 1 11447
2 93851 1 11447
2 93852 1 11447
2 93853 1 11448
2 93854 1 11448
2 93855 1 11448
2 93856 1 11448
2 93857 1 11449
2 93858 1 11449
2 93859 1 11450
2 93860 1 11450
2 93861 1 11453
2 93862 1 11453
2 93863 1 11453
2 93864 1 11453
2 93865 1 11453
2 93866 1 11453
2 93867 1 11453
2 93868 1 11455
2 93869 1 11455
2 93870 1 11458
2 93871 1 11458
2 93872 1 11472
2 93873 1 11472
2 93874 1 11477
2 93875 1 11477
2 93876 1 11477
2 93877 1 11477
2 93878 1 11477
2 93879 1 11477
2 93880 1 11482
2 93881 1 11482
2 93882 1 11482
2 93883 1 11482
2 93884 1 11482
2 93885 1 11482
2 93886 1 11482
2 93887 1 11482
2 93888 1 11483
2 93889 1 11483
2 93890 1 11487
2 93891 1 11487
2 93892 1 11503
2 93893 1 11503
2 93894 1 11503
2 93895 1 11503
2 93896 1 11503
2 93897 1 11504
2 93898 1 11504
2 93899 1 11504
2 93900 1 11516
2 93901 1 11516
2 93902 1 11517
2 93903 1 11517
2 93904 1 11518
2 93905 1 11518
2 93906 1 11518
2 93907 1 11518
2 93908 1 11519
2 93909 1 11519
2 93910 1 11525
2 93911 1 11525
2 93912 1 11531
2 93913 1 11531
2 93914 1 11534
2 93915 1 11534
2 93916 1 11534
2 93917 1 11546
2 93918 1 11546
2 93919 1 11547
2 93920 1 11547
2 93921 1 11567
2 93922 1 11567
2 93923 1 11568
2 93924 1 11568
2 93925 1 11568
2 93926 1 11568
2 93927 1 11569
2 93928 1 11569
2 93929 1 11570
2 93930 1 11570
2 93931 1 11570
2 93932 1 11570
2 93933 1 11570
2 93934 1 11570
2 93935 1 11570
2 93936 1 11571
2 93937 1 11571
2 93938 1 11571
2 93939 1 11582
2 93940 1 11582
2 93941 1 11582
2 93942 1 11582
2 93943 1 11584
2 93944 1 11584
2 93945 1 11585
2 93946 1 11585
2 93947 1 11585
2 93948 1 11587
2 93949 1 11587
2 93950 1 11589
2 93951 1 11589
2 93952 1 11589
2 93953 1 11591
2 93954 1 11591
2 93955 1 11600
2 93956 1 11600
2 93957 1 11600
2 93958 1 11600
2 93959 1 11601
2 93960 1 11601
2 93961 1 11602
2 93962 1 11602
2 93963 1 11603
2 93964 1 11603
2 93965 1 11610
2 93966 1 11610
2 93967 1 11610
2 93968 1 11610
2 93969 1 11610
2 93970 1 11610
2 93971 1 11611
2 93972 1 11611
2 93973 1 11612
2 93974 1 11612
2 93975 1 11634
2 93976 1 11634
2 93977 1 11635
2 93978 1 11635
2 93979 1 11635
2 93980 1 11635
2 93981 1 11635
2 93982 1 11637
2 93983 1 11637
2 93984 1 11637
2 93985 1 11637
2 93986 1 11646
2 93987 1 11646
2 93988 1 11659
2 93989 1 11659
2 93990 1 11659
2 93991 1 11660
2 93992 1 11660
2 93993 1 11674
2 93994 1 11674
2 93995 1 11682
2 93996 1 11682
2 93997 1 11690
2 93998 1 11690
2 93999 1 11690
2 94000 1 11690
2 94001 1 11691
2 94002 1 11691
2 94003 1 11692
2 94004 1 11692
2 94005 1 11692
2 94006 1 11703
2 94007 1 11703
2 94008 1 11711
2 94009 1 11711
2 94010 1 11711
2 94011 1 11711
2 94012 1 11711
2 94013 1 11719
2 94014 1 11719
2 94015 1 11721
2 94016 1 11721
2 94017 1 11721
2 94018 1 11737
2 94019 1 11737
2 94020 1 11737
2 94021 1 11739
2 94022 1 11739
2 94023 1 11739
2 94024 1 11754
2 94025 1 11754
2 94026 1 11760
2 94027 1 11760
2 94028 1 11768
2 94029 1 11768
2 94030 1 11768
2 94031 1 11768
2 94032 1 11768
2 94033 1 11768
2 94034 1 11769
2 94035 1 11769
2 94036 1 11769
2 94037 1 11774
2 94038 1 11774
2 94039 1 11781
2 94040 1 11781
2 94041 1 11790
2 94042 1 11790
2 94043 1 11791
2 94044 1 11791
2 94045 1 11791
2 94046 1 11808
2 94047 1 11808
2 94048 1 11808
2 94049 1 11811
2 94050 1 11811
2 94051 1 11816
2 94052 1 11816
2 94053 1 11836
2 94054 1 11836
2 94055 1 11836
2 94056 1 11836
2 94057 1 11836
2 94058 1 11868
2 94059 1 11868
2 94060 1 11868
2 94061 1 11869
2 94062 1 11869
2 94063 1 11869
2 94064 1 11869
2 94065 1 11869
2 94066 1 11870
2 94067 1 11870
2 94068 1 11870
2 94069 1 11878
2 94070 1 11878
2 94071 1 11878
2 94072 1 11878
2 94073 1 11878
2 94074 1 11878
2 94075 1 11878
2 94076 1 11879
2 94077 1 11879
2 94078 1 11882
2 94079 1 11882
2 94080 1 11882
2 94081 1 11882
2 94082 1 11882
2 94083 1 11882
2 94084 1 11882
2 94085 1 11882
2 94086 1 11882
2 94087 1 11882
2 94088 1 11882
2 94089 1 11890
2 94090 1 11890
2 94091 1 11899
2 94092 1 11899
2 94093 1 11899
2 94094 1 11921
2 94095 1 11921
2 94096 1 11921
2 94097 1 11921
2 94098 1 11928
2 94099 1 11928
2 94100 1 11928
2 94101 1 11967
2 94102 1 11967
2 94103 1 11968
2 94104 1 11968
2 94105 1 11968
2 94106 1 11968
2 94107 1 11969
2 94108 1 11969
2 94109 1 11978
2 94110 1 11978
2 94111 1 11978
2 94112 1 11979
2 94113 1 11979
2 94114 1 11979
2 94115 1 11982
2 94116 1 11982
2 94117 1 11983
2 94118 1 11983
2 94119 1 11998
2 94120 1 11998
2 94121 1 11999
2 94122 1 11999
2 94123 1 12001
2 94124 1 12001
2 94125 1 12001
2 94126 1 12002
2 94127 1 12002
2 94128 1 12002
2 94129 1 12011
2 94130 1 12011
2 94131 1 12012
2 94132 1 12012
2 94133 1 12013
2 94134 1 12013
2 94135 1 12013
2 94136 1 12013
2 94137 1 12013
2 94138 1 12013
2 94139 1 12013
2 94140 1 12013
2 94141 1 12013
2 94142 1 12024
2 94143 1 12024
2 94144 1 12024
2 94145 1 12025
2 94146 1 12025
2 94147 1 12030
2 94148 1 12030
2 94149 1 12030
2 94150 1 12030
2 94151 1 12044
2 94152 1 12044
2 94153 1 12045
2 94154 1 12045
2 94155 1 12052
2 94156 1 12052
2 94157 1 12052
2 94158 1 12054
2 94159 1 12054
2 94160 1 12055
2 94161 1 12055
2 94162 1 12056
2 94163 1 12056
2 94164 1 12083
2 94165 1 12083
2 94166 1 12098
2 94167 1 12098
2 94168 1 12098
2 94169 1 12098
2 94170 1 12104
2 94171 1 12104
2 94172 1 12107
2 94173 1 12107
2 94174 1 12107
2 94175 1 12107
2 94176 1 12107
2 94177 1 12108
2 94178 1 12108
2 94179 1 12109
2 94180 1 12109
2 94181 1 12116
2 94182 1 12116
2 94183 1 12117
2 94184 1 12117
2 94185 1 12117
2 94186 1 12117
2 94187 1 12117
2 94188 1 12119
2 94189 1 12119
2 94190 1 12119
2 94191 1 12120
2 94192 1 12120
2 94193 1 12121
2 94194 1 12121
2 94195 1 12122
2 94196 1 12122
2 94197 1 12134
2 94198 1 12134
2 94199 1 12149
2 94200 1 12149
2 94201 1 12150
2 94202 1 12150
2 94203 1 12155
2 94204 1 12155
2 94205 1 12157
2 94206 1 12157
2 94207 1 12157
2 94208 1 12157
2 94209 1 12157
2 94210 1 12157
2 94211 1 12191
2 94212 1 12191
2 94213 1 12194
2 94214 1 12194
2 94215 1 12200
2 94216 1 12200
2 94217 1 12200
2 94218 1 12200
2 94219 1 12200
2 94220 1 12200
2 94221 1 12202
2 94222 1 12202
2 94223 1 12209
2 94224 1 12209
2 94225 1 12209
2 94226 1 12209
2 94227 1 12209
2 94228 1 12217
2 94229 1 12217
2 94230 1 12217
2 94231 1 12231
2 94232 1 12231
2 94233 1 12231
2 94234 1 12231
2 94235 1 12231
2 94236 1 12231
2 94237 1 12231
2 94238 1 12231
2 94239 1 12232
2 94240 1 12232
2 94241 1 12232
2 94242 1 12232
2 94243 1 12232
2 94244 1 12233
2 94245 1 12233
2 94246 1 12233
2 94247 1 12233
2 94248 1 12233
2 94249 1 12237
2 94250 1 12237
2 94251 1 12237
2 94252 1 12245
2 94253 1 12245
2 94254 1 12246
2 94255 1 12246
2 94256 1 12247
2 94257 1 12247
2 94258 1 12248
2 94259 1 12248
2 94260 1 12248
2 94261 1 12248
2 94262 1 12249
2 94263 1 12249
2 94264 1 12249
2 94265 1 12249
2 94266 1 12249
2 94267 1 12249
2 94268 1 12249
2 94269 1 12249
2 94270 1 12249
2 94271 1 12249
2 94272 1 12250
2 94273 1 12250
2 94274 1 12250
2 94275 1 12250
2 94276 1 12251
2 94277 1 12251
2 94278 1 12251
2 94279 1 12252
2 94280 1 12252
2 94281 1 12252
2 94282 1 12252
2 94283 1 12252
2 94284 1 12252
2 94285 1 12252
2 94286 1 12252
2 94287 1 12253
2 94288 1 12253
2 94289 1 12253
2 94290 1 12253
2 94291 1 12253
2 94292 1 12253
2 94293 1 12253
2 94294 1 12264
2 94295 1 12264
2 94296 1 12265
2 94297 1 12265
2 94298 1 12265
2 94299 1 12267
2 94300 1 12267
2 94301 1 12273
2 94302 1 12273
2 94303 1 12277
2 94304 1 12277
2 94305 1 12280
2 94306 1 12280
2 94307 1 12280
2 94308 1 12280
2 94309 1 12317
2 94310 1 12317
2 94311 1 12317
2 94312 1 12317
2 94313 1 12317
2 94314 1 12319
2 94315 1 12319
2 94316 1 12321
2 94317 1 12321
2 94318 1 12321
2 94319 1 12321
2 94320 1 12323
2 94321 1 12323
2 94322 1 12323
2 94323 1 12323
2 94324 1 12323
2 94325 1 12323
2 94326 1 12324
2 94327 1 12324
2 94328 1 12324
2 94329 1 12324
2 94330 1 12324
2 94331 1 12341
2 94332 1 12341
2 94333 1 12350
2 94334 1 12350
2 94335 1 12351
2 94336 1 12351
2 94337 1 12359
2 94338 1 12359
2 94339 1 12359
2 94340 1 12359
2 94341 1 12360
2 94342 1 12360
2 94343 1 12360
2 94344 1 12361
2 94345 1 12361
2 94346 1 12371
2 94347 1 12371
2 94348 1 12380
2 94349 1 12380
2 94350 1 12386
2 94351 1 12386
2 94352 1 12398
2 94353 1 12398
2 94354 1 12398
2 94355 1 12398
2 94356 1 12399
2 94357 1 12399
2 94358 1 12399
2 94359 1 12400
2 94360 1 12400
2 94361 1 12400
2 94362 1 12400
2 94363 1 12403
2 94364 1 12403
2 94365 1 12410
2 94366 1 12410
2 94367 1 12410
2 94368 1 12412
2 94369 1 12412
2 94370 1 12426
2 94371 1 12426
2 94372 1 12426
2 94373 1 12426
2 94374 1 12426
2 94375 1 12440
2 94376 1 12440
2 94377 1 12443
2 94378 1 12443
2 94379 1 12443
2 94380 1 12451
2 94381 1 12451
2 94382 1 12451
2 94383 1 12452
2 94384 1 12452
2 94385 1 12452
2 94386 1 12453
2 94387 1 12453
2 94388 1 12453
2 94389 1 12454
2 94390 1 12454
2 94391 1 12454
2 94392 1 12458
2 94393 1 12458
2 94394 1 12474
2 94395 1 12474
2 94396 1 12474
2 94397 1 12474
2 94398 1 12474
2 94399 1 12474
2 94400 1 12476
2 94401 1 12476
2 94402 1 12486
2 94403 1 12486
2 94404 1 12494
2 94405 1 12494
2 94406 1 12495
2 94407 1 12495
2 94408 1 12496
2 94409 1 12496
2 94410 1 12496
2 94411 1 12504
2 94412 1 12504
2 94413 1 12504
2 94414 1 12505
2 94415 1 12505
2 94416 1 12506
2 94417 1 12506
2 94418 1 12519
2 94419 1 12519
2 94420 1 12521
2 94421 1 12521
2 94422 1 12532
2 94423 1 12532
2 94424 1 12536
2 94425 1 12536
2 94426 1 12537
2 94427 1 12537
2 94428 1 12539
2 94429 1 12539
2 94430 1 12540
2 94431 1 12540
2 94432 1 12540
2 94433 1 12540
2 94434 1 12549
2 94435 1 12549
2 94436 1 12549
2 94437 1 12549
2 94438 1 12549
2 94439 1 12550
2 94440 1 12550
2 94441 1 12550
2 94442 1 12550
2 94443 1 12550
2 94444 1 12551
2 94445 1 12551
2 94446 1 12551
2 94447 1 12551
2 94448 1 12551
2 94449 1 12552
2 94450 1 12552
2 94451 1 12556
2 94452 1 12556
2 94453 1 12557
2 94454 1 12557
2 94455 1 12569
2 94456 1 12569
2 94457 1 12569
2 94458 1 12591
2 94459 1 12591
2 94460 1 12604
2 94461 1 12604
2 94462 1 12607
2 94463 1 12607
2 94464 1 12625
2 94465 1 12625
2 94466 1 12625
2 94467 1 12626
2 94468 1 12626
2 94469 1 12626
2 94470 1 12626
2 94471 1 12626
2 94472 1 12626
2 94473 1 12626
2 94474 1 12626
2 94475 1 12626
2 94476 1 12626
2 94477 1 12626
2 94478 1 12626
2 94479 1 12626
2 94480 1 12634
2 94481 1 12634
2 94482 1 12634
2 94483 1 12634
2 94484 1 12634
2 94485 1 12634
2 94486 1 12634
2 94487 1 12634
2 94488 1 12635
2 94489 1 12635
2 94490 1 12638
2 94491 1 12638
2 94492 1 12645
2 94493 1 12645
2 94494 1 12656
2 94495 1 12656
2 94496 1 12656
2 94497 1 12656
2 94498 1 12656
2 94499 1 12657
2 94500 1 12657
2 94501 1 12657
2 94502 1 12657
2 94503 1 12663
2 94504 1 12663
2 94505 1 12664
2 94506 1 12664
2 94507 1 12675
2 94508 1 12675
2 94509 1 12675
2 94510 1 12675
2 94511 1 12675
2 94512 1 12675
2 94513 1 12675
2 94514 1 12684
2 94515 1 12684
2 94516 1 12692
2 94517 1 12692
2 94518 1 12701
2 94519 1 12701
2 94520 1 12715
2 94521 1 12715
2 94522 1 12716
2 94523 1 12716
2 94524 1 12716
2 94525 1 12725
2 94526 1 12725
2 94527 1 12725
2 94528 1 12725
2 94529 1 12725
2 94530 1 12731
2 94531 1 12731
2 94532 1 12731
2 94533 1 12731
2 94534 1 12731
2 94535 1 12731
2 94536 1 12735
2 94537 1 12735
2 94538 1 12765
2 94539 1 12765
2 94540 1 12766
2 94541 1 12766
2 94542 1 12771
2 94543 1 12771
2 94544 1 12794
2 94545 1 12794
2 94546 1 12794
2 94547 1 12794
2 94548 1 12794
2 94549 1 12795
2 94550 1 12795
2 94551 1 12795
2 94552 1 12795
2 94553 1 12795
2 94554 1 12798
2 94555 1 12798
2 94556 1 12807
2 94557 1 12807
2 94558 1 12821
2 94559 1 12821
2 94560 1 12822
2 94561 1 12822
2 94562 1 12822
2 94563 1 12822
2 94564 1 12822
2 94565 1 12822
2 94566 1 12822
2 94567 1 12822
2 94568 1 12822
2 94569 1 12823
2 94570 1 12823
2 94571 1 12823
2 94572 1 12823
2 94573 1 12823
2 94574 1 12824
2 94575 1 12824
2 94576 1 12832
2 94577 1 12832
2 94578 1 12832
2 94579 1 12832
2 94580 1 12835
2 94581 1 12835
2 94582 1 12835
2 94583 1 12843
2 94584 1 12843
2 94585 1 12843
2 94586 1 12843
2 94587 1 12843
2 94588 1 12843
2 94589 1 12843
2 94590 1 12843
2 94591 1 12843
2 94592 1 12843
2 94593 1 12843
2 94594 1 12843
2 94595 1 12843
2 94596 1 12843
2 94597 1 12844
2 94598 1 12844
2 94599 1 12844
2 94600 1 12844
2 94601 1 12844
2 94602 1 12845
2 94603 1 12845
2 94604 1 12846
2 94605 1 12846
2 94606 1 12846
2 94607 1 12848
2 94608 1 12848
2 94609 1 12866
2 94610 1 12866
2 94611 1 12866
2 94612 1 12866
2 94613 1 12866
2 94614 1 12868
2 94615 1 12868
2 94616 1 12876
2 94617 1 12876
2 94618 1 12876
2 94619 1 12876
2 94620 1 12877
2 94621 1 12877
2 94622 1 12899
2 94623 1 12899
2 94624 1 12899
2 94625 1 12899
2 94626 1 12907
2 94627 1 12907
2 94628 1 12907
2 94629 1 12908
2 94630 1 12908
2 94631 1 12908
2 94632 1 12908
2 94633 1 12919
2 94634 1 12919
2 94635 1 12932
2 94636 1 12932
2 94637 1 12932
2 94638 1 12955
2 94639 1 12955
2 94640 1 12969
2 94641 1 12969
2 94642 1 12969
2 94643 1 12987
2 94644 1 12987
2 94645 1 12988
2 94646 1 12988
2 94647 1 12988
2 94648 1 12988
2 94649 1 12988
2 94650 1 12990
2 94651 1 12990
2 94652 1 13006
2 94653 1 13006
2 94654 1 13021
2 94655 1 13021
2 94656 1 13021
2 94657 1 13021
2 94658 1 13021
2 94659 1 13021
2 94660 1 13021
2 94661 1 13021
2 94662 1 13058
2 94663 1 13058
2 94664 1 13058
2 94665 1 13059
2 94666 1 13059
2 94667 1 13060
2 94668 1 13060
2 94669 1 13060
2 94670 1 13060
2 94671 1 13060
2 94672 1 13062
2 94673 1 13062
2 94674 1 13062
2 94675 1 13075
2 94676 1 13075
2 94677 1 13075
2 94678 1 13082
2 94679 1 13082
2 94680 1 13084
2 94681 1 13084
2 94682 1 13118
2 94683 1 13118
2 94684 1 13118
2 94685 1 13118
2 94686 1 13118
2 94687 1 13118
2 94688 1 13119
2 94689 1 13119
2 94690 1 13119
2 94691 1 13119
2 94692 1 13119
2 94693 1 13119
2 94694 1 13120
2 94695 1 13120
2 94696 1 13120
2 94697 1 13121
2 94698 1 13121
2 94699 1 13122
2 94700 1 13122
2 94701 1 13122
2 94702 1 13122
2 94703 1 13130
2 94704 1 13130
2 94705 1 13141
2 94706 1 13141
2 94707 1 13182
2 94708 1 13182
2 94709 1 13193
2 94710 1 13193
2 94711 1 13195
2 94712 1 13195
2 94713 1 13196
2 94714 1 13196
2 94715 1 13207
2 94716 1 13207
2 94717 1 13207
2 94718 1 13207
2 94719 1 13207
2 94720 1 13208
2 94721 1 13208
2 94722 1 13208
2 94723 1 13210
2 94724 1 13210
2 94725 1 13210
2 94726 1 13210
2 94727 1 13210
2 94728 1 13210
2 94729 1 13211
2 94730 1 13211
2 94731 1 13211
2 94732 1 13211
2 94733 1 13222
2 94734 1 13222
2 94735 1 13222
2 94736 1 13222
2 94737 1 13222
2 94738 1 13224
2 94739 1 13224
2 94740 1 13226
2 94741 1 13226
2 94742 1 13228
2 94743 1 13228
2 94744 1 13243
2 94745 1 13243
2 94746 1 13243
2 94747 1 13244
2 94748 1 13244
2 94749 1 13246
2 94750 1 13246
2 94751 1 13246
2 94752 1 13246
2 94753 1 13246
2 94754 1 13246
2 94755 1 13247
2 94756 1 13247
2 94757 1 13247
2 94758 1 13247
2 94759 1 13247
2 94760 1 13247
2 94761 1 13247
2 94762 1 13248
2 94763 1 13248
2 94764 1 13250
2 94765 1 13250
2 94766 1 13250
2 94767 1 13250
2 94768 1 13255
2 94769 1 13255
2 94770 1 13255
2 94771 1 13258
2 94772 1 13258
2 94773 1 13263
2 94774 1 13263
2 94775 1 13263
2 94776 1 13263
2 94777 1 13263
2 94778 1 13263
2 94779 1 13263
2 94780 1 13263
2 94781 1 13263
2 94782 1 13263
2 94783 1 13263
2 94784 1 13263
2 94785 1 13264
2 94786 1 13264
2 94787 1 13264
2 94788 1 13265
2 94789 1 13265
2 94790 1 13273
2 94791 1 13273
2 94792 1 13275
2 94793 1 13275
2 94794 1 13281
2 94795 1 13281
2 94796 1 13281
2 94797 1 13288
2 94798 1 13288
2 94799 1 13288
2 94800 1 13288
2 94801 1 13288
2 94802 1 13288
2 94803 1 13288
2 94804 1 13288
2 94805 1 13288
2 94806 1 13289
2 94807 1 13289
2 94808 1 13289
2 94809 1 13289
2 94810 1 13294
2 94811 1 13294
2 94812 1 13294
2 94813 1 13295
2 94814 1 13295
2 94815 1 13295
2 94816 1 13295
2 94817 1 13295
2 94818 1 13295
2 94819 1 13295
2 94820 1 13309
2 94821 1 13309
2 94822 1 13309
2 94823 1 13310
2 94824 1 13310
2 94825 1 13311
2 94826 1 13311
2 94827 1 13312
2 94828 1 13312
2 94829 1 13319
2 94830 1 13319
2 94831 1 13319
2 94832 1 13319
2 94833 1 13319
2 94834 1 13327
2 94835 1 13327
2 94836 1 13327
2 94837 1 13327
2 94838 1 13327
2 94839 1 13327
2 94840 1 13327
2 94841 1 13327
2 94842 1 13328
2 94843 1 13328
2 94844 1 13331
2 94845 1 13331
2 94846 1 13332
2 94847 1 13332
2 94848 1 13335
2 94849 1 13335
2 94850 1 13335
2 94851 1 13345
2 94852 1 13345
2 94853 1 13345
2 94854 1 13347
2 94855 1 13347
2 94856 1 13352
2 94857 1 13352
2 94858 1 13353
2 94859 1 13353
2 94860 1 13353
2 94861 1 13353
2 94862 1 13353
2 94863 1 13353
2 94864 1 13353
2 94865 1 13353
2 94866 1 13353
2 94867 1 13354
2 94868 1 13354
2 94869 1 13354
2 94870 1 13369
2 94871 1 13369
2 94872 1 13372
2 94873 1 13372
2 94874 1 13385
2 94875 1 13385
2 94876 1 13397
2 94877 1 13397
2 94878 1 13400
2 94879 1 13400
2 94880 1 13400
2 94881 1 13429
2 94882 1 13429
2 94883 1 13441
2 94884 1 13441
2 94885 1 13442
2 94886 1 13442
2 94887 1 13450
2 94888 1 13450
2 94889 1 13450
2 94890 1 13460
2 94891 1 13460
2 94892 1 13470
2 94893 1 13470
2 94894 1 13472
2 94895 1 13472
2 94896 1 13472
2 94897 1 13472
2 94898 1 13473
2 94899 1 13473
2 94900 1 13473
2 94901 1 13480
2 94902 1 13480
2 94903 1 13480
2 94904 1 13480
2 94905 1 13480
2 94906 1 13480
2 94907 1 13487
2 94908 1 13487
2 94909 1 13503
2 94910 1 13503
2 94911 1 13504
2 94912 1 13504
2 94913 1 13504
2 94914 1 13504
2 94915 1 13513
2 94916 1 13513
2 94917 1 13514
2 94918 1 13514
2 94919 1 13526
2 94920 1 13526
2 94921 1 13526
2 94922 1 13536
2 94923 1 13536
2 94924 1 13549
2 94925 1 13549
2 94926 1 13550
2 94927 1 13550
2 94928 1 13550
2 94929 1 13550
2 94930 1 13550
2 94931 1 13552
2 94932 1 13552
2 94933 1 13552
2 94934 1 13552
2 94935 1 13552
2 94936 1 13553
2 94937 1 13553
2 94938 1 13555
2 94939 1 13555
2 94940 1 13555
2 94941 1 13613
2 94942 1 13613
2 94943 1 13614
2 94944 1 13614
2 94945 1 13614
2 94946 1 13615
2 94947 1 13615
2 94948 1 13616
2 94949 1 13616
2 94950 1 13617
2 94951 1 13617
2 94952 1 13617
2 94953 1 13618
2 94954 1 13618
2 94955 1 13632
2 94956 1 13632
2 94957 1 13646
2 94958 1 13646
2 94959 1 13647
2 94960 1 13647
2 94961 1 13665
2 94962 1 13665
2 94963 1 13665
2 94964 1 13666
2 94965 1 13666
2 94966 1 13666
2 94967 1 13667
2 94968 1 13667
2 94969 1 13674
2 94970 1 13674
2 94971 1 13674
2 94972 1 13674
2 94973 1 13674
2 94974 1 13686
2 94975 1 13686
2 94976 1 13686
2 94977 1 13686
2 94978 1 13687
2 94979 1 13687
2 94980 1 13698
2 94981 1 13698
2 94982 1 13698
2 94983 1 13698
2 94984 1 13699
2 94985 1 13699
2 94986 1 13700
2 94987 1 13700
2 94988 1 13701
2 94989 1 13701
2 94990 1 13709
2 94991 1 13709
2 94992 1 13709
2 94993 1 13709
2 94994 1 13723
2 94995 1 13723
2 94996 1 13725
2 94997 1 13725
2 94998 1 13725
2 94999 1 13725
2 95000 1 13725
2 95001 1 13725
2 95002 1 13726
2 95003 1 13726
2 95004 1 13736
2 95005 1 13736
2 95006 1 13737
2 95007 1 13737
2 95008 1 13756
2 95009 1 13756
2 95010 1 13757
2 95011 1 13757
2 95012 1 13757
2 95013 1 13760
2 95014 1 13760
2 95015 1 13764
2 95016 1 13764
2 95017 1 13785
2 95018 1 13785
2 95019 1 13786
2 95020 1 13786
2 95021 1 13787
2 95022 1 13787
2 95023 1 13794
2 95024 1 13794
2 95025 1 13794
2 95026 1 13794
2 95027 1 13796
2 95028 1 13796
2 95029 1 13804
2 95030 1 13804
2 95031 1 13804
2 95032 1 13804
2 95033 1 13805
2 95034 1 13805
2 95035 1 13822
2 95036 1 13822
2 95037 1 13822
2 95038 1 13822
2 95039 1 13823
2 95040 1 13823
2 95041 1 13844
2 95042 1 13844
2 95043 1 13852
2 95044 1 13852
2 95045 1 13852
2 95046 1 13852
2 95047 1 13852
2 95048 1 13852
2 95049 1 13852
2 95050 1 13853
2 95051 1 13853
2 95052 1 13853
2 95053 1 13854
2 95054 1 13854
2 95055 1 13874
2 95056 1 13874
2 95057 1 13876
2 95058 1 13876
2 95059 1 13877
2 95060 1 13877
2 95061 1 13877
2 95062 1 13892
2 95063 1 13892
2 95064 1 13895
2 95065 1 13895
2 95066 1 13895
2 95067 1 13895
2 95068 1 13895
2 95069 1 13895
2 95070 1 13895
2 95071 1 13895
2 95072 1 13909
2 95073 1 13909
2 95074 1 13949
2 95075 1 13949
2 95076 1 13958
2 95077 1 13958
2 95078 1 13961
2 95079 1 13961
2 95080 1 13983
2 95081 1 13983
2 95082 1 13985
2 95083 1 13985
2 95084 1 13985
2 95085 1 13985
2 95086 1 13985
2 95087 1 13985
2 95088 1 13986
2 95089 1 13986
2 95090 1 13986
2 95091 1 13988
2 95092 1 13988
2 95093 1 14001
2 95094 1 14001
2 95095 1 14001
2 95096 1 14002
2 95097 1 14002
2 95098 1 14002
2 95099 1 14015
2 95100 1 14015
2 95101 1 14015
2 95102 1 14015
2 95103 1 14016
2 95104 1 14016
2 95105 1 14027
2 95106 1 14027
2 95107 1 14027
2 95108 1 14034
2 95109 1 14034
2 95110 1 14036
2 95111 1 14036
2 95112 1 14036
2 95113 1 14036
2 95114 1 14036
2 95115 1 14037
2 95116 1 14037
2 95117 1 14037
2 95118 1 14061
2 95119 1 14061
2 95120 1 14068
2 95121 1 14068
2 95122 1 14068
2 95123 1 14068
2 95124 1 14069
2 95125 1 14069
2 95126 1 14069
2 95127 1 14069
2 95128 1 14069
2 95129 1 14087
2 95130 1 14087
2 95131 1 14100
2 95132 1 14100
2 95133 1 14100
2 95134 1 14100
2 95135 1 14100
2 95136 1 14100
2 95137 1 14100
2 95138 1 14100
2 95139 1 14108
2 95140 1 14108
2 95141 1 14113
2 95142 1 14113
2 95143 1 14131
2 95144 1 14131
2 95145 1 14131
2 95146 1 14132
2 95147 1 14132
2 95148 1 14132
2 95149 1 14150
2 95150 1 14150
2 95151 1 14150
2 95152 1 14150
2 95153 1 14150
2 95154 1 14161
2 95155 1 14161
2 95156 1 14161
2 95157 1 14164
2 95158 1 14164
2 95159 1 14175
2 95160 1 14175
2 95161 1 14175
2 95162 1 14175
2 95163 1 14176
2 95164 1 14176
2 95165 1 14176
2 95166 1 14176
2 95167 1 14176
2 95168 1 14176
2 95169 1 14176
2 95170 1 14176
2 95171 1 14184
2 95172 1 14184
2 95173 1 14185
2 95174 1 14185
2 95175 1 14199
2 95176 1 14199
2 95177 1 14199
2 95178 1 14200
2 95179 1 14200
2 95180 1 14202
2 95181 1 14202
2 95182 1 14219
2 95183 1 14219
2 95184 1 14220
2 95185 1 14220
2 95186 1 14236
2 95187 1 14236
2 95188 1 14236
2 95189 1 14236
2 95190 1 14240
2 95191 1 14240
2 95192 1 14240
2 95193 1 14240
2 95194 1 14240
2 95195 1 14241
2 95196 1 14241
2 95197 1 14249
2 95198 1 14249
2 95199 1 14249
2 95200 1 14250
2 95201 1 14250
2 95202 1 14251
2 95203 1 14251
2 95204 1 14251
2 95205 1 14251
2 95206 1 14272
2 95207 1 14272
2 95208 1 14272
2 95209 1 14289
2 95210 1 14289
2 95211 1 14289
2 95212 1 14289
2 95213 1 14289
2 95214 1 14289
2 95215 1 14289
2 95216 1 14289
2 95217 1 14289
2 95218 1 14297
2 95219 1 14297
2 95220 1 14298
2 95221 1 14298
2 95222 1 14298
2 95223 1 14309
2 95224 1 14309
2 95225 1 14309
2 95226 1 14310
2 95227 1 14310
2 95228 1 14321
2 95229 1 14321
2 95230 1 14321
2 95231 1 14321
2 95232 1 14321
2 95233 1 14321
2 95234 1 14321
2 95235 1 14321
2 95236 1 14335
2 95237 1 14335
2 95238 1 14336
2 95239 1 14336
2 95240 1 14344
2 95241 1 14344
2 95242 1 14355
2 95243 1 14355
2 95244 1 14359
2 95245 1 14359
2 95246 1 14401
2 95247 1 14401
2 95248 1 14401
2 95249 1 14410
2 95250 1 14410
2 95251 1 14428
2 95252 1 14428
2 95253 1 14429
2 95254 1 14429
2 95255 1 14429
2 95256 1 14429
2 95257 1 14429
2 95258 1 14429
2 95259 1 14440
2 95260 1 14440
2 95261 1 14441
2 95262 1 14441
2 95263 1 14441
2 95264 1 14441
2 95265 1 14441
2 95266 1 14441
2 95267 1 14441
2 95268 1 14441
2 95269 1 14441
2 95270 1 14441
2 95271 1 14441
2 95272 1 14441
2 95273 1 14442
2 95274 1 14442
2 95275 1 14442
2 95276 1 14442
2 95277 1 14442
2 95278 1 14442
2 95279 1 14443
2 95280 1 14443
2 95281 1 14443
2 95282 1 14443
2 95283 1 14443
2 95284 1 14443
2 95285 1 14443
2 95286 1 14451
2 95287 1 14451
2 95288 1 14451
2 95289 1 14451
2 95290 1 14451
2 95291 1 14451
2 95292 1 14451
2 95293 1 14451
2 95294 1 14451
2 95295 1 14451
2 95296 1 14452
2 95297 1 14452
2 95298 1 14453
2 95299 1 14453
2 95300 1 14453
2 95301 1 14463
2 95302 1 14463
2 95303 1 14463
2 95304 1 14463
2 95305 1 14464
2 95306 1 14464
2 95307 1 14464
2 95308 1 14464
2 95309 1 14464
2 95310 1 14464
2 95311 1 14464
2 95312 1 14464
2 95313 1 14464
2 95314 1 14464
2 95315 1 14464
2 95316 1 14464
2 95317 1 14464
2 95318 1 14464
2 95319 1 14464
2 95320 1 14464
2 95321 1 14464
2 95322 1 14464
2 95323 1 14477
2 95324 1 14477
2 95325 1 14485
2 95326 1 14485
2 95327 1 14499
2 95328 1 14499
2 95329 1 14499
2 95330 1 14499
2 95331 1 14504
2 95332 1 14504
2 95333 1 14504
2 95334 1 14504
2 95335 1 14504
2 95336 1 14504
2 95337 1 14504
2 95338 1 14504
2 95339 1 14504
2 95340 1 14504
2 95341 1 14504
2 95342 1 14504
2 95343 1 14504
2 95344 1 14504
2 95345 1 14504
2 95346 1 14504
2 95347 1 14506
2 95348 1 14506
2 95349 1 14506
2 95350 1 14506
2 95351 1 14506
2 95352 1 14506
2 95353 1 14506
2 95354 1 14508
2 95355 1 14508
2 95356 1 14508
2 95357 1 14516
2 95358 1 14516
2 95359 1 14516
2 95360 1 14517
2 95361 1 14517
2 95362 1 14519
2 95363 1 14519
2 95364 1 14522
2 95365 1 14522
2 95366 1 14522
2 95367 1 14522
2 95368 1 14522
2 95369 1 14522
2 95370 1 14522
2 95371 1 14522
2 95372 1 14522
2 95373 1 14523
2 95374 1 14523
2 95375 1 14523
2 95376 1 14523
2 95377 1 14523
2 95378 1 14524
2 95379 1 14524
2 95380 1 14525
2 95381 1 14525
2 95382 1 14526
2 95383 1 14526
2 95384 1 14526
2 95385 1 14526
2 95386 1 14526
2 95387 1 14526
2 95388 1 14526
2 95389 1 14535
2 95390 1 14535
2 95391 1 14536
2 95392 1 14536
2 95393 1 14536
2 95394 1 14551
2 95395 1 14551
2 95396 1 14553
2 95397 1 14553
2 95398 1 14554
2 95399 1 14554
2 95400 1 14558
2 95401 1 14558
2 95402 1 14559
2 95403 1 14559
2 95404 1 14565
2 95405 1 14565
2 95406 1 14571
2 95407 1 14571
2 95408 1 14573
2 95409 1 14573
2 95410 1 14584
2 95411 1 14584
2 95412 1 14584
2 95413 1 14592
2 95414 1 14592
2 95415 1 14592
2 95416 1 14592
2 95417 1 14592
2 95418 1 14593
2 95419 1 14593
2 95420 1 14593
2 95421 1 14593
2 95422 1 14593
2 95423 1 14593
2 95424 1 14596
2 95425 1 14596
2 95426 1 14597
2 95427 1 14597
2 95428 1 14597
2 95429 1 14597
2 95430 1 14598
2 95431 1 14598
2 95432 1 14599
2 95433 1 14599
2 95434 1 14602
2 95435 1 14602
2 95436 1 14610
2 95437 1 14610
2 95438 1 14611
2 95439 1 14611
2 95440 1 14629
2 95441 1 14629
2 95442 1 14637
2 95443 1 14637
2 95444 1 14637
2 95445 1 14637
2 95446 1 14637
2 95447 1 14639
2 95448 1 14639
2 95449 1 14641
2 95450 1 14641
2 95451 1 14644
2 95452 1 14644
2 95453 1 14653
2 95454 1 14653
2 95455 1 14678
2 95456 1 14678
2 95457 1 14678
2 95458 1 14678
2 95459 1 14678
2 95460 1 14690
2 95461 1 14690
2 95462 1 14702
2 95463 1 14702
2 95464 1 14702
2 95465 1 14703
2 95466 1 14703
2 95467 1 14704
2 95468 1 14704
2 95469 1 14705
2 95470 1 14705
2 95471 1 14705
2 95472 1 14730
2 95473 1 14730
2 95474 1 14730
2 95475 1 14730
2 95476 1 14730
2 95477 1 14730
2 95478 1 14732
2 95479 1 14732
2 95480 1 14741
2 95481 1 14741
2 95482 1 14741
2 95483 1 14741
2 95484 1 14741
2 95485 1 14750
2 95486 1 14750
2 95487 1 14750
2 95488 1 14750
2 95489 1 14750
2 95490 1 14750
2 95491 1 14767
2 95492 1 14767
2 95493 1 14767
2 95494 1 14767
2 95495 1 14767
2 95496 1 14779
2 95497 1 14779
2 95498 1 14787
2 95499 1 14787
2 95500 1 14789
2 95501 1 14789
2 95502 1 14790
2 95503 1 14790
2 95504 1 14790
2 95505 1 14790
2 95506 1 14790
2 95507 1 14790
2 95508 1 14790
2 95509 1 14790
2 95510 1 14790
2 95511 1 14792
2 95512 1 14792
2 95513 1 14792
2 95514 1 14792
2 95515 1 14792
2 95516 1 14794
2 95517 1 14794
2 95518 1 14794
2 95519 1 14794
2 95520 1 14798
2 95521 1 14798
2 95522 1 14798
2 95523 1 14798
2 95524 1 14798
2 95525 1 14798
2 95526 1 14798
2 95527 1 14798
2 95528 1 14799
2 95529 1 14799
2 95530 1 14799
2 95531 1 14800
2 95532 1 14800
2 95533 1 14801
2 95534 1 14801
2 95535 1 14816
2 95536 1 14816
2 95537 1 14823
2 95538 1 14823
2 95539 1 14828
2 95540 1 14828
2 95541 1 14828
2 95542 1 14828
2 95543 1 14829
2 95544 1 14829
2 95545 1 14836
2 95546 1 14836
2 95547 1 14836
2 95548 1 14836
2 95549 1 14836
2 95550 1 14846
2 95551 1 14846
2 95552 1 14846
2 95553 1 14856
2 95554 1 14856
2 95555 1 14882
2 95556 1 14882
2 95557 1 14882
2 95558 1 14882
2 95559 1 14894
2 95560 1 14894
2 95561 1 14913
2 95562 1 14913
2 95563 1 14913
2 95564 1 14913
2 95565 1 14913
2 95566 1 14914
2 95567 1 14914
2 95568 1 14915
2 95569 1 14915
2 95570 1 14916
2 95571 1 14916
2 95572 1 14916
2 95573 1 14925
2 95574 1 14925
2 95575 1 14925
2 95576 1 14925
2 95577 1 14925
2 95578 1 14926
2 95579 1 14926
2 95580 1 14927
2 95581 1 14927
2 95582 1 14927
2 95583 1 14927
2 95584 1 14932
2 95585 1 14932
2 95586 1 14932
2 95587 1 14932
2 95588 1 14932
2 95589 1 14932
2 95590 1 14935
2 95591 1 14935
2 95592 1 14935
2 95593 1 14935
2 95594 1 14936
2 95595 1 14936
2 95596 1 14944
2 95597 1 14944
2 95598 1 14945
2 95599 1 14945
2 95600 1 14950
2 95601 1 14950
2 95602 1 14950
2 95603 1 14951
2 95604 1 14951
2 95605 1 14952
2 95606 1 14952
2 95607 1 14952
2 95608 1 14970
2 95609 1 14970
2 95610 1 14971
2 95611 1 14971
2 95612 1 14979
2 95613 1 14979
2 95614 1 14979
2 95615 1 14979
2 95616 1 14980
2 95617 1 14980
2 95618 1 14980
2 95619 1 14980
2 95620 1 14980
2 95621 1 14980
2 95622 1 14980
2 95623 1 14980
2 95624 1 14980
2 95625 1 14990
2 95626 1 14990
2 95627 1 14991
2 95628 1 14991
2 95629 1 14991
2 95630 1 14992
2 95631 1 14992
2 95632 1 14992
2 95633 1 14993
2 95634 1 14993
2 95635 1 14993
2 95636 1 14993
2 95637 1 14993
2 95638 1 14993
2 95639 1 14993
2 95640 1 14993
2 95641 1 14993
2 95642 1 14993
2 95643 1 14993
2 95644 1 14993
2 95645 1 14993
2 95646 1 14993
2 95647 1 15009
2 95648 1 15009
2 95649 1 15009
2 95650 1 15009
2 95651 1 15009
2 95652 1 15009
2 95653 1 15010
2 95654 1 15010
2 95655 1 15025
2 95656 1 15025
2 95657 1 15025
2 95658 1 15025
2 95659 1 15044
2 95660 1 15044
2 95661 1 15044
2 95662 1 15044
2 95663 1 15046
2 95664 1 15046
2 95665 1 15053
2 95666 1 15053
2 95667 1 15053
2 95668 1 15067
2 95669 1 15067
2 95670 1 15067
2 95671 1 15067
2 95672 1 15067
2 95673 1 15067
2 95674 1 15069
2 95675 1 15069
2 95676 1 15069
2 95677 1 15069
2 95678 1 15085
2 95679 1 15085
2 95680 1 15085
2 95681 1 15085
2 95682 1 15099
2 95683 1 15099
2 95684 1 15104
2 95685 1 15104
2 95686 1 15104
2 95687 1 15104
2 95688 1 15112
2 95689 1 15112
2 95690 1 15112
2 95691 1 15112
2 95692 1 15112
2 95693 1 15113
2 95694 1 15113
2 95695 1 15120
2 95696 1 15120
2 95697 1 15120
2 95698 1 15123
2 95699 1 15123
2 95700 1 15123
2 95701 1 15123
2 95702 1 15123
2 95703 1 15124
2 95704 1 15124
2 95705 1 15124
2 95706 1 15124
2 95707 1 15124
2 95708 1 15124
2 95709 1 15124
2 95710 1 15141
2 95711 1 15141
2 95712 1 15150
2 95713 1 15150
2 95714 1 15150
2 95715 1 15162
2 95716 1 15162
2 95717 1 15165
2 95718 1 15165
2 95719 1 15165
2 95720 1 15165
2 95721 1 15165
2 95722 1 15165
2 95723 1 15165
2 95724 1 15165
2 95725 1 15165
2 95726 1 15166
2 95727 1 15166
2 95728 1 15166
2 95729 1 15175
2 95730 1 15175
2 95731 1 15175
2 95732 1 15175
2 95733 1 15176
2 95734 1 15176
2 95735 1 15176
2 95736 1 15176
2 95737 1 15184
2 95738 1 15184
2 95739 1 15184
2 95740 1 15184
2 95741 1 15184
2 95742 1 15184
2 95743 1 15184
2 95744 1 15184
2 95745 1 15184
2 95746 1 15185
2 95747 1 15185
2 95748 1 15195
2 95749 1 15195
2 95750 1 15195
2 95751 1 15210
2 95752 1 15210
2 95753 1 15210
2 95754 1 15212
2 95755 1 15212
2 95756 1 15213
2 95757 1 15213
2 95758 1 15214
2 95759 1 15214
2 95760 1 15214
2 95761 1 15215
2 95762 1 15215
2 95763 1 15215
2 95764 1 15225
2 95765 1 15225
2 95766 1 15227
2 95767 1 15227
2 95768 1 15236
2 95769 1 15236
2 95770 1 15251
2 95771 1 15251
2 95772 1 15251
2 95773 1 15251
2 95774 1 15251
2 95775 1 15269
2 95776 1 15269
2 95777 1 15269
2 95778 1 15269
2 95779 1 15269
2 95780 1 15269
2 95781 1 15269
2 95782 1 15269
2 95783 1 15270
2 95784 1 15270
2 95785 1 15270
2 95786 1 15270
2 95787 1 15270
2 95788 1 15287
2 95789 1 15287
2 95790 1 15287
2 95791 1 15288
2 95792 1 15288
2 95793 1 15288
2 95794 1 15289
2 95795 1 15289
2 95796 1 15296
2 95797 1 15296
2 95798 1 15296
2 95799 1 15296
2 95800 1 15296
2 95801 1 15296
2 95802 1 15297
2 95803 1 15297
2 95804 1 15297
2 95805 1 15305
2 95806 1 15305
2 95807 1 15326
2 95808 1 15326
2 95809 1 15339
2 95810 1 15339
2 95811 1 15343
2 95812 1 15343
2 95813 1 15344
2 95814 1 15344
2 95815 1 15346
2 95816 1 15346
2 95817 1 15346
2 95818 1 15346
2 95819 1 15346
2 95820 1 15361
2 95821 1 15361
2 95822 1 15362
2 95823 1 15362
2 95824 1 15362
2 95825 1 15362
2 95826 1 15362
2 95827 1 15362
2 95828 1 15365
2 95829 1 15365
2 95830 1 15375
2 95831 1 15375
2 95832 1 15382
2 95833 1 15382
2 95834 1 15382
2 95835 1 15414
2 95836 1 15414
2 95837 1 15429
2 95838 1 15429
2 95839 1 15444
2 95840 1 15444
2 95841 1 15444
2 95842 1 15448
2 95843 1 15448
2 95844 1 15448
2 95845 1 15448
2 95846 1 15449
2 95847 1 15449
2 95848 1 15450
2 95849 1 15450
2 95850 1 15450
2 95851 1 15458
2 95852 1 15458
2 95853 1 15459
2 95854 1 15459
2 95855 1 15460
2 95856 1 15460
2 95857 1 15476
2 95858 1 15476
2 95859 1 15476
2 95860 1 15481
2 95861 1 15481
2 95862 1 15500
2 95863 1 15500
2 95864 1 15500
2 95865 1 15504
2 95866 1 15504
2 95867 1 15515
2 95868 1 15515
2 95869 1 15516
2 95870 1 15516
2 95871 1 15516
2 95872 1 15538
2 95873 1 15538
2 95874 1 15546
2 95875 1 15546
2 95876 1 15546
2 95877 1 15546
2 95878 1 15569
2 95879 1 15569
2 95880 1 15571
2 95881 1 15571
2 95882 1 15571
2 95883 1 15572
2 95884 1 15572
2 95885 1 15634
2 95886 1 15634
2 95887 1 15634
2 95888 1 15634
2 95889 1 15634
2 95890 1 15634
2 95891 1 15634
2 95892 1 15660
2 95893 1 15660
2 95894 1 15660
2 95895 1 15661
2 95896 1 15661
2 95897 1 15663
2 95898 1 15663
2 95899 1 15669
2 95900 1 15669
2 95901 1 15669
2 95902 1 15687
2 95903 1 15687
2 95904 1 15687
2 95905 1 15694
2 95906 1 15694
2 95907 1 15694
2 95908 1 15701
2 95909 1 15701
2 95910 1 15701
2 95911 1 15701
2 95912 1 15702
2 95913 1 15702
2 95914 1 15702
2 95915 1 15722
2 95916 1 15722
2 95917 1 15722
2 95918 1 15724
2 95919 1 15724
2 95920 1 15729
2 95921 1 15729
2 95922 1 15737
2 95923 1 15737
2 95924 1 15750
2 95925 1 15750
2 95926 1 15754
2 95927 1 15754
2 95928 1 15774
2 95929 1 15774
2 95930 1 15777
2 95931 1 15777
2 95932 1 15789
2 95933 1 15789
2 95934 1 15789
2 95935 1 15789
2 95936 1 15789
2 95937 1 15791
2 95938 1 15791
2 95939 1 15795
2 95940 1 15795
2 95941 1 15795
2 95942 1 15795
2 95943 1 15795
2 95944 1 15796
2 95945 1 15796
2 95946 1 15796
2 95947 1 15796
2 95948 1 15797
2 95949 1 15797
2 95950 1 15805
2 95951 1 15805
2 95952 1 15813
2 95953 1 15813
2 95954 1 15816
2 95955 1 15816
2 95956 1 15816
2 95957 1 15816
2 95958 1 15824
2 95959 1 15824
2 95960 1 15827
2 95961 1 15827
2 95962 1 15827
2 95963 1 15834
2 95964 1 15834
2 95965 1 15834
2 95966 1 15856
2 95967 1 15856
2 95968 1 15856
2 95969 1 15880
2 95970 1 15880
2 95971 1 15880
2 95972 1 15880
2 95973 1 15880
2 95974 1 15880
2 95975 1 15880
2 95976 1 15881
2 95977 1 15881
2 95978 1 15890
2 95979 1 15890
2 95980 1 15898
2 95981 1 15898
2 95982 1 15968
2 95983 1 15968
2 95984 1 15968
2 95985 1 15983
2 95986 1 15983
2 95987 1 15984
2 95988 1 15984
2 95989 1 15984
2 95990 1 15999
2 95991 1 15999
2 95992 1 16015
2 95993 1 16015
2 95994 1 16034
2 95995 1 16034
2 95996 1 16035
2 95997 1 16035
2 95998 1 16035
2 95999 1 16035
2 96000 1 16035
2 96001 1 16035
2 96002 1 16035
2 96003 1 16035
2 96004 1 16035
2 96005 1 16035
2 96006 1 16035
2 96007 1 16035
2 96008 1 16037
2 96009 1 16037
2 96010 1 16044
2 96011 1 16044
2 96012 1 16047
2 96013 1 16047
2 96014 1 16057
2 96015 1 16057
2 96016 1 16057
2 96017 1 16070
2 96018 1 16070
2 96019 1 16070
2 96020 1 16070
2 96021 1 16070
2 96022 1 16070
2 96023 1 16070
2 96024 1 16078
2 96025 1 16078
2 96026 1 16078
2 96027 1 16078
2 96028 1 16078
2 96029 1 16078
2 96030 1 16091
2 96031 1 16091
2 96032 1 16091
2 96033 1 16091
2 96034 1 16091
2 96035 1 16091
2 96036 1 16091
2 96037 1 16100
2 96038 1 16100
2 96039 1 16100
2 96040 1 16100
2 96041 1 16111
2 96042 1 16111
2 96043 1 16111
2 96044 1 16112
2 96045 1 16112
2 96046 1 16119
2 96047 1 16119
2 96048 1 16119
2 96049 1 16119
2 96050 1 16119
2 96051 1 16130
2 96052 1 16130
2 96053 1 16144
2 96054 1 16144
2 96055 1 16159
2 96056 1 16159
2 96057 1 16159
2 96058 1 16159
2 96059 1 16160
2 96060 1 16160
2 96061 1 16184
2 96062 1 16184
2 96063 1 16197
2 96064 1 16197
2 96065 1 16197
2 96066 1 16198
2 96067 1 16198
2 96068 1 16209
2 96069 1 16209
2 96070 1 16209
2 96071 1 16209
2 96072 1 16211
2 96073 1 16211
2 96074 1 16211
2 96075 1 16211
2 96076 1 16211
2 96077 1 16211
2 96078 1 16227
2 96079 1 16227
2 96080 1 16227
2 96081 1 16227
2 96082 1 16227
2 96083 1 16227
2 96084 1 16227
2 96085 1 16227
2 96086 1 16227
2 96087 1 16228
2 96088 1 16228
2 96089 1 16228
2 96090 1 16228
2 96091 1 16230
2 96092 1 16230
2 96093 1 16238
2 96094 1 16238
2 96095 1 16238
2 96096 1 16245
2 96097 1 16245
2 96098 1 16246
2 96099 1 16246
2 96100 1 16246
2 96101 1 16246
2 96102 1 16246
2 96103 1 16246
2 96104 1 16246
2 96105 1 16246
2 96106 1 16246
2 96107 1 16246
2 96108 1 16246
2 96109 1 16246
2 96110 1 16246
2 96111 1 16246
2 96112 1 16255
2 96113 1 16255
2 96114 1 16273
2 96115 1 16273
2 96116 1 16273
2 96117 1 16274
2 96118 1 16274
2 96119 1 16274
2 96120 1 16277
2 96121 1 16277
2 96122 1 16278
2 96123 1 16278
2 96124 1 16278
2 96125 1 16278
2 96126 1 16279
2 96127 1 16279
2 96128 1 16280
2 96129 1 16280
2 96130 1 16297
2 96131 1 16297
2 96132 1 16297
2 96133 1 16297
2 96134 1 16297
2 96135 1 16298
2 96136 1 16298
2 96137 1 16315
2 96138 1 16315
2 96139 1 16320
2 96140 1 16320
2 96141 1 16343
2 96142 1 16343
2 96143 1 16353
2 96144 1 16353
2 96145 1 16353
2 96146 1 16365
2 96147 1 16365
2 96148 1 16373
2 96149 1 16373
2 96150 1 16374
2 96151 1 16374
2 96152 1 16410
2 96153 1 16410
2 96154 1 16410
2 96155 1 16410
2 96156 1 16411
2 96157 1 16411
2 96158 1 16419
2 96159 1 16419
2 96160 1 16420
2 96161 1 16420
2 96162 1 16420
2 96163 1 16428
2 96164 1 16428
2 96165 1 16429
2 96166 1 16429
2 96167 1 16429
2 96168 1 16451
2 96169 1 16451
2 96170 1 16452
2 96171 1 16452
2 96172 1 16452
2 96173 1 16452
2 96174 1 16453
2 96175 1 16453
2 96176 1 16453
2 96177 1 16453
2 96178 1 16466
2 96179 1 16466
2 96180 1 16504
2 96181 1 16504
2 96182 1 16504
2 96183 1 16516
2 96184 1 16516
2 96185 1 16516
2 96186 1 16529
2 96187 1 16529
2 96188 1 16529
2 96189 1 16530
2 96190 1 16530
2 96191 1 16545
2 96192 1 16545
2 96193 1 16545
2 96194 1 16553
2 96195 1 16553
2 96196 1 16554
2 96197 1 16554
2 96198 1 16554
2 96199 1 16554
2 96200 1 16554
2 96201 1 16554
2 96202 1 16583
2 96203 1 16583
2 96204 1 16583
2 96205 1 16607
2 96206 1 16607
2 96207 1 16607
2 96208 1 16638
2 96209 1 16638
2 96210 1 16638
2 96211 1 16640
2 96212 1 16640
2 96213 1 16645
2 96214 1 16645
2 96215 1 16657
2 96216 1 16657
2 96217 1 16658
2 96218 1 16658
2 96219 1 16658
2 96220 1 16677
2 96221 1 16677
2 96222 1 16688
2 96223 1 16688
2 96224 1 16688
2 96225 1 16688
2 96226 1 16688
2 96227 1 16688
2 96228 1 16711
2 96229 1 16711
2 96230 1 16712
2 96231 1 16712
2 96232 1 16721
2 96233 1 16721
2 96234 1 16733
2 96235 1 16733
2 96236 1 16733
2 96237 1 16733
2 96238 1 16781
2 96239 1 16781
2 96240 1 16783
2 96241 1 16783
2 96242 1 16783
2 96243 1 16783
2 96244 1 16783
2 96245 1 16784
2 96246 1 16784
2 96247 1 16789
2 96248 1 16789
2 96249 1 16791
2 96250 1 16791
2 96251 1 16791
2 96252 1 16791
2 96253 1 16791
2 96254 1 16791
2 96255 1 16791
2 96256 1 16791
2 96257 1 16806
2 96258 1 16806
2 96259 1 16806
2 96260 1 16806
2 96261 1 16807
2 96262 1 16807
2 96263 1 16807
2 96264 1 16807
2 96265 1 16807
2 96266 1 16807
2 96267 1 16807
2 96268 1 16809
2 96269 1 16809
2 96270 1 16809
2 96271 1 16809
2 96272 1 16809
2 96273 1 16809
2 96274 1 16809
2 96275 1 16809
2 96276 1 16809
2 96277 1 16809
2 96278 1 16809
2 96279 1 16809
2 96280 1 16809
2 96281 1 16809
2 96282 1 16809
2 96283 1 16810
2 96284 1 16810
2 96285 1 16810
2 96286 1 16810
2 96287 1 16810
2 96288 1 16810
2 96289 1 16811
2 96290 1 16811
2 96291 1 16812
2 96292 1 16812
2 96293 1 16812
2 96294 1 16812
2 96295 1 16815
2 96296 1 16815
2 96297 1 16815
2 96298 1 16815
2 96299 1 16815
2 96300 1 16815
2 96301 1 16815
2 96302 1 16815
2 96303 1 16815
2 96304 1 16815
2 96305 1 16816
2 96306 1 16816
2 96307 1 16824
2 96308 1 16824
2 96309 1 16825
2 96310 1 16825
2 96311 1 16825
2 96312 1 16825
2 96313 1 16825
2 96314 1 16825
2 96315 1 16825
2 96316 1 16825
2 96317 1 16825
2 96318 1 16835
2 96319 1 16835
2 96320 1 16851
2 96321 1 16851
2 96322 1 16854
2 96323 1 16854
2 96324 1 16854
2 96325 1 16854
2 96326 1 16854
2 96327 1 16854
2 96328 1 16854
2 96329 1 16854
2 96330 1 16854
2 96331 1 16854
2 96332 1 16854
2 96333 1 16854
2 96334 1 16854
2 96335 1 16855
2 96336 1 16855
2 96337 1 16855
2 96338 1 16855
2 96339 1 16855
2 96340 1 16855
2 96341 1 16856
2 96342 1 16856
2 96343 1 16856
2 96344 1 16856
2 96345 1 16857
2 96346 1 16857
2 96347 1 16875
2 96348 1 16875
2 96349 1 16875
2 96350 1 16875
2 96351 1 16875
2 96352 1 16879
2 96353 1 16879
2 96354 1 16879
2 96355 1 16881
2 96356 1 16881
2 96357 1 16881
2 96358 1 16883
2 96359 1 16883
2 96360 1 16884
2 96361 1 16884
2 96362 1 16884
2 96363 1 16884
2 96364 1 16884
2 96365 1 16884
2 96366 1 16884
2 96367 1 16884
2 96368 1 16884
2 96369 1 16884
2 96370 1 16884
2 96371 1 16884
2 96372 1 16884
2 96373 1 16884
2 96374 1 16884
2 96375 1 16884
2 96376 1 16884
2 96377 1 16884
2 96378 1 16884
2 96379 1 16884
2 96380 1 16884
2 96381 1 16884
2 96382 1 16887
2 96383 1 16887
2 96384 1 16887
2 96385 1 16887
2 96386 1 16887
2 96387 1 16887
2 96388 1 16891
2 96389 1 16891
2 96390 1 16891
2 96391 1 16892
2 96392 1 16892
2 96393 1 16893
2 96394 1 16893
2 96395 1 16893
2 96396 1 16893
2 96397 1 16893
2 96398 1 16893
2 96399 1 16893
2 96400 1 16893
2 96401 1 16893
2 96402 1 16893
2 96403 1 16893
2 96404 1 16899
2 96405 1 16899
2 96406 1 16900
2 96407 1 16900
2 96408 1 16900
2 96409 1 16900
2 96410 1 16900
2 96411 1 16900
2 96412 1 16900
2 96413 1 16900
2 96414 1 16900
2 96415 1 16902
2 96416 1 16902
2 96417 1 16908
2 96418 1 16908
2 96419 1 16925
2 96420 1 16925
2 96421 1 16925
2 96422 1 16925
2 96423 1 16925
2 96424 1 16925
2 96425 1 16925
2 96426 1 16925
2 96427 1 16925
2 96428 1 16925
2 96429 1 16925
2 96430 1 16925
2 96431 1 16925
2 96432 1 16925
2 96433 1 16925
2 96434 1 16925
2 96435 1 16925
2 96436 1 16925
2 96437 1 16925
2 96438 1 16925
2 96439 1 16925
2 96440 1 16925
2 96441 1 16925
2 96442 1 16927
2 96443 1 16927
2 96444 1 16927
2 96445 1 16927
2 96446 1 16927
2 96447 1 16927
2 96448 1 16927
2 96449 1 16928
2 96450 1 16928
2 96451 1 16928
2 96452 1 16928
2 96453 1 16928
2 96454 1 16929
2 96455 1 16929
2 96456 1 16929
2 96457 1 16929
2 96458 1 16929
2 96459 1 16931
2 96460 1 16931
2 96461 1 16931
2 96462 1 16931
2 96463 1 16931
2 96464 1 16932
2 96465 1 16932
2 96466 1 16934
2 96467 1 16934
2 96468 1 16943
2 96469 1 16943
2 96470 1 16944
2 96471 1 16944
2 96472 1 16945
2 96473 1 16945
2 96474 1 16946
2 96475 1 16946
2 96476 1 16948
2 96477 1 16948
2 96478 1 16962
2 96479 1 16962
2 96480 1 16962
2 96481 1 16977
2 96482 1 16977
2 96483 1 16977
2 96484 1 16977
2 96485 1 16977
2 96486 1 16984
2 96487 1 16984
2 96488 1 16984
2 96489 1 16984
2 96490 1 16991
2 96491 1 16991
2 96492 1 16996
2 96493 1 16996
2 96494 1 16997
2 96495 1 16997
2 96496 1 17024
2 96497 1 17024
2 96498 1 17038
2 96499 1 17038
2 96500 1 17038
2 96501 1 17038
2 96502 1 17039
2 96503 1 17039
2 96504 1 17039
2 96505 1 17039
2 96506 1 17041
2 96507 1 17041
2 96508 1 17042
2 96509 1 17042
2 96510 1 17042
2 96511 1 17042
2 96512 1 17042
2 96513 1 17042
2 96514 1 17042
2 96515 1 17042
2 96516 1 17042
2 96517 1 17054
2 96518 1 17054
2 96519 1 17054
2 96520 1 17054
2 96521 1 17054
2 96522 1 17064
2 96523 1 17064
2 96524 1 17064
2 96525 1 17064
2 96526 1 17064
2 96527 1 17064
2 96528 1 17064
2 96529 1 17064
2 96530 1 17064
2 96531 1 17064
2 96532 1 17066
2 96533 1 17066
2 96534 1 17079
2 96535 1 17079
2 96536 1 17087
2 96537 1 17087
2 96538 1 17096
2 96539 1 17096
2 96540 1 17096
2 96541 1 17096
2 96542 1 17105
2 96543 1 17105
2 96544 1 17108
2 96545 1 17108
2 96546 1 17117
2 96547 1 17117
2 96548 1 17117
2 96549 1 17117
2 96550 1 17117
2 96551 1 17117
2 96552 1 17131
2 96553 1 17131
2 96554 1 17131
2 96555 1 17131
2 96556 1 17132
2 96557 1 17132
2 96558 1 17132
2 96559 1 17133
2 96560 1 17133
2 96561 1 17133
2 96562 1 17133
2 96563 1 17133
2 96564 1 17133
2 96565 1 17133
2 96566 1 17133
2 96567 1 17136
2 96568 1 17136
2 96569 1 17136
2 96570 1 17136
2 96571 1 17136
2 96572 1 17136
2 96573 1 17136
2 96574 1 17136
2 96575 1 17136
2 96576 1 17136
2 96577 1 17137
2 96578 1 17137
2 96579 1 17138
2 96580 1 17138
2 96581 1 17166
2 96582 1 17166
2 96583 1 17166
2 96584 1 17166
2 96585 1 17166
2 96586 1 17174
2 96587 1 17174
2 96588 1 17175
2 96589 1 17175
2 96590 1 17175
2 96591 1 17183
2 96592 1 17183
2 96593 1 17183
2 96594 1 17184
2 96595 1 17184
2 96596 1 17184
2 96597 1 17192
2 96598 1 17192
2 96599 1 17193
2 96600 1 17193
2 96601 1 17194
2 96602 1 17194
2 96603 1 17208
2 96604 1 17208
2 96605 1 17208
2 96606 1 17211
2 96607 1 17211
2 96608 1 17215
2 96609 1 17215
2 96610 1 17223
2 96611 1 17223
2 96612 1 17223
2 96613 1 17223
2 96614 1 17223
2 96615 1 17223
2 96616 1 17223
2 96617 1 17223
2 96618 1 17223
2 96619 1 17223
2 96620 1 17223
2 96621 1 17223
2 96622 1 17224
2 96623 1 17224
2 96624 1 17226
2 96625 1 17226
2 96626 1 17226
2 96627 1 17233
2 96628 1 17233
2 96629 1 17234
2 96630 1 17234
2 96631 1 17244
2 96632 1 17244
2 96633 1 17245
2 96634 1 17245
2 96635 1 17246
2 96636 1 17246
2 96637 1 17256
2 96638 1 17256
2 96639 1 17256
2 96640 1 17256
2 96641 1 17284
2 96642 1 17284
2 96643 1 17286
2 96644 1 17286
2 96645 1 17286
2 96646 1 17286
2 96647 1 17286
2 96648 1 17286
2 96649 1 17286
2 96650 1 17286
2 96651 1 17286
2 96652 1 17286
2 96653 1 17287
2 96654 1 17287
2 96655 1 17288
2 96656 1 17288
2 96657 1 17288
2 96658 1 17288
2 96659 1 17289
2 96660 1 17289
2 96661 1 17289
2 96662 1 17291
2 96663 1 17291
2 96664 1 17298
2 96665 1 17298
2 96666 1 17315
2 96667 1 17315
2 96668 1 17315
2 96669 1 17318
2 96670 1 17318
2 96671 1 17318
2 96672 1 17318
2 96673 1 17318
2 96674 1 17319
2 96675 1 17319
2 96676 1 17319
2 96677 1 17320
2 96678 1 17320
2 96679 1 17320
2 96680 1 17325
2 96681 1 17325
2 96682 1 17325
2 96683 1 17326
2 96684 1 17326
2 96685 1 17327
2 96686 1 17327
2 96687 1 17338
2 96688 1 17338
2 96689 1 17340
2 96690 1 17340
2 96691 1 17359
2 96692 1 17359
2 96693 1 17359
2 96694 1 17361
2 96695 1 17361
2 96696 1 17368
2 96697 1 17368
2 96698 1 17368
2 96699 1 17368
2 96700 1 17368
2 96701 1 17368
2 96702 1 17369
2 96703 1 17369
2 96704 1 17369
2 96705 1 17373
2 96706 1 17373
2 96707 1 17373
2 96708 1 17376
2 96709 1 17376
2 96710 1 17380
2 96711 1 17380
2 96712 1 17381
2 96713 1 17381
2 96714 1 17384
2 96715 1 17384
2 96716 1 17393
2 96717 1 17393
2 96718 1 17393
2 96719 1 17442
2 96720 1 17442
2 96721 1 17447
2 96722 1 17447
2 96723 1 17448
2 96724 1 17448
2 96725 1 17448
2 96726 1 17448
2 96727 1 17448
2 96728 1 17448
2 96729 1 17448
2 96730 1 17448
2 96731 1 17448
2 96732 1 17457
2 96733 1 17457
2 96734 1 17457
2 96735 1 17457
2 96736 1 17457
2 96737 1 17457
2 96738 1 17457
2 96739 1 17457
2 96740 1 17457
2 96741 1 17457
2 96742 1 17457
2 96743 1 17457
2 96744 1 17457
2 96745 1 17457
2 96746 1 17457
2 96747 1 17457
2 96748 1 17457
2 96749 1 17457
2 96750 1 17457
2 96751 1 17457
2 96752 1 17457
2 96753 1 17457
2 96754 1 17457
2 96755 1 17457
2 96756 1 17457
2 96757 1 17457
2 96758 1 17457
2 96759 1 17457
2 96760 1 17457
2 96761 1 17457
2 96762 1 17457
2 96763 1 17457
2 96764 1 17457
2 96765 1 17457
2 96766 1 17457
2 96767 1 17457
2 96768 1 17457
2 96769 1 17457
2 96770 1 17457
2 96771 1 17457
2 96772 1 17457
2 96773 1 17457
2 96774 1 17457
2 96775 1 17457
2 96776 1 17457
2 96777 1 17457
2 96778 1 17457
2 96779 1 17457
2 96780 1 17457
2 96781 1 17457
2 96782 1 17457
2 96783 1 17457
2 96784 1 17457
2 96785 1 17458
2 96786 1 17458
2 96787 1 17459
2 96788 1 17459
2 96789 1 17459
2 96790 1 17459
2 96791 1 17459
2 96792 1 17460
2 96793 1 17460
2 96794 1 17460
2 96795 1 17475
2 96796 1 17475
2 96797 1 17475
2 96798 1 17476
2 96799 1 17476
2 96800 1 17476
2 96801 1 17476
2 96802 1 17476
2 96803 1 17476
2 96804 1 17476
2 96805 1 17476
2 96806 1 17478
2 96807 1 17478
2 96808 1 17478
2 96809 1 17480
2 96810 1 17480
2 96811 1 17480
2 96812 1 17481
2 96813 1 17481
2 96814 1 17482
2 96815 1 17482
2 96816 1 17484
2 96817 1 17484
2 96818 1 17507
2 96819 1 17507
2 96820 1 17529
2 96821 1 17529
2 96822 1 17529
2 96823 1 17530
2 96824 1 17530
2 96825 1 17530
2 96826 1 17537
2 96827 1 17537
2 96828 1 17537
2 96829 1 17548
2 96830 1 17548
2 96831 1 17548
2 96832 1 17551
2 96833 1 17551
2 96834 1 17583
2 96835 1 17583
2 96836 1 17583
2 96837 1 17583
2 96838 1 17584
2 96839 1 17584
2 96840 1 17585
2 96841 1 17585
2 96842 1 17585
2 96843 1 17595
2 96844 1 17595
2 96845 1 17595
2 96846 1 17606
2 96847 1 17606
2 96848 1 17606
2 96849 1 17608
2 96850 1 17608
2 96851 1 17642
2 96852 1 17642
2 96853 1 17645
2 96854 1 17645
2 96855 1 17658
2 96856 1 17658
2 96857 1 17666
2 96858 1 17666
2 96859 1 17666
2 96860 1 17667
2 96861 1 17667
2 96862 1 17685
2 96863 1 17685
2 96864 1 17685
2 96865 1 17685
2 96866 1 17685
2 96867 1 17685
2 96868 1 17685
2 96869 1 17685
2 96870 1 17686
2 96871 1 17686
2 96872 1 17691
2 96873 1 17691
2 96874 1 17694
2 96875 1 17694
2 96876 1 17695
2 96877 1 17695
2 96878 1 17702
2 96879 1 17702
2 96880 1 17719
2 96881 1 17719
2 96882 1 17720
2 96883 1 17720
2 96884 1 17732
2 96885 1 17732
2 96886 1 17734
2 96887 1 17734
2 96888 1 17747
2 96889 1 17747
2 96890 1 17748
2 96891 1 17748
2 96892 1 17750
2 96893 1 17750
2 96894 1 17750
2 96895 1 17755
2 96896 1 17755
2 96897 1 17755
2 96898 1 17755
2 96899 1 17756
2 96900 1 17756
2 96901 1 17756
2 96902 1 17757
2 96903 1 17757
2 96904 1 17764
2 96905 1 17764
2 96906 1 17773
2 96907 1 17773
2 96908 1 17794
2 96909 1 17794
2 96910 1 17808
2 96911 1 17808
2 96912 1 17865
2 96913 1 17865
2 96914 1 17879
2 96915 1 17879
2 96916 1 17879
2 96917 1 17879
2 96918 1 17879
2 96919 1 17879
2 96920 1 17879
2 96921 1 17879
2 96922 1 17879
2 96923 1 17879
2 96924 1 17879
2 96925 1 17879
2 96926 1 17879
2 96927 1 17879
2 96928 1 17879
2 96929 1 17879
2 96930 1 17879
2 96931 1 17879
2 96932 1 17879
2 96933 1 17879
2 96934 1 17879
2 96935 1 17879
2 96936 1 17879
2 96937 1 17879
2 96938 1 17879
2 96939 1 17879
2 96940 1 17879
2 96941 1 17879
2 96942 1 17879
2 96943 1 17879
2 96944 1 17879
2 96945 1 17879
2 96946 1 17879
2 96947 1 17879
2 96948 1 17879
2 96949 1 17879
2 96950 1 17879
2 96951 1 17880
2 96952 1 17880
2 96953 1 17881
2 96954 1 17881
2 96955 1 17881
2 96956 1 17881
2 96957 1 17881
2 96958 1 17881
2 96959 1 17881
2 96960 1 17881
2 96961 1 17881
2 96962 1 17881
2 96963 1 17881
2 96964 1 17881
2 96965 1 17881
2 96966 1 17881
2 96967 1 17881
2 96968 1 17881
2 96969 1 17881
2 96970 1 17881
2 96971 1 17881
2 96972 1 17881
2 96973 1 17881
2 96974 1 17881
2 96975 1 17881
2 96976 1 17881
2 96977 1 17881
2 96978 1 17881
2 96979 1 17881
2 96980 1 17881
2 96981 1 17881
2 96982 1 17881
2 96983 1 17881
2 96984 1 17881
2 96985 1 17881
2 96986 1 17881
2 96987 1 17881
2 96988 1 17881
2 96989 1 17881
2 96990 1 17881
2 96991 1 17882
2 96992 1 17882
2 96993 1 17883
2 96994 1 17883
2 96995 1 17884
2 96996 1 17884
2 96997 1 17884
2 96998 1 17884
2 96999 1 17884
2 97000 1 17884
2 97001 1 17884
2 97002 1 17884
2 97003 1 17884
2 97004 1 17886
2 97005 1 17886
2 97006 1 17886
2 97007 1 17887
2 97008 1 17887
2 97009 1 17887
2 97010 1 17888
2 97011 1 17888
2 97012 1 17913
2 97013 1 17913
2 97014 1 17913
2 97015 1 17913
2 97016 1 17913
2 97017 1 17913
2 97018 1 17913
2 97019 1 17916
2 97020 1 17916
2 97021 1 17917
2 97022 1 17917
2 97023 1 17917
2 97024 1 17917
2 97025 1 17917
2 97026 1 17917
2 97027 1 17917
2 97028 1 17917
2 97029 1 17917
2 97030 1 17917
2 97031 1 17917
2 97032 1 17917
2 97033 1 17917
2 97034 1 17917
2 97035 1 17917
2 97036 1 17917
2 97037 1 17917
2 97038 1 17917
2 97039 1 17917
2 97040 1 17917
2 97041 1 17917
2 97042 1 17917
2 97043 1 17917
2 97044 1 17917
2 97045 1 17917
2 97046 1 17917
2 97047 1 17917
2 97048 1 17917
2 97049 1 17917
2 97050 1 17917
2 97051 1 17917
2 97052 1 17917
2 97053 1 17917
2 97054 1 17917
2 97055 1 17917
2 97056 1 17917
2 97057 1 17917
2 97058 1 17917
2 97059 1 17917
2 97060 1 17917
2 97061 1 17917
2 97062 1 17917
2 97063 1 17917
2 97064 1 17917
2 97065 1 17917
2 97066 1 17917
2 97067 1 17917
2 97068 1 17917
2 97069 1 17917
2 97070 1 17919
2 97071 1 17919
2 97072 1 17919
2 97073 1 17919
2 97074 1 17919
2 97075 1 17919
2 97076 1 17919
2 97077 1 17919
2 97078 1 17920
2 97079 1 17920
2 97080 1 17933
2 97081 1 17933
2 97082 1 17933
2 97083 1 17933
2 97084 1 17933
2 97085 1 17933
2 97086 1 17933
2 97087 1 17933
2 97088 1 17933
2 97089 1 17933
2 97090 1 17933
2 97091 1 17968
2 97092 1 17968
2 97093 1 17968
2 97094 1 17968
2 97095 1 17972
2 97096 1 17972
2 97097 1 17972
2 97098 1 17990
2 97099 1 17990
2 97100 1 17990
2 97101 1 17990
2 97102 1 17990
2 97103 1 17990
2 97104 1 17990
2 97105 1 17990
2 97106 1 17990
2 97107 1 17990
2 97108 1 17990
2 97109 1 17990
2 97110 1 17998
2 97111 1 17998
2 97112 1 17998
2 97113 1 17999
2 97114 1 17999
2 97115 1 18002
2 97116 1 18002
2 97117 1 18002
2 97118 1 18002
2 97119 1 18002
2 97120 1 18002
2 97121 1 18002
2 97122 1 18002
2 97123 1 18002
2 97124 1 18002
2 97125 1 18002
2 97126 1 18002
2 97127 1 18002
2 97128 1 18002
2 97129 1 18002
2 97130 1 18002
2 97131 1 18002
2 97132 1 18002
2 97133 1 18002
2 97134 1 18002
2 97135 1 18002
2 97136 1 18002
2 97137 1 18002
2 97138 1 18003
2 97139 1 18003
2 97140 1 18004
2 97141 1 18004
2 97142 1 18016
2 97143 1 18016
2 97144 1 18023
2 97145 1 18023
2 97146 1 18023
2 97147 1 18023
2 97148 1 18025
2 97149 1 18025
2 97150 1 18025
2 97151 1 18025
2 97152 1 18025
2 97153 1 18025
2 97154 1 18026
2 97155 1 18026
2 97156 1 18033
2 97157 1 18033
2 97158 1 18036
2 97159 1 18036
2 97160 1 18036
2 97161 1 18044
2 97162 1 18044
2 97163 1 18044
2 97164 1 18044
2 97165 1 18044
2 97166 1 18044
2 97167 1 18044
2 97168 1 18044
2 97169 1 18060
2 97170 1 18060
2 97171 1 18060
2 97172 1 18060
2 97173 1 18061
2 97174 1 18061
2 97175 1 18061
2 97176 1 18062
2 97177 1 18062
2 97178 1 18062
2 97179 1 18076
2 97180 1 18076
2 97181 1 18076
2 97182 1 18077
2 97183 1 18077
2 97184 1 18077
2 97185 1 18077
2 97186 1 18081
2 97187 1 18081
2 97188 1 18084
2 97189 1 18084
2 97190 1 18086
2 97191 1 18086
2 97192 1 18093
2 97193 1 18093
2 97194 1 18107
2 97195 1 18107
2 97196 1 18115
2 97197 1 18115
2 97198 1 18115
2 97199 1 18115
2 97200 1 18115
2 97201 1 18123
2 97202 1 18123
2 97203 1 18123
2 97204 1 18123
2 97205 1 18123
2 97206 1 18123
2 97207 1 18123
2 97208 1 18123
2 97209 1 18123
2 97210 1 18123
2 97211 1 18123
2 97212 1 18123
2 97213 1 18127
2 97214 1 18127
2 97215 1 18127
2 97216 1 18127
2 97217 1 18128
2 97218 1 18128
2 97219 1 18128
2 97220 1 18128
2 97221 1 18133
2 97222 1 18133
2 97223 1 18136
2 97224 1 18136
2 97225 1 18136
2 97226 1 18136
2 97227 1 18148
2 97228 1 18148
2 97229 1 18148
2 97230 1 18148
2 97231 1 18165
2 97232 1 18165
2 97233 1 18165
2 97234 1 18165
2 97235 1 18165
2 97236 1 18166
2 97237 1 18166
2 97238 1 18166
2 97239 1 18166
2 97240 1 18167
2 97241 1 18167
2 97242 1 18176
2 97243 1 18176
2 97244 1 18196
2 97245 1 18196
2 97246 1 18197
2 97247 1 18197
2 97248 1 18197
2 97249 1 18197
2 97250 1 18201
2 97251 1 18201
2 97252 1 18201
2 97253 1 18202
2 97254 1 18202
2 97255 1 18203
2 97256 1 18203
2 97257 1 18203
2 97258 1 18203
2 97259 1 18203
2 97260 1 18212
2 97261 1 18212
2 97262 1 18225
2 97263 1 18225
2 97264 1 18225
2 97265 1 18225
2 97266 1 18225
2 97267 1 18225
2 97268 1 18225
2 97269 1 18225
2 97270 1 18226
2 97271 1 18226
2 97272 1 18227
2 97273 1 18227
2 97274 1 18230
2 97275 1 18230
2 97276 1 18237
2 97277 1 18237
2 97278 1 18237
2 97279 1 18237
2 97280 1 18237
2 97281 1 18237
2 97282 1 18237
2 97283 1 18237
2 97284 1 18237
2 97285 1 18237
2 97286 1 18239
2 97287 1 18239
2 97288 1 18239
2 97289 1 18239
2 97290 1 18241
2 97291 1 18241
2 97292 1 18242
2 97293 1 18242
2 97294 1 18250
2 97295 1 18250
2 97296 1 18250
2 97297 1 18250
2 97298 1 18250
2 97299 1 18261
2 97300 1 18261
2 97301 1 18261
2 97302 1 18270
2 97303 1 18270
2 97304 1 18282
2 97305 1 18282
2 97306 1 18291
2 97307 1 18291
2 97308 1 18291
2 97309 1 18300
2 97310 1 18300
2 97311 1 18309
2 97312 1 18309
2 97313 1 18309
2 97314 1 18309
2 97315 1 18309
2 97316 1 18311
2 97317 1 18311
2 97318 1 18312
2 97319 1 18312
2 97320 1 18312
2 97321 1 18358
2 97322 1 18358
2 97323 1 18358
2 97324 1 18358
2 97325 1 18359
2 97326 1 18359
2 97327 1 18367
2 97328 1 18367
2 97329 1 18367
2 97330 1 18367
2 97331 1 18367
2 97332 1 18367
2 97333 1 18375
2 97334 1 18375
2 97335 1 18384
2 97336 1 18384
2 97337 1 18384
2 97338 1 18384
2 97339 1 18384
2 97340 1 18384
2 97341 1 18385
2 97342 1 18385
2 97343 1 18385
2 97344 1 18385
2 97345 1 18385
2 97346 1 18393
2 97347 1 18393
2 97348 1 18416
2 97349 1 18416
2 97350 1 18422
2 97351 1 18422
2 97352 1 18430
2 97353 1 18430
2 97354 1 18455
2 97355 1 18455
2 97356 1 18475
2 97357 1 18475
2 97358 1 18475
2 97359 1 18475
2 97360 1 18475
2 97361 1 18475
2 97362 1 18475
2 97363 1 18475
2 97364 1 18475
2 97365 1 18475
2 97366 1 18476
2 97367 1 18476
2 97368 1 18476
2 97369 1 18476
2 97370 1 18476
2 97371 1 18476
2 97372 1 18477
2 97373 1 18477
2 97374 1 18478
2 97375 1 18478
2 97376 1 18478
2 97377 1 18478
2 97378 1 18478
2 97379 1 18478
2 97380 1 18478
2 97381 1 18478
2 97382 1 18478
2 97383 1 18478
2 97384 1 18478
2 97385 1 18478
2 97386 1 18478
2 97387 1 18478
2 97388 1 18478
2 97389 1 18478
2 97390 1 18478
2 97391 1 18478
2 97392 1 18478
2 97393 1 18478
2 97394 1 18478
2 97395 1 18478
2 97396 1 18478
2 97397 1 18478
2 97398 1 18478
2 97399 1 18478
2 97400 1 18478
2 97401 1 18478
2 97402 1 18478
2 97403 1 18478
2 97404 1 18478
2 97405 1 18478
2 97406 1 18478
2 97407 1 18478
2 97408 1 18478
2 97409 1 18478
2 97410 1 18478
2 97411 1 18478
2 97412 1 18478
2 97413 1 18478
2 97414 1 18478
2 97415 1 18478
2 97416 1 18478
2 97417 1 18478
2 97418 1 18478
2 97419 1 18478
2 97420 1 18478
2 97421 1 18478
2 97422 1 18478
2 97423 1 18478
2 97424 1 18478
2 97425 1 18478
2 97426 1 18478
2 97427 1 18478
2 97428 1 18478
2 97429 1 18478
2 97430 1 18478
2 97431 1 18478
2 97432 1 18481
2 97433 1 18481
2 97434 1 18488
2 97435 1 18488
2 97436 1 18489
2 97437 1 18489
2 97438 1 18489
2 97439 1 18489
2 97440 1 18489
2 97441 1 18489
2 97442 1 18489
2 97443 1 18489
2 97444 1 18489
2 97445 1 18489
2 97446 1 18489
2 97447 1 18490
2 97448 1 18490
2 97449 1 18491
2 97450 1 18491
2 97451 1 18498
2 97452 1 18498
2 97453 1 18499
2 97454 1 18499
2 97455 1 18507
2 97456 1 18507
2 97457 1 18508
2 97458 1 18508
2 97459 1 18509
2 97460 1 18509
2 97461 1 18525
2 97462 1 18525
2 97463 1 18525
2 97464 1 18525
2 97465 1 18525
2 97466 1 18525
2 97467 1 18525
2 97468 1 18533
2 97469 1 18533
2 97470 1 18536
2 97471 1 18536
2 97472 1 18536
2 97473 1 18536
2 97474 1 18536
2 97475 1 18536
2 97476 1 18536
2 97477 1 18536
2 97478 1 18536
2 97479 1 18536
2 97480 1 18536
2 97481 1 18536
2 97482 1 18536
2 97483 1 18536
2 97484 1 18536
2 97485 1 18536
2 97486 1 18536
2 97487 1 18537
2 97488 1 18537
2 97489 1 18537
2 97490 1 18537
2 97491 1 18537
2 97492 1 18538
2 97493 1 18538
2 97494 1 18538
2 97495 1 18538
2 97496 1 18538
2 97497 1 18546
2 97498 1 18546
2 97499 1 18547
2 97500 1 18547
2 97501 1 18547
2 97502 1 18547
2 97503 1 18551
2 97504 1 18551
2 97505 1 18551
2 97506 1 18564
2 97507 1 18564
2 97508 1 18565
2 97509 1 18565
2 97510 1 18565
2 97511 1 18566
2 97512 1 18566
2 97513 1 18567
2 97514 1 18567
2 97515 1 18567
2 97516 1 18575
2 97517 1 18575
2 97518 1 18575
2 97519 1 18575
2 97520 1 18585
2 97521 1 18585
2 97522 1 18589
2 97523 1 18589
2 97524 1 18597
2 97525 1 18597
2 97526 1 18598
2 97527 1 18598
2 97528 1 18618
2 97529 1 18618
2 97530 1 18618
2 97531 1 18618
2 97532 1 18618
2 97533 1 18618
2 97534 1 18618
2 97535 1 18619
2 97536 1 18619
2 97537 1 18621
2 97538 1 18621
2 97539 1 18622
2 97540 1 18622
2 97541 1 18622
2 97542 1 18622
2 97543 1 18622
2 97544 1 18622
2 97545 1 18622
2 97546 1 18623
2 97547 1 18623
2 97548 1 18623
2 97549 1 18623
2 97550 1 18625
2 97551 1 18625
2 97552 1 18626
2 97553 1 18626
2 97554 1 18626
2 97555 1 18626
2 97556 1 18626
2 97557 1 18626
2 97558 1 18626
2 97559 1 18628
2 97560 1 18628
2 97561 1 18628
2 97562 1 18628
2 97563 1 18628
2 97564 1 18628
2 97565 1 18648
2 97566 1 18648
2 97567 1 18648
2 97568 1 18648
2 97569 1 18648
2 97570 1 18650
2 97571 1 18650
2 97572 1 18653
2 97573 1 18653
2 97574 1 18660
2 97575 1 18660
2 97576 1 18670
2 97577 1 18670
2 97578 1 18670
2 97579 1 18679
2 97580 1 18679
2 97581 1 18691
2 97582 1 18691
2 97583 1 18692
2 97584 1 18692
2 97585 1 18695
2 97586 1 18695
2 97587 1 18695
2 97588 1 18695
2 97589 1 18695
2 97590 1 18695
2 97591 1 18695
2 97592 1 18695
2 97593 1 18696
2 97594 1 18696
2 97595 1 18696
2 97596 1 18703
2 97597 1 18703
2 97598 1 18703
2 97599 1 18715
2 97600 1 18715
2 97601 1 18715
2 97602 1 18715
2 97603 1 18715
2 97604 1 18716
2 97605 1 18716
2 97606 1 18719
2 97607 1 18719
2 97608 1 18720
2 97609 1 18720
2 97610 1 18720
2 97611 1 18721
2 97612 1 18721
2 97613 1 18730
2 97614 1 18730
2 97615 1 18734
2 97616 1 18734
2 97617 1 18734
2 97618 1 18734
2 97619 1 18735
2 97620 1 18735
2 97621 1 18741
2 97622 1 18741
2 97623 1 18756
2 97624 1 18756
2 97625 1 18756
2 97626 1 18756
2 97627 1 18756
2 97628 1 18756
2 97629 1 18758
2 97630 1 18758
2 97631 1 18759
2 97632 1 18759
2 97633 1 18810
2 97634 1 18810
2 97635 1 18811
2 97636 1 18811
2 97637 1 18812
2 97638 1 18812
2 97639 1 18824
2 97640 1 18824
2 97641 1 18832
2 97642 1 18832
2 97643 1 18835
2 97644 1 18835
2 97645 1 18843
2 97646 1 18843
2 97647 1 18851
2 97648 1 18851
2 97649 1 18851
2 97650 1 18864
2 97651 1 18864
2 97652 1 18865
2 97653 1 18865
2 97654 1 18866
2 97655 1 18866
2 97656 1 18867
2 97657 1 18867
2 97658 1 18869
2 97659 1 18869
2 97660 1 18873
2 97661 1 18873
2 97662 1 18873
2 97663 1 18873
2 97664 1 18873
2 97665 1 18881
2 97666 1 18881
2 97667 1 18893
2 97668 1 18893
2 97669 1 18893
2 97670 1 18893
2 97671 1 18893
2 97672 1 18894
2 97673 1 18894
2 97674 1 18897
2 97675 1 18897
2 97676 1 18904
2 97677 1 18904
2 97678 1 18906
2 97679 1 18906
2 97680 1 18906
2 97681 1 18906
2 97682 1 18906
2 97683 1 18906
2 97684 1 18907
2 97685 1 18907
2 97686 1 18907
2 97687 1 18907
2 97688 1 18908
2 97689 1 18908
2 97690 1 18913
2 97691 1 18913
2 97692 1 18913
2 97693 1 18921
2 97694 1 18921
2 97695 1 18921
2 97696 1 18921
2 97697 1 18921
2 97698 1 18921
2 97699 1 18921
2 97700 1 18921
2 97701 1 18922
2 97702 1 18922
2 97703 1 18923
2 97704 1 18923
2 97705 1 18923
2 97706 1 18923
2 97707 1 18926
2 97708 1 18926
2 97709 1 18946
2 97710 1 18946
2 97711 1 18964
2 97712 1 18964
2 97713 1 18966
2 97714 1 18966
2 97715 1 18967
2 97716 1 18967
2 97717 1 18967
2 97718 1 18967
2 97719 1 18967
2 97720 1 18967
2 97721 1 18967
2 97722 1 18967
2 97723 1 18967
2 97724 1 18967
2 97725 1 18967
2 97726 1 18967
2 97727 1 18967
2 97728 1 18968
2 97729 1 18968
2 97730 1 18984
2 97731 1 18984
2 97732 1 18984
2 97733 1 18984
2 97734 1 18984
2 97735 1 18984
2 97736 1 18984
2 97737 1 18984
2 97738 1 18984
2 97739 1 18984
2 97740 1 18984
2 97741 1 18984
2 97742 1 18984
2 97743 1 18984
2 97744 1 18984
2 97745 1 18984
2 97746 1 18984
2 97747 1 18984
2 97748 1 18984
2 97749 1 18986
2 97750 1 18986
2 97751 1 18986
2 97752 1 18986
2 97753 1 18986
2 97754 1 18986
2 97755 1 18986
2 97756 1 18986
2 97757 1 18986
2 97758 1 18995
2 97759 1 18995
2 97760 1 19016
2 97761 1 19016
2 97762 1 19017
2 97763 1 19017
2 97764 1 19034
2 97765 1 19034
2 97766 1 19037
2 97767 1 19037
2 97768 1 19037
2 97769 1 19037
2 97770 1 19037
2 97771 1 19037
2 97772 1 19037
2 97773 1 19053
2 97774 1 19053
2 97775 1 19053
2 97776 1 19053
2 97777 1 19053
2 97778 1 19054
2 97779 1 19054
2 97780 1 19054
2 97781 1 19054
2 97782 1 19055
2 97783 1 19055
2 97784 1 19057
2 97785 1 19057
2 97786 1 19058
2 97787 1 19058
2 97788 1 19062
2 97789 1 19062
2 97790 1 19062
2 97791 1 19062
2 97792 1 19066
2 97793 1 19066
2 97794 1 19077
2 97795 1 19077
2 97796 1 19083
2 97797 1 19083
2 97798 1 19090
2 97799 1 19090
2 97800 1 19102
2 97801 1 19102
2 97802 1 19102
2 97803 1 19102
2 97804 1 19102
2 97805 1 19104
2 97806 1 19104
2 97807 1 19105
2 97808 1 19105
2 97809 1 19117
2 97810 1 19117
2 97811 1 19131
2 97812 1 19131
2 97813 1 19132
2 97814 1 19132
2 97815 1 19133
2 97816 1 19133
2 97817 1 19136
2 97818 1 19136
2 97819 1 19136
2 97820 1 19140
2 97821 1 19140
2 97822 1 19140
2 97823 1 19143
2 97824 1 19143
2 97825 1 19143
2 97826 1 19144
2 97827 1 19144
2 97828 1 19144
2 97829 1 19144
2 97830 1 19146
2 97831 1 19146
2 97832 1 19147
2 97833 1 19147
2 97834 1 19147
2 97835 1 19147
2 97836 1 19148
2 97837 1 19148
2 97838 1 19152
2 97839 1 19152
2 97840 1 19155
2 97841 1 19155
2 97842 1 19156
2 97843 1 19156
2 97844 1 19162
2 97845 1 19162
2 97846 1 19169
2 97847 1 19169
2 97848 1 19177
2 97849 1 19177
2 97850 1 19177
2 97851 1 19178
2 97852 1 19178
2 97853 1 19197
2 97854 1 19197
2 97855 1 19197
2 97856 1 19197
2 97857 1 19198
2 97858 1 19198
2 97859 1 19198
2 97860 1 19198
2 97861 1 19198
2 97862 1 19199
2 97863 1 19199
2 97864 1 19199
2 97865 1 19200
2 97866 1 19200
2 97867 1 19200
2 97868 1 19200
2 97869 1 19200
2 97870 1 19200
2 97871 1 19201
2 97872 1 19201
2 97873 1 19201
2 97874 1 19201
2 97875 1 19201
2 97876 1 19201
2 97877 1 19201
2 97878 1 19201
2 97879 1 19201
2 97880 1 19201
2 97881 1 19201
2 97882 1 19201
2 97883 1 19201
2 97884 1 19201
2 97885 1 19201
2 97886 1 19201
2 97887 1 19201
2 97888 1 19201
2 97889 1 19202
2 97890 1 19202
2 97891 1 19202
2 97892 1 19205
2 97893 1 19205
2 97894 1 19205
2 97895 1 19205
2 97896 1 19205
2 97897 1 19205
2 97898 1 19205
2 97899 1 19205
2 97900 1 19205
2 97901 1 19205
2 97902 1 19205
2 97903 1 19205
2 97904 1 19205
2 97905 1 19205
2 97906 1 19205
2 97907 1 19205
2 97908 1 19205
2 97909 1 19205
2 97910 1 19205
2 97911 1 19205
2 97912 1 19205
2 97913 1 19205
2 97914 1 19205
2 97915 1 19205
2 97916 1 19205
2 97917 1 19206
2 97918 1 19206
2 97919 1 19206
2 97920 1 19206
2 97921 1 19206
2 97922 1 19206
2 97923 1 19206
2 97924 1 19206
2 97925 1 19206
2 97926 1 19207
2 97927 1 19207
2 97928 1 19207
2 97929 1 19208
2 97930 1 19208
2 97931 1 19208
2 97932 1 19208
2 97933 1 19208
2 97934 1 19208
2 97935 1 19208
2 97936 1 19208
2 97937 1 19209
2 97938 1 19209
2 97939 1 19209
2 97940 1 19209
2 97941 1 19210
2 97942 1 19210
2 97943 1 19210
2 97944 1 19210
2 97945 1 19211
2 97946 1 19211
2 97947 1 19218
2 97948 1 19218
2 97949 1 19224
2 97950 1 19224
2 97951 1 19224
2 97952 1 19224
2 97953 1 19224
2 97954 1 19224
2 97955 1 19224
2 97956 1 19224
2 97957 1 19224
2 97958 1 19224
2 97959 1 19237
2 97960 1 19237
2 97961 1 19237
2 97962 1 19237
2 97963 1 19237
2 97964 1 19237
2 97965 1 19237
2 97966 1 19237
2 97967 1 19237
2 97968 1 19237
2 97969 1 19239
2 97970 1 19239
2 97971 1 19239
2 97972 1 19246
2 97973 1 19246
2 97974 1 19260
2 97975 1 19260
2 97976 1 19263
2 97977 1 19263
2 97978 1 19270
2 97979 1 19270
2 97980 1 19270
2 97981 1 19270
2 97982 1 19271
2 97983 1 19271
2 97984 1 19279
2 97985 1 19279
2 97986 1 19288
2 97987 1 19288
2 97988 1 19298
2 97989 1 19298
2 97990 1 19298
2 97991 1 19298
2 97992 1 19321
2 97993 1 19321
2 97994 1 19333
2 97995 1 19333
2 97996 1 19335
2 97997 1 19335
2 97998 1 19337
2 97999 1 19337
2 98000 1 19337
2 98001 1 19337
2 98002 1 19337
2 98003 1 19340
2 98004 1 19340
2 98005 1 19340
2 98006 1 19340
2 98007 1 19340
2 98008 1 19343
2 98009 1 19343
2 98010 1 19352
2 98011 1 19352
2 98012 1 19352
2 98013 1 19352
2 98014 1 19352
2 98015 1 19352
2 98016 1 19352
2 98017 1 19362
2 98018 1 19362
2 98019 1 19362
2 98020 1 19362
2 98021 1 19362
2 98022 1 19362
2 98023 1 19362
2 98024 1 19362
2 98025 1 19362
2 98026 1 19362
2 98027 1 19362
2 98028 1 19362
2 98029 1 19362
2 98030 1 19362
2 98031 1 19362
2 98032 1 19362
2 98033 1 19362
2 98034 1 19362
2 98035 1 19362
2 98036 1 19362
2 98037 1 19362
2 98038 1 19362
2 98039 1 19362
2 98040 1 19362
2 98041 1 19362
2 98042 1 19363
2 98043 1 19363
2 98044 1 19369
2 98045 1 19369
2 98046 1 19369
2 98047 1 19369
2 98048 1 19370
2 98049 1 19370
2 98050 1 19370
2 98051 1 19371
2 98052 1 19371
2 98053 1 19374
2 98054 1 19374
2 98055 1 19374
2 98056 1 19383
2 98057 1 19383
2 98058 1 19383
2 98059 1 19401
2 98060 1 19401
2 98061 1 19410
2 98062 1 19410
2 98063 1 19411
2 98064 1 19411
2 98065 1 19414
2 98066 1 19414
2 98067 1 19421
2 98068 1 19421
2 98069 1 19422
2 98070 1 19422
2 98071 1 19422
2 98072 1 19426
2 98073 1 19426
2 98074 1 19426
2 98075 1 19441
2 98076 1 19441
2 98077 1 19450
2 98078 1 19450
2 98079 1 19454
2 98080 1 19454
2 98081 1 19454
2 98082 1 19454
2 98083 1 19454
2 98084 1 19454
2 98085 1 19466
2 98086 1 19466
2 98087 1 19466
2 98088 1 19466
2 98089 1 19481
2 98090 1 19481
2 98091 1 19482
2 98092 1 19482
2 98093 1 19482
2 98094 1 19482
2 98095 1 19483
2 98096 1 19483
2 98097 1 19483
2 98098 1 19483
2 98099 1 19483
2 98100 1 19491
2 98101 1 19491
2 98102 1 19491
2 98103 1 19491
2 98104 1 19491
2 98105 1 19500
2 98106 1 19500
2 98107 1 19523
2 98108 1 19523
2 98109 1 19523
2 98110 1 19528
2 98111 1 19528
2 98112 1 19528
2 98113 1 19528
2 98114 1 19528
2 98115 1 19528
2 98116 1 19528
2 98117 1 19528
2 98118 1 19529
2 98119 1 19529
2 98120 1 19529
2 98121 1 19529
2 98122 1 19533
2 98123 1 19533
2 98124 1 19533
2 98125 1 19533
2 98126 1 19534
2 98127 1 19534
2 98128 1 19534
2 98129 1 19534
2 98130 1 19534
2 98131 1 19535
2 98132 1 19535
2 98133 1 19545
2 98134 1 19545
2 98135 1 19546
2 98136 1 19546
2 98137 1 19546
2 98138 1 19546
2 98139 1 19546
2 98140 1 19546
2 98141 1 19547
2 98142 1 19547
2 98143 1 19548
2 98144 1 19548
2 98145 1 19552
2 98146 1 19552
2 98147 1 19552
2 98148 1 19552
2 98149 1 19552
2 98150 1 19552
2 98151 1 19553
2 98152 1 19553
2 98153 1 19553
2 98154 1 19553
2 98155 1 19561
2 98156 1 19561
2 98157 1 19561
2 98158 1 19561
2 98159 1 19561
2 98160 1 19561
2 98161 1 19561
2 98162 1 19562
2 98163 1 19562
2 98164 1 19565
2 98165 1 19565
2 98166 1 19565
2 98167 1 19566
2 98168 1 19566
2 98169 1 19571
2 98170 1 19571
2 98171 1 19601
2 98172 1 19601
2 98173 1 19601
2 98174 1 19601
2 98175 1 19601
2 98176 1 19601
2 98177 1 19601
2 98178 1 19601
2 98179 1 19601
2 98180 1 19601
2 98181 1 19601
2 98182 1 19601
2 98183 1 19602
2 98184 1 19602
2 98185 1 19614
2 98186 1 19614
2 98187 1 19614
2 98188 1 19614
2 98189 1 19614
2 98190 1 19614
2 98191 1 19614
2 98192 1 19614
2 98193 1 19614
2 98194 1 19614
2 98195 1 19615
2 98196 1 19615
2 98197 1 19615
2 98198 1 19615
2 98199 1 19615
2 98200 1 19616
2 98201 1 19616
2 98202 1 19616
2 98203 1 19616
2 98204 1 19616
2 98205 1 19616
2 98206 1 19616
2 98207 1 19616
2 98208 1 19617
2 98209 1 19617
2 98210 1 19628
2 98211 1 19628
2 98212 1 19628
2 98213 1 19628
2 98214 1 19628
2 98215 1 19628
2 98216 1 19628
2 98217 1 19628
2 98218 1 19640
2 98219 1 19640
2 98220 1 19640
2 98221 1 19640
2 98222 1 19640
2 98223 1 19640
2 98224 1 19640
2 98225 1 19640
2 98226 1 19641
2 98227 1 19641
2 98228 1 19641
2 98229 1 19641
2 98230 1 19641
2 98231 1 19641
2 98232 1 19642
2 98233 1 19642
2 98234 1 19642
2 98235 1 19642
2 98236 1 19642
2 98237 1 19642
2 98238 1 19642
2 98239 1 19642
2 98240 1 19642
2 98241 1 19642
2 98242 1 19642
2 98243 1 19642
2 98244 1 19642
2 98245 1 19642
2 98246 1 19643
2 98247 1 19643
2 98248 1 19643
2 98249 1 19643
2 98250 1 19643
2 98251 1 19644
2 98252 1 19644
2 98253 1 19644
2 98254 1 19646
2 98255 1 19646
2 98256 1 19646
2 98257 1 19646
2 98258 1 19646
2 98259 1 19646
2 98260 1 19646
2 98261 1 19646
2 98262 1 19646
2 98263 1 19646
2 98264 1 19647
2 98265 1 19647
2 98266 1 19649
2 98267 1 19649
2 98268 1 19649
2 98269 1 19649
2 98270 1 19649
2 98271 1 19649
2 98272 1 19649
2 98273 1 19649
2 98274 1 19649
2 98275 1 19649
2 98276 1 19649
2 98277 1 19649
2 98278 1 19649
2 98279 1 19649
2 98280 1 19649
2 98281 1 19649
2 98282 1 19649
2 98283 1 19650
2 98284 1 19650
2 98285 1 19651
2 98286 1 19651
2 98287 1 19651
2 98288 1 19651
2 98289 1 19651
2 98290 1 19651
2 98291 1 19651
2 98292 1 19651
2 98293 1 19651
2 98294 1 19658
2 98295 1 19658
2 98296 1 19671
2 98297 1 19671
2 98298 1 19716
2 98299 1 19716
2 98300 1 19729
2 98301 1 19729
2 98302 1 19729
2 98303 1 19729
2 98304 1 19729
2 98305 1 19730
2 98306 1 19730
2 98307 1 19742
2 98308 1 19742
2 98309 1 19742
2 98310 1 19743
2 98311 1 19743
2 98312 1 19757
2 98313 1 19757
2 98314 1 19774
2 98315 1 19774
2 98316 1 19784
2 98317 1 19784
2 98318 1 19784
2 98319 1 19786
2 98320 1 19786
2 98321 1 19786
2 98322 1 19792
2 98323 1 19792
2 98324 1 19792
2 98325 1 19807
2 98326 1 19807
2 98327 1 19807
2 98328 1 19807
2 98329 1 19807
2 98330 1 19808
2 98331 1 19808
2 98332 1 19808
2 98333 1 19810
2 98334 1 19810
2 98335 1 19810
2 98336 1 19810
2 98337 1 19820
2 98338 1 19820
2 98339 1 19820
2 98340 1 19820
2 98341 1 19820
2 98342 1 19820
2 98343 1 19820
2 98344 1 19820
2 98345 1 19820
2 98346 1 19820
2 98347 1 19820
2 98348 1 19820
2 98349 1 19820
2 98350 1 19828
2 98351 1 19828
2 98352 1 19833
2 98353 1 19833
2 98354 1 19874
2 98355 1 19874
2 98356 1 19884
2 98357 1 19884
2 98358 1 19884
2 98359 1 19884
2 98360 1 19884
2 98361 1 19892
2 98362 1 19892
2 98363 1 19892
2 98364 1 19892
2 98365 1 19900
2 98366 1 19900
2 98367 1 19900
2 98368 1 19902
2 98369 1 19902
2 98370 1 19915
2 98371 1 19915
2 98372 1 19915
2 98373 1 19915
2 98374 1 19915
2 98375 1 19915
2 98376 1 19915
2 98377 1 19915
2 98378 1 19915
2 98379 1 19915
2 98380 1 19915
2 98381 1 19919
2 98382 1 19919
2 98383 1 19919
2 98384 1 19919
2 98385 1 19919
2 98386 1 19919
2 98387 1 19919
2 98388 1 19919
2 98389 1 19946
2 98390 1 19946
2 98391 1 19946
2 98392 1 19947
2 98393 1 19947
2 98394 1 19947
2 98395 1 19947
2 98396 1 19948
2 98397 1 19948
2 98398 1 19948
2 98399 1 19948
2 98400 1 19948
2 98401 1 19949
2 98402 1 19949
2 98403 1 19951
2 98404 1 19951
2 98405 1 19951
2 98406 1 19951
2 98407 1 19951
2 98408 1 19951
2 98409 1 19951
2 98410 1 19951
2 98411 1 19951
2 98412 1 19951
2 98413 1 19951
2 98414 1 19951
2 98415 1 19951
2 98416 1 19951
2 98417 1 19951
2 98418 1 19954
2 98419 1 19954
2 98420 1 19954
2 98421 1 19954
2 98422 1 19954
2 98423 1 19954
2 98424 1 19954
2 98425 1 19954
2 98426 1 19954
2 98427 1 19954
2 98428 1 19954
2 98429 1 19954
2 98430 1 19954
2 98431 1 19954
2 98432 1 19954
2 98433 1 19954
2 98434 1 19954
2 98435 1 19954
2 98436 1 19954
2 98437 1 19954
2 98438 1 19954
2 98439 1 19954
2 98440 1 19954
2 98441 1 19954
2 98442 1 19954
2 98443 1 19954
2 98444 1 19954
2 98445 1 19954
2 98446 1 19955
2 98447 1 19955
2 98448 1 19956
2 98449 1 19956
2 98450 1 19956
2 98451 1 19956
2 98452 1 19956
2 98453 1 19956
2 98454 1 19956
2 98455 1 19964
2 98456 1 19964
2 98457 1 19964
2 98458 1 19964
2 98459 1 19964
2 98460 1 19964
2 98461 1 19964
2 98462 1 19964
2 98463 1 19964
2 98464 1 19964
2 98465 1 19964
2 98466 1 19964
2 98467 1 19965
2 98468 1 19965
2 98469 1 19967
2 98470 1 19967
2 98471 1 19972
2 98472 1 19972
2 98473 1 19972
2 98474 1 19972
2 98475 1 19972
2 98476 1 19972
2 98477 1 19972
2 98478 1 19979
2 98479 1 19979
2 98480 1 19979
2 98481 1 19979
2 98482 1 19979
2 98483 1 19983
2 98484 1 19983
2 98485 1 19983
2 98486 1 19983
2 98487 1 19983
2 98488 1 19983
2 98489 1 19983
2 98490 1 19983
2 98491 1 19983
2 98492 1 19983
2 98493 1 19983
2 98494 1 19983
2 98495 1 19983
2 98496 1 19983
2 98497 1 19983
2 98498 1 19983
2 98499 1 19983
2 98500 1 19983
2 98501 1 19983
2 98502 1 19983
2 98503 1 19983
2 98504 1 19983
2 98505 1 19983
2 98506 1 19983
2 98507 1 19983
2 98508 1 19983
2 98509 1 19983
2 98510 1 19983
2 98511 1 19983
2 98512 1 19983
2 98513 1 19983
2 98514 1 19983
2 98515 1 19983
2 98516 1 19994
2 98517 1 19994
2 98518 1 20019
2 98519 1 20019
2 98520 1 20019
2 98521 1 20019
2 98522 1 20019
2 98523 1 20019
2 98524 1 20019
2 98525 1 20019
2 98526 1 20019
2 98527 1 20019
2 98528 1 20024
2 98529 1 20024
2 98530 1 20024
2 98531 1 20033
2 98532 1 20033
2 98533 1 20033
2 98534 1 20040
2 98535 1 20040
2 98536 1 20054
2 98537 1 20054
2 98538 1 20071
2 98539 1 20071
2 98540 1 20072
2 98541 1 20072
2 98542 1 20072
2 98543 1 20072
2 98544 1 20072
2 98545 1 20072
2 98546 1 20072
2 98547 1 20090
2 98548 1 20090
2 98549 1 20097
2 98550 1 20097
2 98551 1 20097
2 98552 1 20097
2 98553 1 20097
2 98554 1 20097
2 98555 1 20097
2 98556 1 20098
2 98557 1 20098
2 98558 1 20098
2 98559 1 20098
2 98560 1 20098
2 98561 1 20116
2 98562 1 20116
2 98563 1 20127
2 98564 1 20127
2 98565 1 20128
2 98566 1 20128
2 98567 1 20199
2 98568 1 20199
2 98569 1 20210
2 98570 1 20210
2 98571 1 20232
2 98572 1 20232
2 98573 1 20247
2 98574 1 20247
2 98575 1 20264
2 98576 1 20264
2 98577 1 20264
2 98578 1 20264
2 98579 1 20264
2 98580 1 20264
2 98581 1 20264
2 98582 1 20264
2 98583 1 20265
2 98584 1 20265
2 98585 1 20267
2 98586 1 20267
2 98587 1 20268
2 98588 1 20268
2 98589 1 20268
2 98590 1 20268
2 98591 1 20268
2 98592 1 20268
2 98593 1 20268
2 98594 1 20268
2 98595 1 20268
2 98596 1 20268
2 98597 1 20268
2 98598 1 20268
2 98599 1 20268
2 98600 1 20268
2 98601 1 20272
2 98602 1 20272
2 98603 1 20272
2 98604 1 20272
2 98605 1 20272
2 98606 1 20279
2 98607 1 20279
2 98608 1 20279
2 98609 1 20279
2 98610 1 20279
2 98611 1 20279
2 98612 1 20279
2 98613 1 20279
2 98614 1 20279
2 98615 1 20279
2 98616 1 20279
2 98617 1 20279
2 98618 1 20279
2 98619 1 20279
2 98620 1 20279
2 98621 1 20279
2 98622 1 20280
2 98623 1 20280
2 98624 1 20283
2 98625 1 20283
2 98626 1 20308
2 98627 1 20308
2 98628 1 20308
2 98629 1 20308
2 98630 1 20308
2 98631 1 20308
2 98632 1 20323
2 98633 1 20323
2 98634 1 20334
2 98635 1 20334
2 98636 1 20361
2 98637 1 20361
2 98638 1 20361
2 98639 1 20361
2 98640 1 20362
2 98641 1 20362
2 98642 1 20362
2 98643 1 20404
2 98644 1 20404
2 98645 1 20404
2 98646 1 20406
2 98647 1 20406
2 98648 1 20411
2 98649 1 20411
2 98650 1 20411
2 98651 1 20411
2 98652 1 20411
2 98653 1 20416
2 98654 1 20416
2 98655 1 20426
2 98656 1 20426
2 98657 1 20426
2 98658 1 20426
2 98659 1 20426
2 98660 1 20426
2 98661 1 20427
2 98662 1 20427
2 98663 1 20435
2 98664 1 20435
2 98665 1 20443
2 98666 1 20443
2 98667 1 20462
2 98668 1 20462
2 98669 1 20462
2 98670 1 20463
2 98671 1 20463
2 98672 1 20463
2 98673 1 20467
2 98674 1 20467
2 98675 1 20467
2 98676 1 20467
2 98677 1 20472
2 98678 1 20472
2 98679 1 20472
2 98680 1 20481
2 98681 1 20481
2 98682 1 20481
2 98683 1 20481
2 98684 1 20481
2 98685 1 20481
2 98686 1 20487
2 98687 1 20487
2 98688 1 20487
2 98689 1 20487
2 98690 1 20487
2 98691 1 20487
2 98692 1 20487
2 98693 1 20487
2 98694 1 20487
2 98695 1 20487
2 98696 1 20487
2 98697 1 20487
2 98698 1 20487
2 98699 1 20487
2 98700 1 20487
2 98701 1 20487
2 98702 1 20488
2 98703 1 20488
2 98704 1 20492
2 98705 1 20492
2 98706 1 20492
2 98707 1 20492
2 98708 1 20492
2 98709 1 20492
2 98710 1 20492
2 98711 1 20492
2 98712 1 20492
2 98713 1 20492
2 98714 1 20492
2 98715 1 20492
2 98716 1 20493
2 98717 1 20493
2 98718 1 20493
2 98719 1 20496
2 98720 1 20496
2 98721 1 20497
2 98722 1 20497
2 98723 1 20500
2 98724 1 20500
2 98725 1 20503
2 98726 1 20503
2 98727 1 20507
2 98728 1 20507
2 98729 1 20519
2 98730 1 20519
2 98731 1 20519
2 98732 1 20519
2 98733 1 20519
2 98734 1 20519
2 98735 1 20520
2 98736 1 20520
2 98737 1 20521
2 98738 1 20521
2 98739 1 20524
2 98740 1 20524
2 98741 1 20524
2 98742 1 20524
2 98743 1 20524
2 98744 1 20524
2 98745 1 20524
2 98746 1 20524
2 98747 1 20524
2 98748 1 20524
2 98749 1 20524
2 98750 1 20539
2 98751 1 20539
2 98752 1 20547
2 98753 1 20547
2 98754 1 20547
2 98755 1 20547
2 98756 1 20547
2 98757 1 20547
2 98758 1 20547
2 98759 1 20547
2 98760 1 20547
2 98761 1 20547
2 98762 1 20547
2 98763 1 20547
2 98764 1 20547
2 98765 1 20547
2 98766 1 20547
2 98767 1 20547
2 98768 1 20547
2 98769 1 20547
2 98770 1 20547
2 98771 1 20547
2 98772 1 20547
2 98773 1 20547
2 98774 1 20547
2 98775 1 20547
2 98776 1 20547
2 98777 1 20547
2 98778 1 20547
2 98779 1 20547
2 98780 1 20548
2 98781 1 20548
2 98782 1 20574
2 98783 1 20574
2 98784 1 20575
2 98785 1 20575
2 98786 1 20601
2 98787 1 20601
2 98788 1 20619
2 98789 1 20619
2 98790 1 20622
2 98791 1 20622
2 98792 1 20622
2 98793 1 20622
2 98794 1 20624
2 98795 1 20624
2 98796 1 20624
2 98797 1 20624
2 98798 1 20647
2 98799 1 20647
2 98800 1 20648
2 98801 1 20648
2 98802 1 20648
2 98803 1 20648
2 98804 1 20650
2 98805 1 20650
2 98806 1 20650
2 98807 1 20650
2 98808 1 20650
2 98809 1 20650
2 98810 1 20650
2 98811 1 20658
2 98812 1 20658
2 98813 1 20661
2 98814 1 20661
2 98815 1 20661
2 98816 1 20661
2 98817 1 20661
2 98818 1 20663
2 98819 1 20663
2 98820 1 20663
2 98821 1 20663
2 98822 1 20663
2 98823 1 20663
2 98824 1 20672
2 98825 1 20672
2 98826 1 20673
2 98827 1 20673
2 98828 1 20673
2 98829 1 20673
2 98830 1 20673
2 98831 1 20673
2 98832 1 20674
2 98833 1 20674
2 98834 1 20676
2 98835 1 20676
2 98836 1 20676
2 98837 1 20685
2 98838 1 20685
2 98839 1 20685
2 98840 1 20685
2 98841 1 20685
2 98842 1 20685
2 98843 1 20688
2 98844 1 20688
2 98845 1 20688
2 98846 1 20711
2 98847 1 20711
2 98848 1 20725
2 98849 1 20725
2 98850 1 20725
2 98851 1 20725
2 98852 1 20726
2 98853 1 20726
2 98854 1 20734
2 98855 1 20734
2 98856 1 20734
2 98857 1 20735
2 98858 1 20735
2 98859 1 20735
2 98860 1 20735
2 98861 1 20735
2 98862 1 20763
2 98863 1 20763
2 98864 1 20764
2 98865 1 20764
2 98866 1 20773
2 98867 1 20773
2 98868 1 20773
2 98869 1 20773
2 98870 1 20809
2 98871 1 20809
2 98872 1 20810
2 98873 1 20810
2 98874 1 20810
2 98875 1 20818
2 98876 1 20818
2 98877 1 20818
2 98878 1 20818
2 98879 1 20818
2 98880 1 20818
2 98881 1 20819
2 98882 1 20819
2 98883 1 20819
2 98884 1 20820
2 98885 1 20820
2 98886 1 20830
2 98887 1 20830
2 98888 1 20838
2 98889 1 20838
2 98890 1 20838
2 98891 1 20839
2 98892 1 20839
2 98893 1 20839
2 98894 1 20839
2 98895 1 20839
2 98896 1 20839
2 98897 1 20839
2 98898 1 20840
2 98899 1 20840
2 98900 1 20841
2 98901 1 20841
2 98902 1 20841
2 98903 1 20841
2 98904 1 20854
2 98905 1 20854
2 98906 1 20865
2 98907 1 20865
2 98908 1 20865
2 98909 1 20867
2 98910 1 20867
2 98911 1 20897
2 98912 1 20897
2 98913 1 20897
2 98914 1 20897
2 98915 1 20897
2 98916 1 20897
2 98917 1 20897
2 98918 1 20897
2 98919 1 20897
2 98920 1 20897
2 98921 1 20897
2 98922 1 20897
2 98923 1 20897
2 98924 1 20897
2 98925 1 20897
2 98926 1 20898
2 98927 1 20898
2 98928 1 20901
2 98929 1 20901
2 98930 1 20903
2 98931 1 20903
2 98932 1 20913
2 98933 1 20913
2 98934 1 20920
2 98935 1 20920
2 98936 1 20920
2 98937 1 20921
2 98938 1 20921
2 98939 1 20921
2 98940 1 20921
2 98941 1 20921
2 98942 1 20921
2 98943 1 20921
2 98944 1 20921
2 98945 1 20921
2 98946 1 20933
2 98947 1 20933
2 98948 1 20943
2 98949 1 20943
2 98950 1 20944
2 98951 1 20944
2 98952 1 20952
2 98953 1 20952
2 98954 1 20952
2 98955 1 20968
2 98956 1 20968
2 98957 1 20997
2 98958 1 20997
2 98959 1 21000
2 98960 1 21000
2 98961 1 21000
2 98962 1 21044
2 98963 1 21044
2 98964 1 21044
2 98965 1 21044
2 98966 1 21044
2 98967 1 21044
2 98968 1 21053
2 98969 1 21053
2 98970 1 21054
2 98971 1 21054
2 98972 1 21054
2 98973 1 21055
2 98974 1 21055
2 98975 1 21055
2 98976 1 21055
2 98977 1 21055
2 98978 1 21055
2 98979 1 21055
2 98980 1 21055
2 98981 1 21059
2 98982 1 21059
2 98983 1 21059
2 98984 1 21060
2 98985 1 21060
2 98986 1 21060
2 98987 1 21096
2 98988 1 21096
2 98989 1 21103
2 98990 1 21103
2 98991 1 21103
2 98992 1 21103
2 98993 1 21105
2 98994 1 21105
2 98995 1 21116
2 98996 1 21116
2 98997 1 21117
2 98998 1 21117
2 98999 1 21119
2 99000 1 21119
2 99001 1 21121
2 99002 1 21121
2 99003 1 21121
2 99004 1 21141
2 99005 1 21141
2 99006 1 21150
2 99007 1 21150
2 99008 1 21165
2 99009 1 21165
2 99010 1 21165
2 99011 1 21166
2 99012 1 21166
2 99013 1 21184
2 99014 1 21184
2 99015 1 21195
2 99016 1 21195
2 99017 1 21219
2 99018 1 21219
2 99019 1 21219
2 99020 1 21219
2 99021 1 21219
2 99022 1 21219
2 99023 1 21243
2 99024 1 21243
2 99025 1 21243
2 99026 1 21268
2 99027 1 21268
2 99028 1 21268
2 99029 1 21268
2 99030 1 21268
2 99031 1 21268
2 99032 1 21268
2 99033 1 21268
2 99034 1 21268
2 99035 1 21268
2 99036 1 21269
2 99037 1 21269
2 99038 1 21269
2 99039 1 21276
2 99040 1 21276
2 99041 1 21276
2 99042 1 21281
2 99043 1 21281
2 99044 1 21288
2 99045 1 21288
2 99046 1 21291
2 99047 1 21291
2 99048 1 21294
2 99049 1 21294
2 99050 1 21294
2 99051 1 21294
2 99052 1 21316
2 99053 1 21316
2 99054 1 21329
2 99055 1 21329
2 99056 1 21340
2 99057 1 21340
2 99058 1 21345
2 99059 1 21345
2 99060 1 21345
2 99061 1 21346
2 99062 1 21346
2 99063 1 21347
2 99064 1 21347
2 99065 1 21348
2 99066 1 21348
2 99067 1 21348
2 99068 1 21348
2 99069 1 21348
2 99070 1 21350
2 99071 1 21350
2 99072 1 21354
2 99073 1 21354
2 99074 1 21355
2 99075 1 21355
2 99076 1 21356
2 99077 1 21356
2 99078 1 21356
2 99079 1 21356
2 99080 1 21356
2 99081 1 21356
2 99082 1 21357
2 99083 1 21357
2 99084 1 21357
2 99085 1 21403
2 99086 1 21403
2 99087 1 21403
2 99088 1 21403
2 99089 1 21403
2 99090 1 21404
2 99091 1 21404
2 99092 1 21404
2 99093 1 21404
2 99094 1 21404
2 99095 1 21416
2 99096 1 21416
2 99097 1 21417
2 99098 1 21417
2 99099 1 21417
2 99100 1 21418
2 99101 1 21418
2 99102 1 21419
2 99103 1 21419
2 99104 1 21419
2 99105 1 21420
2 99106 1 21420
2 99107 1 21427
2 99108 1 21427
2 99109 1 21434
2 99110 1 21434
2 99111 1 21437
2 99112 1 21437
2 99113 1 21437
2 99114 1 21478
2 99115 1 21478
2 99116 1 21486
2 99117 1 21486
2 99118 1 21497
2 99119 1 21497
2 99120 1 21497
2 99121 1 21499
2 99122 1 21499
2 99123 1 21514
2 99124 1 21514
2 99125 1 21515
2 99126 1 21515
2 99127 1 21524
2 99128 1 21524
2 99129 1 21536
2 99130 1 21536
2 99131 1 21536
2 99132 1 21536
2 99133 1 21536
2 99134 1 21536
2 99135 1 21536
2 99136 1 21537
2 99137 1 21537
2 99138 1 21537
2 99139 1 21546
2 99140 1 21546
2 99141 1 21546
2 99142 1 21546
2 99143 1 21546
2 99144 1 21547
2 99145 1 21547
2 99146 1 21547
2 99147 1 21558
2 99148 1 21558
2 99149 1 21558
2 99150 1 21570
2 99151 1 21570
2 99152 1 21570
2 99153 1 21570
2 99154 1 21570
2 99155 1 21570
2 99156 1 21570
2 99157 1 21570
2 99158 1 21570
2 99159 1 21570
2 99160 1 21571
2 99161 1 21571
2 99162 1 21571
2 99163 1 21572
2 99164 1 21572
2 99165 1 21578
2 99166 1 21578
2 99167 1 21581
2 99168 1 21581
2 99169 1 21581
2 99170 1 21581
2 99171 1 21583
2 99172 1 21583
2 99173 1 21583
2 99174 1 21583
2 99175 1 21583
2 99176 1 21583
2 99177 1 21583
2 99178 1 21583
2 99179 1 21600
2 99180 1 21600
2 99181 1 21601
2 99182 1 21601
2 99183 1 21601
2 99184 1 21601
2 99185 1 21601
2 99186 1 21601
2 99187 1 21601
2 99188 1 21601
2 99189 1 21601
2 99190 1 21601
2 99191 1 21609
2 99192 1 21609
2 99193 1 21609
2 99194 1 21610
2 99195 1 21610
2 99196 1 21610
2 99197 1 21611
2 99198 1 21611
2 99199 1 21612
2 99200 1 21612
2 99201 1 21617
2 99202 1 21617
2 99203 1 21619
2 99204 1 21619
2 99205 1 21621
2 99206 1 21621
2 99207 1 21621
2 99208 1 21621
2 99209 1 21621
2 99210 1 21621
2 99211 1 21621
2 99212 1 21621
2 99213 1 21621
2 99214 1 21632
2 99215 1 21632
2 99216 1 21668
2 99217 1 21668
2 99218 1 21668
2 99219 1 21668
2 99220 1 21668
2 99221 1 21688
2 99222 1 21688
2 99223 1 21688
2 99224 1 21697
2 99225 1 21697
2 99226 1 21697
2 99227 1 21720
2 99228 1 21720
2 99229 1 21720
2 99230 1 21721
2 99231 1 21721
2 99232 1 21721
2 99233 1 21721
2 99234 1 21721
2 99235 1 21733
2 99236 1 21733
2 99237 1 21740
2 99238 1 21740
2 99239 1 21748
2 99240 1 21748
2 99241 1 21748
2 99242 1 21748
2 99243 1 21749
2 99244 1 21749
2 99245 1 21749
2 99246 1 21767
2 99247 1 21767
2 99248 1 21773
2 99249 1 21773
2 99250 1 21773
2 99251 1 21774
2 99252 1 21774
2 99253 1 21775
2 99254 1 21775
2 99255 1 21775
2 99256 1 21775
2 99257 1 21788
2 99258 1 21788
2 99259 1 21788
2 99260 1 21794
2 99261 1 21794
2 99262 1 21794
2 99263 1 21794
2 99264 1 21794
2 99265 1 21794
2 99266 1 21794
2 99267 1 21794
2 99268 1 21794
2 99269 1 21794
2 99270 1 21794
2 99271 1 21818
2 99272 1 21818
2 99273 1 21818
2 99274 1 21818
2 99275 1 21818
2 99276 1 21818
2 99277 1 21818
2 99278 1 21819
2 99279 1 21819
2 99280 1 21844
2 99281 1 21844
2 99282 1 21852
2 99283 1 21852
2 99284 1 21852
2 99285 1 21881
2 99286 1 21881
2 99287 1 21901
2 99288 1 21901
2 99289 1 21901
2 99290 1 21902
2 99291 1 21902
2 99292 1 21907
2 99293 1 21907
2 99294 1 21907
2 99295 1 21907
2 99296 1 21907
2 99297 1 21907
2 99298 1 21907
2 99299 1 21907
2 99300 1 21907
2 99301 1 21907
2 99302 1 21908
2 99303 1 21908
2 99304 1 21908
2 99305 1 21909
2 99306 1 21909
2 99307 1 21909
2 99308 1 21931
2 99309 1 21931
2 99310 1 21931
2 99311 1 21938
2 99312 1 21938
2 99313 1 21945
2 99314 1 21945
2 99315 1 21945
2 99316 1 21945
2 99317 1 21947
2 99318 1 21947
2 99319 1 21947
2 99320 1 21947
2 99321 1 21953
2 99322 1 21953
2 99323 1 21953
2 99324 1 21963
2 99325 1 21963
2 99326 1 21963
2 99327 1 21963
2 99328 1 21963
2 99329 1 21963
2 99330 1 21967
2 99331 1 21967
2 99332 1 21971
2 99333 1 21971
2 99334 1 21972
2 99335 1 21972
2 99336 1 21975
2 99337 1 21975
2 99338 1 21991
2 99339 1 21991
2 99340 1 21991
2 99341 1 22011
2 99342 1 22011
2 99343 1 22011
2 99344 1 22011
2 99345 1 22011
2 99346 1 22011
2 99347 1 22013
2 99348 1 22013
2 99349 1 22013
2 99350 1 22013
2 99351 1 22013
2 99352 1 22013
2 99353 1 22015
2 99354 1 22015
2 99355 1 22015
2 99356 1 22015
2 99357 1 22015
2 99358 1 22016
2 99359 1 22016
2 99360 1 22016
2 99361 1 22016
2 99362 1 22016
2 99363 1 22016
2 99364 1 22016
2 99365 1 22016
2 99366 1 22016
2 99367 1 22016
2 99368 1 22016
2 99369 1 22016
2 99370 1 22016
2 99371 1 22016
2 99372 1 22016
2 99373 1 22016
2 99374 1 22016
2 99375 1 22016
2 99376 1 22016
2 99377 1 22016
2 99378 1 22016
2 99379 1 22016
2 99380 1 22017
2 99381 1 22017
2 99382 1 22017
2 99383 1 22017
2 99384 1 22017
2 99385 1 22017
2 99386 1 22017
2 99387 1 22017
2 99388 1 22017
2 99389 1 22017
2 99390 1 22017
2 99391 1 22017
2 99392 1 22017
2 99393 1 22017
2 99394 1 22017
2 99395 1 22017
2 99396 1 22017
2 99397 1 22017
2 99398 1 22017
2 99399 1 22019
2 99400 1 22019
2 99401 1 22019
2 99402 1 22019
2 99403 1 22019
2 99404 1 22019
2 99405 1 22019
2 99406 1 22019
2 99407 1 22019
2 99408 1 22019
2 99409 1 22019
2 99410 1 22019
2 99411 1 22019
2 99412 1 22019
2 99413 1 22019
2 99414 1 22019
2 99415 1 22019
2 99416 1 22019
2 99417 1 22019
2 99418 1 22020
2 99419 1 22020
2 99420 1 22020
2 99421 1 22026
2 99422 1 22026
2 99423 1 22026
2 99424 1 22026
2 99425 1 22026
2 99426 1 22034
2 99427 1 22034
2 99428 1 22034
2 99429 1 22035
2 99430 1 22035
2 99431 1 22035
2 99432 1 22036
2 99433 1 22036
2 99434 1 22036
2 99435 1 22036
2 99436 1 22036
2 99437 1 22037
2 99438 1 22037
2 99439 1 22037
2 99440 1 22037
2 99441 1 22047
2 99442 1 22047
2 99443 1 22047
2 99444 1 22047
2 99445 1 22047
2 99446 1 22047
2 99447 1 22047
2 99448 1 22047
2 99449 1 22047
2 99450 1 22047
2 99451 1 22047
2 99452 1 22047
2 99453 1 22047
2 99454 1 22047
2 99455 1 22047
2 99456 1 22048
2 99457 1 22048
2 99458 1 22049
2 99459 1 22049
2 99460 1 22049
2 99461 1 22049
2 99462 1 22049
2 99463 1 22049
2 99464 1 22049
2 99465 1 22049
2 99466 1 22049
2 99467 1 22050
2 99468 1 22050
2 99469 1 22050
2 99470 1 22051
2 99471 1 22051
2 99472 1 22052
2 99473 1 22052
2 99474 1 22054
2 99475 1 22054
2 99476 1 22054
2 99477 1 22054
2 99478 1 22054
2 99479 1 22054
2 99480 1 22054
2 99481 1 22054
2 99482 1 22054
2 99483 1 22054
2 99484 1 22054
2 99485 1 22054
2 99486 1 22054
2 99487 1 22054
2 99488 1 22054
2 99489 1 22055
2 99490 1 22055
2 99491 1 22055
2 99492 1 22056
2 99493 1 22056
2 99494 1 22065
2 99495 1 22065
2 99496 1 22067
2 99497 1 22067
2 99498 1 22068
2 99499 1 22068
2 99500 1 22076
2 99501 1 22076
2 99502 1 22077
2 99503 1 22077
2 99504 1 22079
2 99505 1 22079
2 99506 1 22082
2 99507 1 22082
2 99508 1 22082
2 99509 1 22083
2 99510 1 22083
2 99511 1 22099
2 99512 1 22099
2 99513 1 22102
2 99514 1 22102
2 99515 1 22102
2 99516 1 22119
2 99517 1 22119
2 99518 1 22125
2 99519 1 22125
2 99520 1 22131
2 99521 1 22131
2 99522 1 22131
2 99523 1 22131
2 99524 1 22131
2 99525 1 22131
2 99526 1 22132
2 99527 1 22132
2 99528 1 22139
2 99529 1 22139
2 99530 1 22139
2 99531 1 22140
2 99532 1 22140
2 99533 1 22140
2 99534 1 22140
2 99535 1 22141
2 99536 1 22141
2 99537 1 22155
2 99538 1 22155
2 99539 1 22155
2 99540 1 22155
2 99541 1 22155
2 99542 1 22156
2 99543 1 22156
2 99544 1 22157
2 99545 1 22157
2 99546 1 22165
2 99547 1 22165
2 99548 1 22183
2 99549 1 22183
2 99550 1 22183
2 99551 1 22183
2 99552 1 22183
2 99553 1 22183
2 99554 1 22183
2 99555 1 22183
2 99556 1 22183
2 99557 1 22193
2 99558 1 22193
2 99559 1 22193
2 99560 1 22193
2 99561 1 22200
2 99562 1 22200
2 99563 1 22207
2 99564 1 22207
2 99565 1 22207
2 99566 1 22207
2 99567 1 22207
2 99568 1 22207
2 99569 1 22207
2 99570 1 22207
2 99571 1 22207
2 99572 1 22208
2 99573 1 22208
2 99574 1 22208
2 99575 1 22227
2 99576 1 22227
2 99577 1 22227
2 99578 1 22238
2 99579 1 22238
2 99580 1 22242
2 99581 1 22242
2 99582 1 22255
2 99583 1 22255
2 99584 1 22263
2 99585 1 22263
2 99586 1 22265
2 99587 1 22265
2 99588 1 22267
2 99589 1 22267
2 99590 1 22278
2 99591 1 22278
2 99592 1 22278
2 99593 1 22278
2 99594 1 22279
2 99595 1 22279
2 99596 1 22281
2 99597 1 22281
2 99598 1 22292
2 99599 1 22292
2 99600 1 22306
2 99601 1 22306
2 99602 1 22306
2 99603 1 22328
2 99604 1 22328
2 99605 1 22337
2 99606 1 22337
2 99607 1 22345
2 99608 1 22345
2 99609 1 22352
2 99610 1 22352
2 99611 1 22354
2 99612 1 22354
2 99613 1 22355
2 99614 1 22355
2 99615 1 22355
2 99616 1 22367
2 99617 1 22367
2 99618 1 22367
2 99619 1 22371
2 99620 1 22371
2 99621 1 22371
2 99622 1 22372
2 99623 1 22372
2 99624 1 22372
2 99625 1 22373
2 99626 1 22373
2 99627 1 22382
2 99628 1 22382
2 99629 1 22382
2 99630 1 22382
2 99631 1 22382
2 99632 1 22382
2 99633 1 22382
2 99634 1 22382
2 99635 1 22382
2 99636 1 22384
2 99637 1 22384
2 99638 1 22384
2 99639 1 22384
2 99640 1 22384
2 99641 1 22386
2 99642 1 22386
2 99643 1 22386
2 99644 1 22386
2 99645 1 22386
2 99646 1 22386
2 99647 1 22386
2 99648 1 22386
2 99649 1 22386
2 99650 1 22386
2 99651 1 22386
2 99652 1 22386
2 99653 1 22386
2 99654 1 22386
2 99655 1 22386
2 99656 1 22386
2 99657 1 22386
2 99658 1 22386
2 99659 1 22386
2 99660 1 22386
2 99661 1 22386
2 99662 1 22386
2 99663 1 22386
2 99664 1 22390
2 99665 1 22390
2 99666 1 22400
2 99667 1 22400
2 99668 1 22400
2 99669 1 22401
2 99670 1 22401
2 99671 1 22401
2 99672 1 22401
2 99673 1 22401
2 99674 1 22401
2 99675 1 22401
2 99676 1 22401
2 99677 1 22401
2 99678 1 22403
2 99679 1 22403
2 99680 1 22403
2 99681 1 22408
2 99682 1 22408
2 99683 1 22408
2 99684 1 22408
2 99685 1 22408
2 99686 1 22408
2 99687 1 22422
2 99688 1 22422
2 99689 1 22422
2 99690 1 22429
2 99691 1 22429
2 99692 1 22429
2 99693 1 22429
2 99694 1 22429
2 99695 1 22429
2 99696 1 22429
2 99697 1 22442
2 99698 1 22442
2 99699 1 22442
2 99700 1 22442
2 99701 1 22443
2 99702 1 22443
2 99703 1 22461
2 99704 1 22461
2 99705 1 22461
2 99706 1 22462
2 99707 1 22462
2 99708 1 22465
2 99709 1 22465
2 99710 1 22472
2 99711 1 22472
2 99712 1 22472
2 99713 1 22472
2 99714 1 22472
2 99715 1 22473
2 99716 1 22473
2 99717 1 22476
2 99718 1 22476
2 99719 1 22476
2 99720 1 22477
2 99721 1 22477
2 99722 1 22486
2 99723 1 22486
2 99724 1 22509
2 99725 1 22509
2 99726 1 22509
2 99727 1 22516
2 99728 1 22516
2 99729 1 22516
2 99730 1 22524
2 99731 1 22524
2 99732 1 22524
2 99733 1 22525
2 99734 1 22525
2 99735 1 22526
2 99736 1 22526
2 99737 1 22528
2 99738 1 22528
2 99739 1 22531
2 99740 1 22531
2 99741 1 22538
2 99742 1 22538
2 99743 1 22538
2 99744 1 22538
2 99745 1 22538
2 99746 1 22544
2 99747 1 22544
2 99748 1 22544
2 99749 1 22563
2 99750 1 22563
2 99751 1 22563
2 99752 1 22563
2 99753 1 22563
2 99754 1 22563
2 99755 1 22563
2 99756 1 22563
2 99757 1 22563
2 99758 1 22563
2 99759 1 22563
2 99760 1 22564
2 99761 1 22564
2 99762 1 22565
2 99763 1 22565
2 99764 1 22569
2 99765 1 22569
2 99766 1 22578
2 99767 1 22578
2 99768 1 22578
2 99769 1 22587
2 99770 1 22587
2 99771 1 22587
2 99772 1 22587
2 99773 1 22596
2 99774 1 22596
2 99775 1 22596
2 99776 1 22596
2 99777 1 22596
2 99778 1 22596
2 99779 1 22596
2 99780 1 22596
2 99781 1 22626
2 99782 1 22626
2 99783 1 22626
2 99784 1 22637
2 99785 1 22637
2 99786 1 22640
2 99787 1 22640
2 99788 1 22644
2 99789 1 22644
2 99790 1 22644
2 99791 1 22649
2 99792 1 22649
2 99793 1 22657
2 99794 1 22657
2 99795 1 22657
2 99796 1 22657
2 99797 1 22657
2 99798 1 22657
2 99799 1 22657
2 99800 1 22659
2 99801 1 22659
2 99802 1 22659
2 99803 1 22660
2 99804 1 22660
2 99805 1 22660
2 99806 1 22661
2 99807 1 22661
2 99808 1 22661
2 99809 1 22661
2 99810 1 22661
2 99811 1 22661
2 99812 1 22661
2 99813 1 22661
2 99814 1 22668
2 99815 1 22668
2 99816 1 22668
2 99817 1 22668
2 99818 1 22669
2 99819 1 22669
2 99820 1 22670
2 99821 1 22670
2 99822 1 22670
2 99823 1 22671
2 99824 1 22671
2 99825 1 22671
2 99826 1 22692
2 99827 1 22692
2 99828 1 22695
2 99829 1 22695
2 99830 1 22695
2 99831 1 22695
2 99832 1 22702
2 99833 1 22702
2 99834 1 22702
2 99835 1 22712
2 99836 1 22712
2 99837 1 22715
2 99838 1 22715
2 99839 1 22731
2 99840 1 22731
2 99841 1 22731
2 99842 1 22732
2 99843 1 22732
2 99844 1 22742
2 99845 1 22742
2 99846 1 22758
2 99847 1 22758
2 99848 1 22758
2 99849 1 22758
2 99850 1 22758
2 99851 1 22758
2 99852 1 22759
2 99853 1 22759
2 99854 1 22759
2 99855 1 22760
2 99856 1 22760
2 99857 1 22761
2 99858 1 22761
2 99859 1 22761
2 99860 1 22761
2 99861 1 22761
2 99862 1 22761
2 99863 1 22761
2 99864 1 22761
2 99865 1 22761
2 99866 1 22761
2 99867 1 22761
2 99868 1 22764
2 99869 1 22764
2 99870 1 22764
2 99871 1 22773
2 99872 1 22773
2 99873 1 22774
2 99874 1 22774
2 99875 1 22774
2 99876 1 22774
2 99877 1 22777
2 99878 1 22777
2 99879 1 22777
2 99880 1 22778
2 99881 1 22778
2 99882 1 22779
2 99883 1 22779
2 99884 1 22801
2 99885 1 22801
2 99886 1 22805
2 99887 1 22805
2 99888 1 22805
2 99889 1 22832
2 99890 1 22832
2 99891 1 22834
2 99892 1 22834
2 99893 1 22836
2 99894 1 22836
2 99895 1 22841
2 99896 1 22841
2 99897 1 22845
2 99898 1 22845
2 99899 1 22859
2 99900 1 22859
2 99901 1 22870
2 99902 1 22870
2 99903 1 22873
2 99904 1 22873
2 99905 1 22873
2 99906 1 22874
2 99907 1 22874
2 99908 1 22890
2 99909 1 22890
2 99910 1 22896
2 99911 1 22896
2 99912 1 22911
2 99913 1 22911
2 99914 1 22923
2 99915 1 22923
2 99916 1 22931
2 99917 1 22931
2 99918 1 22931
2 99919 1 22931
2 99920 1 22933
2 99921 1 22933
2 99922 1 22953
2 99923 1 22953
2 99924 1 22956
2 99925 1 22956
2 99926 1 22956
2 99927 1 22956
2 99928 1 22956
2 99929 1 22956
2 99930 1 22956
2 99931 1 22957
2 99932 1 22957
2 99933 1 22957
2 99934 1 22957
2 99935 1 22957
2 99936 1 22957
2 99937 1 22966
2 99938 1 22966
2 99939 1 22967
2 99940 1 22967
2 99941 1 22979
2 99942 1 22979
2 99943 1 22993
2 99944 1 22993
2 99945 1 22993
2 99946 1 22993
2 99947 1 23008
2 99948 1 23008
2 99949 1 23008
2 99950 1 23008
2 99951 1 23009
2 99952 1 23009
2 99953 1 23011
2 99954 1 23011
2 99955 1 23011
2 99956 1 23011
2 99957 1 23011
2 99958 1 23011
2 99959 1 23011
2 99960 1 23011
2 99961 1 23011
2 99962 1 23011
2 99963 1 23011
2 99964 1 23011
2 99965 1 23011
2 99966 1 23025
2 99967 1 23025
2 99968 1 23025
2 99969 1 23025
2 99970 1 23025
2 99971 1 23025
2 99972 1 23025
2 99973 1 23025
2 99974 1 23025
2 99975 1 23025
2 99976 1 23026
2 99977 1 23026
2 99978 1 23047
2 99979 1 23047
2 99980 1 23062
2 99981 1 23062
2 99982 1 23068
2 99983 1 23068
2 99984 1 23076
2 99985 1 23076
2 99986 1 23076
2 99987 1 23076
2 99988 1 23092
2 99989 1 23092
2 99990 1 23098
2 99991 1 23098
2 99992 1 23109
2 99993 1 23109
2 99994 1 23109
2 99995 1 23112
2 99996 1 23112
2 99997 1 23112
2 99998 1 23112
2 99999 1 23112
2 100000 1 23125
2 100001 1 23125
2 100002 1 23140
2 100003 1 23140
2 100004 1 23140
2 100005 1 23140
2 100006 1 23141
2 100007 1 23141
2 100008 1 23141
2 100009 1 23143
2 100010 1 23143
2 100011 1 23145
2 100012 1 23145
2 100013 1 23151
2 100014 1 23151
2 100015 1 23173
2 100016 1 23173
2 100017 1 23182
2 100018 1 23182
2 100019 1 23182
2 100020 1 23182
2 100021 1 23182
2 100022 1 23182
2 100023 1 23182
2 100024 1 23182
2 100025 1 23182
2 100026 1 23182
2 100027 1 23182
2 100028 1 23182
2 100029 1 23182
2 100030 1 23182
2 100031 1 23182
2 100032 1 23182
2 100033 1 23182
2 100034 1 23191
2 100035 1 23191
2 100036 1 23192
2 100037 1 23192
2 100038 1 23199
2 100039 1 23199
2 100040 1 23199
2 100041 1 23219
2 100042 1 23219
2 100043 1 23219
2 100044 1 23219
2 100045 1 23219
2 100046 1 23219
2 100047 1 23219
2 100048 1 23219
2 100049 1 23229
2 100050 1 23229
2 100051 1 23231
2 100052 1 23231
2 100053 1 23232
2 100054 1 23232
2 100055 1 23233
2 100056 1 23233
2 100057 1 23233
2 100058 1 23233
2 100059 1 23250
2 100060 1 23250
2 100061 1 23250
2 100062 1 23251
2 100063 1 23251
2 100064 1 23263
2 100065 1 23263
2 100066 1 23271
2 100067 1 23271
2 100068 1 23298
2 100069 1 23298
2 100070 1 23300
2 100071 1 23300
2 100072 1 23313
2 100073 1 23313
2 100074 1 23313
2 100075 1 23347
2 100076 1 23347
2 100077 1 23347
2 100078 1 23347
2 100079 1 23347
2 100080 1 23347
2 100081 1 23347
2 100082 1 23347
2 100083 1 23347
2 100084 1 23347
2 100085 1 23347
2 100086 1 23347
2 100087 1 23347
2 100088 1 23347
2 100089 1 23347
2 100090 1 23348
2 100091 1 23348
2 100092 1 23348
2 100093 1 23348
2 100094 1 23350
2 100095 1 23350
2 100096 1 23354
2 100097 1 23354
2 100098 1 23355
2 100099 1 23355
2 100100 1 23355
2 100101 1 23358
2 100102 1 23358
2 100103 1 23358
2 100104 1 23358
2 100105 1 23358
2 100106 1 23359
2 100107 1 23359
2 100108 1 23366
2 100109 1 23366
2 100110 1 23366
2 100111 1 23366
2 100112 1 23366
2 100113 1 23366
2 100114 1 23367
2 100115 1 23367
2 100116 1 23367
2 100117 1 23371
2 100118 1 23371
2 100119 1 23371
2 100120 1 23371
2 100121 1 23380
2 100122 1 23380
2 100123 1 23380
2 100124 1 23380
2 100125 1 23381
2 100126 1 23381
2 100127 1 23392
2 100128 1 23392
2 100129 1 23395
2 100130 1 23395
2 100131 1 23396
2 100132 1 23396
2 100133 1 23418
2 100134 1 23418
2 100135 1 23419
2 100136 1 23419
2 100137 1 23419
2 100138 1 23419
2 100139 1 23419
2 100140 1 23419
2 100141 1 23419
2 100142 1 23419
2 100143 1 23419
2 100144 1 23419
2 100145 1 23419
2 100146 1 23419
2 100147 1 23419
2 100148 1 23420
2 100149 1 23420
2 100150 1 23420
2 100151 1 23430
2 100152 1 23430
2 100153 1 23430
2 100154 1 23430
2 100155 1 23430
2 100156 1 23430
2 100157 1 23430
2 100158 1 23432
2 100159 1 23432
2 100160 1 23433
2 100161 1 23433
2 100162 1 23434
2 100163 1 23434
2 100164 1 23434
2 100165 1 23434
2 100166 1 23434
2 100167 1 23434
2 100168 1 23444
2 100169 1 23444
2 100170 1 23444
2 100171 1 23444
2 100172 1 23444
2 100173 1 23444
2 100174 1 23444
2 100175 1 23444
2 100176 1 23444
2 100177 1 23444
2 100178 1 23444
2 100179 1 23444
2 100180 1 23444
2 100181 1 23444
2 100182 1 23444
2 100183 1 23444
2 100184 1 23444
2 100185 1 23444
2 100186 1 23444
2 100187 1 23444
2 100188 1 23444
2 100189 1 23444
2 100190 1 23444
2 100191 1 23444
2 100192 1 23444
2 100193 1 23444
2 100194 1 23444
2 100195 1 23444
2 100196 1 23444
2 100197 1 23444
2 100198 1 23444
2 100199 1 23444
2 100200 1 23444
2 100201 1 23444
2 100202 1 23444
2 100203 1 23444
2 100204 1 23444
2 100205 1 23444
2 100206 1 23444
2 100207 1 23444
2 100208 1 23444
2 100209 1 23444
2 100210 1 23444
2 100211 1 23444
2 100212 1 23444
2 100213 1 23444
2 100214 1 23444
2 100215 1 23444
2 100216 1 23444
2 100217 1 23444
2 100218 1 23444
2 100219 1 23444
2 100220 1 23444
2 100221 1 23444
2 100222 1 23445
2 100223 1 23445
2 100224 1 23445
2 100225 1 23445
2 100226 1 23450
2 100227 1 23450
2 100228 1 23457
2 100229 1 23457
2 100230 1 23470
2 100231 1 23470
2 100232 1 23470
2 100233 1 23470
2 100234 1 23470
2 100235 1 23470
2 100236 1 23471
2 100237 1 23471
2 100238 1 23471
2 100239 1 23473
2 100240 1 23473
2 100241 1 23474
2 100242 1 23474
2 100243 1 23474
2 100244 1 23474
2 100245 1 23475
2 100246 1 23475
2 100247 1 23484
2 100248 1 23484
2 100249 1 23484
2 100250 1 23487
2 100251 1 23487
2 100252 1 23487
2 100253 1 23487
2 100254 1 23487
2 100255 1 23490
2 100256 1 23490
2 100257 1 23490
2 100258 1 23491
2 100259 1 23491
2 100260 1 23495
2 100261 1 23495
2 100262 1 23495
2 100263 1 23495
2 100264 1 23495
2 100265 1 23495
2 100266 1 23495
2 100267 1 23495
2 100268 1 23495
2 100269 1 23495
2 100270 1 23495
2 100271 1 23495
2 100272 1 23495
2 100273 1 23495
2 100274 1 23495
2 100275 1 23495
2 100276 1 23495
2 100277 1 23495
2 100278 1 23495
2 100279 1 23495
2 100280 1 23495
2 100281 1 23495
2 100282 1 23495
2 100283 1 23495
2 100284 1 23495
2 100285 1 23495
2 100286 1 23495
2 100287 1 23495
2 100288 1 23495
2 100289 1 23495
2 100290 1 23495
2 100291 1 23495
2 100292 1 23495
2 100293 1 23503
2 100294 1 23503
2 100295 1 23503
2 100296 1 23503
2 100297 1 23503
2 100298 1 23503
2 100299 1 23503
2 100300 1 23514
2 100301 1 23514
2 100302 1 23514
2 100303 1 23514
2 100304 1 23514
2 100305 1 23523
2 100306 1 23523
2 100307 1 23523
2 100308 1 23526
2 100309 1 23526
2 100310 1 23527
2 100311 1 23527
2 100312 1 23528
2 100313 1 23528
2 100314 1 23528
2 100315 1 23529
2 100316 1 23529
2 100317 1 23529
2 100318 1 23533
2 100319 1 23533
2 100320 1 23533
2 100321 1 23543
2 100322 1 23543
2 100323 1 23544
2 100324 1 23544
2 100325 1 23545
2 100326 1 23545
2 100327 1 23547
2 100328 1 23547
2 100329 1 23547
2 100330 1 23547
2 100331 1 23551
2 100332 1 23551
2 100333 1 23552
2 100334 1 23552
2 100335 1 23553
2 100336 1 23553
2 100337 1 23553
2 100338 1 23553
2 100339 1 23554
2 100340 1 23554
2 100341 1 23554
2 100342 1 23554
2 100343 1 23554
2 100344 1 23554
2 100345 1 23554
2 100346 1 23554
2 100347 1 23554
2 100348 1 23555
2 100349 1 23555
2 100350 1 23555
2 100351 1 23555
2 100352 1 23566
2 100353 1 23566
2 100354 1 23583
2 100355 1 23583
2 100356 1 23591
2 100357 1 23591
2 100358 1 23592
2 100359 1 23592
2 100360 1 23598
2 100361 1 23598
2 100362 1 23599
2 100363 1 23599
2 100364 1 23599
2 100365 1 23608
2 100366 1 23608
2 100367 1 23609
2 100368 1 23609
2 100369 1 23609
2 100370 1 23627
2 100371 1 23627
2 100372 1 23628
2 100373 1 23628
2 100374 1 23628
2 100375 1 23642
2 100376 1 23642
2 100377 1 23650
2 100378 1 23650
2 100379 1 23650
2 100380 1 23650
2 100381 1 23650
2 100382 1 23650
2 100383 1 23650
2 100384 1 23650
2 100385 1 23651
2 100386 1 23651
2 100387 1 23651
2 100388 1 23651
2 100389 1 23652
2 100390 1 23652
2 100391 1 23652
2 100392 1 23666
2 100393 1 23666
2 100394 1 23666
2 100395 1 23666
2 100396 1 23666
2 100397 1 23666
2 100398 1 23667
2 100399 1 23667
2 100400 1 23670
2 100401 1 23670
2 100402 1 23670
2 100403 1 23670
2 100404 1 23670
2 100405 1 23672
2 100406 1 23672
2 100407 1 23672
2 100408 1 23681
2 100409 1 23681
2 100410 1 23681
2 100411 1 23696
2 100412 1 23696
2 100413 1 23697
2 100414 1 23697
2 100415 1 23698
2 100416 1 23698
2 100417 1 23698
2 100418 1 23698
2 100419 1 23698
2 100420 1 23698
2 100421 1 23707
2 100422 1 23707
2 100423 1 23707
2 100424 1 23707
2 100425 1 23707
2 100426 1 23707
2 100427 1 23707
2 100428 1 23707
2 100429 1 23707
2 100430 1 23707
2 100431 1 23707
2 100432 1 23707
2 100433 1 23707
2 100434 1 23707
2 100435 1 23707
2 100436 1 23707
2 100437 1 23707
2 100438 1 23707
2 100439 1 23707
2 100440 1 23707
2 100441 1 23707
2 100442 1 23707
2 100443 1 23711
2 100444 1 23711
2 100445 1 23720
2 100446 1 23720
2 100447 1 23720
2 100448 1 23720
2 100449 1 23720
2 100450 1 23724
2 100451 1 23724
2 100452 1 23724
2 100453 1 23735
2 100454 1 23735
2 100455 1 23736
2 100456 1 23736
2 100457 1 23736
2 100458 1 23738
2 100459 1 23738
2 100460 1 23748
2 100461 1 23748
2 100462 1 23755
2 100463 1 23755
2 100464 1 23756
2 100465 1 23756
2 100466 1 23777
2 100467 1 23777
2 100468 1 23778
2 100469 1 23778
2 100470 1 23795
2 100471 1 23795
2 100472 1 23795
2 100473 1 23795
2 100474 1 23795
2 100475 1 23797
2 100476 1 23797
2 100477 1 23805
2 100478 1 23805
2 100479 1 23810
2 100480 1 23810
2 100481 1 23810
2 100482 1 23810
2 100483 1 23845
2 100484 1 23845
2 100485 1 23853
2 100486 1 23853
2 100487 1 23862
2 100488 1 23862
2 100489 1 23862
2 100490 1 23883
2 100491 1 23883
2 100492 1 23899
2 100493 1 23899
2 100494 1 23899
2 100495 1 23899
2 100496 1 23906
2 100497 1 23906
2 100498 1 23906
2 100499 1 23906
2 100500 1 23906
2 100501 1 23906
2 100502 1 23906
2 100503 1 23906
2 100504 1 23906
2 100505 1 23906
2 100506 1 23907
2 100507 1 23907
2 100508 1 23907
2 100509 1 23908
2 100510 1 23908
2 100511 1 23909
2 100512 1 23909
2 100513 1 23909
2 100514 1 23909
2 100515 1 23909
2 100516 1 23909
2 100517 1 23909
2 100518 1 23909
2 100519 1 23909
2 100520 1 23909
2 100521 1 23909
2 100522 1 23909
2 100523 1 23909
2 100524 1 23909
2 100525 1 23910
2 100526 1 23910
2 100527 1 23910
2 100528 1 23910
2 100529 1 23910
2 100530 1 23910
2 100531 1 23910
2 100532 1 23910
2 100533 1 23913
2 100534 1 23913
2 100535 1 23916
2 100536 1 23916
2 100537 1 23925
2 100538 1 23925
2 100539 1 23936
2 100540 1 23936
2 100541 1 23936
2 100542 1 23936
2 100543 1 23936
2 100544 1 23936
2 100545 1 23961
2 100546 1 23961
2 100547 1 23961
2 100548 1 23962
2 100549 1 23962
2 100550 1 23963
2 100551 1 23963
2 100552 1 23968
2 100553 1 23968
2 100554 1 23975
2 100555 1 23975
2 100556 1 23983
2 100557 1 23983
2 100558 1 23984
2 100559 1 23984
2 100560 1 23984
2 100561 1 23986
2 100562 1 23986
2 100563 1 23994
2 100564 1 23994
2 100565 1 23994
2 100566 1 24017
2 100567 1 24017
2 100568 1 24017
2 100569 1 24018
2 100570 1 24018
2 100571 1 24034
2 100572 1 24034
2 100573 1 24048
2 100574 1 24048
2 100575 1 24048
2 100576 1 24048
2 100577 1 24048
2 100578 1 24048
2 100579 1 24048
2 100580 1 24048
2 100581 1 24048
2 100582 1 24048
2 100583 1 24048
2 100584 1 24048
2 100585 1 24051
2 100586 1 24051
2 100587 1 24059
2 100588 1 24059
2 100589 1 24061
2 100590 1 24061
2 100591 1 24062
2 100592 1 24062
2 100593 1 24063
2 100594 1 24063
2 100595 1 24063
2 100596 1 24064
2 100597 1 24064
2 100598 1 24064
2 100599 1 24065
2 100600 1 24065
2 100601 1 24065
2 100602 1 24065
2 100603 1 24065
2 100604 1 24073
2 100605 1 24073
2 100606 1 24080
2 100607 1 24080
2 100608 1 24081
2 100609 1 24081
2 100610 1 24104
2 100611 1 24104
2 100612 1 24112
2 100613 1 24112
2 100614 1 24117
2 100615 1 24117
2 100616 1 24117
2 100617 1 24118
2 100618 1 24118
2 100619 1 24131
2 100620 1 24131
2 100621 1 24132
2 100622 1 24132
2 100623 1 24156
2 100624 1 24156
2 100625 1 24160
2 100626 1 24160
2 100627 1 24168
2 100628 1 24168
2 100629 1 24168
2 100630 1 24168
2 100631 1 24168
2 100632 1 24173
2 100633 1 24173
2 100634 1 24173
2 100635 1 24174
2 100636 1 24174
2 100637 1 24174
2 100638 1 24174
2 100639 1 24174
2 100640 1 24174
2 100641 1 24174
2 100642 1 24174
2 100643 1 24175
2 100644 1 24175
2 100645 1 24175
2 100646 1 24175
2 100647 1 24189
2 100648 1 24189
2 100649 1 24218
2 100650 1 24218
2 100651 1 24218
2 100652 1 24218
2 100653 1 24218
2 100654 1 24228
2 100655 1 24228
2 100656 1 24243
2 100657 1 24243
2 100658 1 24243
2 100659 1 24259
2 100660 1 24259
2 100661 1 24259
2 100662 1 24259
2 100663 1 24259
2 100664 1 24260
2 100665 1 24260
2 100666 1 24277
2 100667 1 24277
2 100668 1 24285
2 100669 1 24285
2 100670 1 24285
2 100671 1 24285
2 100672 1 24285
2 100673 1 24285
2 100674 1 24286
2 100675 1 24286
2 100676 1 24287
2 100677 1 24287
2 100678 1 24294
2 100679 1 24294
2 100680 1 24294
2 100681 1 24294
2 100682 1 24316
2 100683 1 24316
2 100684 1 24316
2 100685 1 24329
2 100686 1 24329
2 100687 1 24330
2 100688 1 24330
2 100689 1 24341
2 100690 1 24341
2 100691 1 24346
2 100692 1 24346
2 100693 1 24352
2 100694 1 24352
2 100695 1 24362
2 100696 1 24362
2 100697 1 24431
2 100698 1 24431
2 100699 1 24473
2 100700 1 24473
2 100701 1 24473
2 100702 1 24473
2 100703 1 24473
2 100704 1 24474
2 100705 1 24474
2 100706 1 24490
2 100707 1 24490
2 100708 1 24495
2 100709 1 24495
2 100710 1 24495
2 100711 1 24500
2 100712 1 24500
2 100713 1 24510
2 100714 1 24510
2 100715 1 24533
2 100716 1 24533
2 100717 1 24547
2 100718 1 24547
2 100719 1 24555
2 100720 1 24555
2 100721 1 24595
2 100722 1 24595
2 100723 1 24599
2 100724 1 24599
2 100725 1 24613
2 100726 1 24613
2 100727 1 24613
2 100728 1 24652
2 100729 1 24652
2 100730 1 24652
2 100731 1 24652
2 100732 1 24660
2 100733 1 24660
2 100734 1 24660
2 100735 1 24661
2 100736 1 24661
2 100737 1 24661
2 100738 1 24661
2 100739 1 24661
2 100740 1 24661
2 100741 1 24661
2 100742 1 24669
2 100743 1 24669
2 100744 1 24676
2 100745 1 24676
2 100746 1 24677
2 100747 1 24677
2 100748 1 24679
2 100749 1 24679
2 100750 1 24719
2 100751 1 24719
2 100752 1 24719
2 100753 1 24719
2 100754 1 24719
2 100755 1 24719
2 100756 1 24720
2 100757 1 24720
2 100758 1 24720
2 100759 1 24721
2 100760 1 24721
2 100761 1 24721
2 100762 1 24745
2 100763 1 24745
2 100764 1 24745
2 100765 1 24745
2 100766 1 24745
2 100767 1 24746
2 100768 1 24746
2 100769 1 24746
2 100770 1 24749
2 100771 1 24749
2 100772 1 24749
2 100773 1 24749
2 100774 1 24752
2 100775 1 24752
2 100776 1 24761
2 100777 1 24761
2 100778 1 24761
2 100779 1 24762
2 100780 1 24762
2 100781 1 24763
2 100782 1 24763
2 100783 1 24763
2 100784 1 24766
2 100785 1 24766
2 100786 1 24778
2 100787 1 24778
2 100788 1 24778
2 100789 1 24778
2 100790 1 24778
2 100791 1 24796
2 100792 1 24796
2 100793 1 24796
2 100794 1 24832
2 100795 1 24832
2 100796 1 24850
2 100797 1 24850
2 100798 1 24850
2 100799 1 24854
2 100800 1 24854
2 100801 1 24854
2 100802 1 24854
2 100803 1 24854
2 100804 1 24872
2 100805 1 24872
2 100806 1 24872
2 100807 1 24872
2 100808 1 24872
2 100809 1 24872
2 100810 1 24872
2 100811 1 24872
2 100812 1 24872
2 100813 1 24872
2 100814 1 24872
2 100815 1 24874
2 100816 1 24874
2 100817 1 24881
2 100818 1 24881
2 100819 1 24905
2 100820 1 24905
2 100821 1 24905
2 100822 1 24907
2 100823 1 24907
2 100824 1 24907
2 100825 1 24918
2 100826 1 24918
2 100827 1 24932
2 100828 1 24932
2 100829 1 24932
2 100830 1 24938
2 100831 1 24938
2 100832 1 24967
2 100833 1 24967
2 100834 1 24974
2 100835 1 24974
2 100836 1 25020
2 100837 1 25020
2 100838 1 25022
2 100839 1 25022
2 100840 1 25022
2 100841 1 25022
2 100842 1 25022
2 100843 1 25023
2 100844 1 25023
2 100845 1 25023
2 100846 1 25023
2 100847 1 25025
2 100848 1 25025
2 100849 1 25025
2 100850 1 25029
2 100851 1 25029
2 100852 1 25042
2 100853 1 25042
2 100854 1 25046
2 100855 1 25046
2 100856 1 25053
2 100857 1 25053
2 100858 1 25053
2 100859 1 25054
2 100860 1 25054
2 100861 1 25054
2 100862 1 25129
2 100863 1 25129
2 100864 1 25139
2 100865 1 25139
2 100866 1 25164
2 100867 1 25164
2 100868 1 25181
2 100869 1 25181
2 100870 1 25181
2 100871 1 25181
2 100872 1 25184
2 100873 1 25184
2 100874 1 25217
2 100875 1 25217
2 100876 1 25233
2 100877 1 25233
2 100878 1 25233
2 100879 1 25233
2 100880 1 25233
2 100881 1 25234
2 100882 1 25234
2 100883 1 25265
2 100884 1 25265
2 100885 1 25271
2 100886 1 25271
2 100887 1 25272
2 100888 1 25272
2 100889 1 25279
2 100890 1 25279
2 100891 1 25279
2 100892 1 25292
2 100893 1 25292
2 100894 1 25300
2 100895 1 25300
2 100896 1 25314
2 100897 1 25314
2 100898 1 25344
2 100899 1 25344
2 100900 1 25347
2 100901 1 25347
2 100902 1 25380
2 100903 1 25380
2 100904 1 25380
2 100905 1 25380
2 100906 1 25381
2 100907 1 25381
2 100908 1 25381
2 100909 1 25381
2 100910 1 25381
2 100911 1 25381
2 100912 1 25381
2 100913 1 25394
2 100914 1 25394
2 100915 1 25394
2 100916 1 25395
2 100917 1 25395
2 100918 1 25396
2 100919 1 25396
2 100920 1 25426
2 100921 1 25426
2 100922 1 25428
2 100923 1 25428
2 100924 1 25431
2 100925 1 25431
2 100926 1 25433
2 100927 1 25433
2 100928 1 25434
2 100929 1 25434
2 100930 1 25444
2 100931 1 25444
2 100932 1 25444
2 100933 1 25444
2 100934 1 25447
2 100935 1 25447
2 100936 1 25460
2 100937 1 25460
2 100938 1 25463
2 100939 1 25463
2 100940 1 25489
2 100941 1 25489
2 100942 1 25489
2 100943 1 25490
2 100944 1 25490
2 100945 1 25490
2 100946 1 25504
2 100947 1 25504
2 100948 1 25504
2 100949 1 25505
2 100950 1 25505
2 100951 1 25506
2 100952 1 25506
2 100953 1 25506
2 100954 1 25506
2 100955 1 25506
2 100956 1 25516
2 100957 1 25516
2 100958 1 25517
2 100959 1 25517
2 100960 1 25517
2 100961 1 25517
2 100962 1 25518
2 100963 1 25518
2 100964 1 25518
2 100965 1 25518
2 100966 1 25529
2 100967 1 25529
2 100968 1 25529
2 100969 1 25539
2 100970 1 25539
2 100971 1 25539
2 100972 1 25540
2 100973 1 25540
2 100974 1 25549
2 100975 1 25549
2 100976 1 25549
2 100977 1 25550
2 100978 1 25550
2 100979 1 25561
2 100980 1 25561
2 100981 1 25561
2 100982 1 25581
2 100983 1 25581
2 100984 1 25581
2 100985 1 25582
2 100986 1 25582
2 100987 1 25582
2 100988 1 25582
2 100989 1 25596
2 100990 1 25596
2 100991 1 25598
2 100992 1 25598
2 100993 1 25598
2 100994 1 25598
2 100995 1 25599
2 100996 1 25599
2 100997 1 25599
2 100998 1 25602
2 100999 1 25602
2 101000 1 25602
2 101001 1 25602
2 101002 1 25619
2 101003 1 25619
2 101004 1 25619
2 101005 1 25619
2 101006 1 25619
2 101007 1 25619
2 101008 1 25619
2 101009 1 25619
2 101010 1 25619
2 101011 1 25619
2 101012 1 25630
2 101013 1 25630
2 101014 1 25630
2 101015 1 25630
2 101016 1 25630
2 101017 1 25630
2 101018 1 25630
2 101019 1 25630
2 101020 1 25630
2 101021 1 25630
2 101022 1 25630
2 101023 1 25630
2 101024 1 25630
2 101025 1 25630
2 101026 1 25630
2 101027 1 25630
2 101028 1 25630
2 101029 1 25630
2 101030 1 25636
2 101031 1 25636
2 101032 1 25639
2 101033 1 25639
2 101034 1 25639
2 101035 1 25652
2 101036 1 25652
2 101037 1 25652
2 101038 1 25652
2 101039 1 25652
2 101040 1 25660
2 101041 1 25660
2 101042 1 25660
2 101043 1 25660
2 101044 1 25660
2 101045 1 25662
2 101046 1 25662
2 101047 1 25662
2 101048 1 25663
2 101049 1 25663
2 101050 1 25663
2 101051 1 25668
2 101052 1 25668
2 101053 1 25668
2 101054 1 25668
2 101055 1 25668
2 101056 1 25668
2 101057 1 25668
2 101058 1 25668
2 101059 1 25668
2 101060 1 25676
2 101061 1 25676
2 101062 1 25676
2 101063 1 25677
2 101064 1 25677
2 101065 1 25679
2 101066 1 25679
2 101067 1 25679
2 101068 1 25693
2 101069 1 25693
2 101070 1 25696
2 101071 1 25696
2 101072 1 25696
2 101073 1 25696
2 101074 1 25698
2 101075 1 25698
2 101076 1 25698
2 101077 1 25698
2 101078 1 25698
2 101079 1 25698
2 101080 1 25707
2 101081 1 25707
2 101082 1 25711
2 101083 1 25711
2 101084 1 25711
2 101085 1 25712
2 101086 1 25712
2 101087 1 25712
2 101088 1 25714
2 101089 1 25714
2 101090 1 25724
2 101091 1 25724
2 101092 1 25727
2 101093 1 25727
2 101094 1 25727
2 101095 1 25727
2 101096 1 25727
2 101097 1 25727
2 101098 1 25747
2 101099 1 25747
2 101100 1 25748
2 101101 1 25748
2 101102 1 25748
2 101103 1 25748
2 101104 1 25748
2 101105 1 25755
2 101106 1 25755
2 101107 1 25757
2 101108 1 25757
2 101109 1 25764
2 101110 1 25764
2 101111 1 25774
2 101112 1 25774
2 101113 1 25788
2 101114 1 25788
2 101115 1 25800
2 101116 1 25800
2 101117 1 25806
2 101118 1 25806
2 101119 1 25806
2 101120 1 25807
2 101121 1 25807
2 101122 1 25807
2 101123 1 25807
2 101124 1 25807
2 101125 1 25807
2 101126 1 25807
2 101127 1 25807
2 101128 1 25807
2 101129 1 25807
2 101130 1 25807
2 101131 1 25807
2 101132 1 25807
2 101133 1 25807
2 101134 1 25807
2 101135 1 25808
2 101136 1 25808
2 101137 1 25809
2 101138 1 25809
2 101139 1 25809
2 101140 1 25812
2 101141 1 25812
2 101142 1 25812
2 101143 1 25812
2 101144 1 25812
2 101145 1 25812
2 101146 1 25812
2 101147 1 25812
2 101148 1 25812
2 101149 1 25812
2 101150 1 25812
2 101151 1 25812
2 101152 1 25815
2 101153 1 25815
2 101154 1 25816
2 101155 1 25816
2 101156 1 25816
2 101157 1 25816
2 101158 1 25818
2 101159 1 25818
2 101160 1 25822
2 101161 1 25822
2 101162 1 25829
2 101163 1 25829
2 101164 1 25829
2 101165 1 25829
2 101166 1 25875
2 101167 1 25875
2 101168 1 25875
2 101169 1 25875
2 101170 1 25875
2 101171 1 25875
2 101172 1 25880
2 101173 1 25880
2 101174 1 25880
2 101175 1 25881
2 101176 1 25881
2 101177 1 25891
2 101178 1 25891
2 101179 1 25891
2 101180 1 25892
2 101181 1 25892
2 101182 1 25892
2 101183 1 25899
2 101184 1 25899
2 101185 1 25930
2 101186 1 25930
2 101187 1 25931
2 101188 1 25931
2 101189 1 25931
2 101190 1 25934
2 101191 1 25934
2 101192 1 25974
2 101193 1 25974
2 101194 1 25974
2 101195 1 25974
2 101196 1 25974
2 101197 1 25974
2 101198 1 25974
2 101199 1 25974
2 101200 1 25974
2 101201 1 25974
2 101202 1 25975
2 101203 1 25975
2 101204 1 25975
2 101205 1 25996
2 101206 1 25996
2 101207 1 25996
2 101208 1 25996
2 101209 1 26005
2 101210 1 26005
2 101211 1 26006
2 101212 1 26006
2 101213 1 26008
2 101214 1 26008
2 101215 1 26031
2 101216 1 26031
2 101217 1 26033
2 101218 1 26033
2 101219 1 26038
2 101220 1 26038
2 101221 1 26039
2 101222 1 26039
2 101223 1 26049
2 101224 1 26049
2 101225 1 26049
2 101226 1 26054
2 101227 1 26054
2 101228 1 26063
2 101229 1 26063
2 101230 1 26063
2 101231 1 26078
2 101232 1 26078
2 101233 1 26091
2 101234 1 26091
2 101235 1 26091
2 101236 1 26092
2 101237 1 26092
2 101238 1 26092
2 101239 1 26092
2 101240 1 26092
2 101241 1 26093
2 101242 1 26093
2 101243 1 26094
2 101244 1 26094
2 101245 1 26113
2 101246 1 26113
2 101247 1 26113
2 101248 1 26118
2 101249 1 26118
2 101250 1 26118
2 101251 1 26118
2 101252 1 26118
2 101253 1 26119
2 101254 1 26119
2 101255 1 26126
2 101256 1 26126
2 101257 1 26126
2 101258 1 26126
2 101259 1 26128
2 101260 1 26128
2 101261 1 26135
2 101262 1 26135
2 101263 1 26135
2 101264 1 26135
2 101265 1 26137
2 101266 1 26137
2 101267 1 26148
2 101268 1 26148
2 101269 1 26177
2 101270 1 26177
2 101271 1 26177
2 101272 1 26177
2 101273 1 26177
2 101274 1 26178
2 101275 1 26178
2 101276 1 26185
2 101277 1 26185
2 101278 1 26195
2 101279 1 26195
2 101280 1 26201
2 101281 1 26201
2 101282 1 26201
2 101283 1 26201
2 101284 1 26201
2 101285 1 26201
2 101286 1 26205
2 101287 1 26205
2 101288 1 26218
2 101289 1 26218
2 101290 1 26218
2 101291 1 26218
2 101292 1 26219
2 101293 1 26219
2 101294 1 26219
2 101295 1 26232
2 101296 1 26232
2 101297 1 26236
2 101298 1 26236
2 101299 1 26237
2 101300 1 26237
2 101301 1 26246
2 101302 1 26246
2 101303 1 26249
2 101304 1 26249
2 101305 1 26249
2 101306 1 26249
2 101307 1 26257
2 101308 1 26257
2 101309 1 26259
2 101310 1 26259
2 101311 1 26259
2 101312 1 26260
2 101313 1 26260
2 101314 1 26263
2 101315 1 26263
2 101316 1 26291
2 101317 1 26291
2 101318 1 26291
2 101319 1 26291
2 101320 1 26291
2 101321 1 26291
2 101322 1 26298
2 101323 1 26298
2 101324 1 26298
2 101325 1 26309
2 101326 1 26309
2 101327 1 26318
2 101328 1 26318
2 101329 1 26318
2 101330 1 26320
2 101331 1 26320
2 101332 1 26325
2 101333 1 26325
2 101334 1 26331
2 101335 1 26331
2 101336 1 26332
2 101337 1 26332
2 101338 1 26359
2 101339 1 26359
2 101340 1 26382
2 101341 1 26382
2 101342 1 26382
2 101343 1 26409
2 101344 1 26409
2 101345 1 26410
2 101346 1 26410
2 101347 1 26420
2 101348 1 26420
2 101349 1 26423
2 101350 1 26423
2 101351 1 26441
2 101352 1 26441
2 101353 1 26448
2 101354 1 26448
2 101355 1 26503
2 101356 1 26503
2 101357 1 26503
2 101358 1 26504
2 101359 1 26504
2 101360 1 26513
2 101361 1 26513
2 101362 1 26513
2 101363 1 26514
2 101364 1 26514
2 101365 1 26514
2 101366 1 26526
2 101367 1 26526
2 101368 1 26529
2 101369 1 26529
2 101370 1 26532
2 101371 1 26532
2 101372 1 26532
2 101373 1 26533
2 101374 1 26533
2 101375 1 26539
2 101376 1 26539
2 101377 1 26540
2 101378 1 26540
2 101379 1 26540
2 101380 1 26540
2 101381 1 26540
2 101382 1 26554
2 101383 1 26554
2 101384 1 26578
2 101385 1 26578
2 101386 1 26587
2 101387 1 26587
2 101388 1 26587
2 101389 1 26587
2 101390 1 26587
2 101391 1 26605
2 101392 1 26605
2 101393 1 26605
2 101394 1 26605
2 101395 1 26606
2 101396 1 26606
2 101397 1 26606
2 101398 1 26606
2 101399 1 26606
2 101400 1 26609
2 101401 1 26609
2 101402 1 26624
2 101403 1 26624
2 101404 1 26624
2 101405 1 26624
2 101406 1 26624
2 101407 1 26631
2 101408 1 26631
2 101409 1 26643
2 101410 1 26643
2 101411 1 26646
2 101412 1 26646
2 101413 1 26668
2 101414 1 26668
2 101415 1 26683
2 101416 1 26683
2 101417 1 26734
2 101418 1 26734
2 101419 1 26773
2 101420 1 26773
2 101421 1 26774
2 101422 1 26774
2 101423 1 26816
2 101424 1 26816
2 101425 1 26817
2 101426 1 26817
2 101427 1 26820
2 101428 1 26820
2 101429 1 26820
2 101430 1 26820
2 101431 1 26820
2 101432 1 26820
2 101433 1 26820
2 101434 1 26820
2 101435 1 26820
2 101436 1 26820
2 101437 1 26820
2 101438 1 26820
2 101439 1 26837
2 101440 1 26837
2 101441 1 26858
2 101442 1 26858
2 101443 1 26858
2 101444 1 26858
2 101445 1 26858
2 101446 1 26882
2 101447 1 26882
2 101448 1 26891
2 101449 1 26891
2 101450 1 26930
2 101451 1 26930
2 101452 1 26930
2 101453 1 26949
2 101454 1 26949
2 101455 1 26950
2 101456 1 26950
2 101457 1 26952
2 101458 1 26952
2 101459 1 26955
2 101460 1 26955
2 101461 1 26969
2 101462 1 26969
2 101463 1 26988
2 101464 1 26988
2 101465 1 26992
2 101466 1 26992
2 101467 1 26996
2 101468 1 26996
2 101469 1 27030
2 101470 1 27030
2 101471 1 27030
2 101472 1 27030
2 101473 1 27030
2 101474 1 27030
2 101475 1 27030
2 101476 1 27030
2 101477 1 27030
2 101478 1 27030
2 101479 1 27030
2 101480 1 27030
2 101481 1 27046
2 101482 1 27046
2 101483 1 27046
2 101484 1 27047
2 101485 1 27047
2 101486 1 27047
2 101487 1 27064
2 101488 1 27064
2 101489 1 27064
2 101490 1 27064
2 101491 1 27081
2 101492 1 27081
2 101493 1 27092
2 101494 1 27092
2 101495 1 27103
2 101496 1 27103
2 101497 1 27103
2 101498 1 27103
2 101499 1 27103
2 101500 1 27103
2 101501 1 27104
2 101502 1 27104
2 101503 1 27105
2 101504 1 27105
2 101505 1 27106
2 101506 1 27106
2 101507 1 27121
2 101508 1 27121
2 101509 1 27121
2 101510 1 27122
2 101511 1 27122
2 101512 1 27122
2 101513 1 27122
2 101514 1 27123
2 101515 1 27123
2 101516 1 27123
2 101517 1 27123
2 101518 1 27123
2 101519 1 27123
2 101520 1 27123
2 101521 1 27140
2 101522 1 27140
2 101523 1 27147
2 101524 1 27147
2 101525 1 27167
2 101526 1 27167
2 101527 1 27169
2 101528 1 27169
2 101529 1 27179
2 101530 1 27179
2 101531 1 27180
2 101532 1 27180
2 101533 1 27181
2 101534 1 27181
2 101535 1 27181
2 101536 1 27210
2 101537 1 27210
2 101538 1 27220
2 101539 1 27220
2 101540 1 27220
2 101541 1 27220
2 101542 1 27228
2 101543 1 27228
2 101544 1 27232
2 101545 1 27232
2 101546 1 27254
2 101547 1 27254
2 101548 1 27271
2 101549 1 27271
2 101550 1 27271
2 101551 1 27271
2 101552 1 27271
2 101553 1 27271
2 101554 1 27271
2 101555 1 27271
2 101556 1 27271
2 101557 1 27271
2 101558 1 27291
2 101559 1 27291
2 101560 1 27291
2 101561 1 27291
2 101562 1 27291
2 101563 1 27291
2 101564 1 27291
2 101565 1 27291
2 101566 1 27291
2 101567 1 27294
2 101568 1 27294
2 101569 1 27297
2 101570 1 27297
2 101571 1 27297
2 101572 1 27305
2 101573 1 27305
2 101574 1 27305
2 101575 1 27305
2 101576 1 27305
2 101577 1 27305
2 101578 1 27306
2 101579 1 27306
2 101580 1 27306
2 101581 1 27310
2 101582 1 27310
2 101583 1 27322
2 101584 1 27322
2 101585 1 27322
2 101586 1 27333
2 101587 1 27333
2 101588 1 27333
2 101589 1 27334
2 101590 1 27334
2 101591 1 27334
2 101592 1 27345
2 101593 1 27345
2 101594 1 27359
2 101595 1 27359
2 101596 1 27421
2 101597 1 27421
2 101598 1 27422
2 101599 1 27422
2 101600 1 27423
2 101601 1 27423
2 101602 1 27423
2 101603 1 27432
2 101604 1 27432
2 101605 1 27432
2 101606 1 27432
2 101607 1 27432
2 101608 1 27432
2 101609 1 27432
2 101610 1 27436
2 101611 1 27436
2 101612 1 27437
2 101613 1 27437
2 101614 1 27438
2 101615 1 27438
2 101616 1 27438
2 101617 1 27441
2 101618 1 27441
2 101619 1 27444
2 101620 1 27444
2 101621 1 27449
2 101622 1 27449
2 101623 1 27450
2 101624 1 27450
2 101625 1 27451
2 101626 1 27451
2 101627 1 27454
2 101628 1 27454
2 101629 1 27460
2 101630 1 27460
2 101631 1 27523
2 101632 1 27523
2 101633 1 27523
2 101634 1 27531
2 101635 1 27531
2 101636 1 27534
2 101637 1 27534
2 101638 1 27539
2 101639 1 27539
2 101640 1 27554
2 101641 1 27554
2 101642 1 27554
2 101643 1 27578
2 101644 1 27578
2 101645 1 27578
2 101646 1 27616
2 101647 1 27616
2 101648 1 27617
2 101649 1 27617
2 101650 1 27627
2 101651 1 27627
2 101652 1 27630
2 101653 1 27630
2 101654 1 27631
2 101655 1 27631
2 101656 1 27634
2 101657 1 27634
2 101658 1 27661
2 101659 1 27661
2 101660 1 27681
2 101661 1 27681
2 101662 1 27687
2 101663 1 27687
2 101664 1 27691
2 101665 1 27691
2 101666 1 27692
2 101667 1 27692
2 101668 1 27697
2 101669 1 27697
2 101670 1 27732
2 101671 1 27732
2 101672 1 27732
2 101673 1 27735
2 101674 1 27735
2 101675 1 27757
2 101676 1 27757
2 101677 1 27757
2 101678 1 27757
2 101679 1 27757
2 101680 1 27760
2 101681 1 27760
2 101682 1 27762
2 101683 1 27762
2 101684 1 27762
2 101685 1 27777
2 101686 1 27777
2 101687 1 27806
2 101688 1 27806
2 101689 1 27807
2 101690 1 27807
2 101691 1 27813
2 101692 1 27813
2 101693 1 27815
2 101694 1 27815
2 101695 1 27828
2 101696 1 27828
2 101697 1 27849
2 101698 1 27849
2 101699 1 27849
2 101700 1 27938
2 101701 1 27938
2 101702 1 27953
2 101703 1 27953
2 101704 1 27953
2 101705 1 27953
2 101706 1 27956
2 101707 1 27956
2 101708 1 27962
2 101709 1 27962
2 101710 1 27962
2 101711 1 27972
2 101712 1 27972
2 101713 1 27972
2 101714 1 27972
2 101715 1 27981
2 101716 1 27981
2 101717 1 27984
2 101718 1 27984
2 101719 1 27984
2 101720 1 27984
2 101721 1 27984
2 101722 1 27984
2 101723 1 27984
2 101724 1 27984
2 101725 1 27988
2 101726 1 27988
2 101727 1 27988
2 101728 1 28002
2 101729 1 28002
2 101730 1 28004
2 101731 1 28004
2 101732 1 28004
2 101733 1 28004
2 101734 1 28004
2 101735 1 28032
2 101736 1 28032
2 101737 1 28032
2 101738 1 28048
2 101739 1 28048
2 101740 1 28089
2 101741 1 28089
2 101742 1 28089
2 101743 1 28089
2 101744 1 28097
2 101745 1 28097
2 101746 1 28097
2 101747 1 28099
2 101748 1 28099
2 101749 1 28100
2 101750 1 28100
2 101751 1 28107
2 101752 1 28107
2 101753 1 28121
2 101754 1 28121
2 101755 1 28121
2 101756 1 28122
2 101757 1 28122
2 101758 1 28132
2 101759 1 28132
2 101760 1 28142
2 101761 1 28142
2 101762 1 28143
2 101763 1 28143
2 101764 1 28143
2 101765 1 28147
2 101766 1 28147
2 101767 1 28147
2 101768 1 28147
2 101769 1 28147
2 101770 1 28148
2 101771 1 28148
2 101772 1 28148
2 101773 1 28149
2 101774 1 28149
2 101775 1 28152
2 101776 1 28152
2 101777 1 28152
2 101778 1 28160
2 101779 1 28160
2 101780 1 28161
2 101781 1 28161
2 101782 1 28178
2 101783 1 28178
2 101784 1 28178
2 101785 1 28178
2 101786 1 28178
2 101787 1 28178
2 101788 1 28179
2 101789 1 28179
2 101790 1 28188
2 101791 1 28188
2 101792 1 28194
2 101793 1 28194
2 101794 1 28194
2 101795 1 28194
2 101796 1 28194
2 101797 1 28266
2 101798 1 28266
2 101799 1 28266
2 101800 1 28298
2 101801 1 28298
2 101802 1 28307
2 101803 1 28307
2 101804 1 28312
2 101805 1 28312
2 101806 1 28326
2 101807 1 28326
2 101808 1 28329
2 101809 1 28329
2 101810 1 28329
2 101811 1 28373
2 101812 1 28373
2 101813 1 28374
2 101814 1 28374
2 101815 1 28382
2 101816 1 28382
2 101817 1 28400
2 101818 1 28400
2 101819 1 28413
2 101820 1 28413
2 101821 1 28416
2 101822 1 28416
2 101823 1 28430
2 101824 1 28430
2 101825 1 28431
2 101826 1 28431
2 101827 1 28436
2 101828 1 28436
2 101829 1 28436
2 101830 1 28436
2 101831 1 28436
2 101832 1 28447
2 101833 1 28447
2 101834 1 28461
2 101835 1 28461
2 101836 1 28465
2 101837 1 28465
2 101838 1 28487
2 101839 1 28487
2 101840 1 28505
2 101841 1 28505
2 101842 1 28548
2 101843 1 28548
2 101844 1 28556
2 101845 1 28556
2 101846 1 28556
2 101847 1 28556
2 101848 1 28557
2 101849 1 28557
2 101850 1 28558
2 101851 1 28558
2 101852 1 28558
2 101853 1 28567
2 101854 1 28567
2 101855 1 28568
2 101856 1 28568
2 101857 1 28568
2 101858 1 28603
2 101859 1 28603
2 101860 1 28606
2 101861 1 28606
2 101862 1 28606
2 101863 1 28606
2 101864 1 28606
2 101865 1 28606
2 101866 1 28606
2 101867 1 28606
2 101868 1 28626
2 101869 1 28626
2 101870 1 28626
2 101871 1 28626
2 101872 1 28658
2 101873 1 28658
2 101874 1 28658
2 101875 1 28673
2 101876 1 28673
2 101877 1 28679
2 101878 1 28679
2 101879 1 28679
2 101880 1 28687
2 101881 1 28687
2 101882 1 28700
2 101883 1 28700
2 101884 1 28725
2 101885 1 28725
2 101886 1 28726
2 101887 1 28726
2 101888 1 28727
2 101889 1 28727
2 101890 1 28735
2 101891 1 28735
2 101892 1 28744
2 101893 1 28744
2 101894 1 28769
2 101895 1 28769
2 101896 1 28770
2 101897 1 28770
2 101898 1 28791
2 101899 1 28791
2 101900 1 28791
2 101901 1 28792
2 101902 1 28792
2 101903 1 28822
2 101904 1 28822
2 101905 1 28832
2 101906 1 28832
2 101907 1 28839
2 101908 1 28839
2 101909 1 28848
2 101910 1 28848
2 101911 1 28858
2 101912 1 28858
2 101913 1 28869
2 101914 1 28869
2 101915 1 28869
2 101916 1 28874
2 101917 1 28874
2 101918 1 28874
2 101919 1 28878
2 101920 1 28878
2 101921 1 28878
2 101922 1 28879
2 101923 1 28879
2 101924 1 28879
2 101925 1 28879
2 101926 1 28879
2 101927 1 28885
2 101928 1 28885
2 101929 1 28918
2 101930 1 28918
2 101931 1 28918
2 101932 1 28918
2 101933 1 28918
2 101934 1 28918
2 101935 1 28920
2 101936 1 28920
2 101937 1 28920
2 101938 1 28920
2 101939 1 28920
2 101940 1 28920
2 101941 1 28920
2 101942 1 28920
2 101943 1 28920
2 101944 1 28920
2 101945 1 28920
2 101946 1 28922
2 101947 1 28922
2 101948 1 28944
2 101949 1 28944
2 101950 1 28945
2 101951 1 28945
2 101952 1 28960
2 101953 1 28960
2 101954 1 28960
2 101955 1 28980
2 101956 1 28980
2 101957 1 28980
2 101958 1 29023
2 101959 1 29023
2 101960 1 29023
2 101961 1 29023
2 101962 1 29035
2 101963 1 29035
2 101964 1 29035
2 101965 1 29049
2 101966 1 29049
2 101967 1 29050
2 101968 1 29050
2 101969 1 29050
2 101970 1 29060
2 101971 1 29060
2 101972 1 29064
2 101973 1 29064
2 101974 1 29064
2 101975 1 29082
2 101976 1 29082
2 101977 1 29082
2 101978 1 29082
2 101979 1 29082
2 101980 1 29082
2 101981 1 29091
2 101982 1 29091
2 101983 1 29101
2 101984 1 29101
2 101985 1 29101
2 101986 1 29101
2 101987 1 29124
2 101988 1 29124
2 101989 1 29124
2 101990 1 29124
2 101991 1 29138
2 101992 1 29138
2 101993 1 29147
2 101994 1 29147
2 101995 1 29147
2 101996 1 29161
2 101997 1 29161
2 101998 1 29161
2 101999 1 29161
2 102000 1 29161
2 102001 1 29161
2 102002 1 29162
2 102003 1 29162
2 102004 1 29162
2 102005 1 29162
2 102006 1 29171
2 102007 1 29171
2 102008 1 29173
2 102009 1 29173
2 102010 1 29174
2 102011 1 29174
2 102012 1 29182
2 102013 1 29182
2 102014 1 29182
2 102015 1 29182
2 102016 1 29182
2 102017 1 29183
2 102018 1 29183
2 102019 1 29193
2 102020 1 29193
2 102021 1 29201
2 102022 1 29201
2 102023 1 29205
2 102024 1 29205
2 102025 1 29206
2 102026 1 29206
2 102027 1 29206
2 102028 1 29206
2 102029 1 29207
2 102030 1 29207
2 102031 1 29218
2 102032 1 29218
2 102033 1 29233
2 102034 1 29233
2 102035 1 29234
2 102036 1 29234
2 102037 1 29234
2 102038 1 29235
2 102039 1 29235
2 102040 1 29235
2 102041 1 29235
2 102042 1 29235
2 102043 1 29236
2 102044 1 29236
2 102045 1 29244
2 102046 1 29244
2 102047 1 29264
2 102048 1 29264
2 102049 1 29264
2 102050 1 29264
2 102051 1 29264
2 102052 1 29264
2 102053 1 29264
2 102054 1 29264
2 102055 1 29264
2 102056 1 29264
2 102057 1 29264
2 102058 1 29265
2 102059 1 29265
2 102060 1 29284
2 102061 1 29284
2 102062 1 29299
2 102063 1 29299
2 102064 1 29311
2 102065 1 29311
2 102066 1 29319
2 102067 1 29319
2 102068 1 29319
2 102069 1 29332
2 102070 1 29332
2 102071 1 29332
2 102072 1 29332
2 102073 1 29348
2 102074 1 29348
2 102075 1 29367
2 102076 1 29367
2 102077 1 29389
2 102078 1 29389
2 102079 1 29389
2 102080 1 29390
2 102081 1 29390
2 102082 1 29398
2 102083 1 29398
2 102084 1 29399
2 102085 1 29399
2 102086 1 29424
2 102087 1 29424
2 102088 1 29428
2 102089 1 29428
2 102090 1 29437
2 102091 1 29437
2 102092 1 29437
2 102093 1 29437
2 102094 1 29438
2 102095 1 29438
2 102096 1 29442
2 102097 1 29442
2 102098 1 29442
2 102099 1 29442
2 102100 1 29443
2 102101 1 29443
2 102102 1 29454
2 102103 1 29454
2 102104 1 29455
2 102105 1 29455
2 102106 1 29456
2 102107 1 29456
2 102108 1 29465
2 102109 1 29465
2 102110 1 29468
2 102111 1 29468
2 102112 1 29476
2 102113 1 29476
2 102114 1 29512
2 102115 1 29512
2 102116 1 29515
2 102117 1 29515
2 102118 1 29527
2 102119 1 29527
2 102120 1 29527
2 102121 1 29527
2 102122 1 29528
2 102123 1 29528
2 102124 1 29529
2 102125 1 29529
2 102126 1 29540
2 102127 1 29540
2 102128 1 29540
2 102129 1 29540
2 102130 1 29540
2 102131 1 29540
2 102132 1 29541
2 102133 1 29541
2 102134 1 29541
2 102135 1 29541
2 102136 1 29541
2 102137 1 29541
2 102138 1 29544
2 102139 1 29544
2 102140 1 29558
2 102141 1 29558
2 102142 1 29568
2 102143 1 29568
2 102144 1 29568
2 102145 1 29570
2 102146 1 29570
2 102147 1 29573
2 102148 1 29573
2 102149 1 29573
2 102150 1 29573
2 102151 1 29589
2 102152 1 29589
2 102153 1 29611
2 102154 1 29611
2 102155 1 29636
2 102156 1 29636
2 102157 1 29655
2 102158 1 29655
2 102159 1 29659
2 102160 1 29659
2 102161 1 29659
2 102162 1 29694
2 102163 1 29694
2 102164 1 29694
2 102165 1 29694
2 102166 1 29694
2 102167 1 29694
2 102168 1 29695
2 102169 1 29695
2 102170 1 29712
2 102171 1 29712
2 102172 1 29712
2 102173 1 29712
2 102174 1 29723
2 102175 1 29723
2 102176 1 29736
2 102177 1 29736
2 102178 1 29742
2 102179 1 29742
2 102180 1 29743
2 102181 1 29743
2 102182 1 29743
2 102183 1 29743
2 102184 1 29757
2 102185 1 29757
2 102186 1 29770
2 102187 1 29770
2 102188 1 29770
2 102189 1 29770
2 102190 1 29770
2 102191 1 29771
2 102192 1 29771
2 102193 1 29772
2 102194 1 29772
2 102195 1 29773
2 102196 1 29773
2 102197 1 29774
2 102198 1 29774
2 102199 1 29785
2 102200 1 29785
2 102201 1 29818
2 102202 1 29818
2 102203 1 29824
2 102204 1 29824
2 102205 1 29838
2 102206 1 29838
2 102207 1 29842
2 102208 1 29842
2 102209 1 29883
2 102210 1 29883
2 102211 1 29895
2 102212 1 29895
2 102213 1 29910
2 102214 1 29910
2 102215 1 29943
2 102216 1 29943
2 102217 1 29950
2 102218 1 29950
2 102219 1 29950
2 102220 1 29950
2 102221 1 29958
2 102222 1 29958
2 102223 1 29960
2 102224 1 29960
2 102225 1 29960
2 102226 1 29960
2 102227 1 29960
2 102228 1 29960
2 102229 1 29960
2 102230 1 29971
2 102231 1 29971
2 102232 1 29971
2 102233 1 29972
2 102234 1 29972
2 102235 1 29972
2 102236 1 29972
2 102237 1 29981
2 102238 1 29981
2 102239 1 29987
2 102240 1 29987
2 102241 1 30015
2 102242 1 30015
2 102243 1 30038
2 102244 1 30038
2 102245 1 30040
2 102246 1 30040
2 102247 1 30040
2 102248 1 30040
2 102249 1 30040
2 102250 1 30040
2 102251 1 30040
2 102252 1 30040
2 102253 1 30040
2 102254 1 30056
2 102255 1 30056
2 102256 1 30056
2 102257 1 30056
2 102258 1 30056
2 102259 1 30056
2 102260 1 30056
2 102261 1 30056
2 102262 1 30056
2 102263 1 30056
2 102264 1 30056
2 102265 1 30056
2 102266 1 30056
2 102267 1 30056
2 102268 1 30056
2 102269 1 30056
2 102270 1 30056
2 102271 1 30056
2 102272 1 30056
2 102273 1 30056
2 102274 1 30056
2 102275 1 30056
2 102276 1 30056
2 102277 1 30056
2 102278 1 30056
2 102279 1 30056
2 102280 1 30056
2 102281 1 30057
2 102282 1 30057
2 102283 1 30057
2 102284 1 30071
2 102285 1 30071
2 102286 1 30084
2 102287 1 30084
2 102288 1 30092
2 102289 1 30092
2 102290 1 30095
2 102291 1 30095
2 102292 1 30098
2 102293 1 30098
2 102294 1 30101
2 102295 1 30101
2 102296 1 30110
2 102297 1 30110
2 102298 1 30121
2 102299 1 30121
2 102300 1 30121
2 102301 1 30121
2 102302 1 30121
2 102303 1 30136
2 102304 1 30136
2 102305 1 30176
2 102306 1 30176
2 102307 1 30198
2 102308 1 30198
2 102309 1 30198
2 102310 1 30199
2 102311 1 30199
2 102312 1 30212
2 102313 1 30212
2 102314 1 30236
2 102315 1 30236
2 102316 1 30243
2 102317 1 30243
2 102318 1 30243
2 102319 1 30243
2 102320 1 30243
2 102321 1 30243
2 102322 1 30243
2 102323 1 30243
2 102324 1 30243
2 102325 1 30243
2 102326 1 30243
2 102327 1 30244
2 102328 1 30244
2 102329 1 30245
2 102330 1 30245
2 102331 1 30246
2 102332 1 30246
2 102333 1 30277
2 102334 1 30277
2 102335 1 30280
2 102336 1 30280
2 102337 1 30289
2 102338 1 30289
2 102339 1 30290
2 102340 1 30290
2 102341 1 30308
2 102342 1 30308
2 102343 1 30309
2 102344 1 30309
2 102345 1 30310
2 102346 1 30310
2 102347 1 30319
2 102348 1 30319
2 102349 1 30319
2 102350 1 30330
2 102351 1 30330
2 102352 1 30332
2 102353 1 30332
2 102354 1 30332
2 102355 1 30332
2 102356 1 30332
2 102357 1 30332
2 102358 1 30333
2 102359 1 30333
2 102360 1 30365
2 102361 1 30365
2 102362 1 30365
2 102363 1 30366
2 102364 1 30366
2 102365 1 30366
2 102366 1 30366
2 102367 1 30369
2 102368 1 30369
2 102369 1 30376
2 102370 1 30376
2 102371 1 30376
2 102372 1 30376
2 102373 1 30377
2 102374 1 30377
2 102375 1 30377
2 102376 1 30377
2 102377 1 30379
2 102378 1 30379
2 102379 1 30386
2 102380 1 30386
2 102381 1 30395
2 102382 1 30395
2 102383 1 30414
2 102384 1 30414
2 102385 1 30414
2 102386 1 30414
2 102387 1 30462
2 102388 1 30462
2 102389 1 30462
2 102390 1 30462
2 102391 1 30462
2 102392 1 30462
2 102393 1 30462
2 102394 1 30462
2 102395 1 30462
2 102396 1 30462
2 102397 1 30470
2 102398 1 30470
2 102399 1 30470
2 102400 1 30471
2 102401 1 30471
2 102402 1 30472
2 102403 1 30472
2 102404 1 30474
2 102405 1 30474
2 102406 1 30474
2 102407 1 30474
2 102408 1 30474
2 102409 1 30474
2 102410 1 30475
2 102411 1 30475
2 102412 1 30475
2 102413 1 30476
2 102414 1 30476
2 102415 1 30476
2 102416 1 30484
2 102417 1 30484
2 102418 1 30484
2 102419 1 30484
2 102420 1 30485
2 102421 1 30485
2 102422 1 30486
2 102423 1 30486
2 102424 1 30486
2 102425 1 30487
2 102426 1 30487
2 102427 1 30489
2 102428 1 30489
2 102429 1 30499
2 102430 1 30499
2 102431 1 30500
2 102432 1 30500
2 102433 1 30500
2 102434 1 30501
2 102435 1 30501
2 102436 1 30501
2 102437 1 30501
2 102438 1 30518
2 102439 1 30518
2 102440 1 30518
2 102441 1 30518
2 102442 1 30518
2 102443 1 30519
2 102444 1 30519
2 102445 1 30543
2 102446 1 30543
2 102447 1 30543
2 102448 1 30543
2 102449 1 30543
2 102450 1 30543
2 102451 1 30543
2 102452 1 30544
2 102453 1 30544
2 102454 1 30544
2 102455 1 30546
2 102456 1 30546
2 102457 1 30554
2 102458 1 30554
2 102459 1 30554
2 102460 1 30555
2 102461 1 30555
2 102462 1 30613
2 102463 1 30613
2 102464 1 30620
2 102465 1 30620
2 102466 1 30620
2 102467 1 30620
2 102468 1 30621
2 102469 1 30621
2 102470 1 30621
2 102471 1 30621
2 102472 1 30636
2 102473 1 30636
2 102474 1 30637
2 102475 1 30637
2 102476 1 30647
2 102477 1 30647
2 102478 1 30648
2 102479 1 30648
2 102480 1 30648
2 102481 1 30662
2 102482 1 30662
2 102483 1 30662
2 102484 1 30676
2 102485 1 30676
2 102486 1 30676
2 102487 1 30676
2 102488 1 30676
2 102489 1 30677
2 102490 1 30677
2 102491 1 30677
2 102492 1 30679
2 102493 1 30679
2 102494 1 30680
2 102495 1 30680
2 102496 1 30690
2 102497 1 30690
2 102498 1 30690
2 102499 1 30690
2 102500 1 30690
2 102501 1 30691
2 102502 1 30691
2 102503 1 30701
2 102504 1 30701
2 102505 1 30702
2 102506 1 30702
2 102507 1 30702
2 102508 1 30702
2 102509 1 30702
2 102510 1 30702
2 102511 1 30702
2 102512 1 30703
2 102513 1 30703
2 102514 1 30712
2 102515 1 30712
2 102516 1 30712
2 102517 1 30713
2 102518 1 30713
2 102519 1 30713
2 102520 1 30716
2 102521 1 30716
2 102522 1 30716
2 102523 1 30716
2 102524 1 30732
2 102525 1 30732
2 102526 1 30734
2 102527 1 30734
2 102528 1 30738
2 102529 1 30738
2 102530 1 30741
2 102531 1 30741
2 102532 1 30751
2 102533 1 30751
2 102534 1 30754
2 102535 1 30754
2 102536 1 30754
2 102537 1 30777
2 102538 1 30777
2 102539 1 30777
2 102540 1 30781
2 102541 1 30781
2 102542 1 30781
2 102543 1 30781
2 102544 1 30781
2 102545 1 30781
2 102546 1 30781
2 102547 1 30781
2 102548 1 30781
2 102549 1 30781
2 102550 1 30781
2 102551 1 30781
2 102552 1 30781
2 102553 1 30781
2 102554 1 30781
2 102555 1 30781
2 102556 1 30782
2 102557 1 30782
2 102558 1 30782
2 102559 1 30783
2 102560 1 30783
2 102561 1 30783
2 102562 1 30784
2 102563 1 30784
2 102564 1 30785
2 102565 1 30785
2 102566 1 30796
2 102567 1 30796
2 102568 1 30797
2 102569 1 30797
2 102570 1 30797
2 102571 1 30825
2 102572 1 30825
2 102573 1 30825
2 102574 1 30825
2 102575 1 30825
2 102576 1 30825
2 102577 1 30825
2 102578 1 30825
2 102579 1 30826
2 102580 1 30826
2 102581 1 30827
2 102582 1 30827
2 102583 1 30827
2 102584 1 30838
2 102585 1 30838
2 102586 1 30846
2 102587 1 30846
2 102588 1 30870
2 102589 1 30870
2 102590 1 30871
2 102591 1 30871
2 102592 1 30872
2 102593 1 30872
2 102594 1 30874
2 102595 1 30874
2 102596 1 30874
2 102597 1 30877
2 102598 1 30877
2 102599 1 30880
2 102600 1 30880
2 102601 1 30880
2 102602 1 30897
2 102603 1 30897
2 102604 1 30897
2 102605 1 30897
2 102606 1 30939
2 102607 1 30939
2 102608 1 30950
2 102609 1 30950
2 102610 1 30950
2 102611 1 30950
2 102612 1 30950
2 102613 1 30951
2 102614 1 30951
2 102615 1 30951
2 102616 1 30955
2 102617 1 30955
2 102618 1 30955
2 102619 1 30955
2 102620 1 30955
2 102621 1 30955
2 102622 1 30955
2 102623 1 30955
2 102624 1 30955
2 102625 1 30955
2 102626 1 30955
2 102627 1 30955
2 102628 1 30955
2 102629 1 30955
2 102630 1 30955
2 102631 1 30955
2 102632 1 30955
2 102633 1 30955
2 102634 1 30955
2 102635 1 30955
2 102636 1 30955
2 102637 1 30955
2 102638 1 30955
2 102639 1 30955
2 102640 1 30955
2 102641 1 30955
2 102642 1 30955
2 102643 1 30955
2 102644 1 30955
2 102645 1 30955
2 102646 1 30955
2 102647 1 30955
2 102648 1 30955
2 102649 1 30955
2 102650 1 30955
2 102651 1 30956
2 102652 1 30956
2 102653 1 30956
2 102654 1 30956
2 102655 1 30956
2 102656 1 30956
2 102657 1 30956
2 102658 1 30956
2 102659 1 30957
2 102660 1 30957
2 102661 1 30963
2 102662 1 30963
2 102663 1 30963
2 102664 1 30963
2 102665 1 30963
2 102666 1 30963
2 102667 1 30963
2 102668 1 30963
2 102669 1 30964
2 102670 1 30964
2 102671 1 30964
2 102672 1 30964
2 102673 1 30964
2 102674 1 30965
2 102675 1 30965
2 102676 1 30965
2 102677 1 30965
2 102678 1 30965
2 102679 1 30965
2 102680 1 30965
2 102681 1 30965
2 102682 1 30965
2 102683 1 30965
2 102684 1 30965
2 102685 1 30965
2 102686 1 30965
2 102687 1 30965
2 102688 1 30965
2 102689 1 30965
2 102690 1 30965
2 102691 1 30965
2 102692 1 30965
2 102693 1 30965
2 102694 1 30965
2 102695 1 30965
2 102696 1 30965
2 102697 1 30965
2 102698 1 30965
2 102699 1 30965
2 102700 1 30965
2 102701 1 30965
2 102702 1 30965
2 102703 1 30966
2 102704 1 30966
2 102705 1 30966
2 102706 1 30966
2 102707 1 30966
2 102708 1 30966
2 102709 1 30966
2 102710 1 30966
2 102711 1 30966
2 102712 1 30967
2 102713 1 30967
2 102714 1 30967
2 102715 1 30967
2 102716 1 30972
2 102717 1 30972
2 102718 1 30986
2 102719 1 30986
2 102720 1 30986
2 102721 1 30986
2 102722 1 30995
2 102723 1 30995
2 102724 1 30996
2 102725 1 30996
2 102726 1 31008
2 102727 1 31008
2 102728 1 31009
2 102729 1 31009
2 102730 1 31009
2 102731 1 31009
2 102732 1 31022
2 102733 1 31022
2 102734 1 31022
2 102735 1 31022
2 102736 1 31022
2 102737 1 31022
2 102738 1 31022
2 102739 1 31022
2 102740 1 31022
2 102741 1 31023
2 102742 1 31023
2 102743 1 31023
2 102744 1 31024
2 102745 1 31024
2 102746 1 31024
2 102747 1 31024
2 102748 1 31024
2 102749 1 31024
2 102750 1 31024
2 102751 1 31024
2 102752 1 31024
2 102753 1 31024
2 102754 1 31024
2 102755 1 31024
2 102756 1 31024
2 102757 1 31025
2 102758 1 31025
2 102759 1 31025
2 102760 1 31025
2 102761 1 31028
2 102762 1 31028
2 102763 1 31028
2 102764 1 31028
2 102765 1 31028
2 102766 1 31030
2 102767 1 31030
2 102768 1 31031
2 102769 1 31031
2 102770 1 31031
2 102771 1 31031
2 102772 1 31031
2 102773 1 31031
2 102774 1 31031
2 102775 1 31031
2 102776 1 31031
2 102777 1 31031
2 102778 1 31035
2 102779 1 31035
2 102780 1 31035
2 102781 1 31038
2 102782 1 31038
2 102783 1 31046
2 102784 1 31046
2 102785 1 31061
2 102786 1 31061
2 102787 1 31062
2 102788 1 31062
2 102789 1 31062
2 102790 1 31071
2 102791 1 31071
2 102792 1 31071
2 102793 1 31071
2 102794 1 31071
2 102795 1 31071
2 102796 1 31071
2 102797 1 31072
2 102798 1 31072
2 102799 1 31072
2 102800 1 31072
2 102801 1 31072
2 102802 1 31088
2 102803 1 31088
2 102804 1 31088
2 102805 1 31088
2 102806 1 31088
2 102807 1 31089
2 102808 1 31089
2 102809 1 31090
2 102810 1 31090
2 102811 1 31092
2 102812 1 31092
2 102813 1 31092
2 102814 1 31092
2 102815 1 31100
2 102816 1 31100
2 102817 1 31100
2 102818 1 31100
2 102819 1 31100
2 102820 1 31100
2 102821 1 31107
2 102822 1 31107
2 102823 1 31107
2 102824 1 31107
2 102825 1 31107
2 102826 1 31108
2 102827 1 31108
2 102828 1 31113
2 102829 1 31113
2 102830 1 31113
2 102831 1 31119
2 102832 1 31119
2 102833 1 31128
2 102834 1 31128
2 102835 1 31129
2 102836 1 31129
2 102837 1 31129
2 102838 1 31129
2 102839 1 31135
2 102840 1 31135
2 102841 1 31141
2 102842 1 31141
2 102843 1 31141
2 102844 1 31141
2 102845 1 31146
2 102846 1 31146
2 102847 1 31154
2 102848 1 31154
2 102849 1 31154
2 102850 1 31154
2 102851 1 31154
2 102852 1 31173
2 102853 1 31173
2 102854 1 31201
2 102855 1 31201
2 102856 1 31201
2 102857 1 31201
2 102858 1 31201
2 102859 1 31201
2 102860 1 31201
2 102861 1 31201
2 102862 1 31201
2 102863 1 31217
2 102864 1 31217
2 102865 1 31217
2 102866 1 31217
2 102867 1 31217
2 102868 1 31227
2 102869 1 31227
2 102870 1 31252
2 102871 1 31252
2 102872 1 31252
2 102873 1 31253
2 102874 1 31253
2 102875 1 31255
2 102876 1 31255
2 102877 1 31271
2 102878 1 31271
2 102879 1 31271
2 102880 1 31272
2 102881 1 31272
2 102882 1 31282
2 102883 1 31282
2 102884 1 31285
2 102885 1 31285
2 102886 1 31287
2 102887 1 31287
2 102888 1 31287
2 102889 1 31290
2 102890 1 31290
2 102891 1 31291
2 102892 1 31291
2 102893 1 31291
2 102894 1 31291
2 102895 1 31299
2 102896 1 31299
2 102897 1 31307
2 102898 1 31307
2 102899 1 31307
2 102900 1 31307
2 102901 1 31308
2 102902 1 31308
2 102903 1 31308
2 102904 1 31308
2 102905 1 31308
2 102906 1 31308
2 102907 1 31308
2 102908 1 31308
2 102909 1 31308
2 102910 1 31312
2 102911 1 31312
2 102912 1 31322
2 102913 1 31322
2 102914 1 31340
2 102915 1 31340
2 102916 1 31348
2 102917 1 31348
2 102918 1 31356
2 102919 1 31356
2 102920 1 31356
2 102921 1 31359
2 102922 1 31359
2 102923 1 31360
2 102924 1 31360
2 102925 1 31360
2 102926 1 31360
2 102927 1 31360
2 102928 1 31360
2 102929 1 31361
2 102930 1 31361
2 102931 1 31364
2 102932 1 31364
2 102933 1 31364
2 102934 1 31364
2 102935 1 31364
2 102936 1 31364
2 102937 1 31364
2 102938 1 31364
2 102939 1 31366
2 102940 1 31366
2 102941 1 31367
2 102942 1 31367
2 102943 1 31382
2 102944 1 31382
2 102945 1 31383
2 102946 1 31383
2 102947 1 31388
2 102948 1 31388
2 102949 1 31388
2 102950 1 31389
2 102951 1 31389
2 102952 1 31392
2 102953 1 31392
2 102954 1 31392
2 102955 1 31392
2 102956 1 31396
2 102957 1 31396
2 102958 1 31396
2 102959 1 31405
2 102960 1 31405
2 102961 1 31406
2 102962 1 31406
2 102963 1 31415
2 102964 1 31415
2 102965 1 31424
2 102966 1 31424
2 102967 1 31470
2 102968 1 31470
2 102969 1 31470
2 102970 1 31475
2 102971 1 31475
2 102972 1 31479
2 102973 1 31479
2 102974 1 31480
2 102975 1 31480
2 102976 1 31490
2 102977 1 31490
2 102978 1 31512
2 102979 1 31512
2 102980 1 31512
2 102981 1 31513
2 102982 1 31513
2 102983 1 31516
2 102984 1 31516
2 102985 1 31516
2 102986 1 31516
2 102987 1 31523
2 102988 1 31523
2 102989 1 31532
2 102990 1 31532
2 102991 1 31532
2 102992 1 31547
2 102993 1 31547
2 102994 1 31547
2 102995 1 31563
2 102996 1 31563
2 102997 1 31564
2 102998 1 31564
2 102999 1 31564
2 103000 1 31564
2 103001 1 31568
2 103002 1 31568
2 103003 1 31569
2 103004 1 31569
2 103005 1 31569
2 103006 1 31591
2 103007 1 31591
2 103008 1 31604
2 103009 1 31604
2 103010 1 31604
2 103011 1 31604
2 103012 1 31640
2 103013 1 31640
2 103014 1 31640
2 103015 1 31640
2 103016 1 31640
2 103017 1 31640
2 103018 1 31640
2 103019 1 31641
2 103020 1 31641
2 103021 1 31655
2 103022 1 31655
2 103023 1 31656
2 103024 1 31656
2 103025 1 31689
2 103026 1 31689
2 103027 1 31729
2 103028 1 31729
2 103029 1 31730
2 103030 1 31730
2 103031 1 31750
2 103032 1 31750
2 103033 1 31756
2 103034 1 31756
2 103035 1 31760
2 103036 1 31760
2 103037 1 31778
2 103038 1 31778
2 103039 1 31778
2 103040 1 31778
2 103041 1 31779
2 103042 1 31779
2 103043 1 31780
2 103044 1 31780
2 103045 1 31784
2 103046 1 31784
2 103047 1 31788
2 103048 1 31788
2 103049 1 31788
2 103050 1 31788
2 103051 1 31788
2 103052 1 31788
2 103053 1 31789
2 103054 1 31789
2 103055 1 31801
2 103056 1 31801
2 103057 1 31801
2 103058 1 31824
2 103059 1 31824
2 103060 1 31824
2 103061 1 31827
2 103062 1 31827
2 103063 1 31827
2 103064 1 31835
2 103065 1 31835
2 103066 1 31835
2 103067 1 31839
2 103068 1 31839
2 103069 1 31839
2 103070 1 31855
2 103071 1 31855
2 103072 1 31855
2 103073 1 31855
2 103074 1 31857
2 103075 1 31857
2 103076 1 31864
2 103077 1 31864
2 103078 1 31873
2 103079 1 31873
2 103080 1 31873
2 103081 1 31885
2 103082 1 31885
2 103083 1 31887
2 103084 1 31887
2 103085 1 31887
2 103086 1 31888
2 103087 1 31888
2 103088 1 31899
2 103089 1 31899
2 103090 1 31924
2 103091 1 31924
2 103092 1 31926
2 103093 1 31926
2 103094 1 31927
2 103095 1 31927
2 103096 1 31928
2 103097 1 31928
2 103098 1 31928
2 103099 1 31928
2 103100 1 31946
2 103101 1 31946
2 103102 1 31946
2 103103 1 31946
2 103104 1 31949
2 103105 1 31949
2 103106 1 31949
2 103107 1 31989
2 103108 1 31989
2 103109 1 32000
2 103110 1 32000
2 103111 1 32007
2 103112 1 32007
2 103113 1 32026
2 103114 1 32026
2 103115 1 32034
2 103116 1 32034
2 103117 1 32036
2 103118 1 32036
2 103119 1 32037
2 103120 1 32037
2 103121 1 32037
2 103122 1 32037
2 103123 1 32038
2 103124 1 32038
2 103125 1 32038
2 103126 1 32058
2 103127 1 32058
2 103128 1 32102
2 103129 1 32102
2 103130 1 32102
2 103131 1 32108
2 103132 1 32108
2 103133 1 32118
2 103134 1 32118
2 103135 1 32118
2 103136 1 32118
2 103137 1 32118
2 103138 1 32118
2 103139 1 32118
2 103140 1 32118
2 103141 1 32118
2 103142 1 32118
2 103143 1 32119
2 103144 1 32119
2 103145 1 32119
2 103146 1 32119
2 103147 1 32119
2 103148 1 32131
2 103149 1 32131
2 103150 1 32131
2 103151 1 32136
2 103152 1 32136
2 103153 1 32137
2 103154 1 32137
2 103155 1 32146
2 103156 1 32146
2 103157 1 32147
2 103158 1 32147
2 103159 1 32154
2 103160 1 32154
2 103161 1 32184
2 103162 1 32184
2 103163 1 32194
2 103164 1 32194
2 103165 1 32198
2 103166 1 32198
2 103167 1 32198
2 103168 1 32198
2 103169 1 32198
2 103170 1 32206
2 103171 1 32206
2 103172 1 32208
2 103173 1 32208
2 103174 1 32208
2 103175 1 32222
2 103176 1 32222
2 103177 1 32223
2 103178 1 32223
2 103179 1 32223
2 103180 1 32232
2 103181 1 32232
2 103182 1 32258
2 103183 1 32258
2 103184 1 32266
2 103185 1 32266
2 103186 1 32268
2 103187 1 32268
2 103188 1 32268
2 103189 1 32285
2 103190 1 32285
2 103191 1 32292
2 103192 1 32292
2 103193 1 32315
2 103194 1 32315
2 103195 1 32315
2 103196 1 32316
2 103197 1 32316
2 103198 1 32317
2 103199 1 32317
2 103200 1 32339
2 103201 1 32339
2 103202 1 32339
2 103203 1 32339
2 103204 1 32339
2 103205 1 32339
2 103206 1 32339
2 103207 1 32341
2 103208 1 32341
2 103209 1 32369
2 103210 1 32369
2 103211 1 32410
2 103212 1 32410
2 103213 1 32418
2 103214 1 32418
2 103215 1 32433
2 103216 1 32433
2 103217 1 32454
2 103218 1 32454
2 103219 1 32454
2 103220 1 32479
2 103221 1 32479
2 103222 1 32481
2 103223 1 32481
2 103224 1 32487
2 103225 1 32487
2 103226 1 32496
2 103227 1 32496
2 103228 1 32565
2 103229 1 32565
2 103230 1 32566
2 103231 1 32566
2 103232 1 32566
2 103233 1 32567
2 103234 1 32567
2 103235 1 32573
2 103236 1 32573
2 103237 1 32573
2 103238 1 32592
2 103239 1 32592
2 103240 1 32592
2 103241 1 32609
2 103242 1 32609
2 103243 1 32619
2 103244 1 32619
2 103245 1 32619
2 103246 1 32627
2 103247 1 32627
2 103248 1 32627
2 103249 1 32639
2 103250 1 32639
2 103251 1 32640
2 103252 1 32640
2 103253 1 32656
2 103254 1 32656
2 103255 1 32657
2 103256 1 32657
2 103257 1 32657
2 103258 1 32657
2 103259 1 32657
2 103260 1 32657
2 103261 1 32657
2 103262 1 32657
2 103263 1 32658
2 103264 1 32658
2 103265 1 32675
2 103266 1 32675
2 103267 1 32675
2 103268 1 32675
2 103269 1 32675
2 103270 1 32675
2 103271 1 32675
2 103272 1 32675
2 103273 1 32675
2 103274 1 32676
2 103275 1 32676
2 103276 1 32676
2 103277 1 32677
2 103278 1 32677
2 103279 1 32677
2 103280 1 32687
2 103281 1 32687
2 103282 1 32688
2 103283 1 32688
2 103284 1 32688
2 103285 1 32700
2 103286 1 32700
2 103287 1 32700
2 103288 1 32703
2 103289 1 32703
2 103290 1 32730
2 103291 1 32730
2 103292 1 32746
2 103293 1 32746
2 103294 1 32746
2 103295 1 32746
2 103296 1 32746
2 103297 1 32746
2 103298 1 32746
2 103299 1 32746
2 103300 1 32746
2 103301 1 32756
2 103302 1 32756
2 103303 1 32757
2 103304 1 32757
2 103305 1 32775
2 103306 1 32775
2 103307 1 32778
2 103308 1 32778
2 103309 1 32778
2 103310 1 32778
2 103311 1 32778
2 103312 1 32778
2 103313 1 32778
2 103314 1 32778
2 103315 1 32778
2 103316 1 32788
2 103317 1 32788
2 103318 1 32788
2 103319 1 32801
2 103320 1 32801
2 103321 1 32809
2 103322 1 32809
2 103323 1 32814
2 103324 1 32814
2 103325 1 32827
2 103326 1 32827
2 103327 1 32836
2 103328 1 32836
2 103329 1 32836
2 103330 1 32837
2 103331 1 32837
2 103332 1 32848
2 103333 1 32848
2 103334 1 32855
2 103335 1 32855
2 103336 1 32855
2 103337 1 32862
2 103338 1 32862
2 103339 1 32862
2 103340 1 32862
2 103341 1 32862
2 103342 1 32862
2 103343 1 32862
2 103344 1 32862
2 103345 1 32862
2 103346 1 32886
2 103347 1 32886
2 103348 1 32886
2 103349 1 32886
2 103350 1 32910
2 103351 1 32910
2 103352 1 32910
2 103353 1 32930
2 103354 1 32930
2 103355 1 32930
2 103356 1 32930
2 103357 1 32930
2 103358 1 32930
2 103359 1 32930
2 103360 1 32947
2 103361 1 32947
2 103362 1 32947
2 103363 1 32947
2 103364 1 32950
2 103365 1 32950
2 103366 1 32969
2 103367 1 32969
2 103368 1 32969
2 103369 1 32970
2 103370 1 32970
2 103371 1 32998
2 103372 1 32998
2 103373 1 32999
2 103374 1 32999
2 103375 1 33012
2 103376 1 33012
2 103377 1 33012
2 103378 1 33013
2 103379 1 33013
2 103380 1 33014
2 103381 1 33014
2 103382 1 33041
2 103383 1 33041
2 103384 1 33041
2 103385 1 33056
2 103386 1 33056
2 103387 1 33057
2 103388 1 33057
2 103389 1 33057
2 103390 1 33069
2 103391 1 33069
2 103392 1 33069
2 103393 1 33073
2 103394 1 33073
2 103395 1 33116
2 103396 1 33116
2 103397 1 33133
2 103398 1 33133
2 103399 1 33135
2 103400 1 33135
2 103401 1 33143
2 103402 1 33143
2 103403 1 33168
2 103404 1 33168
2 103405 1 33179
2 103406 1 33179
2 103407 1 33220
2 103408 1 33220
2 103409 1 33220
2 103410 1 33220
2 103411 1 33220
2 103412 1 33247
2 103413 1 33247
2 103414 1 33248
2 103415 1 33248
2 103416 1 33250
2 103417 1 33250
2 103418 1 33252
2 103419 1 33252
2 103420 1 33268
2 103421 1 33268
2 103422 1 33275
2 103423 1 33275
2 103424 1 33304
2 103425 1 33304
2 103426 1 33305
2 103427 1 33305
2 103428 1 33305
2 103429 1 33305
2 103430 1 33307
2 103431 1 33307
2 103432 1 33307
2 103433 1 33320
2 103434 1 33320
2 103435 1 33325
2 103436 1 33325
2 103437 1 33339
2 103438 1 33339
2 103439 1 33339
2 103440 1 33341
2 103441 1 33341
2 103442 1 33342
2 103443 1 33342
2 103444 1 33342
2 103445 1 33342
2 103446 1 33342
2 103447 1 33342
2 103448 1 33355
2 103449 1 33355
2 103450 1 33355
2 103451 1 33355
2 103452 1 33355
2 103453 1 33364
2 103454 1 33364
2 103455 1 33364
2 103456 1 33364
2 103457 1 33366
2 103458 1 33366
2 103459 1 33371
2 103460 1 33371
2 103461 1 33372
2 103462 1 33372
2 103463 1 33396
2 103464 1 33396
2 103465 1 33396
2 103466 1 33404
2 103467 1 33404
2 103468 1 33420
2 103469 1 33420
2 103470 1 33422
2 103471 1 33422
2 103472 1 33434
2 103473 1 33434
2 103474 1 33436
2 103475 1 33436
2 103476 1 33457
2 103477 1 33457
2 103478 1 33465
2 103479 1 33465
2 103480 1 33475
2 103481 1 33475
2 103482 1 33487
2 103483 1 33487
2 103484 1 33502
2 103485 1 33502
2 103486 1 33503
2 103487 1 33503
2 103488 1 33503
2 103489 1 33503
2 103490 1 33503
2 103491 1 33543
2 103492 1 33543
2 103493 1 33543
2 103494 1 33543
2 103495 1 33543
2 103496 1 33556
2 103497 1 33556
2 103498 1 33566
2 103499 1 33566
2 103500 1 33576
2 103501 1 33576
2 103502 1 33585
2 103503 1 33585
2 103504 1 33585
2 103505 1 33585
2 103506 1 33587
2 103507 1 33587
2 103508 1 33587
2 103509 1 33598
2 103510 1 33598
2 103511 1 33599
2 103512 1 33599
2 103513 1 33625
2 103514 1 33625
2 103515 1 33625
2 103516 1 33640
2 103517 1 33640
2 103518 1 33659
2 103519 1 33659
2 103520 1 33662
2 103521 1 33662
2 103522 1 33662
2 103523 1 33668
2 103524 1 33668
2 103525 1 33668
2 103526 1 33668
2 103527 1 33726
2 103528 1 33726
2 103529 1 33740
2 103530 1 33740
2 103531 1 33807
2 103532 1 33807
2 103533 1 33847
2 103534 1 33847
2 103535 1 33848
2 103536 1 33848
2 103537 1 33850
2 103538 1 33850
2 103539 1 33861
2 103540 1 33861
2 103541 1 33861
2 103542 1 33865
2 103543 1 33865
2 103544 1 33865
2 103545 1 33873
2 103546 1 33873
2 103547 1 33882
2 103548 1 33882
2 103549 1 33892
2 103550 1 33892
2 103551 1 33919
2 103552 1 33919
2 103553 1 33941
2 103554 1 33941
2 103555 1 33941
2 103556 1 33943
2 103557 1 33943
2 103558 1 33944
2 103559 1 33944
2 103560 1 33963
2 103561 1 33963
2 103562 1 33963
2 103563 1 33963
2 103564 1 33963
2 103565 1 33963
2 103566 1 33964
2 103567 1 33964
2 103568 1 33965
2 103569 1 33965
2 103570 1 33967
2 103571 1 33967
2 103572 1 33985
2 103573 1 33985
2 103574 1 33985
2 103575 1 33985
2 103576 1 33986
2 103577 1 33986
2 103578 1 33986
2 103579 1 33992
2 103580 1 33992
2 103581 1 33994
2 103582 1 33994
2 103583 1 33997
2 103584 1 33997
2 103585 1 33997
2 103586 1 34036
2 103587 1 34036
2 103588 1 34036
2 103589 1 34040
2 103590 1 34040
2 103591 1 34060
2 103592 1 34060
2 103593 1 34070
2 103594 1 34070
2 103595 1 34071
2 103596 1 34071
2 103597 1 34071
2 103598 1 34073
2 103599 1 34073
2 103600 1 34077
2 103601 1 34077
2 103602 1 34078
2 103603 1 34078
2 103604 1 34079
2 103605 1 34079
2 103606 1 34079
2 103607 1 34079
2 103608 1 34080
2 103609 1 34080
2 103610 1 34084
2 103611 1 34084
2 103612 1 34112
2 103613 1 34112
2 103614 1 34112
2 103615 1 34112
2 103616 1 34112
2 103617 1 34113
2 103618 1 34113
2 103619 1 34113
2 103620 1 34113
2 103621 1 34113
2 103622 1 34123
2 103623 1 34123
2 103624 1 34123
2 103625 1 34123
2 103626 1 34139
2 103627 1 34139
2 103628 1 34168
2 103629 1 34168
2 103630 1 34199
2 103631 1 34199
2 103632 1 34199
2 103633 1 34199
2 103634 1 34202
2 103635 1 34202
2 103636 1 34237
2 103637 1 34237
2 103638 1 34238
2 103639 1 34238
2 103640 1 34238
2 103641 1 34238
2 103642 1 34238
2 103643 1 34252
2 103644 1 34252
2 103645 1 34254
2 103646 1 34254
2 103647 1 34254
2 103648 1 34263
2 103649 1 34263
2 103650 1 34266
2 103651 1 34266
2 103652 1 34266
2 103653 1 34267
2 103654 1 34267
2 103655 1 34268
2 103656 1 34268
2 103657 1 34268
2 103658 1 34271
2 103659 1 34271
2 103660 1 34306
2 103661 1 34306
2 103662 1 34306
2 103663 1 34307
2 103664 1 34307
2 103665 1 34319
2 103666 1 34319
2 103667 1 34319
2 103668 1 34319
2 103669 1 34319
2 103670 1 34319
2 103671 1 34320
2 103672 1 34320
2 103673 1 34320
2 103674 1 34321
2 103675 1 34321
2 103676 1 34328
2 103677 1 34328
2 103678 1 34381
2 103679 1 34381
2 103680 1 34394
2 103681 1 34394
2 103682 1 34394
2 103683 1 34395
2 103684 1 34395
2 103685 1 34406
2 103686 1 34406
2 103687 1 34428
2 103688 1 34428
2 103689 1 34428
2 103690 1 34428
2 103691 1 34429
2 103692 1 34429
2 103693 1 34441
2 103694 1 34441
2 103695 1 34444
2 103696 1 34444
2 103697 1 34447
2 103698 1 34447
2 103699 1 34447
2 103700 1 34471
2 103701 1 34471
2 103702 1 34471
2 103703 1 34471
2 103704 1 34490
2 103705 1 34490
2 103706 1 34491
2 103707 1 34491
2 103708 1 34506
2 103709 1 34506
2 103710 1 34523
2 103711 1 34523
2 103712 1 34523
2 103713 1 34532
2 103714 1 34532
2 103715 1 34544
2 103716 1 34544
2 103717 1 34544
2 103718 1 34573
2 103719 1 34573
2 103720 1 34596
2 103721 1 34596
2 103722 1 34638
2 103723 1 34638
2 103724 1 34687
2 103725 1 34687
2 103726 1 34687
2 103727 1 34697
2 103728 1 34697
2 103729 1 34719
2 103730 1 34719
2 103731 1 34719
2 103732 1 34719
2 103733 1 34720
2 103734 1 34720
2 103735 1 34747
2 103736 1 34747
2 103737 1 34758
2 103738 1 34758
2 103739 1 34766
2 103740 1 34766
2 103741 1 34774
2 103742 1 34774
2 103743 1 34774
2 103744 1 34774
2 103745 1 34775
2 103746 1 34775
2 103747 1 34783
2 103748 1 34783
2 103749 1 34783
2 103750 1 34783
2 103751 1 34796
2 103752 1 34796
2 103753 1 34796
2 103754 1 34803
2 103755 1 34803
2 103756 1 34813
2 103757 1 34813
2 103758 1 34813
2 103759 1 34813
2 103760 1 34814
2 103761 1 34814
2 103762 1 34815
2 103763 1 34815
2 103764 1 34825
2 103765 1 34825
2 103766 1 34826
2 103767 1 34826
2 103768 1 34826
2 103769 1 34831
2 103770 1 34831
2 103771 1 34857
2 103772 1 34857
2 103773 1 34872
2 103774 1 34872
2 103775 1 34875
2 103776 1 34875
2 103777 1 34876
2 103778 1 34876
2 103779 1 34876
2 103780 1 34879
2 103781 1 34879
2 103782 1 34893
2 103783 1 34893
2 103784 1 34893
2 103785 1 34901
2 103786 1 34901
2 103787 1 34901
2 103788 1 34902
2 103789 1 34902
2 103790 1 34904
2 103791 1 34904
2 103792 1 34904
2 103793 1 34905
2 103794 1 34905
2 103795 1 34916
2 103796 1 34916
2 103797 1 34917
2 103798 1 34917
2 103799 1 34930
2 103800 1 34930
2 103801 1 34930
2 103802 1 34930
2 103803 1 34955
2 103804 1 34955
2 103805 1 34987
2 103806 1 34987
2 103807 1 34990
2 103808 1 34990
2 103809 1 35002
2 103810 1 35002
2 103811 1 35012
2 103812 1 35012
2 103813 1 35012
2 103814 1 35013
2 103815 1 35013
2 103816 1 35023
2 103817 1 35023
2 103818 1 35023
2 103819 1 35025
2 103820 1 35025
2 103821 1 35026
2 103822 1 35026
2 103823 1 35026
2 103824 1 35027
2 103825 1 35027
2 103826 1 35027
2 103827 1 35027
2 103828 1 35027
2 103829 1 35027
2 103830 1 35036
2 103831 1 35036
2 103832 1 35036
2 103833 1 35041
2 103834 1 35041
2 103835 1 35041
2 103836 1 35076
2 103837 1 35076
2 103838 1 35108
2 103839 1 35108
2 103840 1 35125
2 103841 1 35125
2 103842 1 35125
2 103843 1 35140
2 103844 1 35140
2 103845 1 35140
2 103846 1 35140
2 103847 1 35141
2 103848 1 35141
2 103849 1 35155
2 103850 1 35155
2 103851 1 35164
2 103852 1 35164
2 103853 1 35164
2 103854 1 35166
2 103855 1 35166
2 103856 1 35166
2 103857 1 35166
2 103858 1 35172
2 103859 1 35172
2 103860 1 35184
2 103861 1 35184
2 103862 1 35184
2 103863 1 35199
2 103864 1 35199
2 103865 1 35199
2 103866 1 35199
2 103867 1 35214
2 103868 1 35214
2 103869 1 35214
2 103870 1 35221
2 103871 1 35221
2 103872 1 35267
2 103873 1 35267
2 103874 1 35276
2 103875 1 35276
2 103876 1 35277
2 103877 1 35277
2 103878 1 35277
2 103879 1 35287
2 103880 1 35287
2 103881 1 35294
2 103882 1 35294
2 103883 1 35294
2 103884 1 35294
2 103885 1 35294
2 103886 1 35295
2 103887 1 35295
2 103888 1 35295
2 103889 1 35295
2 103890 1 35295
2 103891 1 35295
2 103892 1 35295
2 103893 1 35295
2 103894 1 35295
2 103895 1 35298
2 103896 1 35298
2 103897 1 35305
2 103898 1 35305
2 103899 1 35305
2 103900 1 35305
2 103901 1 35305
2 103902 1 35306
2 103903 1 35306
2 103904 1 35319
2 103905 1 35319
2 103906 1 35319
2 103907 1 35319
2 103908 1 35319
2 103909 1 35319
2 103910 1 35319
2 103911 1 35328
2 103912 1 35328
2 103913 1 35360
2 103914 1 35360
2 103915 1 35369
2 103916 1 35369
2 103917 1 35369
2 103918 1 35374
2 103919 1 35374
2 103920 1 35405
2 103921 1 35405
2 103922 1 35431
2 103923 1 35431
2 103924 1 35431
2 103925 1 35434
2 103926 1 35434
2 103927 1 35434
2 103928 1 35434
2 103929 1 35434
2 103930 1 35434
2 103931 1 35434
2 103932 1 35434
2 103933 1 35434
2 103934 1 35435
2 103935 1 35435
2 103936 1 35435
2 103937 1 35435
2 103938 1 35435
2 103939 1 35435
2 103940 1 35435
2 103941 1 35435
2 103942 1 35435
2 103943 1 35435
2 103944 1 35436
2 103945 1 35436
2 103946 1 35438
2 103947 1 35438
2 103948 1 35438
2 103949 1 35438
2 103950 1 35438
2 103951 1 35438
2 103952 1 35438
2 103953 1 35438
2 103954 1 35438
2 103955 1 35438
2 103956 1 35438
2 103957 1 35438
2 103958 1 35438
2 103959 1 35438
2 103960 1 35438
2 103961 1 35438
2 103962 1 35438
2 103963 1 35438
2 103964 1 35438
2 103965 1 35445
2 103966 1 35445
2 103967 1 35449
2 103968 1 35449
2 103969 1 35466
2 103970 1 35466
2 103971 1 35466
2 103972 1 35466
2 103973 1 35466
2 103974 1 35466
2 103975 1 35475
2 103976 1 35475
2 103977 1 35476
2 103978 1 35476
2 103979 1 35485
2 103980 1 35485
2 103981 1 35485
2 103982 1 35505
2 103983 1 35505
2 103984 1 35506
2 103985 1 35506
2 103986 1 35531
2 103987 1 35531
2 103988 1 35565
2 103989 1 35565
2 103990 1 35565
2 103991 1 35565
2 103992 1 35573
2 103993 1 35573
2 103994 1 35582
2 103995 1 35582
2 103996 1 35583
2 103997 1 35583
2 103998 1 35587
2 103999 1 35587
2 104000 1 35587
2 104001 1 35587
2 104002 1 35589
2 104003 1 35589
2 104004 1 35597
2 104005 1 35597
2 104006 1 35616
2 104007 1 35616
2 104008 1 35638
2 104009 1 35638
2 104010 1 35647
2 104011 1 35647
2 104012 1 35655
2 104013 1 35655
2 104014 1 35655
2 104015 1 35658
2 104016 1 35658
2 104017 1 35659
2 104018 1 35659
2 104019 1 35664
2 104020 1 35664
2 104021 1 35690
2 104022 1 35690
2 104023 1 35697
2 104024 1 35697
2 104025 1 35717
2 104026 1 35717
2 104027 1 35735
2 104028 1 35735
2 104029 1 35736
2 104030 1 35736
2 104031 1 35785
2 104032 1 35785
2 104033 1 35786
2 104034 1 35786
2 104035 1 35795
2 104036 1 35795
2 104037 1 35796
2 104038 1 35796
2 104039 1 35799
2 104040 1 35799
2 104041 1 35808
2 104042 1 35808
2 104043 1 35848
2 104044 1 35848
2 104045 1 35866
2 104046 1 35866
2 104047 1 35869
2 104048 1 35869
2 104049 1 35883
2 104050 1 35883
2 104051 1 35883
2 104052 1 35884
2 104053 1 35884
2 104054 1 35885
2 104055 1 35885
2 104056 1 35885
2 104057 1 35910
2 104058 1 35910
2 104059 1 35910
2 104060 1 35910
2 104061 1 35910
2 104062 1 35910
2 104063 1 35910
2 104064 1 35910
2 104065 1 35911
2 104066 1 35911
2 104067 1 35911
2 104068 1 35911
2 104069 1 35913
2 104070 1 35913
2 104071 1 35927
2 104072 1 35927
2 104073 1 35944
2 104074 1 35944
2 104075 1 35944
2 104076 1 35985
2 104077 1 35985
2 104078 1 35989
2 104079 1 35989
2 104080 1 35997
2 104081 1 35997
2 104082 1 36017
2 104083 1 36017
2 104084 1 36020
2 104085 1 36020
2 104086 1 36026
2 104087 1 36026
2 104088 1 36070
2 104089 1 36070
2 104090 1 36072
2 104091 1 36072
2 104092 1 36073
2 104093 1 36073
2 104094 1 36121
2 104095 1 36121
2 104096 1 36128
2 104097 1 36128
2 104098 1 36128
2 104099 1 36135
2 104100 1 36135
2 104101 1 36135
2 104102 1 36135
2 104103 1 36135
2 104104 1 36160
2 104105 1 36160
2 104106 1 36214
2 104107 1 36214
2 104108 1 36294
2 104109 1 36294
2 104110 1 36314
2 104111 1 36314
2 104112 1 36314
2 104113 1 36314
2 104114 1 36316
2 104115 1 36316
2 104116 1 36326
2 104117 1 36326
2 104118 1 36329
2 104119 1 36329
2 104120 1 36329
2 104121 1 36360
2 104122 1 36360
2 104123 1 36363
2 104124 1 36363
2 104125 1 36363
2 104126 1 36363
2 104127 1 36363
2 104128 1 36363
2 104129 1 36363
2 104130 1 36363
2 104131 1 36363
2 104132 1 36363
2 104133 1 36372
2 104134 1 36372
2 104135 1 36379
2 104136 1 36379
2 104137 1 36419
2 104138 1 36419
2 104139 1 36419
2 104140 1 36419
2 104141 1 36419
2 104142 1 36419
2 104143 1 36437
2 104144 1 36437
2 104145 1 36442
2 104146 1 36442
2 104147 1 36447
2 104148 1 36447
2 104149 1 36461
2 104150 1 36461
2 104151 1 36493
2 104152 1 36493
2 104153 1 36493
2 104154 1 36493
2 104155 1 36493
2 104156 1 36493
2 104157 1 36493
2 104158 1 36493
2 104159 1 36493
2 104160 1 36493
2 104161 1 36494
2 104162 1 36494
2 104163 1 36495
2 104164 1 36495
2 104165 1 36498
2 104166 1 36498
2 104167 1 36553
2 104168 1 36553
2 104169 1 36553
2 104170 1 36592
2 104171 1 36592
2 104172 1 36617
2 104173 1 36617
2 104174 1 36634
2 104175 1 36634
2 104176 1 36649
2 104177 1 36649
2 104178 1 36662
2 104179 1 36662
2 104180 1 36662
2 104181 1 36695
2 104182 1 36695
2 104183 1 36739
2 104184 1 36739
2 104185 1 36758
2 104186 1 36758
2 104187 1 36758
2 104188 1 36771
2 104189 1 36771
2 104190 1 36782
2 104191 1 36782
2 104192 1 36822
2 104193 1 36822
2 104194 1 36829
2 104195 1 36829
2 104196 1 36868
2 104197 1 36868
2 104198 1 36868
2 104199 1 36868
2 104200 1 36870
2 104201 1 36870
2 104202 1 36877
2 104203 1 36877
2 104204 1 36884
2 104205 1 36884
2 104206 1 36895
2 104207 1 36895
2 104208 1 36895
2 104209 1 36895
2 104210 1 36896
2 104211 1 36896
2 104212 1 36941
2 104213 1 36941
2 104214 1 36945
2 104215 1 36945
2 104216 1 36980
2 104217 1 36980
2 104218 1 36981
2 104219 1 36981
2 104220 1 36982
2 104221 1 36982
2 104222 1 36982
2 104223 1 36983
2 104224 1 36983
2 104225 1 36993
2 104226 1 36993
2 104227 1 36993
2 104228 1 37001
2 104229 1 37001
2 104230 1 37001
2 104231 1 37006
2 104232 1 37006
2 104233 1 37030
2 104234 1 37030
2 104235 1 37150
2 104236 1 37150
2 104237 1 37163
2 104238 1 37163
2 104239 1 37163
2 104240 1 37182
2 104241 1 37182
2 104242 1 37215
2 104243 1 37215
2 104244 1 37215
2 104245 1 37225
2 104246 1 37225
2 104247 1 37247
2 104248 1 37247
2 104249 1 37279
2 104250 1 37279
2 104251 1 37286
2 104252 1 37286
2 104253 1 37296
2 104254 1 37296
2 104255 1 37297
2 104256 1 37297
2 104257 1 37310
2 104258 1 37310
2 104259 1 37310
2 104260 1 37310
2 104261 1 37310
2 104262 1 37310
2 104263 1 37322
2 104264 1 37322
2 104265 1 37334
2 104266 1 37334
2 104267 1 37335
2 104268 1 37335
2 104269 1 37335
2 104270 1 37335
2 104271 1 37335
2 104272 1 37336
2 104273 1 37336
2 104274 1 37359
2 104275 1 37359
2 104276 1 37359
2 104277 1 37359
2 104278 1 37363
2 104279 1 37363
2 104280 1 37363
2 104281 1 37363
2 104282 1 37365
2 104283 1 37365
2 104284 1 37368
2 104285 1 37368
2 104286 1 37368
2 104287 1 37392
2 104288 1 37392
2 104289 1 37392
2 104290 1 37426
2 104291 1 37426
2 104292 1 37447
2 104293 1 37447
2 104294 1 37447
2 104295 1 37447
2 104296 1 37447
2 104297 1 37467
2 104298 1 37467
2 104299 1 37483
2 104300 1 37483
2 104301 1 37504
2 104302 1 37504
2 104303 1 37507
2 104304 1 37507
2 104305 1 37526
2 104306 1 37526
2 104307 1 37527
2 104308 1 37527
2 104309 1 37535
2 104310 1 37535
2 104311 1 37548
2 104312 1 37548
2 104313 1 37548
2 104314 1 37564
2 104315 1 37564
2 104316 1 37564
2 104317 1 37564
2 104318 1 37582
2 104319 1 37582
2 104320 1 37630
2 104321 1 37630
2 104322 1 37630
2 104323 1 37630
2 104324 1 37630
2 104325 1 37630
2 104326 1 37630
2 104327 1 37630
2 104328 1 37635
2 104329 1 37635
2 104330 1 37635
2 104331 1 37638
2 104332 1 37638
2 104333 1 37647
2 104334 1 37647
2 104335 1 37662
2 104336 1 37662
2 104337 1 37662
2 104338 1 37671
2 104339 1 37671
2 104340 1 37676
2 104341 1 37676
2 104342 1 37679
2 104343 1 37679
2 104344 1 37679
2 104345 1 37690
2 104346 1 37690
2 104347 1 37713
2 104348 1 37713
2 104349 1 37734
2 104350 1 37734
2 104351 1 37734
2 104352 1 37754
2 104353 1 37754
2 104354 1 37758
2 104355 1 37758
2 104356 1 37799
2 104357 1 37799
2 104358 1 37806
2 104359 1 37806
2 104360 1 37819
2 104361 1 37819
2 104362 1 37822
2 104363 1 37822
2 104364 1 37823
2 104365 1 37823
2 104366 1 37867
2 104367 1 37867
2 104368 1 37867
2 104369 1 37867
2 104370 1 37867
2 104371 1 37867
2 104372 1 37868
2 104373 1 37868
2 104374 1 37905
2 104375 1 37905
2 104376 1 37906
2 104377 1 37906
2 104378 1 37913
2 104379 1 37913
2 104380 1 37913
2 104381 1 37915
2 104382 1 37915
2 104383 1 37915
2 104384 1 37916
2 104385 1 37916
2 104386 1 37922
2 104387 1 37922
2 104388 1 37940
2 104389 1 37940
2 104390 1 37940
2 104391 1 37948
2 104392 1 37948
2 104393 1 37948
2 104394 1 37967
2 104395 1 37967
2 104396 1 37973
2 104397 1 37973
2 104398 1 38000
2 104399 1 38000
2 104400 1 38013
2 104401 1 38013
2 104402 1 38026
2 104403 1 38026
2 104404 1 38026
2 104405 1 38050
2 104406 1 38050
2 104407 1 38052
2 104408 1 38052
2 104409 1 38061
2 104410 1 38061
2 104411 1 38129
2 104412 1 38129
2 104413 1 38129
2 104414 1 38142
2 104415 1 38142
2 104416 1 38168
2 104417 1 38168
2 104418 1 38168
2 104419 1 38169
2 104420 1 38169
2 104421 1 38170
2 104422 1 38170
2 104423 1 38179
2 104424 1 38179
2 104425 1 38179
2 104426 1 38179
2 104427 1 38179
2 104428 1 38186
2 104429 1 38186
2 104430 1 38226
2 104431 1 38226
2 104432 1 38226
2 104433 1 38227
2 104434 1 38227
2 104435 1 38227
2 104436 1 38235
2 104437 1 38235
2 104438 1 38235
2 104439 1 38235
2 104440 1 38249
2 104441 1 38249
2 104442 1 38249
2 104443 1 38270
2 104444 1 38270
2 104445 1 38270
2 104446 1 38270
2 104447 1 38298
2 104448 1 38298
2 104449 1 38314
2 104450 1 38314
2 104451 1 38314
2 104452 1 38314
2 104453 1 38324
2 104454 1 38324
2 104455 1 38324
2 104456 1 38337
2 104457 1 38337
2 104458 1 38340
2 104459 1 38340
2 104460 1 38346
2 104461 1 38346
2 104462 1 38346
2 104463 1 38346
2 104464 1 38355
2 104465 1 38355
2 104466 1 38356
2 104467 1 38356
2 104468 1 38363
2 104469 1 38363
2 104470 1 38371
2 104471 1 38371
2 104472 1 38373
2 104473 1 38373
2 104474 1 38420
2 104475 1 38420
2 104476 1 38469
2 104477 1 38469
2 104478 1 38484
2 104479 1 38484
2 104480 1 38494
2 104481 1 38494
2 104482 1 38505
2 104483 1 38505
2 104484 1 38510
2 104485 1 38510
2 104486 1 38517
2 104487 1 38517
2 104488 1 38547
2 104489 1 38547
2 104490 1 38550
2 104491 1 38550
2 104492 1 38551
2 104493 1 38551
2 104494 1 38584
2 104495 1 38584
2 104496 1 38585
2 104497 1 38585
2 104498 1 38585
2 104499 1 38586
2 104500 1 38586
2 104501 1 38599
2 104502 1 38599
2 104503 1 38599
2 104504 1 38602
2 104505 1 38602
2 104506 1 38609
2 104507 1 38609
2 104508 1 38610
2 104509 1 38610
2 104510 1 38610
2 104511 1 38610
2 104512 1 38610
2 104513 1 38610
2 104514 1 38610
2 104515 1 38618
2 104516 1 38618
2 104517 1 38618
2 104518 1 38620
2 104519 1 38620
2 104520 1 38628
2 104521 1 38628
2 104522 1 38628
2 104523 1 38628
2 104524 1 38638
2 104525 1 38638
2 104526 1 38638
2 104527 1 38639
2 104528 1 38639
2 104529 1 38647
2 104530 1 38647
2 104531 1 38647
2 104532 1 38669
2 104533 1 38669
2 104534 1 38669
2 104535 1 38669
2 104536 1 38669
2 104537 1 38670
2 104538 1 38670
2 104539 1 38671
2 104540 1 38671
2 104541 1 38671
2 104542 1 38671
2 104543 1 38671
2 104544 1 38689
2 104545 1 38689
2 104546 1 38689
2 104547 1 38689
2 104548 1 38724
2 104549 1 38724
2 104550 1 38739
2 104551 1 38739
2 104552 1 38800
2 104553 1 38800
2 104554 1 38837
2 104555 1 38837
2 104556 1 38845
2 104557 1 38845
2 104558 1 38863
2 104559 1 38863
2 104560 1 38889
2 104561 1 38889
2 104562 1 38889
2 104563 1 38889
2 104564 1 38890
2 104565 1 38890
2 104566 1 38905
2 104567 1 38905
2 104568 1 38909
2 104569 1 38909
2 104570 1 38913
2 104571 1 38913
2 104572 1 38925
2 104573 1 38925
2 104574 1 38925
2 104575 1 38925
2 104576 1 38925
2 104577 1 38925
2 104578 1 38935
2 104579 1 38935
2 104580 1 38940
2 104581 1 38940
2 104582 1 38960
2 104583 1 38960
2 104584 1 38964
2 104585 1 38964
2 104586 1 38974
2 104587 1 38974
2 104588 1 38996
2 104589 1 38996
2 104590 1 38996
2 104591 1 39002
2 104592 1 39002
2 104593 1 39002
2 104594 1 39004
2 104595 1 39004
2 104596 1 39012
2 104597 1 39012
2 104598 1 39028
2 104599 1 39028
2 104600 1 39043
2 104601 1 39043
2 104602 1 39060
2 104603 1 39060
2 104604 1 39060
2 104605 1 39060
2 104606 1 39068
2 104607 1 39068
2 104608 1 39068
2 104609 1 39068
2 104610 1 39069
2 104611 1 39069
2 104612 1 39078
2 104613 1 39078
2 104614 1 39088
2 104615 1 39088
2 104616 1 39095
2 104617 1 39095
2 104618 1 39095
2 104619 1 39095
2 104620 1 39095
2 104621 1 39096
2 104622 1 39096
2 104623 1 39127
2 104624 1 39127
2 104625 1 39127
2 104626 1 39138
2 104627 1 39138
2 104628 1 39138
2 104629 1 39138
2 104630 1 39147
2 104631 1 39147
2 104632 1 39162
2 104633 1 39162
2 104634 1 39162
2 104635 1 39195
2 104636 1 39195
2 104637 1 39195
2 104638 1 39195
2 104639 1 39208
2 104640 1 39208
2 104641 1 39208
2 104642 1 39208
2 104643 1 39208
2 104644 1 39235
2 104645 1 39235
2 104646 1 39290
2 104647 1 39290
2 104648 1 39315
2 104649 1 39315
2 104650 1 39326
2 104651 1 39326
2 104652 1 39335
2 104653 1 39335
2 104654 1 39408
2 104655 1 39408
2 104656 1 39419
2 104657 1 39419
2 104658 1 39419
2 104659 1 39419
2 104660 1 39433
2 104661 1 39433
2 104662 1 39438
2 104663 1 39438
2 104664 1 39446
2 104665 1 39446
2 104666 1 39446
2 104667 1 39446
2 104668 1 39446
2 104669 1 39458
2 104670 1 39458
2 104671 1 39469
2 104672 1 39469
2 104673 1 39477
2 104674 1 39477
2 104675 1 39478
2 104676 1 39478
2 104677 1 39478
2 104678 1 39533
2 104679 1 39533
2 104680 1 39533
2 104681 1 39540
2 104682 1 39540
2 104683 1 39540
2 104684 1 39540
2 104685 1 39540
2 104686 1 39547
2 104687 1 39547
2 104688 1 39549
2 104689 1 39549
2 104690 1 39560
2 104691 1 39560
2 104692 1 39582
2 104693 1 39582
2 104694 1 39598
2 104695 1 39598
2 104696 1 39628
2 104697 1 39628
2 104698 1 39638
2 104699 1 39638
2 104700 1 39653
2 104701 1 39653
2 104702 1 39659
2 104703 1 39659
2 104704 1 39659
2 104705 1 39659
2 104706 1 39659
2 104707 1 39668
2 104708 1 39668
2 104709 1 39686
2 104710 1 39686
2 104711 1 39687
2 104712 1 39687
2 104713 1 39687
2 104714 1 39687
2 104715 1 39695
2 104716 1 39695
2 104717 1 39726
2 104718 1 39726
2 104719 1 39742
2 104720 1 39742
2 104721 1 39759
2 104722 1 39759
2 104723 1 39759
2 104724 1 39771
2 104725 1 39771
2 104726 1 39790
2 104727 1 39790
2 104728 1 39791
2 104729 1 39791
2 104730 1 39791
2 104731 1 39798
2 104732 1 39798
2 104733 1 39798
2 104734 1 39799
2 104735 1 39799
2 104736 1 39819
2 104737 1 39819
2 104738 1 39881
2 104739 1 39881
2 104740 1 39881
2 104741 1 39925
2 104742 1 39925
2 104743 1 39926
2 104744 1 39926
2 104745 1 39926
2 104746 1 39926
2 104747 1 39955
2 104748 1 39955
2 104749 1 39999
2 104750 1 39999
2 104751 1 40020
2 104752 1 40020
2 104753 1 40025
2 104754 1 40025
2 104755 1 40025
2 104756 1 40026
2 104757 1 40026
2 104758 1 40044
2 104759 1 40044
2 104760 1 40044
2 104761 1 40044
2 104762 1 40044
2 104763 1 40044
2 104764 1 40044
2 104765 1 40061
2 104766 1 40061
2 104767 1 40061
2 104768 1 40063
2 104769 1 40063
2 104770 1 40063
2 104771 1 40063
2 104772 1 40087
2 104773 1 40087
2 104774 1 40095
2 104775 1 40095
2 104776 1 40104
2 104777 1 40104
2 104778 1 40109
2 104779 1 40109
2 104780 1 40137
2 104781 1 40137
2 104782 1 40138
2 104783 1 40138
2 104784 1 40146
2 104785 1 40146
2 104786 1 40149
2 104787 1 40149
2 104788 1 40157
2 104789 1 40157
2 104790 1 40173
2 104791 1 40173
2 104792 1 40195
2 104793 1 40195
2 104794 1 40195
2 104795 1 40196
2 104796 1 40196
2 104797 1 40198
2 104798 1 40198
2 104799 1 40198
2 104800 1 40198
2 104801 1 40198
2 104802 1 40201
2 104803 1 40201
2 104804 1 40228
2 104805 1 40228
2 104806 1 40229
2 104807 1 40229
2 104808 1 40231
2 104809 1 40231
2 104810 1 40237
2 104811 1 40237
2 104812 1 40277
2 104813 1 40277
2 104814 1 40324
2 104815 1 40324
2 104816 1 40352
2 104817 1 40352
2 104818 1 40353
2 104819 1 40353
2 104820 1 40373
2 104821 1 40373
2 104822 1 40373
2 104823 1 40373
2 104824 1 40383
2 104825 1 40383
2 104826 1 40383
2 104827 1 40398
2 104828 1 40398
2 104829 1 40430
2 104830 1 40430
2 104831 1 40437
2 104832 1 40437
2 104833 1 40438
2 104834 1 40438
2 104835 1 40449
2 104836 1 40449
2 104837 1 40457
2 104838 1 40457
2 104839 1 40458
2 104840 1 40458
2 104841 1 40458
2 104842 1 40459
2 104843 1 40459
2 104844 1 40459
2 104845 1 40460
2 104846 1 40460
2 104847 1 40465
2 104848 1 40465
2 104849 1 40521
2 104850 1 40521
2 104851 1 40557
2 104852 1 40557
2 104853 1 40599
2 104854 1 40599
2 104855 1 40600
2 104856 1 40600
2 104857 1 40603
2 104858 1 40603
2 104859 1 40675
2 104860 1 40675
2 104861 1 40718
2 104862 1 40718
2 104863 1 40718
2 104864 1 40751
2 104865 1 40751
2 104866 1 40751
2 104867 1 40761
2 104868 1 40761
2 104869 1 40776
2 104870 1 40776
2 104871 1 40799
2 104872 1 40799
2 104873 1 40800
2 104874 1 40800
2 104875 1 40808
2 104876 1 40808
2 104877 1 40850
2 104878 1 40850
2 104879 1 40858
2 104880 1 40858
2 104881 1 40858
2 104882 1 40858
2 104883 1 40858
2 104884 1 40858
2 104885 1 40858
2 104886 1 40866
2 104887 1 40866
2 104888 1 40894
2 104889 1 40894
2 104890 1 40894
2 104891 1 40894
2 104892 1 40908
2 104893 1 40908
2 104894 1 40922
2 104895 1 40922
2 104896 1 41002
2 104897 1 41002
2 104898 1 41010
2 104899 1 41010
2 104900 1 41023
2 104901 1 41023
2 104902 1 41118
2 104903 1 41118
2 104904 1 41118
2 104905 1 41132
2 104906 1 41132
2 104907 1 41132
2 104908 1 41132
2 104909 1 41132
2 104910 1 41133
2 104911 1 41133
2 104912 1 41158
2 104913 1 41158
2 104914 1 41159
2 104915 1 41159
2 104916 1 41170
2 104917 1 41170
2 104918 1 41184
2 104919 1 41184
2 104920 1 41185
2 104921 1 41185
2 104922 1 41185
2 104923 1 41186
2 104924 1 41186
2 104925 1 41189
2 104926 1 41189
2 104927 1 41208
2 104928 1 41208
2 104929 1 41227
2 104930 1 41227
2 104931 1 41237
2 104932 1 41237
2 104933 1 41245
2 104934 1 41245
2 104935 1 41321
2 104936 1 41321
2 104937 1 41321
2 104938 1 41321
2 104939 1 41321
2 104940 1 41359
2 104941 1 41359
2 104942 1 41367
2 104943 1 41367
2 104944 1 41375
2 104945 1 41375
2 104946 1 41375
2 104947 1 41375
2 104948 1 41416
2 104949 1 41416
2 104950 1 41422
2 104951 1 41422
2 104952 1 41422
2 104953 1 41474
2 104954 1 41474
2 104955 1 41587
2 104956 1 41587
2 104957 1 41599
2 104958 1 41599
2 104959 1 41599
2 104960 1 41612
2 104961 1 41612
2 104962 1 41616
2 104963 1 41616
2 104964 1 41619
2 104965 1 41619
2 104966 1 41651
2 104967 1 41651
2 104968 1 41662
2 104969 1 41662
2 104970 1 41696
2 104971 1 41696
2 104972 1 41696
2 104973 1 41717
2 104974 1 41717
2 104975 1 41717
2 104976 1 41717
2 104977 1 41788
2 104978 1 41788
2 104979 1 41853
2 104980 1 41853
2 104981 1 41864
2 104982 1 41864
2 104983 1 41866
2 104984 1 41866
2 104985 1 41902
2 104986 1 41902
2 104987 1 41929
2 104988 1 41929
2 104989 1 42025
2 104990 1 42025
2 104991 1 42073
2 104992 1 42073
2 104993 1 42090
2 104994 1 42090
2 104995 1 42091
2 104996 1 42091
2 104997 1 42102
2 104998 1 42102
2 104999 1 42102
2 105000 1 42102
2 105001 1 42141
2 105002 1 42141
2 105003 1 42141
2 105004 1 42234
2 105005 1 42234
2 105006 1 42235
2 105007 1 42235
2 105008 1 42237
2 105009 1 42237
2 105010 1 42237
2 105011 1 42237
2 105012 1 42237
2 105013 1 42237
2 105014 1 42254
2 105015 1 42254
2 105016 1 42254
2 105017 1 42261
2 105018 1 42261
2 105019 1 42261
2 105020 1 42262
2 105021 1 42262
2 105022 1 42306
2 105023 1 42306
2 105024 1 42342
2 105025 1 42342
2 105026 1 42345
2 105027 1 42345
2 105028 1 42345
2 105029 1 42345
2 105030 1 42372
2 105031 1 42372
2 105032 1 42386
2 105033 1 42386
2 105034 1 42389
2 105035 1 42389
2 105036 1 42397
2 105037 1 42397
2 105038 1 42397
2 105039 1 42417
2 105040 1 42417
2 105041 1 42417
2 105042 1 42433
2 105043 1 42433
2 105044 1 42434
2 105045 1 42434
2 105046 1 42434
2 105047 1 42436
2 105048 1 42436
2 105049 1 42439
2 105050 1 42439
2 105051 1 42446
2 105052 1 42446
2 105053 1 42447
2 105054 1 42447
2 105055 1 42456
2 105056 1 42456
2 105057 1 42463
2 105058 1 42463
2 105059 1 42464
2 105060 1 42464
2 105061 1 42471
2 105062 1 42471
2 105063 1 42471
2 105064 1 42525
2 105065 1 42525
2 105066 1 42532
2 105067 1 42532
2 105068 1 42532
2 105069 1 42532
2 105070 1 42532
2 105071 1 42533
2 105072 1 42533
2 105073 1 42533
2 105074 1 42533
2 105075 1 42538
2 105076 1 42538
2 105077 1 42539
2 105078 1 42539
2 105079 1 42558
2 105080 1 42558
2 105081 1 42558
2 105082 1 42558
2 105083 1 42558
2 105084 1 42558
2 105085 1 42558
2 105086 1 42558
2 105087 1 42558
2 105088 1 42558
2 105089 1 42559
2 105090 1 42559
2 105091 1 42587
2 105092 1 42587
2 105093 1 42590
2 105094 1 42590
2 105095 1 42617
2 105096 1 42617
2 105097 1 42617
2 105098 1 42627
2 105099 1 42627
2 105100 1 42627
2 105101 1 42643
2 105102 1 42643
2 105103 1 42651
2 105104 1 42651
2 105105 1 42651
2 105106 1 42685
2 105107 1 42685
2 105108 1 42685
2 105109 1 42693
2 105110 1 42693
2 105111 1 42695
2 105112 1 42695
2 105113 1 42748
2 105114 1 42748
2 105115 1 42773
2 105116 1 42773
2 105117 1 42788
2 105118 1 42788
2 105119 1 42792
2 105120 1 42792
2 105121 1 42855
2 105122 1 42855
2 105123 1 42863
2 105124 1 42863
2 105125 1 42868
2 105126 1 42868
2 105127 1 42871
2 105128 1 42871
2 105129 1 42871
2 105130 1 42884
2 105131 1 42884
2 105132 1 42884
2 105133 1 42893
2 105134 1 42893
2 105135 1 42916
2 105136 1 42916
2 105137 1 42916
2 105138 1 42916
2 105139 1 42916
2 105140 1 42916
2 105141 1 42918
2 105142 1 42918
2 105143 1 42934
2 105144 1 42934
2 105145 1 42934
2 105146 1 42934
2 105147 1 42934
2 105148 1 42953
2 105149 1 42953
2 105150 1 42958
2 105151 1 42958
2 105152 1 42958
2 105153 1 42958
2 105154 1 42981
2 105155 1 42981
2 105156 1 42982
2 105157 1 42982
2 105158 1 42982
2 105159 1 42983
2 105160 1 42983
2 105161 1 42983
2 105162 1 42983
2 105163 1 43001
2 105164 1 43001
2 105165 1 43001
2 105166 1 43001
2 105167 1 43026
2 105168 1 43026
2 105169 1 43056
2 105170 1 43056
2 105171 1 43076
2 105172 1 43076
2 105173 1 43079
2 105174 1 43079
2 105175 1 43092
2 105176 1 43092
2 105177 1 43095
2 105178 1 43095
2 105179 1 43129
2 105180 1 43129
2 105181 1 43157
2 105182 1 43157
2 105183 1 43175
2 105184 1 43175
2 105185 1 43175
2 105186 1 43252
2 105187 1 43252
2 105188 1 43254
2 105189 1 43254
2 105190 1 43254
2 105191 1 43298
2 105192 1 43298
2 105193 1 43298
2 105194 1 43298
2 105195 1 43298
2 105196 1 43341
2 105197 1 43341
2 105198 1 43344
2 105199 1 43344
2 105200 1 43344
2 105201 1 43346
2 105202 1 43346
2 105203 1 43368
2 105204 1 43368
2 105205 1 43368
2 105206 1 43368
2 105207 1 43369
2 105208 1 43369
2 105209 1 43382
2 105210 1 43382
2 105211 1 43390
2 105212 1 43390
2 105213 1 43497
2 105214 1 43497
2 105215 1 43508
2 105216 1 43508
2 105217 1 43532
2 105218 1 43532
2 105219 1 43552
2 105220 1 43552
2 105221 1 43552
2 105222 1 43572
2 105223 1 43572
2 105224 1 43617
2 105225 1 43617
2 105226 1 43617
2 105227 1 43645
2 105228 1 43645
2 105229 1 43648
2 105230 1 43648
2 105231 1 43651
2 105232 1 43651
2 105233 1 43651
2 105234 1 43652
2 105235 1 43652
2 105236 1 43652
2 105237 1 43653
2 105238 1 43653
2 105239 1 43653
2 105240 1 43667
2 105241 1 43667
2 105242 1 43694
2 105243 1 43694
2 105244 1 43761
2 105245 1 43761
2 105246 1 43761
2 105247 1 43761
2 105248 1 43761
2 105249 1 43763
2 105250 1 43763
2 105251 1 43766
2 105252 1 43766
2 105253 1 43766
2 105254 1 43776
2 105255 1 43776
2 105256 1 43817
2 105257 1 43817
2 105258 1 43817
2 105259 1 43819
2 105260 1 43819
2 105261 1 43831
2 105262 1 43831
2 105263 1 43832
2 105264 1 43832
2 105265 1 43853
2 105266 1 43853
2 105267 1 43862
2 105268 1 43862
2 105269 1 43862
2 105270 1 43862
2 105271 1 43862
2 105272 1 43862
2 105273 1 43863
2 105274 1 43863
2 105275 1 43872
2 105276 1 43872
2 105277 1 43873
2 105278 1 43873
2 105279 1 43877
2 105280 1 43877
2 105281 1 43897
2 105282 1 43897
2 105283 1 43898
2 105284 1 43898
2 105285 1 43907
2 105286 1 43907
2 105287 1 43910
2 105288 1 43910
2 105289 1 43934
2 105290 1 43934
2 105291 1 43935
2 105292 1 43935
2 105293 1 43945
2 105294 1 43945
2 105295 1 43950
2 105296 1 43950
2 105297 1 43993
2 105298 1 43993
2 105299 1 44046
2 105300 1 44046
2 105301 1 44059
2 105302 1 44059
2 105303 1 44059
2 105304 1 44086
2 105305 1 44086
2 105306 1 44086
2 105307 1 44086
2 105308 1 44087
2 105309 1 44087
2 105310 1 44096
2 105311 1 44096
2 105312 1 44099
2 105313 1 44099
2 105314 1 44099
2 105315 1 44108
2 105316 1 44108
2 105317 1 44108
2 105318 1 44109
2 105319 1 44109
2 105320 1 44134
2 105321 1 44134
2 105322 1 44136
2 105323 1 44136
2 105324 1 44140
2 105325 1 44140
2 105326 1 44141
2 105327 1 44141
2 105328 1 44141
2 105329 1 44141
2 105330 1 44144
2 105331 1 44144
2 105332 1 44166
2 105333 1 44166
2 105334 1 44166
2 105335 1 44204
2 105336 1 44204
2 105337 1 44217
2 105338 1 44217
2 105339 1 44217
2 105340 1 44222
2 105341 1 44222
2 105342 1 44246
2 105343 1 44246
2 105344 1 44246
2 105345 1 44247
2 105346 1 44247
2 105347 1 44247
2 105348 1 44250
2 105349 1 44250
2 105350 1 44251
2 105351 1 44251
2 105352 1 44254
2 105353 1 44254
2 105354 1 44277
2 105355 1 44277
2 105356 1 44303
2 105357 1 44303
2 105358 1 44303
2 105359 1 44316
2 105360 1 44316
2 105361 1 44320
2 105362 1 44320
2 105363 1 44330
2 105364 1 44330
2 105365 1 44331
2 105366 1 44331
2 105367 1 44348
2 105368 1 44348
2 105369 1 44356
2 105370 1 44356
2 105371 1 44356
2 105372 1 44391
2 105373 1 44391
2 105374 1 44405
2 105375 1 44405
2 105376 1 44418
2 105377 1 44418
2 105378 1 44418
2 105379 1 44423
2 105380 1 44423
2 105381 1 44443
2 105382 1 44443
2 105383 1 44471
2 105384 1 44471
2 105385 1 44480
2 105386 1 44480
2 105387 1 44480
2 105388 1 44488
2 105389 1 44488
2 105390 1 44507
2 105391 1 44507
2 105392 1 44508
2 105393 1 44508
2 105394 1 44508
2 105395 1 44523
2 105396 1 44523
2 105397 1 44611
2 105398 1 44611
2 105399 1 44623
2 105400 1 44623
2 105401 1 44677
2 105402 1 44677
2 105403 1 44695
2 105404 1 44695
2 105405 1 44703
2 105406 1 44703
2 105407 1 44713
2 105408 1 44713
2 105409 1 44731
2 105410 1 44731
2 105411 1 44807
2 105412 1 44807
2 105413 1 44816
2 105414 1 44816
2 105415 1 44877
2 105416 1 44877
2 105417 1 44894
2 105418 1 44894
2 105419 1 44908
2 105420 1 44908
2 105421 1 44938
2 105422 1 44938
2 105423 1 44972
2 105424 1 44972
2 105425 1 44972
2 105426 1 44975
2 105427 1 44975
2 105428 1 44999
2 105429 1 44999
2 105430 1 45061
2 105431 1 45061
2 105432 1 45073
2 105433 1 45073
2 105434 1 45088
2 105435 1 45088
2 105436 1 45109
2 105437 1 45109
2 105438 1 45117
2 105439 1 45117
2 105440 1 45144
2 105441 1 45144
2 105442 1 45145
2 105443 1 45145
2 105444 1 45187
2 105445 1 45187
2 105446 1 45189
2 105447 1 45189
2 105448 1 45191
2 105449 1 45191
2 105450 1 45191
2 105451 1 45192
2 105452 1 45192
2 105453 1 45230
2 105454 1 45230
2 105455 1 45260
2 105456 1 45260
2 105457 1 45268
2 105458 1 45268
2 105459 1 45282
2 105460 1 45282
2 105461 1 45284
2 105462 1 45284
2 105463 1 45284
2 105464 1 45285
2 105465 1 45285
2 105466 1 45286
2 105467 1 45286
2 105468 1 45286
2 105469 1 45288
2 105470 1 45288
2 105471 1 45298
2 105472 1 45298
2 105473 1 45306
2 105474 1 45306
2 105475 1 45314
2 105476 1 45314
2 105477 1 45316
2 105478 1 45316
2 105479 1 45325
2 105480 1 45325
2 105481 1 45355
2 105482 1 45355
2 105483 1 45355
2 105484 1 45355
2 105485 1 45355
2 105486 1 45365
2 105487 1 45365
2 105488 1 45375
2 105489 1 45375
2 105490 1 45375
2 105491 1 45385
2 105492 1 45385
2 105493 1 45388
2 105494 1 45388
2 105495 1 45390
2 105496 1 45390
2 105497 1 45398
2 105498 1 45398
2 105499 1 45402
2 105500 1 45402
2 105501 1 45410
2 105502 1 45410
2 105503 1 45439
2 105504 1 45439
2 105505 1 45454
2 105506 1 45454
2 105507 1 45457
2 105508 1 45457
2 105509 1 45475
2 105510 1 45475
2 105511 1 45509
2 105512 1 45509
2 105513 1 45519
2 105514 1 45519
2 105515 1 45531
2 105516 1 45531
2 105517 1 45554
2 105518 1 45554
2 105519 1 45554
2 105520 1 45555
2 105521 1 45555
2 105522 1 45564
2 105523 1 45564
2 105524 1 45582
2 105525 1 45582
2 105526 1 45583
2 105527 1 45583
2 105528 1 45583
2 105529 1 45583
2 105530 1 45591
2 105531 1 45591
2 105532 1 45591
2 105533 1 45598
2 105534 1 45598
2 105535 1 45635
2 105536 1 45635
2 105537 1 45636
2 105538 1 45636
2 105539 1 45636
2 105540 1 45656
2 105541 1 45656
2 105542 1 45661
2 105543 1 45661
2 105544 1 45661
2 105545 1 45670
2 105546 1 45670
2 105547 1 45681
2 105548 1 45681
2 105549 1 45700
2 105550 1 45700
2 105551 1 45715
2 105552 1 45715
2 105553 1 45715
2 105554 1 45715
2 105555 1 45722
2 105556 1 45722
2 105557 1 45722
2 105558 1 45723
2 105559 1 45723
2 105560 1 45727
2 105561 1 45727
2 105562 1 45733
2 105563 1 45733
2 105564 1 45761
2 105565 1 45761
2 105566 1 45777
2 105567 1 45777
2 105568 1 45830
2 105569 1 45830
2 105570 1 45837
2 105571 1 45837
2 105572 1 45920
2 105573 1 45920
2 105574 1 45923
2 105575 1 45923
2 105576 1 45932
2 105577 1 45932
2 105578 1 45944
2 105579 1 45944
2 105580 1 46008
2 105581 1 46008
2 105582 1 46051
2 105583 1 46051
2 105584 1 46067
2 105585 1 46067
2 105586 1 46080
2 105587 1 46080
2 105588 1 46092
2 105589 1 46092
2 105590 1 46108
2 105591 1 46108
2 105592 1 46108
2 105593 1 46108
2 105594 1 46109
2 105595 1 46109
2 105596 1 46109
2 105597 1 46143
2 105598 1 46143
2 105599 1 46207
2 105600 1 46207
2 105601 1 46291
2 105602 1 46291
2 105603 1 46322
2 105604 1 46322
2 105605 1 46322
2 105606 1 46360
2 105607 1 46360
2 105608 1 46360
2 105609 1 46360
2 105610 1 46384
2 105611 1 46384
2 105612 1 46418
2 105613 1 46418
2 105614 1 46437
2 105615 1 46437
2 105616 1 46448
2 105617 1 46448
2 105618 1 46448
2 105619 1 46448
2 105620 1 46449
2 105621 1 46449
2 105622 1 46449
2 105623 1 46467
2 105624 1 46467
2 105625 1 46467
2 105626 1 46470
2 105627 1 46470
2 105628 1 46475
2 105629 1 46475
2 105630 1 46479
2 105631 1 46479
2 105632 1 46479
2 105633 1 46492
2 105634 1 46492
2 105635 1 46492
2 105636 1 46502
2 105637 1 46502
2 105638 1 46502
2 105639 1 46502
2 105640 1 46510
2 105641 1 46510
2 105642 1 46510
2 105643 1 46511
2 105644 1 46511
2 105645 1 46520
2 105646 1 46520
2 105647 1 46520
2 105648 1 46520
2 105649 1 46521
2 105650 1 46521
2 105651 1 46537
2 105652 1 46537
2 105653 1 46593
2 105654 1 46593
2 105655 1 46594
2 105656 1 46594
2 105657 1 46594
2 105658 1 46594
2 105659 1 46626
2 105660 1 46626
2 105661 1 46626
2 105662 1 46626
2 105663 1 46664
2 105664 1 46664
2 105665 1 46667
2 105666 1 46667
2 105667 1 46667
2 105668 1 46667
2 105669 1 46667
2 105670 1 46667
2 105671 1 46670
2 105672 1 46670
2 105673 1 46679
2 105674 1 46679
2 105675 1 46707
2 105676 1 46707
2 105677 1 46714
2 105678 1 46714
2 105679 1 46716
2 105680 1 46716
2 105681 1 46716
2 105682 1 46732
2 105683 1 46732
2 105684 1 46745
2 105685 1 46745
2 105686 1 46777
2 105687 1 46777
2 105688 1 46777
2 105689 1 46777
2 105690 1 46810
2 105691 1 46810
2 105692 1 46854
2 105693 1 46854
2 105694 1 46875
2 105695 1 46875
2 105696 1 46887
2 105697 1 46887
2 105698 1 46887
2 105699 1 46914
2 105700 1 46914
2 105701 1 46996
2 105702 1 46996
2 105703 1 47015
2 105704 1 47015
2 105705 1 47016
2 105706 1 47016
2 105707 1 47022
2 105708 1 47022
2 105709 1 47022
2 105710 1 47024
2 105711 1 47024
2 105712 1 47025
2 105713 1 47025
2 105714 1 47044
2 105715 1 47044
2 105716 1 47070
2 105717 1 47070
2 105718 1 47097
2 105719 1 47097
2 105720 1 47111
2 105721 1 47111
2 105722 1 47129
2 105723 1 47129
2 105724 1 47129
2 105725 1 47130
2 105726 1 47130
2 105727 1 47132
2 105728 1 47132
2 105729 1 47142
2 105730 1 47142
2 105731 1 47142
2 105732 1 47186
2 105733 1 47186
2 105734 1 47191
2 105735 1 47191
2 105736 1 47195
2 105737 1 47195
2 105738 1 47208
2 105739 1 47208
2 105740 1 47220
2 105741 1 47220
2 105742 1 47234
2 105743 1 47234
2 105744 1 47238
2 105745 1 47238
2 105746 1 47273
2 105747 1 47273
2 105748 1 47300
2 105749 1 47300
2 105750 1 47324
2 105751 1 47324
2 105752 1 47324
2 105753 1 47327
2 105754 1 47327
2 105755 1 47327
2 105756 1 47331
2 105757 1 47331
2 105758 1 47331
2 105759 1 47366
2 105760 1 47366
2 105761 1 47490
2 105762 1 47490
2 105763 1 47518
2 105764 1 47518
2 105765 1 47518
2 105766 1 47518
2 105767 1 47522
2 105768 1 47522
2 105769 1 47545
2 105770 1 47545
2 105771 1 47545
2 105772 1 47567
2 105773 1 47567
2 105774 1 47568
2 105775 1 47568
2 105776 1 47570
2 105777 1 47570
2 105778 1 47571
2 105779 1 47571
2 105780 1 47571
2 105781 1 47572
2 105782 1 47572
2 105783 1 47600
2 105784 1 47600
2 105785 1 47610
2 105786 1 47610
2 105787 1 47618
2 105788 1 47618
2 105789 1 47618
2 105790 1 47619
2 105791 1 47619
2 105792 1 47620
2 105793 1 47620
2 105794 1 47648
2 105795 1 47648
2 105796 1 47650
2 105797 1 47650
2 105798 1 47671
2 105799 1 47671
2 105800 1 47674
2 105801 1 47674
2 105802 1 47674
2 105803 1 47696
2 105804 1 47696
2 105805 1 47700
2 105806 1 47700
2 105807 1 47701
2 105808 1 47701
2 105809 1 47716
2 105810 1 47716
2 105811 1 47756
2 105812 1 47756
2 105813 1 47756
2 105814 1 47793
2 105815 1 47793
2 105816 1 47795
2 105817 1 47795
2 105818 1 47795
2 105819 1 47795
2 105820 1 47806
2 105821 1 47806
2 105822 1 47806
2 105823 1 47822
2 105824 1 47822
2 105825 1 47832
2 105826 1 47832
2 105827 1 47846
2 105828 1 47846
2 105829 1 47861
2 105830 1 47861
2 105831 1 47862
2 105832 1 47862
2 105833 1 47862
2 105834 1 47862
2 105835 1 47873
2 105836 1 47873
2 105837 1 47874
2 105838 1 47874
2 105839 1 47926
2 105840 1 47926
2 105841 1 47966
2 105842 1 47966
2 105843 1 47976
2 105844 1 47976
2 105845 1 47979
2 105846 1 47979
2 105847 1 47980
2 105848 1 47980
2 105849 1 47980
2 105850 1 47983
2 105851 1 47983
2 105852 1 47994
2 105853 1 47994
2 105854 1 47995
2 105855 1 47995
2 105856 1 47995
2 105857 1 47995
2 105858 1 48015
2 105859 1 48015
2 105860 1 48015
2 105861 1 48021
2 105862 1 48021
2 105863 1 48072
2 105864 1 48072
2 105865 1 48072
2 105866 1 48098
2 105867 1 48098
2 105868 1 48099
2 105869 1 48099
2 105870 1 48123
2 105871 1 48123
2 105872 1 48126
2 105873 1 48126
2 105874 1 48139
2 105875 1 48139
2 105876 1 48159
2 105877 1 48159
2 105878 1 48186
2 105879 1 48186
2 105880 1 48186
2 105881 1 48194
2 105882 1 48194
2 105883 1 48204
2 105884 1 48204
2 105885 1 48237
2 105886 1 48237
2 105887 1 48237
2 105888 1 48237
2 105889 1 48325
2 105890 1 48325
2 105891 1 48366
2 105892 1 48366
2 105893 1 48373
2 105894 1 48373
2 105895 1 48396
2 105896 1 48396
2 105897 1 48396
2 105898 1 48396
2 105899 1 48396
2 105900 1 48396
2 105901 1 48398
2 105902 1 48398
2 105903 1 48398
2 105904 1 48413
2 105905 1 48413
2 105906 1 48427
2 105907 1 48427
2 105908 1 48432
2 105909 1 48432
2 105910 1 48432
2 105911 1 48432
2 105912 1 48438
2 105913 1 48438
2 105914 1 48456
2 105915 1 48456
2 105916 1 48456
2 105917 1 48456
2 105918 1 48457
2 105919 1 48457
2 105920 1 48475
2 105921 1 48475
2 105922 1 48492
2 105923 1 48492
2 105924 1 48499
2 105925 1 48499
2 105926 1 48662
2 105927 1 48662
2 105928 1 48670
2 105929 1 48670
2 105930 1 48670
2 105931 1 48670
2 105932 1 48670
2 105933 1 48671
2 105934 1 48671
2 105935 1 48690
2 105936 1 48690
2 105937 1 48759
2 105938 1 48759
2 105939 1 48788
2 105940 1 48788
2 105941 1 48814
2 105942 1 48814
2 105943 1 48822
2 105944 1 48822
2 105945 1 48857
2 105946 1 48857
2 105947 1 48871
2 105948 1 48871
2 105949 1 48871
2 105950 1 48921
2 105951 1 48921
2 105952 1 48942
2 105953 1 48942
2 105954 1 48951
2 105955 1 48951
2 105956 1 48957
2 105957 1 48957
2 105958 1 48965
2 105959 1 48965
2 105960 1 48965
2 105961 1 48966
2 105962 1 48966
2 105963 1 48975
2 105964 1 48975
2 105965 1 48998
2 105966 1 48998
2 105967 1 49007
2 105968 1 49007
2 105969 1 49008
2 105970 1 49008
2 105971 1 49008
2 105972 1 49010
2 105973 1 49010
2 105974 1 49011
2 105975 1 49011
2 105976 1 49019
2 105977 1 49019
2 105978 1 49020
2 105979 1 49020
2 105980 1 49020
2 105981 1 49021
2 105982 1 49021
2 105983 1 49034
2 105984 1 49034
2 105985 1 49041
2 105986 1 49041
2 105987 1 49042
2 105988 1 49042
2 105989 1 49076
2 105990 1 49076
2 105991 1 49090
2 105992 1 49090
2 105993 1 49126
2 105994 1 49126
2 105995 1 49135
2 105996 1 49135
2 105997 1 49145
2 105998 1 49145
2 105999 1 49151
2 106000 1 49151
2 106001 1 49162
2 106002 1 49162
2 106003 1 49171
2 106004 1 49171
2 106005 1 49181
2 106006 1 49181
2 106007 1 49213
2 106008 1 49213
2 106009 1 49240
2 106010 1 49240
2 106011 1 49250
2 106012 1 49250
2 106013 1 49265
2 106014 1 49265
2 106015 1 49269
2 106016 1 49269
2 106017 1 49280
2 106018 1 49280
2 106019 1 49292
2 106020 1 49292
2 106021 1 49293
2 106022 1 49293
2 106023 1 49320
2 106024 1 49320
2 106025 1 49331
2 106026 1 49331
2 106027 1 49347
2 106028 1 49347
2 106029 1 49360
2 106030 1 49360
2 106031 1 49361
2 106032 1 49361
2 106033 1 49364
2 106034 1 49364
2 106035 1 49388
2 106036 1 49388
2 106037 1 49391
2 106038 1 49391
2 106039 1 49404
2 106040 1 49404
2 106041 1 49417
2 106042 1 49417
2 106043 1 49424
2 106044 1 49424
2 106045 1 49433
2 106046 1 49433
2 106047 1 49434
2 106048 1 49434
2 106049 1 49443
2 106050 1 49443
2 106051 1 49453
2 106052 1 49453
2 106053 1 49465
2 106054 1 49465
2 106055 1 49483
2 106056 1 49483
2 106057 1 49502
2 106058 1 49502
2 106059 1 49509
2 106060 1 49509
2 106061 1 49518
2 106062 1 49518
2 106063 1 49519
2 106064 1 49519
2 106065 1 49526
2 106066 1 49526
2 106067 1 49548
2 106068 1 49548
2 106069 1 49549
2 106070 1 49549
2 106071 1 49552
2 106072 1 49552
2 106073 1 49553
2 106074 1 49553
2 106075 1 49554
2 106076 1 49554
2 106077 1 49561
2 106078 1 49561
2 106079 1 49564
2 106080 1 49564
2 106081 1 49596
2 106082 1 49596
2 106083 1 49599
2 106084 1 49599
2 106085 1 49600
2 106086 1 49600
2 106087 1 49607
2 106088 1 49607
2 106089 1 49616
2 106090 1 49616
2 106091 1 49634
2 106092 1 49634
2 106093 1 49670
2 106094 1 49670
2 106095 1 49686
2 106096 1 49686
2 106097 1 49693
2 106098 1 49693
2 106099 1 49706
2 106100 1 49706
2 106101 1 49722
2 106102 1 49722
2 106103 1 49739
2 106104 1 49739
2 106105 1 49749
2 106106 1 49749
2 106107 1 49758
2 106108 1 49758
2 106109 1 49759
2 106110 1 49759
2 106111 1 49766
2 106112 1 49766
2 106113 1 49771
2 106114 1 49771
2 106115 1 49806
2 106116 1 49806
2 106117 1 49825
2 106118 1 49825
2 106119 1 49826
2 106120 1 49826
2 106121 1 49842
2 106122 1 49842
2 106123 1 49984
2 106124 1 49984
2 106125 1 49991
2 106126 1 49991
2 106127 1 50057
2 106128 1 50057
2 106129 1 50057
2 106130 1 50135
2 106131 1 50135
2 106132 1 50135
2 106133 1 50135
2 106134 1 50135
2 106135 1 50220
2 106136 1 50220
2 106137 1 50327
2 106138 1 50327
2 106139 1 50333
2 106140 1 50333
2 106141 1 50404
2 106142 1 50404
2 106143 1 50445
2 106144 1 50445
2 106145 1 50445
2 106146 1 50522
2 106147 1 50522
2 106148 1 50535
2 106149 1 50535
2 106150 1 50536
2 106151 1 50536
2 106152 1 50541
2 106153 1 50541
2 106154 1 50648
2 106155 1 50648
2 106156 1 50674
2 106157 1 50674
2 106158 1 50678
2 106159 1 50678
2 106160 1 50682
2 106161 1 50682
2 106162 1 50709
2 106163 1 50709
2 106164 1 50726
2 106165 1 50726
2 106166 1 50753
2 106167 1 50753
2 106168 1 50754
2 106169 1 50754
2 106170 1 50784
2 106171 1 50784
2 106172 1 50805
2 106173 1 50805
2 106174 1 50839
2 106175 1 50839
2 106176 1 50856
2 106177 1 50856
2 106178 1 50856
2 106179 1 50889
2 106180 1 50889
2 106181 1 50910
2 106182 1 50910
2 106183 1 50936
2 106184 1 50936
2 106185 1 50939
2 106186 1 50939
2 106187 1 50960
2 106188 1 50960
2 106189 1 50971
2 106190 1 50971
2 106191 1 50973
2 106192 1 50973
2 106193 1 51009
2 106194 1 51009
2 106195 1 51012
2 106196 1 51012
2 106197 1 51012
2 106198 1 51025
2 106199 1 51025
2 106200 1 51059
2 106201 1 51059
2 106202 1 51119
2 106203 1 51119
2 106204 1 51120
2 106205 1 51120
2 106206 1 51122
2 106207 1 51122
2 106208 1 51151
2 106209 1 51151
2 106210 1 51192
2 106211 1 51192
2 106212 1 51193
2 106213 1 51193
2 106214 1 51193
2 106215 1 51193
2 106216 1 51193
2 106217 1 51194
2 106218 1 51194
2 106219 1 51194
2 106220 1 51196
2 106221 1 51196
2 106222 1 51196
2 106223 1 51196
2 106224 1 51196
2 106225 1 51196
2 106226 1 51196
2 106227 1 51226
2 106228 1 51226
2 106229 1 51227
2 106230 1 51227
2 106231 1 51228
2 106232 1 51228
2 106233 1 51245
2 106234 1 51245
2 106235 1 51245
2 106236 1 51245
2 106237 1 51245
2 106238 1 51245
2 106239 1 51248
2 106240 1 51248
2 106241 1 51254
2 106242 1 51254
2 106243 1 51254
2 106244 1 51261
2 106245 1 51261
2 106246 1 51261
2 106247 1 51300
2 106248 1 51300
2 106249 1 51300
2 106250 1 51343
2 106251 1 51343
2 106252 1 51370
2 106253 1 51370
2 106254 1 51410
2 106255 1 51410
2 106256 1 51452
2 106257 1 51452
2 106258 1 51462
2 106259 1 51462
2 106260 1 51485
2 106261 1 51485
2 106262 1 51496
2 106263 1 51496
2 106264 1 51496
2 106265 1 51506
2 106266 1 51506
2 106267 1 51515
2 106268 1 51515
2 106269 1 51527
2 106270 1 51527
2 106271 1 51530
2 106272 1 51530
2 106273 1 51530
2 106274 1 51541
2 106275 1 51541
2 106276 1 51548
2 106277 1 51548
2 106278 1 51548
2 106279 1 51548
2 106280 1 51551
2 106281 1 51551
2 106282 1 51604
2 106283 1 51604
2 106284 1 51612
2 106285 1 51612
2 106286 1 51647
2 106287 1 51647
2 106288 1 51656
2 106289 1 51656
2 106290 1 51677
2 106291 1 51677
2 106292 1 51684
2 106293 1 51684
2 106294 1 51686
2 106295 1 51686
2 106296 1 51738
2 106297 1 51738
2 106298 1 51761
2 106299 1 51761
2 106300 1 51774
2 106301 1 51774
2 106302 1 51774
2 106303 1 51808
2 106304 1 51808
2 106305 1 51827
2 106306 1 51827
2 106307 1 51835
2 106308 1 51835
2 106309 1 51868
2 106310 1 51868
2 106311 1 51875
2 106312 1 51875
2 106313 1 51884
2 106314 1 51884
2 106315 1 51902
2 106316 1 51902
2 106317 1 51938
2 106318 1 51938
2 106319 1 51996
2 106320 1 51996
2 106321 1 52049
2 106322 1 52049
2 106323 1 52059
2 106324 1 52059
2 106325 1 52080
2 106326 1 52080
2 106327 1 52095
2 106328 1 52095
2 106329 1 52102
2 106330 1 52102
2 106331 1 52114
2 106332 1 52114
2 106333 1 52115
2 106334 1 52115
2 106335 1 52123
2 106336 1 52123
2 106337 1 52264
2 106338 1 52264
2 106339 1 52271
2 106340 1 52271
2 106341 1 52280
2 106342 1 52280
2 106343 1 52288
2 106344 1 52288
2 106345 1 52291
2 106346 1 52291
2 106347 1 52306
2 106348 1 52306
2 106349 1 52367
2 106350 1 52367
2 106351 1 52367
2 106352 1 52367
2 106353 1 52367
2 106354 1 52371
2 106355 1 52371
2 106356 1 52371
2 106357 1 52371
2 106358 1 52387
2 106359 1 52387
2 106360 1 52391
2 106361 1 52391
2 106362 1 52460
2 106363 1 52460
2 106364 1 52474
2 106365 1 52474
2 106366 1 52476
2 106367 1 52476
2 106368 1 52476
2 106369 1 52479
2 106370 1 52479
2 106371 1 52482
2 106372 1 52482
2 106373 1 52490
2 106374 1 52490
2 106375 1 52557
2 106376 1 52557
2 106377 1 52558
2 106378 1 52558
2 106379 1 52558
2 106380 1 52558
2 106381 1 52585
2 106382 1 52585
2 106383 1 52611
2 106384 1 52611
2 106385 1 52628
2 106386 1 52628
2 106387 1 52628
2 106388 1 52628
2 106389 1 52645
2 106390 1 52645
2 106391 1 52649
2 106392 1 52649
2 106393 1 52651
2 106394 1 52651
2 106395 1 52661
2 106396 1 52661
2 106397 1 52661
2 106398 1 52672
2 106399 1 52672
2 106400 1 52708
2 106401 1 52708
2 106402 1 52716
2 106403 1 52716
2 106404 1 52725
2 106405 1 52725
2 106406 1 52725
2 106407 1 52725
2 106408 1 52726
2 106409 1 52726
2 106410 1 52734
2 106411 1 52734
2 106412 1 52744
2 106413 1 52744
2 106414 1 52754
2 106415 1 52754
2 106416 1 52754
2 106417 1 52788
2 106418 1 52788
2 106419 1 52818
2 106420 1 52818
2 106421 1 52818
2 106422 1 52851
2 106423 1 52851
2 106424 1 52852
2 106425 1 52852
2 106426 1 52855
2 106427 1 52855
2 106428 1 52856
2 106429 1 52856
2 106430 1 52861
2 106431 1 52861
2 106432 1 52900
2 106433 1 52900
2 106434 1 52914
2 106435 1 52914
2 106436 1 52915
2 106437 1 52915
2 106438 1 52915
2 106439 1 52932
2 106440 1 52932
2 106441 1 52986
2 106442 1 52986
2 106443 1 52987
2 106444 1 52987
2 106445 1 52987
2 106446 1 52987
2 106447 1 52987
2 106448 1 52995
2 106449 1 52995
2 106450 1 52996
2 106451 1 52996
2 106452 1 52996
2 106453 1 53017
2 106454 1 53017
2 106455 1 53019
2 106456 1 53019
2 106457 1 53127
2 106458 1 53127
2 106459 1 53142
2 106460 1 53142
2 106461 1 53151
2 106462 1 53151
2 106463 1 53151
2 106464 1 53151
2 106465 1 53151
2 106466 1 53187
2 106467 1 53187
2 106468 1 53188
2 106469 1 53188
2 106470 1 53198
2 106471 1 53198
2 106472 1 53265
2 106473 1 53265
2 106474 1 53265
2 106475 1 53265
2 106476 1 53275
2 106477 1 53275
2 106478 1 53323
2 106479 1 53323
2 106480 1 53378
2 106481 1 53378
2 106482 1 53379
2 106483 1 53379
2 106484 1 53396
2 106485 1 53396
2 106486 1 53408
2 106487 1 53408
2 106488 1 53408
2 106489 1 53423
2 106490 1 53423
2 106491 1 53424
2 106492 1 53424
2 106493 1 53444
2 106494 1 53444
2 106495 1 53447
2 106496 1 53447
2 106497 1 53468
2 106498 1 53468
2 106499 1 53479
2 106500 1 53479
2 106501 1 53489
2 106502 1 53489
2 106503 1 53542
2 106504 1 53542
2 106505 1 53568
2 106506 1 53568
2 106507 1 53603
2 106508 1 53603
2 106509 1 53660
2 106510 1 53660
2 106511 1 53660
2 106512 1 53682
2 106513 1 53682
2 106514 1 53685
2 106515 1 53685
2 106516 1 53685
2 106517 1 53710
2 106518 1 53710
2 106519 1 53737
2 106520 1 53737
2 106521 1 53745
2 106522 1 53745
2 106523 1 53745
2 106524 1 53771
2 106525 1 53771
2 106526 1 53783
2 106527 1 53783
2 106528 1 53808
2 106529 1 53808
2 106530 1 53814
2 106531 1 53814
2 106532 1 53817
2 106533 1 53817
2 106534 1 53817
2 106535 1 53837
2 106536 1 53837
2 106537 1 53838
2 106538 1 53838
2 106539 1 53840
2 106540 1 53840
2 106541 1 53844
2 106542 1 53844
2 106543 1 53869
2 106544 1 53869
2 106545 1 53872
2 106546 1 53872
2 106547 1 53872
2 106548 1 53904
2 106549 1 53904
2 106550 1 53915
2 106551 1 53915
2 106552 1 53921
2 106553 1 53921
2 106554 1 53939
2 106555 1 53939
2 106556 1 53939
2 106557 1 53939
2 106558 1 53939
2 106559 1 53939
2 106560 1 53941
2 106561 1 53941
2 106562 1 53994
2 106563 1 53994
2 106564 1 54009
2 106565 1 54009
2 106566 1 54018
2 106567 1 54018
2 106568 1 54024
2 106569 1 54024
2 106570 1 54029
2 106571 1 54029
2 106572 1 54139
2 106573 1 54139
2 106574 1 54253
2 106575 1 54253
2 106576 1 54453
2 106577 1 54453
2 106578 1 54541
2 106579 1 54541
2 106580 1 54541
2 106581 1 54558
2 106582 1 54558
2 106583 1 54576
2 106584 1 54576
2 106585 1 54684
2 106586 1 54684
2 106587 1 54701
2 106588 1 54701
2 106589 1 54701
2 106590 1 54767
2 106591 1 54767
2 106592 1 54936
2 106593 1 54936
2 106594 1 55034
2 106595 1 55034
2 106596 1 55046
2 106597 1 55046
2 106598 1 55074
2 106599 1 55074
2 106600 1 55074
2 106601 1 55139
2 106602 1 55139
2 106603 1 55162
2 106604 1 55162
2 106605 1 55162
2 106606 1 55162
2 106607 1 55177
2 106608 1 55177
2 106609 1 55214
2 106610 1 55214
2 106611 1 55244
2 106612 1 55244
2 106613 1 55250
2 106614 1 55250
2 106615 1 55256
2 106616 1 55256
2 106617 1 55263
2 106618 1 55263
2 106619 1 55286
2 106620 1 55286
2 106621 1 55361
2 106622 1 55361
2 106623 1 55361
2 106624 1 55361
2 106625 1 55362
2 106626 1 55362
2 106627 1 55362
2 106628 1 55366
2 106629 1 55366
2 106630 1 55530
2 106631 1 55530
2 106632 1 55530
2 106633 1 55530
2 106634 1 55538
2 106635 1 55538
2 106636 1 55539
2 106637 1 55539
2 106638 1 55681
2 106639 1 55681
2 106640 1 55729
2 106641 1 55729
2 106642 1 55840
2 106643 1 55840
2 106644 1 55840
2 106645 1 55840
2 106646 1 55840
2 106647 1 55840
2 106648 1 55840
2 106649 1 55840
2 106650 1 55840
2 106651 1 55840
2 106652 1 55840
2 106653 1 55840
2 106654 1 55840
2 106655 1 55840
2 106656 1 55840
2 106657 1 55840
2 106658 1 55840
2 106659 1 55840
2 106660 1 55840
2 106661 1 55840
2 106662 1 55840
2 106663 1 55840
2 106664 1 55840
2 106665 1 55840
2 106666 1 55840
2 106667 1 55840
2 106668 1 55840
2 106669 1 55840
2 106670 1 55850
2 106671 1 55850
2 106672 1 55868
2 106673 1 55868
2 106674 1 55878
2 106675 1 55878
2 106676 1 55878
2 106677 1 55878
2 106678 1 55878
2 106679 1 55879
2 106680 1 55879
2 106681 1 55885
2 106682 1 55885
2 106683 1 55907
2 106684 1 55907
2 106685 1 55925
2 106686 1 55925
2 106687 1 55939
2 106688 1 55939
2 106689 1 55970
2 106690 1 55970
2 106691 1 56014
2 106692 1 56014
2 106693 1 56021
2 106694 1 56021
2 106695 1 56030
2 106696 1 56030
2 106697 1 56051
2 106698 1 56051
2 106699 1 56106
2 106700 1 56106
2 106701 1 56113
2 106702 1 56113
2 106703 1 56114
2 106704 1 56114
2 106705 1 56118
2 106706 1 56118
2 106707 1 56150
2 106708 1 56150
2 106709 1 56152
2 106710 1 56152
2 106711 1 56191
2 106712 1 56191
2 106713 1 56225
2 106714 1 56225
2 106715 1 56225
2 106716 1 56225
2 106717 1 56226
2 106718 1 56226
2 106719 1 56229
2 106720 1 56229
2 106721 1 56230
2 106722 1 56230
2 106723 1 56247
2 106724 1 56247
2 106725 1 56248
2 106726 1 56248
2 106727 1 56249
2 106728 1 56249
2 106729 1 56249
2 106730 1 56258
2 106731 1 56258
2 106732 1 56271
2 106733 1 56271
2 106734 1 56271
2 106735 1 56283
2 106736 1 56283
2 106737 1 56287
2 106738 1 56287
2 106739 1 56287
2 106740 1 56287
2 106741 1 56287
2 106742 1 56287
2 106743 1 56287
2 106744 1 56296
2 106745 1 56296
2 106746 1 56298
2 106747 1 56298
2 106748 1 56306
2 106749 1 56306
2 106750 1 56307
2 106751 1 56307
2 106752 1 56343
2 106753 1 56343
2 106754 1 56343
2 106755 1 56354
2 106756 1 56354
2 106757 1 56420
2 106758 1 56420
2 106759 1 56434
2 106760 1 56434
2 106761 1 56435
2 106762 1 56435
2 106763 1 56444
2 106764 1 56444
2 106765 1 56455
2 106766 1 56455
2 106767 1 56455
2 106768 1 56485
2 106769 1 56485
2 106770 1 56506
2 106771 1 56506
2 106772 1 56506
2 106773 1 56519
2 106774 1 56519
2 106775 1 56521
2 106776 1 56521
2 106777 1 56581
2 106778 1 56581
2 106779 1 56581
2 106780 1 56581
2 106781 1 56609
2 106782 1 56609
2 106783 1 56630
2 106784 1 56630
2 106785 1 56630
2 106786 1 56630
2 106787 1 56630
2 106788 1 56630
2 106789 1 56630
2 106790 1 56630
2 106791 1 56630
2 106792 1 56630
2 106793 1 56649
2 106794 1 56649
2 106795 1 56659
2 106796 1 56659
2 106797 1 56662
2 106798 1 56662
2 106799 1 56677
2 106800 1 56677
2 106801 1 56721
2 106802 1 56721
2 106803 1 56741
2 106804 1 56741
2 106805 1 56748
2 106806 1 56748
2 106807 1 56748
2 106808 1 56749
2 106809 1 56749
2 106810 1 56760
2 106811 1 56760
2 106812 1 56771
2 106813 1 56771
2 106814 1 56793
2 106815 1 56793
2 106816 1 56972
2 106817 1 56972
2 106818 1 57012
2 106819 1 57012
2 106820 1 57024
2 106821 1 57024
2 106822 1 57050
2 106823 1 57050
2 106824 1 57146
2 106825 1 57146
2 106826 1 57147
2 106827 1 57147
2 106828 1 57170
2 106829 1 57170
2 106830 1 57178
2 106831 1 57178
2 106832 1 57202
2 106833 1 57202
2 106834 1 57223
2 106835 1 57223
2 106836 1 57223
2 106837 1 57223
2 106838 1 57267
2 106839 1 57267
2 106840 1 57274
2 106841 1 57274
2 106842 1 57276
2 106843 1 57276
2 106844 1 57445
2 106845 1 57445
2 106846 1 57493
2 106847 1 57493
2 106848 1 57527
2 106849 1 57527
2 106850 1 57528
2 106851 1 57528
2 106852 1 57545
2 106853 1 57545
2 106854 1 57559
2 106855 1 57559
2 106856 1 57572
2 106857 1 57572
2 106858 1 57579
2 106859 1 57579
2 106860 1 57580
2 106861 1 57580
2 106862 1 57612
2 106863 1 57612
2 106864 1 57623
2 106865 1 57623
2 106866 1 57634
2 106867 1 57634
2 106868 1 57634
2 106869 1 57647
2 106870 1 57647
2 106871 1 57670
2 106872 1 57670
2 106873 1 57679
2 106874 1 57679
2 106875 1 57690
2 106876 1 57690
2 106877 1 57701
2 106878 1 57701
2 106879 1 57715
2 106880 1 57715
2 106881 1 57722
2 106882 1 57722
2 106883 1 57810
2 106884 1 57810
2 106885 1 57810
2 106886 1 58019
2 106887 1 58019
2 106888 1 58190
2 106889 1 58190
2 106890 1 58278
2 106891 1 58278
2 106892 1 58360
2 106893 1 58360
2 106894 1 58365
2 106895 1 58365
2 106896 1 58377
2 106897 1 58377
2 106898 1 58387
2 106899 1 58387
2 106900 1 58404
2 106901 1 58404
2 106902 1 58434
2 106903 1 58434
2 106904 1 58501
2 106905 1 58501
2 106906 1 58537
2 106907 1 58537
2 106908 1 58540
2 106909 1 58540
2 106910 1 58563
2 106911 1 58563
2 106912 1 58564
2 106913 1 58564
2 106914 1 58566
2 106915 1 58566
2 106916 1 58573
2 106917 1 58573
2 106918 1 58573
2 106919 1 58573
2 106920 1 58573
2 106921 1 58573
2 106922 1 58574
2 106923 1 58574
2 106924 1 58574
2 106925 1 58574
2 106926 1 58581
2 106927 1 58581
2 106928 1 58581
2 106929 1 58581
2 106930 1 58584
2 106931 1 58584
2 106932 1 58584
2 106933 1 58584
2 106934 1 58584
2 106935 1 58584
2 106936 1 58584
2 106937 1 58584
2 106938 1 58584
2 106939 1 58585
2 106940 1 58585
2 106941 1 58585
2 106942 1 58585
2 106943 1 58585
2 106944 1 58639
2 106945 1 58639
2 106946 1 58639
2 106947 1 58639
2 106948 1 58639
2 106949 1 58639
2 106950 1 58639
2 106951 1 58639
2 106952 1 58639
2 106953 1 58639
2 106954 1 58639
2 106955 1 58639
2 106956 1 58639
2 106957 1 58640
2 106958 1 58640
2 106959 1 58640
2 106960 1 58640
2 106961 1 58640
2 106962 1 58640
2 106963 1 58640
2 106964 1 58640
2 106965 1 58640
2 106966 1 58640
2 106967 1 58640
2 106968 1 58675
2 106969 1 58675
2 106970 1 58693
2 106971 1 58693
2 106972 1 58693
2 106973 1 58693
2 106974 1 58693
2 106975 1 58693
2 106976 1 58693
2 106977 1 58693
2 106978 1 58693
2 106979 1 58693
2 106980 1 58693
2 106981 1 58693
2 106982 1 58694
2 106983 1 58694
2 106984 1 58711
2 106985 1 58711
2 106986 1 58711
2 106987 1 58733
2 106988 1 58733
2 106989 1 58741
2 106990 1 58741
2 106991 1 58748
2 106992 1 58748
2 106993 1 58748
2 106994 1 58748
2 106995 1 58750
2 106996 1 58750
2 106997 1 58758
2 106998 1 58758
2 106999 1 58758
2 107000 1 58758
2 107001 1 58758
2 107002 1 58758
2 107003 1 58758
2 107004 1 58758
2 107005 1 58759
2 107006 1 58759
2 107007 1 58767
2 107008 1 58767
2 107009 1 58781
2 107010 1 58781
2 107011 1 58824
2 107012 1 58824
2 107013 1 58835
2 107014 1 58835
2 107015 1 58850
2 107016 1 58850
2 107017 1 58850
2 107018 1 58862
2 107019 1 58862
2 107020 1 58862
2 107021 1 58863
2 107022 1 58863
2 107023 1 58908
2 107024 1 58908
2 107025 1 58926
2 107026 1 58926
2 107027 1 58927
2 107028 1 58927
2 107029 1 58934
2 107030 1 58934
2 107031 1 58958
2 107032 1 58958
2 107033 1 58958
2 107034 1 58973
2 107035 1 58973
2 107036 1 58973
2 107037 1 58973
2 107038 1 58973
2 107039 1 59041
2 107040 1 59041
2 107041 1 59042
2 107042 1 59042
2 107043 1 59042
2 107044 1 59108
2 107045 1 59108
2 107046 1 59156
2 107047 1 59156
2 107048 1 59156
2 107049 1 59156
2 107050 1 59167
2 107051 1 59167
2 107052 1 59167
2 107053 1 59191
2 107054 1 59191
2 107055 1 59191
2 107056 1 59191
2 107057 1 59191
2 107058 1 59192
2 107059 1 59192
2 107060 1 59193
2 107061 1 59193
2 107062 1 59193
2 107063 1 59195
2 107064 1 59195
2 107065 1 59196
2 107066 1 59196
2 107067 1 59196
2 107068 1 59196
2 107069 1 59198
2 107070 1 59198
2 107071 1 59199
2 107072 1 59199
2 107073 1 59203
2 107074 1 59203
2 107075 1 59205
2 107076 1 59205
2 107077 1 59216
2 107078 1 59216
2 107079 1 59221
2 107080 1 59221
2 107081 1 59221
2 107082 1 59221
2 107083 1 59221
2 107084 1 59223
2 107085 1 59223
2 107086 1 59230
2 107087 1 59230
2 107088 1 59233
2 107089 1 59233
2 107090 1 59233
2 107091 1 59245
2 107092 1 59245
2 107093 1 59246
2 107094 1 59246
2 107095 1 59250
2 107096 1 59250
2 107097 1 59274
2 107098 1 59274
2 107099 1 59274
2 107100 1 59281
2 107101 1 59281
2 107102 1 59300
2 107103 1 59300
2 107104 1 59300
2 107105 1 59300
2 107106 1 59300
2 107107 1 59300
2 107108 1 59300
2 107109 1 59300
2 107110 1 59301
2 107111 1 59301
2 107112 1 59308
2 107113 1 59308
2 107114 1 59311
2 107115 1 59311
2 107116 1 59312
2 107117 1 59312
2 107118 1 59321
2 107119 1 59321
2 107120 1 59321
2 107121 1 59323
2 107122 1 59323
2 107123 1 59328
2 107124 1 59328
2 107125 1 59328
2 107126 1 59328
2 107127 1 59328
2 107128 1 59328
2 107129 1 59328
2 107130 1 59328
2 107131 1 59339
2 107132 1 59339
2 107133 1 59339
2 107134 1 59346
2 107135 1 59346
2 107136 1 59354
2 107137 1 59354
2 107138 1 59354
2 107139 1 59354
2 107140 1 59354
2 107141 1 59357
2 107142 1 59357
2 107143 1 59382
2 107144 1 59382
2 107145 1 59393
2 107146 1 59393
2 107147 1 59426
2 107148 1 59426
2 107149 1 59462
2 107150 1 59462
2 107151 1 59479
2 107152 1 59479
2 107153 1 59481
2 107154 1 59481
2 107155 1 59481
2 107156 1 59493
2 107157 1 59493
2 107158 1 59510
2 107159 1 59510
2 107160 1 59540
2 107161 1 59540
2 107162 1 59540
2 107163 1 59540
2 107164 1 59548
2 107165 1 59548
2 107166 1 59572
2 107167 1 59572
2 107168 1 59587
2 107169 1 59587
2 107170 1 59596
2 107171 1 59596
2 107172 1 59623
2 107173 1 59623
2 107174 1 59634
2 107175 1 59634
2 107176 1 59666
2 107177 1 59666
2 107178 1 59679
2 107179 1 59679
2 107180 1 59743
2 107181 1 59743
2 107182 1 59757
2 107183 1 59757
2 107184 1 59758
2 107185 1 59758
2 107186 1 59777
2 107187 1 59777
2 107188 1 59806
2 107189 1 59806
2 107190 1 59818
2 107191 1 59818
2 107192 1 59820
2 107193 1 59820
2 107194 1 59820
2 107195 1 59829
2 107196 1 59829
2 107197 1 59885
2 107198 1 59885
2 107199 1 59902
2 107200 1 59902
2 107201 1 59912
2 107202 1 59912
2 107203 1 59921
2 107204 1 59921
2 107205 1 59940
2 107206 1 59940
2 107207 1 59951
2 107208 1 59951
2 107209 1 59951
2 107210 1 59951
2 107211 1 59961
2 107212 1 59961
2 107213 1 60072
2 107214 1 60072
2 107215 1 60117
2 107216 1 60117
2 107217 1 60136
2 107218 1 60136
2 107219 1 60151
2 107220 1 60151
2 107221 1 60178
2 107222 1 60178
2 107223 1 60191
2 107224 1 60191
2 107225 1 60191
2 107226 1 60201
2 107227 1 60201
2 107228 1 60209
2 107229 1 60209
2 107230 1 60259
2 107231 1 60259
2 107232 1 60259
2 107233 1 60337
2 107234 1 60337
2 107235 1 60362
2 107236 1 60362
2 107237 1 60389
2 107238 1 60389
2 107239 1 60389
2 107240 1 60447
2 107241 1 60447
2 107242 1 60452
2 107243 1 60452
2 107244 1 60462
2 107245 1 60462
2 107246 1 60462
2 107247 1 60462
2 107248 1 60462
2 107249 1 60487
2 107250 1 60487
2 107251 1 60500
2 107252 1 60500
2 107253 1 60503
2 107254 1 60503
2 107255 1 60506
2 107256 1 60506
2 107257 1 60510
2 107258 1 60510
2 107259 1 60511
2 107260 1 60511
2 107261 1 60525
2 107262 1 60525
2 107263 1 60525
2 107264 1 60526
2 107265 1 60526
2 107266 1 60529
2 107267 1 60529
2 107268 1 60544
2 107269 1 60544
2 107270 1 60546
2 107271 1 60546
2 107272 1 60555
2 107273 1 60555
2 107274 1 60555
2 107275 1 60555
2 107276 1 60571
2 107277 1 60571
2 107278 1 60571
2 107279 1 60571
2 107280 1 60581
2 107281 1 60581
2 107282 1 60581
2 107283 1 60581
2 107284 1 60581
2 107285 1 60582
2 107286 1 60582
2 107287 1 60587
2 107288 1 60587
2 107289 1 60607
2 107290 1 60607
2 107291 1 60617
2 107292 1 60617
2 107293 1 60665
2 107294 1 60665
2 107295 1 60665
2 107296 1 60665
2 107297 1 60665
2 107298 1 60665
2 107299 1 60675
2 107300 1 60675
2 107301 1 60693
2 107302 1 60693
2 107303 1 60694
2 107304 1 60694
2 107305 1 60695
2 107306 1 60695
2 107307 1 60711
2 107308 1 60711
2 107309 1 60745
2 107310 1 60745
2 107311 1 60745
2 107312 1 60746
2 107313 1 60746
2 107314 1 60751
2 107315 1 60751
2 107316 1 60786
2 107317 1 60786
2 107318 1 60795
2 107319 1 60795
2 107320 1 60804
2 107321 1 60804
2 107322 1 60814
2 107323 1 60814
2 107324 1 60815
2 107325 1 60815
2 107326 1 60869
2 107327 1 60869
2 107328 1 60907
2 107329 1 60907
2 107330 1 60921
2 107331 1 60921
2 107332 1 60939
2 107333 1 60939
2 107334 1 60968
2 107335 1 60968
2 107336 1 60968
2 107337 1 60990
2 107338 1 60990
2 107339 1 61025
2 107340 1 61025
2 107341 1 61025
2 107342 1 61025
2 107343 1 61025
2 107344 1 61025
2 107345 1 61025
2 107346 1 61025
2 107347 1 61032
2 107348 1 61032
2 107349 1 61032
2 107350 1 61049
2 107351 1 61049
2 107352 1 61066
2 107353 1 61066
2 107354 1 61095
2 107355 1 61095
2 107356 1 61095
2 107357 1 61112
2 107358 1 61112
2 107359 1 61161
2 107360 1 61161
2 107361 1 61161
2 107362 1 61161
2 107363 1 61172
2 107364 1 61172
2 107365 1 61176
2 107366 1 61176
2 107367 1 61197
2 107368 1 61197
2 107369 1 61206
2 107370 1 61206
2 107371 1 61207
2 107372 1 61207
2 107373 1 61207
2 107374 1 61213
2 107375 1 61213
2 107376 1 61219
2 107377 1 61219
2 107378 1 61219
2 107379 1 61219
2 107380 1 61315
2 107381 1 61315
2 107382 1 61325
2 107383 1 61325
2 107384 1 61325
2 107385 1 61331
2 107386 1 61331
2 107387 1 61343
2 107388 1 61343
2 107389 1 61343
2 107390 1 61343
2 107391 1 61343
2 107392 1 61343
2 107393 1 61343
2 107394 1 61402
2 107395 1 61402
2 107396 1 61410
2 107397 1 61410
2 107398 1 61419
2 107399 1 61419
2 107400 1 61428
2 107401 1 61428
2 107402 1 61439
2 107403 1 61439
2 107404 1 61451
2 107405 1 61451
2 107406 1 61451
2 107407 1 61451
2 107408 1 61462
2 107409 1 61462
2 107410 1 61466
2 107411 1 61466
2 107412 1 61466
2 107413 1 61466
2 107414 1 61481
2 107415 1 61481
2 107416 1 61481
2 107417 1 61481
2 107418 1 61482
2 107419 1 61482
2 107420 1 61549
2 107421 1 61549
2 107422 1 61553
2 107423 1 61553
2 107424 1 61572
2 107425 1 61572
2 107426 1 61604
2 107427 1 61604
2 107428 1 61605
2 107429 1 61605
2 107430 1 61605
2 107431 1 61605
2 107432 1 61605
2 107433 1 61640
2 107434 1 61640
2 107435 1 61640
2 107436 1 61707
2 107437 1 61707
2 107438 1 61725
2 107439 1 61725
2 107440 1 61726
2 107441 1 61726
2 107442 1 61735
2 107443 1 61735
2 107444 1 61742
2 107445 1 61742
2 107446 1 61778
2 107447 1 61778
2 107448 1 61780
2 107449 1 61780
2 107450 1 61782
2 107451 1 61782
2 107452 1 61782
2 107453 1 61783
2 107454 1 61783
2 107455 1 61783
2 107456 1 61785
2 107457 1 61785
2 107458 1 61785
2 107459 1 61798
2 107460 1 61798
2 107461 1 61839
2 107462 1 61839
2 107463 1 61860
2 107464 1 61860
2 107465 1 61891
2 107466 1 61891
2 107467 1 61891
2 107468 1 61891
2 107469 1 61968
2 107470 1 61968
2 107471 1 62000
2 107472 1 62000
2 107473 1 62014
2 107474 1 62014
2 107475 1 62018
2 107476 1 62018
2 107477 1 62061
2 107478 1 62061
2 107479 1 62069
2 107480 1 62069
2 107481 1 62069
2 107482 1 62077
2 107483 1 62077
2 107484 1 62097
2 107485 1 62097
2 107486 1 62131
2 107487 1 62131
2 107488 1 62131
2 107489 1 62164
2 107490 1 62164
2 107491 1 62164
2 107492 1 62164
2 107493 1 62164
2 107494 1 62164
2 107495 1 62164
2 107496 1 62164
2 107497 1 62164
2 107498 1 62167
2 107499 1 62167
2 107500 1 62183
2 107501 1 62183
2 107502 1 62192
2 107503 1 62192
2 107504 1 62201
2 107505 1 62201
2 107506 1 62201
2 107507 1 62204
2 107508 1 62204
2 107509 1 62219
2 107510 1 62219
2 107511 1 62227
2 107512 1 62227
2 107513 1 62236
2 107514 1 62236
2 107515 1 62245
2 107516 1 62245
2 107517 1 62247
2 107518 1 62247
2 107519 1 62249
2 107520 1 62249
2 107521 1 62250
2 107522 1 62250
2 107523 1 62250
2 107524 1 62275
2 107525 1 62275
2 107526 1 62276
2 107527 1 62276
2 107528 1 62316
2 107529 1 62316
2 107530 1 62319
2 107531 1 62319
2 107532 1 62324
2 107533 1 62324
2 107534 1 62356
2 107535 1 62356
2 107536 1 62358
2 107537 1 62358
2 107538 1 62360
2 107539 1 62360
2 107540 1 62388
2 107541 1 62388
2 107542 1 62397
2 107543 1 62397
2 107544 1 62406
2 107545 1 62406
2 107546 1 62446
2 107547 1 62446
2 107548 1 62508
2 107549 1 62508
2 107550 1 62512
2 107551 1 62512
2 107552 1 62527
2 107553 1 62527
2 107554 1 62552
2 107555 1 62552
2 107556 1 62597
2 107557 1 62597
2 107558 1 62605
2 107559 1 62605
2 107560 1 62658
2 107561 1 62658
2 107562 1 62670
2 107563 1 62670
2 107564 1 62674
2 107565 1 62674
2 107566 1 62678
2 107567 1 62678
2 107568 1 62761
2 107569 1 62761
2 107570 1 62761
2 107571 1 62801
2 107572 1 62801
2 107573 1 62876
2 107574 1 62876
2 107575 1 62876
2 107576 1 62876
2 107577 1 62898
2 107578 1 62898
2 107579 1 62916
2 107580 1 62916
2 107581 1 62917
2 107582 1 62917
2 107583 1 62944
2 107584 1 62944
2 107585 1 62953
2 107586 1 62953
2 107587 1 63006
2 107588 1 63006
2 107589 1 63014
2 107590 1 63014
2 107591 1 63017
2 107592 1 63017
2 107593 1 63026
2 107594 1 63026
2 107595 1 63084
2 107596 1 63084
2 107597 1 63084
2 107598 1 63144
2 107599 1 63144
2 107600 1 63168
2 107601 1 63168
2 107602 1 63169
2 107603 1 63169
2 107604 1 63205
2 107605 1 63205
2 107606 1 63310
2 107607 1 63310
2 107608 1 63387
2 107609 1 63387
2 107610 1 63498
2 107611 1 63498
2 107612 1 63605
2 107613 1 63605
0 27 5 165 1 25
0 28 5 132 1 63836
0 29 5 51 1 63950
0 30 5 242 1 64010
0 31 5 344 1 64229
0 32 5 361 1 64536
0 33 5 271 1 64920
0 34 5 278 1 65242
0 35 5 63 1 65548
0 36 5 51 1 65617
0 37 5 55 1 65669
0 38 5 180 1 65708
0 39 5 284 1 65866
0 40 5 301 1 66096
0 41 5 192 1 66415
0 42 5 166 1 66621
0 43 5 98 1 66811
0 44 5 103 1 66909
0 45 5 130 1 67017
0 46 5 87 1 67152
0 47 5 208 1 67251
0 48 5 347 1 67495
0 49 5 455 1 67839
0 50 5 316 1 68231
0 51 5 184 1 68541
0 52 7 9 2 70650 65670
0 53 7 8 2 63951 73807
0 54 5 1 1 73816
0 55 7 5 2 65618 70701
0 56 7 6 2 69040 73824
0 57 5 1 1 73829
0 58 7 1 2 54 57
0 59 5 50 1 58
0 60 7 46 2 71521 68232
0 61 5 66 1 73885
0 62 7 5 2 68743 65549
0 63 5 1 1 73997
0 64 7 8 2 26 70587
0 65 5 1 1 74002
0 66 7 5 2 63 65
0 67 5 34 1 74010
0 68 7 32 2 65709 70936
0 69 5 1 1 74049
0 70 7 2 2 70309 74050
0 71 7 8 2 68908 71879
0 72 7 17 2 66910 67018
0 73 7 17 2 74083 74091
0 74 7 6 2 69333 67840
0 75 5 2 1 74125
0 76 7 5 2 64011 71220
0 77 7 1 2 74126 74133
0 78 7 1 2 74108 77
0 79 7 1 2 74081 78
0 80 5 1 1 79
0 81 7 18 2 65867 66097
0 82 5 2 1 74138
0 83 7 4 2 66812 74139
0 84 7 16 2 64921 70756
0 85 5 1 1 74162
0 86 7 1 2 64537 74163
0 87 7 2 2 74158 86
0 88 7 22 2 69091 64230
0 89 7 2 2 63837 74180
0 90 7 7 2 71977 72852
0 91 7 17 2 72080 73623
0 92 5 1 1 74211
0 93 7 1 2 74204 74212
0 94 7 1 2 74202 93
0 95 7 1 2 74178 94
0 96 5 1 1 95
0 97 7 1 2 80 96
0 98 5 1 1 97
0 99 7 1 2 74015 98
0 100 5 1 1 99
0 101 7 30 2 66911 72081
0 102 7 12 2 63838 74228
0 103 5 7 1 74258
0 104 7 14 2 67019 73624
0 105 7 10 2 68909 71978
0 106 7 2 2 74277 74291
0 107 5 1 1 74301
0 108 7 1 2 74270 107
0 109 5 3 1 108
0 110 7 2 2 72853 74303
0 111 7 14 2 65868 66813
0 112 7 3 2 65243 74308
0 113 7 1 2 65550 74322
0 114 7 14 2 64538 70757
0 115 5 1 1 74325
0 116 7 9 2 66098 74326
0 117 5 1 1 74339
0 118 7 13 2 63719 69092
0 119 7 2 2 64231 74348
0 120 7 1 2 74340 74361
0 121 7 1 2 113 120
0 122 7 1 2 74306 121
0 123 5 1 1 122
0 124 7 1 2 100 123
0 125 5 1 1 124
0 126 7 1 2 73931 125
0 127 5 1 1 126
0 128 7 53 2 64012 65710
0 129 5 30 1 74363
0 130 7 11 2 68910 67020
0 131 7 27 2 70588 71979
0 132 7 8 2 71522 72854
0 133 7 3 2 70038 74484
0 134 5 4 1 74492
0 135 7 82 2 70039 71523
0 136 5 135 1 74499
0 137 7 33 2 67841 73307
0 138 5 7 1 74716
0 139 7 3 2 74581 74717
0 140 5 3 1 74756
0 141 7 2 2 74495 74759
0 142 5 1 1 74762
0 143 7 1 2 73625 142
0 144 5 1 1 143
0 145 7 41 2 72855 68233
0 146 5 5 1 74764
0 147 7 5 2 70040 74765
0 148 5 3 1 74810
0 149 7 7 2 73626 74582
0 150 5 3 1 74818
0 151 7 1 2 67842 74819
0 152 5 1 1 151
0 153 7 1 2 74815 152
0 154 5 1 1 153
0 155 7 1 2 65244 154
0 156 5 1 1 155
0 157 7 1 2 144 156
0 158 5 1 1 157
0 159 7 1 2 71221 158
0 160 5 1 1 159
0 161 7 37 2 68234 68542
0 162 5 19 1 74828
0 163 7 3 2 71524 74829
0 164 5 5 1 74884
0 165 7 22 2 70041 65245
0 166 5 1 1 74892
0 167 7 2 2 72856 74893
0 168 7 1 2 74885 74914
0 169 5 1 1 168
0 170 7 1 2 160 169
0 171 5 1 1 170
0 172 7 1 2 74457 171
0 173 5 1 1 172
0 174 7 7 2 65246 66912
0 175 7 5 2 65551 73627
0 176 7 2 2 74916 74923
0 177 7 56 2 71222 67843
0 178 5 40 1 74930
0 179 7 9 2 70042 73886
0 180 5 19 1 75026
0 181 7 1 2 74986 75035
0 182 5 1 1 181
0 183 7 1 2 74928 182
0 184 5 1 1 183
0 185 7 1 2 173 184
0 186 5 1 1 185
0 187 7 1 2 74446 186
0 188 5 1 1 187
0 189 7 10 2 66099 68235
0 190 5 6 1 75054
0 191 7 18 2 71223 73308
0 192 5 5 1 75070
0 193 7 18 2 65247 73628
0 194 5 25 1 75093
0 195 7 2 2 74500 75111
0 196 5 4 1 75136
0 197 7 1 2 75071 75138
0 198 5 1 1 197
0 199 7 1 2 75064 198
0 200 5 1 1 199
0 201 7 7 2 66913 67844
0 202 7 22 2 63839 70589
0 203 7 18 2 72082 75149
0 204 7 1 2 75142 75171
0 205 7 1 2 200 204
0 206 5 1 1 205
0 207 7 1 2 188 206
0 208 5 1 1 207
0 209 7 1 2 69677 208
0 210 5 1 1 209
0 211 7 11 2 63840 66914
0 212 7 39 2 72083 75189
0 213 5 2 1 75200
0 214 7 62 2 64922 66416
0 215 5 166 1 75241
0 216 7 8 2 68543 75303
0 217 5 2 1 75469
0 218 7 4 2 74583 75477
0 219 5 1 1 75479
0 220 7 7 2 70310 75304
0 221 5 2 1 75483
0 222 7 3 2 75480 75490
0 223 7 1 2 75201 75492
0 224 5 1 1 223
0 225 7 19 2 64923 65248
0 226 5 3 1 75495
0 227 7 4 2 68911 75496
0 228 7 7 2 66417 71980
0 229 7 10 2 67021 68544
0 230 7 1 2 75521 75528
0 231 7 1 2 75517 230
0 232 5 1 1 231
0 233 7 1 2 224 232
0 234 5 1 1 233
0 235 7 47 2 67845 68236
0 236 5 4 1 75538
0 237 7 6 2 70590 71224
0 238 7 1 2 75539 75589
0 239 7 1 2 234 238
0 240 5 1 1 239
0 241 7 1 2 210 240
0 242 5 1 1 241
0 243 7 1 2 71880 242
0 244 5 1 1 243
0 245 7 18 2 64539 72857
0 246 5 19 1 75595
0 247 7 4 2 71525 73629
0 248 5 2 1 75632
0 249 7 2 2 70043 75633
0 250 7 1 2 75613 75638
0 251 5 1 1 250
0 252 7 11 2 65249 67846
0 253 5 4 1 75640
0 254 7 2 2 64540 74865
0 255 5 2 1 75655
0 256 7 1 2 66100 75656
0 257 5 1 1 256
0 258 7 1 2 75641 257
0 259 5 1 1 258
0 260 7 1 2 251 259
0 261 5 1 1 260
0 262 7 13 2 63841 66814
0 263 7 4 2 65552 72084
0 264 7 8 2 75659 75672
0 265 7 2 2 71981 75676
0 266 7 1 2 261 75684
0 267 5 1 1 266
0 268 7 1 2 244 267
0 269 5 1 1 268
0 270 7 1 2 69334 269
0 271 5 1 1 270
0 272 7 11 2 71225 68237
0 273 5 3 1 75686
0 274 7 2 2 64924 75687
0 275 5 2 1 75700
0 276 7 8 2 68912 70311
0 277 7 53 2 71881 66915
0 278 7 11 2 67022 75712
0 279 7 1 2 75704 75765
0 280 7 1 2 75701 279
0 281 5 1 1 280
0 282 7 12 2 71226 73630
0 283 5 4 1 75776
0 284 7 2 2 65250 74830
0 285 5 1 1 75792
0 286 7 1 2 75788 285
0 287 5 2 1 286
0 288 7 15 2 63842 70044
0 289 7 17 2 71982 72085
0 290 7 13 2 66815 75811
0 291 7 1 2 75796 75828
0 292 7 1 2 75794 291
0 293 5 1 1 292
0 294 7 1 2 281 293
0 295 5 1 1 294
0 296 7 13 2 71526 67847
0 297 5 3 1 75841
0 298 7 5 2 69678 65553
0 299 7 1 2 75842 75857
0 300 7 1 2 295 299
0 301 5 1 1 300
0 302 7 1 2 271 301
0 303 5 1 1 302
0 304 7 1 2 70937 303
0 305 5 1 1 304
0 306 7 4 2 70591 72858
0 307 7 19 2 63843 72086
0 308 5 1 1 75866
0 309 7 3 2 70312 74831
0 310 5 4 1 75885
0 311 7 1 2 66101 75888
0 312 5 1 1 311
0 313 7 2 2 75867 312
0 314 7 1 2 75862 75892
0 315 5 1 1 314
0 316 7 52 2 66102 72859
0 317 5 47 1 75894
0 318 7 2 2 73631 75946
0 319 5 1 1 75993
0 320 7 12 2 68913 65251
0 321 5 1 1 75995
0 322 7 6 2 65554 67023
0 323 7 3 2 75996 76007
0 324 7 1 2 75994 76013
0 325 5 1 1 324
0 326 7 1 2 315 325
0 327 5 1 1 326
0 328 7 1 2 69679 327
0 329 5 1 1 328
0 330 7 19 2 66103 67848
0 331 5 6 1 76016
0 332 7 14 2 71227 72860
0 333 5 4 1 76041
0 334 7 3 2 76035 76055
0 335 5 52 1 76059
0 336 7 6 2 68238 76062
0 337 7 4 2 70313 72087
0 338 7 3 2 75150 76120
0 339 7 1 2 68545 76124
0 340 7 1 2 76114 339
0 341 5 1 1 340
0 342 7 10 2 65252 65555
0 343 7 2 2 68914 76127
0 344 7 29 2 67849 73632
0 345 5 1 1 76139
0 346 7 4 2 71228 67024
0 347 7 1 2 76140 76168
0 348 7 1 2 76137 347
0 349 5 1 1 348
0 350 7 1 2 341 349
0 351 7 1 2 329 350
0 352 5 1 1 351
0 353 7 1 2 75713 352
0 354 5 1 1 353
0 355 7 84 2 64541 66104
0 356 5 91 1 76172
0 357 7 2 2 73633 76256
0 358 5 1 1 76347
0 359 7 1 2 75651 358
0 360 5 1 1 359
0 361 7 10 2 71983 68239
0 362 7 1 2 76349 75677
0 363 7 1 2 360 362
0 364 5 1 1 363
0 365 7 1 2 354 364
0 366 5 1 1 365
0 367 7 1 2 70938 366
0 368 5 1 1 367
0 369 7 41 2 66816 71984
0 370 7 2 2 75540 76359
0 371 7 24 2 65253 71229
0 372 5 1 1 76402
0 373 7 1 2 76403 75858
0 374 7 1 2 75868 373
0 375 7 1 2 76400 374
0 376 5 1 1 375
0 377 7 1 2 368 376
0 378 5 1 1 377
0 379 7 1 2 69335 378
0 380 5 1 1 379
0 381 7 5 2 67850 76360
0 382 7 95 2 69680 71230
0 383 5 91 1 76431
0 384 7 8 2 70939 68240
0 385 5 2 1 76617
0 386 7 3 2 76432 76618
0 387 7 1 2 76128 75869
0 388 7 1 2 76627 387
0 389 7 1 2 76426 388
0 390 5 1 1 389
0 391 7 1 2 380 390
0 392 5 1 1 391
0 393 7 1 2 75305 392
0 394 5 1 1 393
0 395 7 4 2 64542 74584
0 396 5 34 1 76630
0 397 7 27 2 68241 73634
0 398 5 3 1 76668
0 399 7 18 2 65254 70940
0 400 7 2 2 76698 74109
0 401 7 1 2 76669 76716
0 402 5 1 1 401
0 403 7 21 2 75660 75812
0 404 5 5 1 76718
0 405 7 4 2 70941 73635
0 406 5 1 1 76744
0 407 7 8 2 68546 75541
0 408 7 1 2 65255 76748
0 409 5 1 1 408
0 410 7 1 2 406 409
0 411 5 1 1 410
0 412 7 1 2 76719 411
0 413 5 1 1 412
0 414 7 1 2 402 413
0 415 5 1 1 414
0 416 7 1 2 65556 415
0 417 5 1 1 416
0 418 7 24 2 67025 74292
0 419 5 1 1 76756
0 420 7 12 2 72861 74832
0 421 5 1 1 76780
0 422 7 25 2 70592 71882
0 423 7 1 2 76792 76699
0 424 7 1 2 76781 423
0 425 7 1 2 76757 424
0 426 5 1 1 425
0 427 7 1 2 417 426
0 428 5 1 1 427
0 429 7 1 2 71231 428
0 430 5 1 1 429
0 431 7 12 2 67851 74833
0 432 5 1 1 76817
0 433 7 1 2 68915 76818
0 434 7 33 2 71985 67026
0 435 7 4 2 71883 76829
0 436 7 11 2 70942 66105
0 437 7 17 2 65256 70593
0 438 7 2 2 76866 76877
0 439 7 1 2 76862 76894
0 440 7 1 2 433 439
0 441 5 1 1 440
0 442 7 1 2 430 441
0 443 5 1 1 442
0 444 7 1 2 69336 443
0 445 5 1 1 444
0 446 7 12 2 72088 76361
0 447 7 2 2 76896 76749
0 448 7 15 2 63844 65557
0 449 7 19 2 70943 71232
0 450 5 1 1 76925
0 451 7 2 2 65257 76926
0 452 7 1 2 76910 76944
0 453 7 1 2 76908 452
0 454 5 1 1 453
0 455 7 1 2 445 454
0 456 5 1 1 455
0 457 7 1 2 76634 456
0 458 5 1 1 457
0 459 7 23 2 69337 69681
0 460 5 2 1 76946
0 461 7 3 2 67852 76947
0 462 7 6 2 65558 71527
0 463 7 2 2 75797 76974
0 464 7 1 2 76897 76980
0 465 7 1 2 76971 464
0 466 7 1 2 75795 465
0 467 5 1 1 466
0 468 7 1 2 458 467
0 469 7 1 2 394 468
0 470 7 1 2 305 469
0 471 5 1 1 470
0 472 7 1 2 74364 471
0 473 5 1 1 472
0 474 7 25 2 72862 73636
0 475 5 3 1 76982
0 476 7 13 2 72089 73309
0 477 7 3 2 76983 77010
0 478 7 5 2 64543 71986
0 479 7 1 2 74181 77026
0 480 7 1 2 77023 479
0 481 7 6 2 66817 76911
0 482 7 17 2 66106 66418
0 483 5 3 1 77037
0 484 7 19 2 70758 65869
0 485 7 2 2 77038 77057
0 486 7 1 2 77031 77076
0 487 7 1 2 480 486
0 488 5 1 1 487
0 489 7 1 2 68744 488
0 490 7 1 2 473 489
0 491 5 1 1 490
0 492 7 14 2 71528 68547
0 493 5 15 1 77078
0 494 7 10 2 70045 77079
0 495 5 13 1 77107
0 496 7 2 2 76257 77108
0 497 5 2 1 77130
0 498 7 64 2 69338 70944
0 499 5 79 1 77134
0 500 7 1 2 76526 77198
0 501 7 1 2 77132 500
0 502 5 1 1 501
0 503 7 12 2 66419 73637
0 504 5 7 1 77277
0 505 7 5 2 64925 77278
0 506 5 13 1 77296
0 507 7 74 2 64232 65870
0 508 5 105 1 77314
0 509 7 1 2 77301 77388
0 510 7 2 2 502 509
0 511 7 10 2 63845 65258
0 512 7 2 2 75829 77495
0 513 7 1 2 77493 77505
0 514 5 1 1 513
0 515 7 4 2 68916 71529
0 516 7 2 2 75766 77507
0 517 5 1 1 77511
0 518 7 4 2 64926 76433
0 519 5 1 1 77513
0 520 7 14 2 70314 70945
0 521 5 1 1 77517
0 522 7 1 2 77514 77518
0 523 7 1 2 77512 522
0 524 5 1 1 523
0 525 7 1 2 514 524
0 526 5 1 1 525
0 527 7 1 2 75542 526
0 528 5 1 1 527
0 529 7 17 2 67853 76434
0 530 5 8 1 77531
0 531 7 6 2 66107 75596
0 532 5 11 1 77556
0 533 7 3 2 70946 77562
0 534 5 1 1 77573
0 535 7 3 2 77548 534
0 536 5 2 1 77576
0 537 7 1 2 71530 77579
0 538 5 1 1 537
0 539 7 3 2 70947 76258
0 540 5 7 1 77581
0 541 7 1 2 68242 77582
0 542 5 1 1 541
0 543 7 1 2 538 542
0 544 5 2 1 543
0 545 7 1 2 76720 77591
0 546 5 1 1 545
0 547 7 10 2 72863 73932
0 548 5 14 1 77593
0 549 7 1 2 76527 77594
0 550 5 2 1 549
0 551 7 2 2 76259 77617
0 552 5 2 1 77619
0 553 7 1 2 77620 76717
0 554 5 1 1 553
0 555 7 1 2 546 554
0 556 5 1 1 555
0 557 7 1 2 70046 556
0 558 5 1 1 557
0 559 7 3 2 66108 73933
0 560 5 7 1 77623
0 561 7 1 2 77626 76721
0 562 5 1 1 561
0 563 7 8 2 67027 74084
0 564 7 4 2 74917 77633
0 565 7 1 2 66109 75854
0 566 5 2 1 565
0 567 7 38 2 72864 73310
0 568 5 9 1 77647
0 569 7 9 2 66420 77648
0 570 5 4 1 77694
0 571 7 1 2 77645 77703
0 572 7 1 2 77641 571
0 573 5 1 1 572
0 574 7 1 2 562 573
0 575 5 1 1 574
0 576 7 1 2 69682 575
0 577 5 1 1 576
0 578 7 11 2 71233 71531
0 579 7 18 2 72090 68243
0 580 7 3 2 63846 76362
0 581 7 2 2 77718 77736
0 582 5 1 1 77739
0 583 7 18 2 67028 67854
0 584 7 3 2 74085 77741
0 585 7 1 2 74918 77759
0 586 5 1 1 585
0 587 7 1 2 582 586
0 588 5 1 1 587
0 589 7 1 2 77707 588
0 590 5 1 1 589
0 591 7 1 2 577 590
0 592 5 1 1 591
0 593 7 1 2 70948 592
0 594 5 1 1 593
0 595 7 1 2 558 594
0 596 5 1 1 595
0 597 7 1 2 69339 596
0 598 5 1 1 597
0 599 7 3 2 71532 71987
0 600 7 17 2 66818 72091
0 601 7 5 2 67855 77765
0 602 7 2 2 77762 77782
0 603 7 6 2 63847 70949
0 604 7 16 2 70047 71234
0 605 5 1 1 77795
0 606 7 5 2 69683 77796
0 607 7 1 2 77789 77811
0 608 7 1 2 77787 607
0 609 5 1 1 608
0 610 7 1 2 598 609
0 611 5 1 1 610
0 612 7 1 2 73638 611
0 613 5 1 1 612
0 614 7 1 2 528 613
0 615 5 1 1 614
0 616 7 1 2 74365 615
0 617 5 1 1 616
0 618 7 21 2 68917 64927
0 619 7 6 2 71884 74092
0 620 7 2 2 77816 77837
0 621 5 2 1 77843
0 622 7 1 2 76739 77845
0 623 5 1 1 622
0 624 7 6 2 74140 74327
0 625 5 3 1 77847
0 626 7 23 2 66421 72865
0 627 5 3 1 77856
0 628 7 6 2 73311 77857
0 629 5 1 1 77882
0 630 7 1 2 77883 74182
0 631 7 1 2 77848 630
0 632 7 2 2 623 631
0 633 5 1 1 77888
0 634 7 1 2 73639 77889
0 635 5 1 1 634
0 636 7 1 2 617 635
0 637 5 1 1 636
0 638 7 1 2 70594 637
0 639 5 1 1 638
0 640 7 25 2 65559 66819
0 641 7 8 2 71533 76260
0 642 5 3 1 77915
0 643 7 4 2 76528 77923
0 644 5 1 1 77926
0 645 7 4 2 68244 76261
0 646 5 7 1 77930
0 647 7 4 2 77927 77934
0 648 5 1 1 77941
0 649 7 1 2 77942 74307
0 650 5 1 1 649
0 651 7 9 2 64544 66422
0 652 5 2 1 77945
0 653 7 11 2 66110 73312
0 654 5 1 1 77956
0 655 7 3 2 77946 77957
0 656 5 1 1 77967
0 657 7 1 2 75239 419
0 658 5 1 1 657
0 659 7 1 2 77968 658
0 660 5 1 1 659
0 661 7 1 2 650 660
0 662 5 1 1 661
0 663 7 10 2 65259 65871
0 664 5 1 1 77970
0 665 7 2 2 64928 77971
0 666 7 17 2 64233 70759
0 667 7 5 2 69093 77982
0 668 7 1 2 77980 77999
0 669 7 1 2 662 668
0 670 5 1 1 669
0 671 7 4 2 76948 76927
0 672 5 1 1 78004
0 673 7 15 2 70315 68548
0 674 5 4 1 78008
0 675 7 7 2 69684 68245
0 676 5 3 1 78027
0 677 7 1 2 78009 78028
0 678 5 2 1 677
0 679 7 1 2 77199 78037
0 680 5 1 1 679
0 681 7 1 2 75947 680
0 682 5 1 1 681
0 683 7 1 2 64545 75889
0 684 5 3 1 683
0 685 7 3 2 66111 77200
0 686 5 1 1 78042
0 687 7 4 2 72866 77201
0 688 5 1 1 78045
0 689 7 2 2 686 688
0 690 7 1 2 78039 78049
0 691 5 1 1 690
0 692 7 1 2 682 691
0 693 5 1 1 692
0 694 7 5 2 70950 75306
0 695 5 2 1 78051
0 696 7 5 2 69340 75307
0 697 5 2 1 78058
0 698 7 2 2 78056 78063
0 699 5 1 1 78065
0 700 7 1 2 693 699
0 701 5 1 1 700
0 702 7 1 2 672 701
0 703 5 1 1 702
0 704 7 1 2 74366 76758
0 705 7 1 2 703 704
0 706 5 1 1 705
0 707 7 1 2 670 706
0 708 5 1 1 707
0 709 7 1 2 77890 708
0 710 5 1 1 709
0 711 7 1 2 63720 710
0 712 7 1 2 639 711
0 713 5 1 1 712
0 714 7 1 2 491 713
0 715 5 1 1 714
0 716 7 1 2 127 715
0 717 5 1 1 716
0 718 7 1 2 72505 717
0 719 5 1 1 718
0 720 7 19 2 68918 65560
0 721 7 16 2 67029 78067
0 722 5 5 1 78086
0 723 7 10 2 65260 72092
0 724 7 3 2 78107 75151
0 725 5 1 1 78117
0 726 7 1 2 78102 725
0 727 5 1 1 726
0 728 7 16 2 64013 69341
0 729 7 6 2 78120 74051
0 730 7 10 2 67496 76529
0 731 5 1 1 78142
0 732 7 37 2 63721 66820
0 733 7 91 2 71988 78152
0 734 5 2 1 78189
0 735 7 2 2 78143 78190
0 736 5 1 1 78282
0 737 7 1 2 78136 78283
0 738 5 1 1 737
0 739 7 8 2 69094 77315
0 740 5 1 1 78284
0 741 7 6 2 70760 73640
0 742 7 4 2 78285 78292
0 743 7 2 2 73313 78298
0 744 5 1 1 78302
0 745 7 23 2 64546 64929
0 746 5 5 1 78304
0 747 7 5 2 68745 78305
0 748 7 17 2 66423 71885
0 749 7 4 2 66112 78337
0 750 7 11 2 66916 72506
0 751 7 1 2 78354 78358
0 752 7 1 2 78332 751
0 753 7 1 2 78303 752
0 754 5 1 1 753
0 755 7 1 2 738 754
0 756 5 1 1 755
0 757 7 1 2 72867 756
0 758 5 1 1 757
0 759 7 19 2 64234 70951
0 760 5 3 1 78369
0 761 7 7 2 67497 76435
0 762 7 1 2 78370 78391
0 763 5 1 1 762
0 764 7 23 2 70952 72507
0 765 5 3 1 78398
0 766 7 18 2 65872 67498
0 767 5 9 1 78424
0 768 7 3 2 78421 78442
0 769 5 10 1 78451
0 770 7 2 2 69342 78454
0 771 5 2 1 78464
0 772 7 26 2 70953 67499
0 773 5 5 1 78468
0 774 7 3 2 64235 78469
0 775 5 2 1 78499
0 776 7 1 2 78466 78502
0 777 5 20 1 776
0 778 7 2 2 76262 78504
0 779 5 1 1 78524
0 780 7 1 2 67856 78525
0 781 5 1 1 780
0 782 7 1 2 763 781
0 783 5 1 1 782
0 784 7 4 2 74367 76363
0 785 7 1 2 63722 78526
0 786 7 1 2 783 785
0 787 5 1 1 786
0 788 7 1 2 758 787
0 789 5 2 1 788
0 790 7 1 2 727 78530
0 791 5 1 1 790
0 792 7 12 2 67500 74368
0 793 7 15 2 68919 76830
0 794 7 2 2 75242 78544
0 795 5 1 1 78559
0 796 7 25 2 73314 73641
0 797 5 14 1 78561
0 798 7 3 2 72093 78562
0 799 7 1 2 75190 78600
0 800 5 1 1 799
0 801 7 1 2 795 800
0 802 5 1 1 801
0 803 7 1 2 69685 802
0 804 5 1 1 803
0 805 7 2 2 75191 77719
0 806 5 1 1 78603
0 807 7 1 2 74820 78604
0 808 5 1 1 807
0 809 7 1 2 804 808
0 810 5 1 1 809
0 811 7 1 2 67857 810
0 812 5 1 1 811
0 813 7 1 2 69686 74834
0 814 5 1 1 813
0 815 7 66 2 66424 73315
0 816 5 43 1 78605
0 817 7 1 2 64547 74887
0 818 5 1 1 817
0 819 7 2 2 70048 818
0 820 7 1 2 78671 78714
0 821 5 1 1 820
0 822 7 1 2 814 821
0 823 5 1 1 822
0 824 7 16 2 67030 72868
0 825 7 1 2 78716 74293
0 826 7 1 2 823 825
0 827 5 1 1 826
0 828 7 1 2 812 827
0 829 5 1 1 828
0 830 7 1 2 71235 829
0 831 5 1 1 830
0 832 7 2 2 74835 78545
0 833 7 17 2 69687 72869
0 834 5 4 1 78734
0 835 7 3 2 76036 78751
0 836 5 7 1 78755
0 837 7 2 2 74501 78758
0 838 5 3 1 78765
0 839 7 1 2 78732 78766
0 840 5 1 1 839
0 841 7 1 2 831 840
0 842 5 1 1 841
0 843 7 1 2 64236 842
0 844 5 1 1 843
0 845 7 2 2 66425 74766
0 846 5 1 1 78770
0 847 7 1 2 66426 74718
0 848 5 5 1 847
0 849 7 1 2 74805 78772
0 850 5 2 1 849
0 851 7 1 2 64930 78777
0 852 5 2 1 851
0 853 7 1 2 846 78779
0 854 5 1 1 853
0 855 7 1 2 76530 854
0 856 5 1 1 855
0 857 7 1 2 66113 76631
0 858 5 6 1 857
0 859 7 4 2 68246 78781
0 860 5 1 1 78787
0 861 7 20 2 64931 71236
0 862 5 1 1 78791
0 863 7 2 2 77858 78792
0 864 5 2 1 78811
0 865 7 1 2 73316 78813
0 866 5 1 1 865
0 867 7 1 2 860 866
0 868 5 1 1 867
0 869 7 1 2 856 868
0 870 5 1 1 869
0 871 7 1 2 69343 73642
0 872 7 1 2 74259 871
0 873 7 1 2 870 872
0 874 5 1 1 873
0 875 7 1 2 844 874
0 876 5 1 1 875
0 877 7 1 2 76793 876
0 878 5 1 1 877
0 879 7 8 2 72870 76531
0 880 5 6 1 78815
0 881 7 9 2 64237 76263
0 882 5 2 1 78829
0 883 7 1 2 78823 78830
0 884 5 2 1 883
0 885 7 6 2 69344 76532
0 886 5 1 1 78842
0 887 7 1 2 72871 78843
0 888 5 1 1 887
0 889 7 1 2 78840 888
0 890 5 1 1 889
0 891 7 1 2 75685 890
0 892 5 1 1 891
0 893 7 1 2 878 892
0 894 5 1 1 893
0 895 7 1 2 68746 894
0 896 5 1 1 895
0 897 7 42 2 65561 78153
0 898 5 1 1 78848
0 899 7 10 2 68247 74585
0 900 5 1 1 78890
0 901 7 8 2 67858 76533
0 902 5 2 1 78900
0 903 7 1 2 76056 78908
0 904 5 6 1 903
0 905 7 2 2 78891 78910
0 906 5 1 1 78916
0 907 7 8 2 66427 67859
0 908 5 1 1 78918
0 909 7 5 2 64932 78919
0 910 5 9 1 78926
0 911 7 1 2 78752 78931
0 912 5 2 1 911
0 913 7 2 2 71237 78940
0 914 5 1 1 78942
0 915 7 2 2 73317 78943
0 916 5 1 1 78944
0 917 7 1 2 906 916
0 918 5 1 1 917
0 919 7 1 2 74302 918
0 920 5 1 1 919
0 921 7 11 2 64933 66114
0 922 5 4 1 78946
0 923 7 2 2 76635 78957
0 924 5 2 1 78961
0 925 7 1 2 67860 78963
0 926 5 1 1 925
0 927 7 1 2 64934 76042
0 928 5 2 1 927
0 929 7 1 2 68248 78965
0 930 7 1 2 926 929
0 931 5 1 1 930
0 932 7 2 2 70049 76063
0 933 5 1 1 78967
0 934 7 3 2 69345 74987
0 935 5 2 1 78969
0 936 7 1 2 73318 78972
0 937 7 1 2 933 936
0 938 7 1 2 914 937
0 939 5 1 1 938
0 940 7 1 2 75202 939
0 941 7 1 2 931 940
0 942 5 1 1 941
0 943 7 1 2 920 942
0 944 5 1 1 943
0 945 7 1 2 78849 944
0 946 5 1 1 945
0 947 7 1 2 896 946
0 948 5 1 1 947
0 949 7 1 2 65261 948
0 950 5 1 1 949
0 951 7 29 2 68747 70595
0 952 5 4 1 78974
0 953 7 5 2 64238 71886
0 954 7 4 2 78975 79007
0 955 7 2 2 66917 76264
0 956 7 1 2 79016 78040
0 957 7 1 2 75893 956
0 958 5 1 1 957
0 959 7 21 2 69688 65262
0 960 5 2 1 79018
0 961 7 5 2 68920 79019
0 962 7 12 2 71989 68549
0 963 7 1 2 79046 76169
0 964 7 1 2 79041 963
0 965 5 1 1 964
0 966 7 1 2 958 965
0 967 5 1 1 966
0 968 7 1 2 79012 967
0 969 5 1 1 968
0 970 7 16 2 70316 66115
0 971 5 2 1 79058
0 972 7 1 2 79059 78733
0 973 5 1 1 972
0 974 7 3 2 66918 77011
0 975 7 16 2 63848 69689
0 976 7 1 2 65263 79079
0 977 7 1 2 79076 976
0 978 5 1 1 977
0 979 7 1 2 973 978
0 980 5 1 1 979
0 981 7 1 2 78850 980
0 982 5 1 1 981
0 983 7 1 2 969 982
0 984 5 1 1 983
0 985 7 1 2 72872 984
0 986 5 1 1 985
0 987 7 2 2 79060 76819
0 988 5 1 1 79095
0 989 7 21 2 68748 64239
0 990 7 8 2 79097 75714
0 991 7 1 2 79118 75172
0 992 7 1 2 79096 991
0 993 5 1 1 992
0 994 7 1 2 986 993
0 995 5 1 1 994
0 996 7 1 2 75308 995
0 997 5 1 1 996
0 998 7 32 2 71887 78976
0 999 7 4 2 71990 74278
0 1000 7 1 2 75705 79158
0 1001 5 1 1 1000
0 1002 7 1 2 74271 1001
0 1003 5 1 1 1002
0 1004 7 10 2 69346 66428
0 1005 5 1 1 79162
0 1006 7 5 2 69690 75948
0 1007 5 5 1 79172
0 1008 7 6 2 68249 74988
0 1009 7 4 2 79177 79182
0 1010 7 1 2 79163 79188
0 1011 7 1 2 1003 1010
0 1012 5 1 1 1011
0 1013 7 11 2 65264 68250
0 1014 5 2 1 79192
0 1015 7 1 2 79193 74272
0 1016 5 1 1 1015
0 1017 7 9 2 69691 73319
0 1018 5 4 1 79205
0 1019 7 18 2 66429 68251
0 1020 5 3 1 79218
0 1021 7 1 2 79214 79236
0 1022 5 5 1 1021
0 1023 7 8 2 64240 71238
0 1024 5 3 1 79244
0 1025 7 9 2 67861 79245
0 1026 5 2 1 79255
0 1027 7 1 2 79239 79256
0 1028 7 1 2 74304 1027
0 1029 7 1 2 1016 1028
0 1030 5 1 1 1029
0 1031 7 1 2 1012 1030
0 1032 5 1 1 1031
0 1033 7 1 2 64935 1032
0 1034 5 1 1 1033
0 1035 7 27 2 64241 69692
0 1036 5 2 1 79266
0 1037 7 5 2 71239 78606
0 1038 5 3 1 79295
0 1039 7 3 2 75065 79300
0 1040 5 3 1 79303
0 1041 7 1 2 79306 75203
0 1042 5 1 1 1041
0 1043 7 7 2 68921 66430
0 1044 7 2 2 76831 79309
0 1045 5 1 1 79316
0 1046 7 2 2 73320 79317
0 1047 5 1 1 79318
0 1048 7 1 2 75777 79319
0 1049 5 1 1 1048
0 1050 7 1 2 1042 1049
0 1051 5 1 1 1050
0 1052 7 1 2 67862 1051
0 1053 5 1 1 1052
0 1054 7 11 2 67031 68252
0 1055 7 4 2 79320 74294
0 1056 5 1 1 79331
0 1057 7 6 2 70317 73643
0 1058 5 5 1 79335
0 1059 7 1 2 76043 79336
0 1060 7 1 2 79332 1059
0 1061 5 1 1 1060
0 1062 7 1 2 1053 1061
0 1063 5 1 1 1062
0 1064 7 1 2 79267 1063
0 1065 5 1 1 1064
0 1066 7 1 2 1034 1065
0 1067 5 1 1 1066
0 1068 7 1 2 79126 1067
0 1069 5 1 1 1068
0 1070 7 11 2 67032 76364
0 1071 7 29 2 63723 68922
0 1072 7 9 2 65562 79357
0 1073 7 8 2 79346 79386
0 1074 5 3 1 79395
0 1075 7 13 2 64548 67863
0 1076 5 8 1 79406
0 1077 7 2 2 76057 79419
0 1078 5 6 1 79427
0 1079 7 1 2 75243 79429
0 1080 5 2 1 1079
0 1081 7 1 2 66116 78941
0 1082 5 1 1 1081
0 1083 7 1 2 79435 1082
0 1084 5 1 1 1083
0 1085 7 1 2 68253 1084
0 1086 5 1 1 1085
0 1087 7 2 2 76436 74586
0 1088 7 1 2 77649 79437
0 1089 5 2 1 1088
0 1090 7 2 2 1086 79439
0 1091 5 1 1 79441
0 1092 7 1 2 79396 1091
0 1093 5 1 1 1092
0 1094 7 1 2 1069 1093
0 1095 7 1 2 997 1094
0 1096 7 1 2 950 1095
0 1097 5 1 1 1096
0 1098 7 1 2 70954 1097
0 1099 5 1 1 1098
0 1100 7 10 2 63724 64549
0 1101 7 5 2 77891 79443
0 1102 5 1 1 79453
0 1103 7 25 2 65873 71240
0 1104 5 2 1 79458
0 1105 7 4 2 73644 79127
0 1106 7 1 2 79459 79485
0 1107 5 1 1 1106
0 1108 7 1 2 1102 1107
0 1109 5 1 1 1108
0 1110 7 1 2 74587 1109
0 1111 5 1 1 1110
0 1112 7 1 2 78947 78851
0 1113 5 1 1 1112
0 1114 7 1 2 1111 1113
0 1115 5 1 1 1114
0 1116 7 1 2 65265 1115
0 1117 5 1 1 1116
0 1118 7 2 2 75309 78010
0 1119 5 2 1 79489
0 1120 7 1 2 76173 79491
0 1121 5 1 1 1120
0 1122 7 3 2 71241 75310
0 1123 5 17 1 79493
0 1124 7 10 2 65874 71888
0 1125 7 4 2 78977 79513
0 1126 7 1 2 79496 79523
0 1127 7 1 2 1121 1126
0 1128 5 1 1 1127
0 1129 7 1 2 67864 1128
0 1130 7 1 2 1117 1129
0 1131 5 1 1 1130
0 1132 7 1 2 76534 79492
0 1133 5 1 1 1132
0 1134 7 1 2 76265 79524
0 1135 7 1 2 1133 1134
0 1136 5 1 1 1135
0 1137 7 3 2 65563 71242
0 1138 7 3 2 78154 79527
0 1139 7 1 2 75497 79530
0 1140 5 1 1 1139
0 1141 7 1 2 72873 1140
0 1142 7 1 2 1136 1141
0 1143 5 1 1 1142
0 1144 7 1 2 68254 1143
0 1145 7 1 2 1131 1144
0 1146 5 1 1 1145
0 1147 7 1 2 64550 605
0 1148 5 3 1 1147
0 1149 7 4 2 66431 78948
0 1150 5 2 1 79536
0 1151 7 5 2 79533 79540
0 1152 7 2 2 72874 79542
0 1153 5 2 1 79547
0 1154 7 12 2 70050 66117
0 1155 5 2 1 79551
0 1156 7 19 2 71243 66432
0 1157 5 1 1 79565
0 1158 7 2 2 64936 79566
0 1159 5 3 1 79584
0 1160 7 1 2 79563 79586
0 1161 5 3 1 1160
0 1162 7 1 2 67865 79589
0 1163 5 1 1 1162
0 1164 7 1 2 79549 1163
0 1165 5 1 1 1164
0 1166 7 7 2 63725 65266
0 1167 7 5 2 66821 73321
0 1168 7 3 2 65564 79599
0 1169 7 1 2 79592 79604
0 1170 7 1 2 1165 1169
0 1171 5 1 1 1170
0 1172 7 1 2 1146 1171
0 1173 5 1 1 1172
0 1174 7 1 2 66919 1173
0 1175 5 1 1 1174
0 1176 7 3 2 68749 65875
0 1177 7 2 2 76129 79607
0 1178 7 6 2 67866 76266
0 1179 5 4 1 79612
0 1180 7 1 2 79613 76365
0 1181 7 1 2 79610 1180
0 1182 5 1 1 1181
0 1183 7 1 2 1175 1182
0 1184 5 1 1 1183
0 1185 7 1 2 75870 1184
0 1186 5 1 1 1185
0 1187 7 29 2 63726 65565
0 1188 7 17 2 66822 79622
0 1189 7 2 2 75311 79651
0 1190 7 2 2 70318 74767
0 1191 5 3 1 79670
0 1192 7 1 2 68550 79671
0 1193 5 1 1 1192
0 1194 7 1 2 79420 1193
0 1195 5 1 1 1194
0 1196 7 1 2 79668 1195
0 1197 5 1 1 1196
0 1198 7 4 2 70596 65876
0 1199 7 6 2 68750 70051
0 1200 7 3 2 79675 79679
0 1201 7 7 2 71889 68255
0 1202 7 3 2 75843 79688
0 1203 7 9 2 65267 68551
0 1204 5 3 1 79698
0 1205 7 1 2 79695 79699
0 1206 7 1 2 79685 1205
0 1207 5 1 1 1206
0 1208 7 1 2 1197 1207
0 1209 5 1 1 1208
0 1210 7 1 2 66118 1209
0 1211 5 1 1 1210
0 1212 7 34 2 72875 68552
0 1213 5 2 1 79710
0 1214 7 2 2 71534 79711
0 1215 7 3 2 74894 79746
0 1216 5 1 1 79748
0 1217 7 1 2 69693 79749
0 1218 5 1 1 1217
0 1219 7 1 2 66119 1218
0 1220 5 1 1 1219
0 1221 7 5 2 66433 76141
0 1222 7 21 2 64937 70319
0 1223 5 1 1 79756
0 1224 7 1 2 79751 79757
0 1225 5 1 1 1224
0 1226 7 1 2 1216 1225
0 1227 5 2 1 1226
0 1228 7 9 2 65877 68256
0 1229 5 1 1 79779
0 1230 7 9 2 68751 76794
0 1231 7 1 2 79780 79788
0 1232 7 1 2 79777 1231
0 1233 7 1 2 1220 1232
0 1234 5 1 1 1233
0 1235 7 1 2 1211 1234
0 1236 5 1 1 1235
0 1237 7 1 2 76759 1236
0 1238 5 1 1 1237
0 1239 7 1 2 1186 1238
0 1240 5 1 1 1239
0 1241 7 1 2 69347 1240
0 1242 5 1 1 1241
0 1243 7 19 2 70320 68257
0 1244 5 7 1 79797
0 1245 7 8 2 69694 75312
0 1246 5 29 1 79823
0 1247 7 4 2 79831 79497
0 1248 5 2 1 79860
0 1249 7 1 2 78901 79861
0 1250 5 3 1 1249
0 1251 7 1 2 79866 78814
0 1252 5 1 1 1251
0 1253 7 1 2 79798 1252
0 1254 5 1 1 1253
0 1255 7 1 2 79440 1254
0 1256 5 1 1 1255
0 1257 7 1 2 76722 1256
0 1258 5 1 1 1257
0 1259 7 3 2 66120 78607
0 1260 5 3 1 79869
0 1261 7 2 2 69348 79872
0 1262 5 2 1 79875
0 1263 7 1 2 71244 78672
0 1264 5 4 1 1263
0 1265 7 1 2 79876 79879
0 1266 5 1 1 1265
0 1267 7 4 2 69695 78608
0 1268 5 4 1 79883
0 1269 7 1 2 71245 79887
0 1270 5 1 1 1269
0 1271 7 4 2 64242 66121
0 1272 5 2 1 79891
0 1273 7 1 2 70052 79895
0 1274 7 1 2 1270 1273
0 1275 5 1 1 1274
0 1276 7 1 2 1266 1275
0 1277 5 1 1 1276
0 1278 7 1 2 72876 1277
0 1279 5 1 1 1278
0 1280 7 6 2 69696 78673
0 1281 5 11 1 79897
0 1282 7 2 2 79898 79246
0 1283 5 1 1 79914
0 1284 7 4 2 66434 76535
0 1285 5 1 1 79916
0 1286 7 1 2 78831 1285
0 1287 5 1 1 1286
0 1288 7 8 2 69349 73322
0 1289 5 4 1 79920
0 1290 7 2 2 79921 79917
0 1291 5 1 1 79932
0 1292 7 1 2 1287 1291
0 1293 5 1 1 1292
0 1294 7 1 2 67867 1293
0 1295 5 1 1 1294
0 1296 7 1 2 1283 1295
0 1297 7 1 2 1279 1296
0 1298 5 1 1 1297
0 1299 7 1 2 77642 1298
0 1300 5 1 1 1299
0 1301 7 1 2 1258 1300
0 1302 5 1 1 1301
0 1303 7 1 2 70955 1302
0 1304 5 1 1 1303
0 1305 7 5 2 69697 75688
0 1306 5 3 1 79934
0 1307 7 7 2 76267 78824
0 1308 5 25 1 79942
0 1309 7 1 2 71535 79943
0 1310 5 1 1 1309
0 1311 7 1 2 79939 1310
0 1312 5 1 1 1311
0 1313 7 1 2 65878 1312
0 1314 5 1 1 1313
0 1315 7 1 2 77695 77812
0 1316 5 2 1 1315
0 1317 7 1 2 1314 79974
0 1318 5 1 1 1317
0 1319 7 10 2 69350 65268
0 1320 5 1 1 79976
0 1321 7 1 2 79977 74110
0 1322 7 1 2 1318 1321
0 1323 5 1 1 1322
0 1324 7 1 2 1304 1323
0 1325 5 1 1 1324
0 1326 7 1 2 73645 1325
0 1327 5 1 1 1326
0 1328 7 5 2 64551 74989
0 1329 5 6 1 79986
0 1330 7 5 2 65879 75949
0 1331 7 2 2 79991 79997
0 1332 5 1 1 80002
0 1333 7 1 2 74836 80003
0 1334 5 2 1 1333
0 1335 7 33 2 69351 64552
0 1336 5 3 1 80006
0 1337 7 1 2 76017 80007
0 1338 5 2 1 1337
0 1339 7 1 2 80004 80042
0 1340 5 1 1 1339
0 1341 7 5 2 67868 76174
0 1342 7 3 2 69352 78586
0 1343 7 2 2 80044 80049
0 1344 5 2 1 80052
0 1345 7 1 2 66435 80054
0 1346 5 1 1 1345
0 1347 7 2 2 70053 1346
0 1348 7 1 2 1340 80056
0 1349 5 1 1 1348
0 1350 7 8 2 68553 77389
0 1351 7 21 2 66122 71536
0 1352 5 1 1 80066
0 1353 7 7 2 70054 68258
0 1354 5 12 1 80087
0 1355 7 4 2 80067 80088
0 1356 5 1 1 80106
0 1357 7 1 2 80058 80107
0 1358 5 1 1 1357
0 1359 7 23 2 64938 70956
0 1360 7 4 2 69698 79567
0 1361 7 3 2 80110 80133
0 1362 5 1 1 80137
0 1363 7 1 2 1358 1362
0 1364 5 1 1 1363
0 1365 7 1 2 72877 1364
0 1366 5 1 1 1365
0 1367 7 4 2 66436 74866
0 1368 5 2 1 80140
0 1369 7 1 2 80144 80053
0 1370 5 2 1 1369
0 1371 7 1 2 1366 80146
0 1372 7 1 2 1349 1371
0 1373 5 1 1 1372
0 1374 7 1 2 77506 1373
0 1375 5 1 1 1374
0 1376 7 1 2 1327 1375
0 1377 5 1 1 1376
0 1378 7 1 2 74016 1377
0 1379 5 1 1 1378
0 1380 7 8 2 69699 74931
0 1381 5 14 1 80148
0 1382 7 12 2 75950 79992
0 1383 7 2 2 75313 80170
0 1384 5 1 1 80182
0 1385 7 1 2 80156 1384
0 1386 5 2 1 1385
0 1387 7 1 2 78023 77549
0 1388 5 1 1 1387
0 1389 7 1 2 79781 79397
0 1390 7 1 2 1388 1389
0 1391 7 1 2 80184 1390
0 1392 5 1 1 1391
0 1393 7 1 2 1379 1392
0 1394 7 1 2 1242 1393
0 1395 7 1 2 1099 1394
0 1396 5 1 1 1395
0 1397 7 1 2 78532 1396
0 1398 5 1 1 1397
0 1399 7 1 2 791 1398
0 1400 7 1 2 719 1399
0 1401 5 1 1 1400
0 1402 7 1 2 66622 1401
0 1403 5 1 1 1402
0 1404 7 10 2 79623 74447
0 1405 7 11 2 65711 71713
0 1406 7 10 2 64014 70321
0 1407 7 2 2 80196 80207
0 1408 7 3 2 76268 77135
0 1409 5 1 1 80219
0 1410 7 17 2 68259 75314
0 1411 5 12 1 80222
0 1412 7 3 2 65880 76536
0 1413 5 4 1 80251
0 1414 7 3 2 64243 76537
0 1415 5 11 1 80258
0 1416 7 4 2 80254 80261
0 1417 5 1 1 80272
0 1418 7 7 2 77390 80273
0 1419 7 1 2 80223 80276
0 1420 5 1 1 1419
0 1421 7 1 2 1409 1420
0 1422 5 1 1 1421
0 1423 7 1 2 80217 1422
0 1424 5 1 1 1423
0 1425 7 23 2 70055 70322
0 1426 5 3 1 80283
0 1427 7 2 2 64553 80306
0 1428 5 1 1 80309
0 1429 7 11 2 65881 66437
0 1430 5 1 1 80311
0 1431 7 2 2 77958 80312
0 1432 7 1 2 80310 80322
0 1433 7 1 2 78000 1432
0 1434 5 1 1 1433
0 1435 7 1 2 1424 1434
0 1436 5 1 1 1435
0 1437 7 1 2 72878 1436
0 1438 5 1 1 1437
0 1439 7 6 2 69353 76700
0 1440 5 1 1 80324
0 1441 7 53 2 71714 68554
0 1442 5 51 1 80330
0 1443 7 5 2 64939 80383
0 1444 5 9 1 80434
0 1445 7 2 2 80435 78609
0 1446 5 5 1 80448
0 1447 7 1 2 80325 80450
0 1448 5 1 1 1447
0 1449 7 5 2 69700 77391
0 1450 5 1 1 80455
0 1451 7 10 2 71537 71715
0 1452 5 4 1 80460
0 1453 7 9 2 70323 73323
0 1454 5 2 1 80474
0 1455 7 1 2 80461 80475
0 1456 5 3 1 1455
0 1457 7 5 2 66438 80384
0 1458 5 9 1 80488
0 1459 7 7 2 73324 80385
0 1460 5 23 1 80502
0 1461 7 2 2 80493 80509
0 1462 7 5 2 78674 80532
0 1463 7 1 2 65269 80534
0 1464 5 1 1 1463
0 1465 7 1 2 80485 1464
0 1466 5 1 1 1465
0 1467 7 1 2 70056 1466
0 1468 5 1 1 1467
0 1469 7 11 2 65270 71716
0 1470 5 1 1 80539
0 1471 7 8 2 68555 80540
0 1472 5 1 1 80550
0 1473 7 1 2 73887 80551
0 1474 5 1 1 1473
0 1475 7 1 2 1440 1474
0 1476 7 1 2 1468 1475
0 1477 5 1 1 1476
0 1478 7 1 2 80456 1477
0 1479 5 1 1 1478
0 1480 7 1 2 1448 1479
0 1481 5 1 1 1480
0 1482 7 1 2 75951 1481
0 1483 5 1 1 1482
0 1484 7 3 2 77392 78050
0 1485 7 108 2 70324 71717
0 1486 5 119 1 80561
0 1487 7 5 2 71538 73325
0 1488 5 1 1 80788
0 1489 7 6 2 70057 80789
0 1490 5 5 1 80793
0 1491 7 1 2 80562 80794
0 1492 5 3 1 1491
0 1493 7 8 2 80331 73888
0 1494 5 2 1 80807
0 1495 7 1 2 70058 80535
0 1496 5 2 1 1495
0 1497 7 2 2 80815 80817
0 1498 5 3 1 80819
0 1499 7 1 2 69701 80451
0 1500 5 1 1 1499
0 1501 7 1 2 80820 1500
0 1502 5 1 1 1501
0 1503 7 1 2 65271 1502
0 1504 5 1 1 1503
0 1505 7 1 2 80804 1504
0 1506 5 1 1 1505
0 1507 7 1 2 80558 1506
0 1508 5 1 1 1507
0 1509 7 18 2 69702 70957
0 1510 5 1 1 80824
0 1511 7 2 2 80563 80825
0 1512 7 15 2 70059 68556
0 1513 5 19 1 80844
0 1514 7 8 2 69354 71539
0 1515 5 3 1 80878
0 1516 7 1 2 80845 80879
0 1517 5 2 1 1516
0 1518 7 1 2 80842 80889
0 1519 5 1 1 1518
0 1520 7 12 2 69703 70325
0 1521 5 2 1 80891
0 1522 7 6 2 71718 80892
0 1523 5 2 1 80905
0 1524 7 1 2 65882 80911
0 1525 5 1 1 1524
0 1526 7 1 2 69355 521
0 1527 7 1 2 1525 1526
0 1528 5 1 1 1527
0 1529 7 1 2 1519 1528
0 1530 5 1 1 1529
0 1531 7 1 2 71246 1530
0 1532 5 1 1 1531
0 1533 7 2 2 80564 77136
0 1534 7 1 2 76538 80913
0 1535 5 1 1 1534
0 1536 7 1 2 1532 1535
0 1537 5 1 1 1536
0 1538 7 1 2 67869 1537
0 1539 5 1 1 1538
0 1540 7 1 2 1508 1539
0 1541 7 1 2 1483 1540
0 1542 5 1 1 1541
0 1543 7 1 2 74369 1542
0 1544 5 1 1 1543
0 1545 7 1 2 1438 1544
0 1546 5 1 1 1545
0 1547 7 1 2 72508 1546
0 1548 5 1 1 1547
0 1549 7 3 2 70060 78675
0 1550 5 11 1 80915
0 1551 7 2 2 73934 80918
0 1552 5 19 1 80929
0 1553 7 3 2 72879 77393
0 1554 7 1 2 66123 80950
0 1555 5 1 1 1554
0 1556 7 1 2 1332 1555
0 1557 5 3 1 1556
0 1558 7 1 2 80931 80953
0 1559 5 1 1 1558
0 1560 7 1 2 80043 1559
0 1561 5 1 1 1560
0 1562 7 1 2 79700 1561
0 1563 5 1 1 1562
0 1564 7 1 2 66439 80859
0 1565 5 5 1 1564
0 1566 7 2 2 69704 80956
0 1567 5 2 1 80961
0 1568 7 1 2 80963 76928
0 1569 5 1 1 1568
0 1570 7 4 2 71540 79552
0 1571 5 1 1 80965
0 1572 7 1 2 80966 77394
0 1573 5 1 1 1572
0 1574 7 1 2 1569 1573
0 1575 5 1 1 1574
0 1576 7 1 2 73326 1575
0 1577 5 1 1 1576
0 1578 7 8 2 66124 75315
0 1579 7 2 2 80008 80969
0 1580 5 1 1 80977
0 1581 7 1 2 68260 80978
0 1582 5 1 1 1581
0 1583 7 18 2 69356 65883
0 1584 5 4 1 80979
0 1585 7 12 2 78388 80997
0 1586 5 74 1 81001
0 1587 7 4 2 69705 81013
0 1588 5 1 1 81087
0 1589 7 4 2 71247 81014
0 1590 5 1 1 81091
0 1591 7 3 2 1588 1590
0 1592 5 1 1 81095
0 1593 7 1 2 72880 81096
0 1594 7 1 2 1582 1593
0 1595 7 1 2 1577 1594
0 1596 5 1 1 1595
0 1597 7 3 2 73327 79164
0 1598 7 1 2 80860 81098
0 1599 5 1 1 1598
0 1600 7 1 2 81002 1599
0 1601 5 1 1 1600
0 1602 7 1 2 76539 1601
0 1603 5 1 1 1602
0 1604 7 1 2 79247 76625
0 1605 5 1 1 1604
0 1606 7 11 2 65884 73328
0 1607 7 5 2 70061 81101
0 1608 5 3 1 81112
0 1609 7 1 2 71541 81113
0 1610 5 1 1 1609
0 1611 7 1 2 1605 1610
0 1612 5 1 1 1611
0 1613 7 1 2 69706 1612
0 1614 5 1 1 1613
0 1615 7 1 2 79460 80795
0 1616 5 1 1 1615
0 1617 7 5 2 64554 76867
0 1618 5 1 1 81120
0 1619 7 1 2 80861 81121
0 1620 5 1 1 1619
0 1621 7 1 2 67870 1620
0 1622 7 1 2 1616 1621
0 1623 7 1 2 1614 1622
0 1624 7 1 2 1603 1623
0 1625 5 1 1 1624
0 1626 7 1 2 1596 1625
0 1627 5 1 1 1626
0 1628 7 20 2 69707 70062
0 1629 5 2 1 81125
0 1630 7 4 2 65885 81126
0 1631 7 1 2 73329 77708
0 1632 7 1 2 81147 1631
0 1633 5 1 1 1632
0 1634 7 1 2 1627 1633
0 1635 5 1 1 1634
0 1636 7 1 2 70326 1635
0 1637 5 1 1 1636
0 1638 7 1 2 1563 1637
0 1639 5 1 1 1638
0 1640 7 1 2 71719 1639
0 1641 5 1 1 1640
0 1642 7 13 2 72881 76175
0 1643 7 1 2 77137 81151
0 1644 5 1 1 1643
0 1645 7 2 2 74811 80068
0 1646 5 2 1 81164
0 1647 7 3 2 64244 75614
0 1648 5 1 1 81168
0 1649 7 8 2 64555 73330
0 1650 5 7 1 81171
0 1651 7 5 2 80919 77595
0 1652 5 6 1 81186
0 1653 7 1 2 81179 81187
0 1654 5 1 1 1653
0 1655 7 1 2 1648 1654
0 1656 5 1 1 1655
0 1657 7 1 2 71248 1656
0 1658 5 1 1 1657
0 1659 7 1 2 66125 74768
0 1660 5 3 1 1659
0 1661 7 19 2 64245 67871
0 1662 5 7 1 81200
0 1663 7 1 2 81197 81219
0 1664 5 1 1 1663
0 1665 7 1 2 69708 1664
0 1666 5 1 1 1665
0 1667 7 18 2 69357 72882
0 1668 5 9 1 81226
0 1669 7 1 2 68261 78927
0 1670 5 1 1 1669
0 1671 7 1 2 81244 1670
0 1672 5 1 1 1671
0 1673 7 1 2 76540 1672
0 1674 5 2 1 1673
0 1675 7 1 2 1666 81253
0 1676 7 2 2 1658 1675
0 1677 5 1 1 81255
0 1678 7 1 2 81166 81256
0 1679 5 1 1 1678
0 1680 7 1 2 70958 1679
0 1681 5 1 1 1680
0 1682 7 8 2 69358 76176
0 1683 5 4 1 81257
0 1684 7 3 2 65886 76269
0 1685 5 2 1 81269
0 1686 7 2 2 66126 74588
0 1687 5 17 1 81274
0 1688 7 2 2 76636 81276
0 1689 5 1 1 81293
0 1690 7 1 2 81270 81294
0 1691 5 1 1 1690
0 1692 7 1 2 81265 1691
0 1693 5 2 1 1692
0 1694 7 1 2 68262 81295
0 1695 5 1 1 1694
0 1696 7 8 2 75244 76177
0 1697 5 1 1 81297
0 1698 7 1 2 69359 77584
0 1699 7 1 2 1697 1698
0 1700 5 1 1 1699
0 1701 7 1 2 1695 1700
0 1702 5 1 1 1701
0 1703 7 1 2 67872 1702
0 1704 5 1 1 1703
0 1705 7 10 2 68263 74502
0 1706 5 8 1 81305
0 1707 7 3 2 69709 79461
0 1708 5 5 1 81323
0 1709 7 1 2 69360 75895
0 1710 5 5 1 1709
0 1711 7 1 2 81326 81331
0 1712 5 2 1 1711
0 1713 7 1 2 81306 81336
0 1714 5 1 1 1713
0 1715 7 1 2 1704 1714
0 1716 7 1 2 1681 1715
0 1717 5 1 1 1716
0 1718 7 1 2 65272 1717
0 1719 5 1 1 1718
0 1720 7 1 2 1644 1719
0 1721 7 1 2 1641 1720
0 1722 5 1 1 1721
0 1723 7 1 2 78533 1722
0 1724 5 1 1 1723
0 1725 7 1 2 1548 1724
0 1726 5 1 1 1725
0 1727 7 1 2 80186 1726
0 1728 5 1 1 1727
0 1729 7 14 2 74017 75871
0 1730 7 3 2 68264 78920
0 1731 5 1 1 81352
0 1732 7 11 2 71542 74769
0 1733 5 5 1 81355
0 1734 7 1 2 81366 74749
0 1735 5 7 1 1734
0 1736 7 2 2 70063 81371
0 1737 5 2 1 81378
0 1738 7 2 2 71543 74719
0 1739 5 1 1 81382
0 1740 7 1 2 81380 1739
0 1741 5 1 1 1740
0 1742 7 1 2 68557 1741
0 1743 5 2 1 1742
0 1744 7 1 2 1731 81384
0 1745 5 1 1 1744
0 1746 7 1 2 70327 1745
0 1747 5 1 1 1746
0 1748 7 1 2 79928 1747
0 1749 5 1 1 1748
0 1750 7 1 2 72509 1749
0 1751 5 1 1 1750
0 1752 7 21 2 67501 73331
0 1753 5 1 1 81386
0 1754 7 18 2 72510 68265
0 1755 7 21 2 70328 67873
0 1756 5 1 1 81425
0 1757 7 1 2 81407 81426
0 1758 5 2 1 1757
0 1759 7 1 2 1753 81446
0 1760 5 1 1 1759
0 1761 7 1 2 64246 1760
0 1762 5 1 1 1761
0 1763 7 2 2 77859 81387
0 1764 5 2 1 81448
0 1765 7 1 2 81450 81447
0 1766 5 1 1 1765
0 1767 7 1 2 64940 1766
0 1768 5 1 1 1767
0 1769 7 1 2 1762 1768
0 1770 7 1 2 1751 1769
0 1771 5 1 1 1770
0 1772 7 1 2 71249 1771
0 1773 5 1 1 1772
0 1774 7 39 2 69361 72511
0 1775 5 5 1 81452
0 1776 7 15 2 73332 75316
0 1777 5 1 1 81496
0 1778 7 1 2 74806 1777
0 1779 5 2 1 1778
0 1780 7 1 2 78011 81511
0 1781 5 1 1 1780
0 1782 7 1 2 74750 1781
0 1783 5 1 1 1782
0 1784 7 1 2 81453 1783
0 1785 5 1 1 1784
0 1786 7 1 2 72883 79816
0 1787 5 2 1 1786
0 1788 7 28 2 64247 67502
0 1789 5 3 1 81515
0 1790 7 1 2 75585 81516
0 1791 7 1 2 81513 1790
0 1792 5 1 1 1791
0 1793 7 1 2 1785 1792
0 1794 7 1 2 1773 1793
0 1795 5 1 1 1794
0 1796 7 1 2 69710 1795
0 1797 5 1 1 1796
0 1798 7 2 2 64248 77550
0 1799 5 1 1 81546
0 1800 7 5 2 77563 1799
0 1801 5 1 1 81548
0 1802 7 7 2 72512 75317
0 1803 7 2 2 81549 81553
0 1804 7 1 2 75112 81560
0 1805 5 1 1 1804
0 1806 7 5 2 70064 79061
0 1807 5 1 1 81562
0 1808 7 1 2 67503 81563
0 1809 7 1 2 79747 1808
0 1810 5 1 1 1809
0 1811 7 1 2 1805 1810
0 1812 5 1 1 1811
0 1813 7 1 2 73333 1812
0 1814 5 1 1 1813
0 1815 7 1 2 76037 79428
0 1816 5 11 1 1815
0 1817 7 11 2 65273 66440
0 1818 5 3 1 81578
0 1819 7 7 2 64941 81579
0 1820 5 1 1 81592
0 1821 7 1 2 73646 81593
0 1822 5 1 1 1821
0 1823 7 1 2 69362 1822
0 1824 5 1 1 1823
0 1825 7 1 2 81567 1824
0 1826 5 1 1 1825
0 1827 7 1 2 70065 75113
0 1828 5 7 1 1827
0 1829 7 1 2 81599 80045
0 1830 5 1 1 1829
0 1831 7 1 2 64249 78735
0 1832 5 1 1 1831
0 1833 7 1 2 67504 1832
0 1834 7 1 2 1830 1833
0 1835 7 1 2 1826 1834
0 1836 5 1 1 1835
0 1837 7 1 2 69363 81277
0 1838 5 1 1 1837
0 1839 7 1 2 64556 1838
0 1840 5 1 1 1839
0 1841 7 10 2 71544 77797
0 1842 5 4 1 81606
0 1843 7 3 2 64250 81616
0 1844 5 3 1 81620
0 1845 7 3 2 72884 75114
0 1846 5 1 1 81626
0 1847 7 1 2 81623 81627
0 1848 7 1 2 1840 1847
0 1849 5 1 1 1848
0 1850 7 2 2 67874 80262
0 1851 7 3 2 71545 76949
0 1852 7 2 2 81631 77798
0 1853 5 1 1 81634
0 1854 7 1 2 81629 1853
0 1855 5 1 1 1854
0 1856 7 1 2 72513 1855
0 1857 7 1 2 1849 1856
0 1858 5 1 1 1857
0 1859 7 1 2 68266 1858
0 1860 7 1 2 1836 1859
0 1861 5 1 1 1860
0 1862 7 1 2 1814 1861
0 1863 5 1 1 1862
0 1864 7 1 2 71720 1863
0 1865 5 1 1 1864
0 1866 7 1 2 77935 78144
0 1867 5 2 1 1866
0 1868 7 3 2 68267 81278
0 1869 5 1 1 81638
0 1870 7 2 2 72514 81639
0 1871 7 1 2 78012 81641
0 1872 5 1 1 1871
0 1873 7 1 2 81636 1872
0 1874 5 1 1 1873
0 1875 7 1 2 72885 1874
0 1876 5 1 1 1875
0 1877 7 8 2 71250 74720
0 1878 5 3 1 81643
0 1879 7 1 2 68268 78902
0 1880 5 4 1 1879
0 1881 7 3 2 68558 75952
0 1882 5 1 1 81658
0 1883 7 2 2 75318 81659
0 1884 7 1 2 73334 81661
0 1885 5 1 1 1884
0 1886 7 1 2 81654 1885
0 1887 5 1 1 1886
0 1888 7 1 2 70329 1887
0 1889 5 1 1 1888
0 1890 7 1 2 81651 1889
0 1891 5 1 1 1890
0 1892 7 1 2 72515 1891
0 1893 5 1 1 1892
0 1894 7 1 2 1876 1893
0 1895 5 1 1 1894
0 1896 7 1 2 69364 1895
0 1897 5 1 1 1896
0 1898 7 6 2 64557 78949
0 1899 5 3 1 81663
0 1900 7 1 2 80263 81669
0 1901 5 1 1 1900
0 1902 7 1 2 67875 1901
0 1903 5 1 1 1902
0 1904 7 1 2 64251 76044
0 1905 5 1 1 1904
0 1906 7 1 2 1903 1905
0 1907 5 1 1 1906
0 1908 7 1 2 79799 1907
0 1909 5 1 1 1908
0 1910 7 1 2 64252 81644
0 1911 5 1 1 1910
0 1912 7 1 2 1909 1911
0 1913 5 1 1 1912
0 1914 7 1 2 67505 1913
0 1915 5 1 1 1914
0 1916 7 1 2 1897 1915
0 1917 7 1 2 1865 1916
0 1918 7 1 2 1797 1917
0 1919 5 1 1 1918
0 1920 7 1 2 70959 1919
0 1921 5 1 1 1920
0 1922 7 137 2 65274 66623
0 1923 5 145 1 81672
0 1924 7 20 2 71251 72516
0 1925 5 1 1 81954
0 1926 7 3 2 76950 81955
0 1927 5 1 1 81974
0 1928 7 2 2 65887 75543
0 1929 5 1 1 81977
0 1930 7 1 2 81385 1929
0 1931 5 1 1 1930
0 1932 7 1 2 81975 1931
0 1933 5 1 1 1932
0 1934 7 1 2 69365 80252
0 1935 5 2 1 1934
0 1936 7 7 2 70960 71546
0 1937 5 4 1 81981
0 1938 7 4 2 64253 81988
0 1939 5 1 1 81992
0 1940 7 1 2 76437 81993
0 1941 5 1 1 1940
0 1942 7 1 2 81979 1941
0 1943 5 2 1 1942
0 1944 7 1 2 67876 81996
0 1945 5 1 1 1944
0 1946 7 19 2 64558 70066
0 1947 7 2 2 81998 80069
0 1948 5 3 1 82017
0 1949 7 1 2 81272 82019
0 1950 5 1 1 1949
0 1951 7 1 2 81227 1950
0 1952 5 1 1 1951
0 1953 7 1 2 68269 1952
0 1954 7 1 2 1945 1953
0 1955 5 1 1 1954
0 1956 7 12 2 67877 75319
0 1957 5 16 1 82022
0 1958 7 10 2 66127 80009
0 1959 5 4 1 82050
0 1960 7 1 2 82023 82051
0 1961 5 2 1 1960
0 1962 7 1 2 73335 82064
0 1963 5 2 1 1962
0 1964 7 1 2 67506 82066
0 1965 7 1 2 1955 1964
0 1966 5 1 1 1965
0 1967 7 1 2 1933 1966
0 1968 5 1 1 1967
0 1969 7 1 2 81809 1968
0 1970 5 1 1 1969
0 1971 7 3 2 67507 76270
0 1972 5 2 1 82068
0 1973 7 2 2 81102 82069
0 1974 5 1 1 82073
0 1975 7 1 2 74127 82074
0 1976 5 1 1 1975
0 1977 7 10 2 72886 74503
0 1978 5 1 1 82075
0 1979 7 3 2 76438 81408
0 1980 5 1 1 82085
0 1981 7 2 2 66128 81388
0 1982 5 2 1 82088
0 1983 7 1 2 68559 82089
0 1984 5 1 1 1983
0 1985 7 1 2 1980 1984
0 1986 5 1 1 1985
0 1987 7 1 2 82076 1986
0 1988 5 1 1 1987
0 1989 7 35 2 73336 68560
0 1990 5 2 1 82092
0 1991 7 21 2 64559 67508
0 1992 7 3 2 76018 82129
0 1993 5 2 1 82150
0 1994 7 1 2 82093 82151
0 1995 5 1 1 1994
0 1996 7 6 2 72517 74721
0 1997 7 1 2 76439 82155
0 1998 5 2 1 1997
0 1999 7 13 2 64560 68270
0 2000 5 7 1 82163
0 2001 7 23 2 66129 67509
0 2002 5 1 1 82183
0 2003 7 3 2 82164 82184
0 2004 5 1 1 82206
0 2005 7 1 2 79712 82207
0 2006 5 1 1 2005
0 2007 7 1 2 82161 2006
0 2008 5 1 1 2007
0 2009 7 1 2 75320 2008
0 2010 5 1 1 2009
0 2011 7 1 2 1995 2010
0 2012 7 1 2 1988 2011
0 2013 5 1 1 2012
0 2014 7 1 2 69366 2013
0 2015 5 1 1 2014
0 2016 7 2 2 68561 80171
0 2017 7 10 2 71547 67510
0 2018 7 1 2 81114 82211
0 2019 7 1 2 82209 2018
0 2020 5 1 1 2019
0 2021 7 1 2 2015 2020
0 2022 5 1 1 2021
0 2023 7 1 2 80565 2022
0 2024 5 1 1 2023
0 2025 7 1 2 1976 2024
0 2026 7 1 2 1970 2025
0 2027 7 1 2 1921 2026
0 2028 5 1 1 2027
0 2029 7 1 2 74370 2028
0 2030 5 1 1 2029
0 2031 7 9 2 73337 77039
0 2032 5 2 1 82221
0 2033 7 2 2 78286 82222
0 2034 5 1 1 82232
0 2035 7 20 2 72518 72887
0 2036 5 1 1 82234
0 2037 7 2 2 70761 82235
0 2038 5 1 1 82254
0 2039 7 1 2 78306 82255
0 2040 7 1 2 82233 2039
0 2041 5 1 1 2040
0 2042 7 1 2 2030 2041
0 2043 5 1 1 2042
0 2044 7 1 2 81338 2043
0 2045 5 1 1 2044
0 2046 7 1 2 1728 2045
0 2047 5 1 1 2046
0 2048 7 1 2 71991 2047
0 2049 5 1 1 2048
0 2050 7 3 2 81810 77395
0 2051 7 1 2 81127 82256
0 2052 5 1 1 2051
0 2053 7 1 2 77202 2052
0 2054 5 1 1 2053
0 2055 7 1 2 78676 2054
0 2056 5 1 1 2055
0 2057 7 4 2 69367 80826
0 2058 5 1 1 82259
0 2059 7 3 2 69711 73889
0 2060 5 2 1 82263
0 2061 7 1 2 77203 82266
0 2062 5 2 1 2061
0 2063 7 10 2 66624 75498
0 2064 5 7 1 82270
0 2065 7 1 2 77396 82280
0 2066 7 1 2 82268 2065
0 2067 5 1 1 2066
0 2068 7 1 2 2058 2067
0 2069 7 1 2 2056 2068
0 2070 5 1 1 2069
0 2071 7 1 2 75953 2070
0 2072 5 1 1 2071
0 2073 7 2 2 69368 74932
0 2074 5 1 1 82287
0 2075 7 1 2 70961 82288
0 2076 5 1 1 2075
0 2077 7 4 2 64561 73935
0 2078 5 10 1 82289
0 2079 7 1 2 79903 82271
0 2080 5 1 1 2079
0 2081 7 1 2 82293 2080
0 2082 5 1 1 2081
0 2083 7 9 2 70067 81811
0 2084 5 22 1 82303
0 2085 7 1 2 82304 78677
0 2086 5 2 1 2085
0 2087 7 1 2 2082 82334
0 2088 5 1 1 2087
0 2089 7 1 2 80559 2088
0 2090 5 1 1 2089
0 2091 7 1 2 2076 2090
0 2092 7 1 2 2072 2091
0 2093 5 1 1 2092
0 2094 7 1 2 64015 2093
0 2095 5 1 1 2094
0 2096 7 25 2 71721 68271
0 2097 5 14 1 82336
0 2098 7 19 2 65888 71548
0 2099 7 3 2 80284 82375
0 2100 7 3 2 82337 82394
0 2101 5 1 1 82397
0 2102 7 6 2 66130 68562
0 2103 5 1 1 82400
0 2104 7 2 2 69369 79407
0 2105 7 1 2 82401 82406
0 2106 7 1 2 82398 2105
0 2107 5 1 1 2106
0 2108 7 1 2 2095 2107
0 2109 5 1 1 2108
0 2110 7 1 2 65712 2109
0 2111 5 1 1 2110
0 2112 7 10 2 70330 65713
0 2113 7 2 2 82408 81128
0 2114 7 2 2 80332 76929
0 2115 7 1 2 82418 82420
0 2116 5 1 1 2115
0 2117 7 61 2 69095 70762
0 2118 5 33 1 82422
0 2119 7 2 2 80333 80285
0 2120 5 4 1 82516
0 2121 7 1 2 82483 82518
0 2122 5 1 1 2121
0 2123 7 11 2 64562 65889
0 2124 5 1 1 82522
0 2125 7 7 2 66131 82523
0 2126 7 1 2 74416 82533
0 2127 7 1 2 2122 2126
0 2128 5 1 1 2127
0 2129 7 1 2 2116 2128
0 2130 5 1 1 2129
0 2131 7 1 2 64254 77884
0 2132 7 1 2 2130 2131
0 2133 5 1 1 2132
0 2134 7 1 2 2111 2133
0 2135 5 1 1 2134
0 2136 7 1 2 72519 2135
0 2137 5 1 1 2136
0 2138 7 15 2 65714 67511
0 2139 5 3 1 82540
0 2140 7 11 2 70962 72888
0 2141 5 1 1 82558
0 2142 7 3 2 69370 82559
0 2143 5 3 1 82569
0 2144 7 9 2 67878 77397
0 2145 5 1 1 82575
0 2146 7 29 2 66625 73338
0 2147 5 15 1 82584
0 2148 7 14 2 65275 82585
0 2149 5 16 1 82628
0 2150 7 3 2 64563 82642
0 2151 5 2 1 82658
0 2152 7 1 2 82576 82659
0 2153 5 1 1 2152
0 2154 7 1 2 82572 2153
0 2155 5 1 1 2154
0 2156 7 1 2 64016 2155
0 2157 5 1 1 2156
0 2158 7 11 2 65890 71722
0 2159 7 2 2 64564 82663
0 2160 7 1 2 68563 74807
0 2161 7 9 2 64255 66441
0 2162 5 2 1 82676
0 2163 7 1 2 74131 1488
0 2164 7 1 2 82685 2163
0 2165 7 3 2 2160 2164
0 2166 7 1 2 82674 82687
0 2167 5 1 1 2166
0 2168 7 11 2 64017 77398
0 2169 5 6 1 82690
0 2170 7 4 2 72889 78678
0 2171 7 1 2 82691 82707
0 2172 5 1 1 2171
0 2173 7 1 2 2167 2172
0 2174 5 1 1 2173
0 2175 7 1 2 70331 2174
0 2176 5 1 1 2175
0 2177 7 3 2 71549 82613
0 2178 5 2 1 82711
0 2179 7 2 2 82361 82714
0 2180 5 2 1 82716
0 2181 7 1 2 64018 80951
0 2182 7 1 2 82718 2181
0 2183 5 1 1 2182
0 2184 7 1 2 2176 2183
0 2185 5 1 1 2184
0 2186 7 1 2 70068 2185
0 2187 5 1 1 2186
0 2188 7 1 2 2157 2187
0 2189 5 1 1 2188
0 2190 7 1 2 66132 2189
0 2191 5 1 1 2190
0 2192 7 9 2 69712 67879
0 2193 5 17 1 82720
0 2194 7 2 2 81812 78610
0 2195 5 2 1 82746
0 2196 7 2 2 82729 82747
0 2197 5 1 1 82750
0 2198 7 1 2 75954 82692
0 2199 7 1 2 82751 2198
0 2200 5 1 1 2199
0 2201 7 1 2 2191 2200
0 2202 5 1 1 2201
0 2203 7 1 2 82541 2202
0 2204 5 1 1 2203
0 2205 7 1 2 2137 2204
0 2206 5 1 1 2205
0 2207 7 15 2 63727 63849
0 2208 7 5 2 66920 82752
0 2209 7 1 2 82767 75673
0 2210 7 1 2 2206 2209
0 2211 5 1 1 2210
0 2212 7 1 2 2049 2211
0 2213 5 1 1 2212
0 2214 7 1 2 66823 2213
0 2215 5 1 1 2214
0 2216 7 9 2 65715 71890
0 2217 7 3 2 64019 82772
0 2218 7 1 2 81600 81099
0 2219 5 1 1 2218
0 2220 7 10 2 64256 68272
0 2221 5 5 1 82784
0 2222 7 4 2 80439 80494
0 2223 5 2 1 82799
0 2224 7 2 2 75484 82800
0 2225 5 1 1 82805
0 2226 7 1 2 82785 82806
0 2227 5 1 1 2226
0 2228 7 1 2 2219 2227
0 2229 5 1 1 2228
0 2230 7 1 2 74458 2229
0 2231 5 1 1 2230
0 2232 7 25 2 65566 66921
0 2233 5 5 1 82807
0 2234 7 8 2 70069 66442
0 2235 5 1 1 82837
0 2236 7 3 2 80566 82094
0 2237 5 9 1 82845
0 2238 7 2 2 82838 82846
0 2239 5 4 1 82857
0 2240 7 2 2 80286 77279
0 2241 5 2 1 82863
0 2242 7 13 2 64942 71550
0 2243 5 1 1 82867
0 2244 7 62 2 66626 73647
0 2245 5 58 1 82880
0 2246 7 9 2 65276 82942
0 2247 5 5 1 83000
0 2248 7 1 2 82868 83001
0 2249 5 1 1 2248
0 2250 7 1 2 82865 2249
0 2251 5 1 1 2250
0 2252 7 1 2 68273 2251
0 2253 5 1 1 2252
0 2254 7 1 2 82859 2253
0 2255 5 1 1 2254
0 2256 7 1 2 82808 2255
0 2257 5 1 1 2256
0 2258 7 1 2 2231 2257
0 2259 5 1 1 2258
0 2260 7 1 2 67880 2259
0 2261 5 1 1 2260
0 2262 7 4 2 75321 82095
0 2263 5 1 1 83014
0 2264 7 1 2 2263 900
0 2265 5 3 1 2264
0 2266 7 1 2 74459 83018
0 2267 5 1 1 2266
0 2268 7 1 2 82832 2267
0 2269 5 1 1 2268
0 2270 7 1 2 81813 2269
0 2271 5 1 1 2270
0 2272 7 2 2 68564 82809
0 2273 5 1 1 83021
0 2274 7 9 2 80567 75322
0 2275 5 1 1 83023
0 2276 7 2 2 73339 74460
0 2277 5 1 1 83032
0 2278 7 1 2 83024 83033
0 2279 5 1 1 2278
0 2280 7 1 2 2273 2279
0 2281 7 1 2 2271 2280
0 2282 5 1 1 2281
0 2283 7 1 2 81228 2282
0 2284 5 1 1 2283
0 2285 7 1 2 2261 2284
0 2286 5 1 1 2285
0 2287 7 1 2 69713 2286
0 2288 5 1 1 2287
0 2289 7 1 2 76142 79758
0 2290 5 1 1 2289
0 2291 7 18 2 65277 73340
0 2292 5 6 1 83034
0 2293 7 1 2 83052 1846
0 2294 5 1 1 2293
0 2295 7 17 2 73648 81673
0 2296 5 6 1 83058
0 2297 7 1 2 80916 83075
0 2298 7 1 2 2294 2297
0 2299 5 1 1 2298
0 2300 7 1 2 2290 2299
0 2301 5 2 1 2300
0 2302 7 1 2 82810 83081
0 2303 5 1 1 2302
0 2304 7 6 2 67881 74461
0 2305 7 6 2 68274 75245
0 2306 5 3 1 83089
0 2307 7 5 2 73649 81814
0 2308 5 1 1 83098
0 2309 7 1 2 83090 83099
0 2310 7 1 2 83083 2309
0 2311 5 1 1 2310
0 2312 7 1 2 2303 2311
0 2313 5 1 1 2312
0 2314 7 1 2 69371 2313
0 2315 5 1 1 2314
0 2316 7 1 2 2288 2315
0 2317 5 1 1 2316
0 2318 7 1 2 68752 2317
0 2319 5 1 1 2318
0 2320 7 5 2 66922 74003
0 2321 7 8 2 65278 71551
0 2322 7 8 2 64943 67882
0 2323 7 2 2 68275 83116
0 2324 5 1 1 83124
0 2325 7 1 2 83108 83125
0 2326 5 2 1 2325
0 2327 7 1 2 83126 81245
0 2328 5 1 1 2327
0 2329 7 1 2 82943 2328
0 2330 5 1 1 2329
0 2331 7 4 2 80141 80510
0 2332 5 1 1 83128
0 2333 7 11 2 70070 67883
0 2334 5 3 1 83132
0 2335 7 1 2 83129 83133
0 2336 5 1 1 2335
0 2337 7 1 2 81246 2336
0 2338 5 1 1 2337
0 2339 7 1 2 70332 2338
0 2340 5 1 1 2339
0 2341 7 1 2 2330 2340
0 2342 5 1 1 2341
0 2343 7 1 2 69714 2342
0 2344 5 1 1 2343
0 2345 7 1 2 69372 83082
0 2346 5 1 1 2345
0 2347 7 1 2 2344 2346
0 2348 5 1 1 2347
0 2349 7 1 2 83103 2348
0 2350 5 1 1 2349
0 2351 7 1 2 2319 2350
0 2352 5 1 1 2351
0 2353 7 1 2 71252 2352
0 2354 5 1 1 2353
0 2355 7 9 2 70333 71552
0 2356 5 6 1 83146
0 2357 7 2 2 68276 75115
0 2358 5 5 1 83161
0 2359 7 1 2 83155 83163
0 2360 5 1 1 2359
0 2361 7 1 2 78759 2360
0 2362 5 1 1 2361
0 2363 7 7 2 73341 82944
0 2364 5 2 1 83168
0 2365 7 1 2 75615 83109
0 2366 7 1 2 83169 2365
0 2367 5 1 1 2366
0 2368 7 1 2 2362 2367
0 2369 5 1 1 2368
0 2370 7 17 2 69373 70071
0 2371 5 1 1 83177
0 2372 7 14 2 66923 74018
0 2373 5 1 1 83194
0 2374 7 1 2 83178 83195
0 2375 7 1 2 2369 2374
0 2376 5 1 1 2375
0 2377 7 1 2 2354 2376
0 2378 5 1 1 2377
0 2379 7 1 2 72520 2378
0 2380 5 1 1 2379
0 2381 7 1 2 79268 74019
0 2382 7 3 2 77799 83147
0 2383 7 15 2 66924 73342
0 2384 5 1 1 83211
0 2385 7 2 2 76143 83212
0 2386 7 1 2 83208 83226
0 2387 7 1 2 2381 2386
0 2388 5 1 1 2387
0 2389 7 1 2 2380 2388
0 2390 5 1 1 2389
0 2391 7 1 2 74448 2390
0 2392 5 1 1 2391
0 2393 7 4 2 64257 74933
0 2394 5 3 1 83228
0 2395 7 1 2 81332 83232
0 2396 5 2 1 2395
0 2397 7 1 2 64565 83235
0 2398 5 1 1 2397
0 2399 7 12 2 72890 76271
0 2400 5 3 1 83237
0 2401 7 1 2 76038 83249
0 2402 5 12 1 2401
0 2403 7 4 2 74504 83252
0 2404 5 1 1 83264
0 2405 7 1 2 64258 83265
0 2406 5 1 1 2405
0 2407 7 1 2 2398 2406
0 2408 5 1 1 2407
0 2409 7 1 2 73343 2408
0 2410 5 1 1 2409
0 2411 7 6 2 71253 79269
0 2412 5 2 1 83268
0 2413 7 4 2 72891 80862
0 2414 5 1 1 83276
0 2415 7 1 2 83269 83277
0 2416 5 1 1 2415
0 2417 7 1 2 2410 2416
0 2418 5 1 1 2417
0 2419 7 1 2 70334 2418
0 2420 5 1 1 2419
0 2421 7 6 2 72892 76440
0 2422 5 2 1 83280
0 2423 7 1 2 83253 80932
0 2424 5 1 1 2423
0 2425 7 1 2 83286 2424
0 2426 5 1 1 2425
0 2427 7 1 2 64259 79701
0 2428 7 1 2 2426 2427
0 2429 5 1 1 2428
0 2430 7 1 2 2420 2429
0 2431 5 1 1 2430
0 2432 7 1 2 71723 2431
0 2433 5 1 1 2432
0 2434 7 15 2 64260 65279
0 2435 7 1 2 74505 76064
0 2436 5 3 1 2435
0 2437 7 3 2 69715 76065
0 2438 5 5 1 83306
0 2439 7 26 2 69716 71553
0 2440 5 1 1 83314
0 2441 7 13 2 70072 72893
0 2442 5 1 1 83340
0 2443 7 1 2 83315 83341
0 2444 5 3 1 2443
0 2445 7 1 2 83309 83353
0 2446 7 1 2 83303 2445
0 2447 5 1 1 2446
0 2448 7 1 2 68277 2447
0 2449 5 2 1 2448
0 2450 7 6 2 64944 77860
0 2451 5 3 1 83358
0 2452 7 12 2 64945 73344
0 2453 5 5 1 83367
0 2454 7 1 2 67884 83379
0 2455 5 3 1 2454
0 2456 7 1 2 76441 83384
0 2457 7 1 2 83364 2456
0 2458 5 1 1 2457
0 2459 7 1 2 83356 2458
0 2460 5 1 1 2459
0 2461 7 1 2 83288 2460
0 2462 5 1 1 2461
0 2463 7 1 2 2433 2462
0 2464 5 1 1 2463
0 2465 7 1 2 74260 2464
0 2466 5 1 1 2465
0 2467 7 2 2 73650 79949
0 2468 7 1 2 82338 79978
0 2469 7 1 2 83387 2468
0 2470 5 1 1 2469
0 2471 7 12 2 66627 68278
0 2472 5 4 1 83389
0 2473 7 1 2 83401 81180
0 2474 7 1 2 83164 2473
0 2475 7 1 2 83229 2474
0 2476 5 1 1 2475
0 2477 7 1 2 2470 2476
0 2478 5 1 1 2477
0 2479 7 1 2 64946 2478
0 2480 5 1 1 2479
0 2481 7 9 2 69717 73651
0 2482 5 1 1 83405
0 2483 7 1 2 83406 83035
0 2484 7 1 2 83230 2483
0 2485 5 1 1 2484
0 2486 7 1 2 2480 2485
0 2487 5 1 1 2486
0 2488 7 1 2 76760 2487
0 2489 5 1 1 2488
0 2490 7 13 2 71724 73652
0 2491 5 2 1 83414
0 2492 7 1 2 83415 80476
0 2493 5 4 1 2492
0 2494 7 9 2 71725 73345
0 2495 5 4 1 83433
0 2496 7 6 2 70335 83434
0 2497 5 8 1 83446
0 2498 7 2 2 79203 83452
0 2499 5 5 1 83460
0 2500 7 1 2 64947 83462
0 2501 5 1 1 2500
0 2502 7 1 2 83429 2501
0 2503 5 1 1 2502
0 2504 7 2 2 79178 78970
0 2505 5 1 1 83467
0 2506 7 1 2 79264 2505
0 2507 5 1 1 2506
0 2508 7 1 2 2503 2507
0 2509 5 1 1 2508
0 2510 7 6 2 71726 72894
0 2511 7 7 2 70336 83469
0 2512 5 3 1 83475
0 2513 7 6 2 65280 74722
0 2514 5 1 1 83485
0 2515 7 1 2 83482 2514
0 2516 5 2 1 2515
0 2517 7 1 2 83270 83491
0 2518 5 1 1 2517
0 2519 7 1 2 2509 2518
0 2520 5 1 1 2519
0 2521 7 1 2 75204 2520
0 2522 5 1 1 2521
0 2523 7 1 2 2489 2522
0 2524 5 1 1 2523
0 2525 7 1 2 66443 2524
0 2526 5 1 1 2525
0 2527 7 15 2 70073 71727
0 2528 5 2 1 83493
0 2529 7 4 2 83494 82096
0 2530 5 3 1 83510
0 2531 7 2 2 83511 83148
0 2532 5 5 1 83517
0 2533 7 12 2 64948 68279
0 2534 5 2 1 83524
0 2535 7 15 2 70074 73346
0 2536 5 1 1 83538
0 2537 7 4 2 83536 2536
0 2538 5 11 1 83553
0 2539 7 3 2 81815 83557
0 2540 5 3 1 83568
0 2541 7 4 2 71728 74867
0 2542 7 1 2 83053 79341
0 2543 7 1 2 83574 2542
0 2544 5 1 1 2543
0 2545 7 1 2 83571 2544
0 2546 5 1 1 2545
0 2547 7 1 2 71254 2546
0 2548 5 1 1 2547
0 2549 7 1 2 83519 2548
0 2550 5 1 1 2549
0 2551 7 1 2 69718 2550
0 2552 5 1 1 2551
0 2553 7 9 2 71729 77080
0 2554 5 2 1 83578
0 2555 7 3 2 80287 83579
0 2556 5 1 1 83589
0 2557 7 2 2 73347 83590
0 2558 7 1 2 71255 83592
0 2559 5 1 1 2558
0 2560 7 1 2 2552 2559
0 2561 5 1 1 2560
0 2562 7 1 2 72895 2561
0 2563 5 1 1 2562
0 2564 7 13 2 71730 67885
0 2565 5 3 1 83594
0 2566 7 4 2 82097 83595
0 2567 7 1 2 80288 80070
0 2568 7 1 2 83610 2567
0 2569 5 1 1 2568
0 2570 7 1 2 2563 2569
0 2571 5 1 1 2570
0 2572 7 12 2 68923 64261
0 2573 7 1 2 83614 76832
0 2574 7 1 2 2571 2573
0 2575 5 1 1 2574
0 2576 7 1 2 2526 2575
0 2577 7 1 2 2466 2576
0 2578 5 1 1 2577
0 2579 7 1 2 78978 2578
0 2580 5 1 1 2579
0 2581 7 1 2 77627 78736
0 2582 5 1 1 2581
0 2583 7 3 2 76019 80495
0 2584 5 1 1 83626
0 2585 7 1 2 68280 83627
0 2586 5 1 1 2585
0 2587 7 1 2 2582 2586
0 2588 5 1 1 2587
0 2589 7 1 2 64262 2588
0 2590 5 1 1 2589
0 2591 7 1 2 79618 79933
0 2592 5 1 1 2591
0 2593 7 1 2 2590 2592
0 2594 5 1 1 2593
0 2595 7 1 2 70337 2594
0 2596 5 1 1 2595
0 2597 7 8 2 64263 71554
0 2598 7 2 2 77564 79183
0 2599 7 2 2 68565 83637
0 2600 7 1 2 83629 83639
0 2601 5 1 1 2600
0 2602 7 3 2 75246 83036
0 2603 5 2 1 83641
0 2604 7 1 2 69374 83644
0 2605 5 1 1 2604
0 2606 7 1 2 83281 2605
0 2607 5 1 1 2606
0 2608 7 4 2 64566 73890
0 2609 5 4 1 83646
0 2610 7 2 2 76020 83647
0 2611 5 2 1 83654
0 2612 7 1 2 75499 83655
0 2613 5 1 1 2612
0 2614 7 1 2 2607 2613
0 2615 5 1 1 2614
0 2616 7 1 2 82945 2615
0 2617 5 1 1 2616
0 2618 7 1 2 2601 2617
0 2619 7 1 2 2596 2618
0 2620 5 1 1 2619
0 2621 7 2 2 68924 74020
0 2622 7 1 2 74093 83658
0 2623 7 1 2 2620 2622
0 2624 5 1 1 2623
0 2625 7 1 2 2580 2624
0 2626 5 1 1 2625
0 2627 7 1 2 67512 2626
0 2628 5 1 1 2627
0 2629 7 12 2 65281 72896
0 2630 5 3 1 83660
0 2631 7 1 2 69375 83661
0 2632 5 2 1 2631
0 2633 7 6 2 68281 80568
0 2634 5 4 1 83677
0 2635 7 1 2 83678 81201
0 2636 5 2 1 2635
0 2637 7 1 2 83675 83687
0 2638 5 1 1 2637
0 2639 7 1 2 75323 2638
0 2640 5 1 1 2639
0 2641 7 1 2 74589 83492
0 2642 5 1 1 2641
0 2643 7 5 2 79707 79342
0 2644 5 15 1 83689
0 2645 7 4 2 72897 83694
0 2646 7 1 2 71731 83709
0 2647 5 1 1 2646
0 2648 7 1 2 2642 2647
0 2649 5 1 1 2648
0 2650 7 1 2 69376 2649
0 2651 5 1 1 2650
0 2652 7 1 2 2640 2651
0 2653 5 1 1 2652
0 2654 7 2 2 81956 74229
0 2655 7 2 2 78979 79080
0 2656 7 1 2 83713 83715
0 2657 7 1 2 2653 2656
0 2658 5 1 1 2657
0 2659 7 1 2 2628 2658
0 2660 7 1 2 2392 2659
0 2661 5 1 1 2660
0 2662 7 1 2 70963 2661
0 2663 5 1 1 2662
0 2664 7 19 2 65891 72521
0 2665 5 4 1 83717
0 2666 7 26 2 78494 83736
0 2667 5 1 1 83740
0 2668 7 2 2 69719 77289
0 2669 5 2 1 83766
0 2670 7 2 2 73348 83768
0 2671 5 1 1 83770
0 2672 7 1 2 81427 83771
0 2673 5 1 1 2672
0 2674 7 5 2 64949 73936
0 2675 5 6 1 83772
0 2676 7 12 2 78679 83777
0 2677 5 1 1 83783
0 2678 7 2 2 72898 83784
0 2679 5 2 1 83795
0 2680 7 1 2 79702 83796
0 2681 5 1 1 2680
0 2682 7 1 2 2673 2681
0 2683 5 1 1 2682
0 2684 7 1 2 71256 2683
0 2685 5 1 1 2684
0 2686 7 1 2 79703 78760
0 2687 7 1 2 80933 2686
0 2688 5 1 1 2687
0 2689 7 1 2 2685 2688
0 2690 5 1 1 2689
0 2691 7 1 2 71732 2690
0 2692 5 1 1 2691
0 2693 7 1 2 79020 76115
0 2694 5 1 1 2693
0 2695 7 1 2 74496 78932
0 2696 5 2 1 2695
0 2697 7 1 2 71257 83799
0 2698 5 1 1 2697
0 2699 7 1 2 78767 2698
0 2700 7 1 2 2694 2699
0 2701 5 1 1 2700
0 2702 7 1 2 83463 2701
0 2703 5 1 1 2702
0 2704 7 1 2 2692 2703
0 2705 5 1 1 2704
0 2706 7 1 2 69377 2705
0 2707 5 1 1 2706
0 2708 7 5 2 68566 81816
0 2709 5 12 1 83801
0 2710 7 2 2 73891 83802
0 2711 5 1 1 83818
0 2712 7 5 2 68567 78680
0 2713 5 5 1 83820
0 2714 7 1 2 71733 83821
0 2715 5 2 1 2714
0 2716 7 2 2 80470 74868
0 2717 5 2 1 83832
0 2718 7 1 2 70338 83834
0 2719 5 1 1 2718
0 2720 7 1 2 83830 2719
0 2721 5 1 1 2720
0 2722 7 1 2 70075 2721
0 2723 5 1 1 2722
0 2724 7 1 2 2711 2723
0 2725 5 1 1 2724
0 2726 7 2 2 74934 79270
0 2727 7 1 2 2725 83836
0 2728 5 1 1 2727
0 2729 7 1 2 2707 2728
0 2730 5 1 1 2729
0 2731 7 1 2 75173 2730
0 2732 5 1 1 2731
0 2733 7 1 2 70339 80496
0 2734 5 2 1 2733
0 2735 7 1 2 77092 83838
0 2736 5 2 1 2735
0 2737 7 9 2 69378 66133
0 2738 5 4 1 83842
0 2739 7 5 2 64264 76442
0 2740 5 2 1 83855
0 2741 7 1 2 83851 83860
0 2742 5 2 1 2741
0 2743 7 1 2 67886 83862
0 2744 7 1 2 83840 2743
0 2745 5 1 1 2744
0 2746 7 4 2 71258 68568
0 2747 5 1 1 83864
0 2748 7 1 2 64567 2747
0 2749 5 2 1 2748
0 2750 7 1 2 80880 83868
0 2751 7 1 2 81628 2750
0 2752 5 1 1 2751
0 2753 7 1 2 2745 2752
0 2754 5 1 1 2753
0 2755 7 2 2 79321 2754
0 2756 7 1 2 78068 83870
0 2757 5 1 1 2756
0 2758 7 1 2 2732 2757
0 2759 5 1 1 2758
0 2760 7 1 2 68753 2759
0 2761 5 1 1 2760
0 2762 7 2 2 70597 79358
0 2763 7 1 2 83872 83871
0 2764 5 1 1 2763
0 2765 7 1 2 2761 2764
0 2766 5 1 1 2765
0 2767 7 1 2 66925 2766
0 2768 5 1 1 2767
0 2769 7 1 2 83843 83447
0 2770 5 1 1 2769
0 2771 7 1 2 64265 79935
0 2772 5 1 1 2771
0 2773 7 1 2 2770 2772
0 2774 5 1 1 2773
0 2775 7 4 2 68925 74506
0 2776 7 9 2 71992 78980
0 2777 7 30 2 67887 68569
0 2778 5 3 1 83887
0 2779 7 2 2 67033 83888
0 2780 7 1 2 83878 83920
0 2781 7 1 2 83874 2780
0 2782 7 1 2 2774 2781
0 2783 5 1 1 2782
0 2784 7 1 2 2768 2783
0 2785 5 1 1 2784
0 2786 7 1 2 83741 2785
0 2787 5 1 1 2786
0 2788 7 1 2 83316 81957
0 2789 5 2 1 2788
0 2790 7 1 2 2004 83922
0 2791 5 1 1 2790
0 2792 7 2 2 79047 74449
0 2793 5 1 1 83924
0 2794 7 1 2 74273 2793
0 2795 5 1 1 2794
0 2796 7 1 2 67888 2795
0 2797 7 1 2 2791 2796
0 2798 5 1 1 2797
0 2799 7 2 2 74485 81389
0 2800 5 1 1 83926
0 2801 7 5 2 68570 76272
0 2802 5 2 1 83928
0 2803 7 1 2 83929 78546
0 2804 7 1 2 83927 2803
0 2805 5 1 1 2804
0 2806 7 1 2 2798 2805
0 2807 5 1 1 2806
0 2808 7 1 2 70340 2807
0 2809 5 1 1 2808
0 2810 7 10 2 67513 76178
0 2811 5 5 1 83935
0 2812 7 8 2 71555 67034
0 2813 7 1 2 68926 83950
0 2814 7 2 2 83936 2813
0 2815 7 1 2 76350 83958
0 2816 5 1 1 2815
0 2817 7 1 2 79081 83822
0 2818 7 1 2 83714 2817
0 2819 5 1 1 2818
0 2820 7 1 2 2816 2819
0 2821 5 1 1 2820
0 2822 7 1 2 67889 2821
0 2823 5 1 1 2822
0 2824 7 1 2 2809 2823
0 2825 5 1 1 2824
0 2826 7 1 2 70076 2825
0 2827 5 1 1 2826
0 2828 7 20 2 64568 70341
0 2829 5 2 1 83960
0 2830 7 1 2 83961 82185
0 2831 5 2 1 2830
0 2832 7 20 2 72522 68571
0 2833 7 2 2 76443 83984
0 2834 5 2 1 84004
0 2835 7 1 2 83982 84006
0 2836 5 2 1 2835
0 2837 7 1 2 75205 84008
0 2838 5 1 1 2837
0 2839 7 3 2 82402 82130
0 2840 7 1 2 75706 76833
0 2841 7 1 2 84010 2840
0 2842 5 1 1 2841
0 2843 7 1 2 2838 2842
0 2844 5 1 1 2843
0 2845 7 1 2 71556 2844
0 2846 5 1 1 2845
0 2847 7 8 2 71993 67514
0 2848 7 3 2 66444 67035
0 2849 7 2 2 84013 84021
0 2850 7 2 2 76404 77817
0 2851 7 1 2 73653 84026
0 2852 7 1 2 84024 2851
0 2853 5 1 1 2852
0 2854 7 1 2 2846 2853
0 2855 5 1 1 2854
0 2856 7 1 2 75544 2855
0 2857 5 1 1 2856
0 2858 7 1 2 2827 2857
0 2859 5 1 1 2858
0 2860 7 1 2 71734 2859
0 2861 5 1 1 2860
0 2862 7 1 2 75485 75206
0 2863 5 1 1 2862
0 2864 7 1 2 74507 78547
0 2865 5 1 1 2864
0 2866 7 1 2 2863 2865
0 2867 5 1 1 2866
0 2868 7 1 2 84005 2867
0 2869 5 1 1 2868
0 2870 7 3 2 71994 80289
0 2871 5 1 1 84028
0 2872 7 1 2 84029 83959
0 2873 5 1 1 2872
0 2874 7 1 2 2869 2873
0 2875 5 1 1 2874
0 2876 7 1 2 75545 2875
0 2877 5 1 1 2876
0 2878 7 1 2 2861 2877
0 2879 5 1 1 2878
0 2880 7 1 2 70598 2879
0 2881 5 1 1 2880
0 2882 7 2 2 68927 75859
0 2883 7 1 2 81409 83841
0 2884 5 1 1 2883
0 2885 7 8 2 70077 73654
0 2886 5 1 1 84033
0 2887 7 2 2 80477 84034
0 2888 5 1 1 84041
0 2889 7 1 2 71557 84042
0 2890 5 1 1 2889
0 2891 7 1 2 2884 2890
0 2892 5 1 1 2891
0 2893 7 4 2 71259 66926
0 2894 7 2 2 84043 77742
0 2895 7 2 2 2892 84047
0 2896 7 1 2 84031 84049
0 2897 5 1 1 2896
0 2898 7 1 2 2881 2897
0 2899 5 1 1 2898
0 2900 7 1 2 68754 2899
0 2901 5 1 1 2900
0 2902 7 9 2 63728 69720
0 2903 7 17 2 68928 70599
0 2904 7 1 2 84051 84060
0 2905 7 1 2 84050 2904
0 2906 5 1 1 2905
0 2907 7 1 2 2901 2906
0 2908 5 1 1 2907
0 2909 7 1 2 65892 2908
0 2910 5 1 1 2909
0 2911 7 10 2 66134 71735
0 2912 7 4 2 64569 84077
0 2913 5 2 1 84087
0 2914 7 3 2 67515 82098
0 2915 7 1 2 84088 84093
0 2916 5 1 1 2915
0 2917 7 12 2 72523 76444
0 2918 5 2 1 84096
0 2919 7 4 2 71736 82099
0 2920 5 5 1 84110
0 2921 7 1 2 76695 84114
0 2922 5 5 1 2921
0 2923 7 1 2 84097 84119
0 2924 5 1 1 2923
0 2925 7 1 2 2916 2924
0 2926 5 1 1 2925
0 2927 7 16 2 70342 66445
0 2928 5 1 1 84124
0 2929 7 5 2 70078 84125
0 2930 7 5 2 68929 77743
0 2931 7 1 2 84140 84145
0 2932 7 1 2 83196 2931
0 2933 7 1 2 2926 2932
0 2934 5 1 1 2933
0 2935 7 1 2 2910 2934
0 2936 5 1 1 2935
0 2937 7 1 2 69379 2936
0 2938 5 1 1 2937
0 2939 7 6 2 68755 83615
0 2940 7 11 2 71260 71737
0 2941 7 2 2 84156 77763
0 2942 7 2 2 84150 84167
0 2943 7 8 2 70079 65893
0 2944 7 11 2 67516 68572
0 2945 5 1 1 84179
0 2946 7 2 2 84171 84180
0 2947 5 1 1 84190
0 2948 7 5 2 70600 67036
0 2949 7 1 2 69721 81428
0 2950 7 1 2 84192 2949
0 2951 7 1 2 84191 2950
0 2952 7 1 2 84169 2951
0 2953 5 1 1 2952
0 2954 7 1 2 2938 2953
0 2955 7 1 2 2787 2954
0 2956 7 1 2 2663 2955
0 2957 5 1 1 2956
0 2958 7 1 2 82781 2957
0 2959 5 1 1 2958
0 2960 7 1 2 70080 77592
0 2961 5 1 1 2960
0 2962 7 2 2 69722 77628
0 2963 5 4 1 84197
0 2964 7 9 2 71261 73892
0 2965 5 1 1 84203
0 2966 7 1 2 84199 2965
0 2967 5 7 1 2966
0 2968 7 1 2 70964 84212
0 2969 5 1 1 2968
0 2970 7 1 2 2961 2969
0 2971 5 1 1 2970
0 2972 7 1 2 69380 2971
0 2973 5 1 1 2972
0 2974 7 3 2 77800 80827
0 2975 5 1 1 84219
0 2976 7 1 2 75844 84220
0 2977 5 1 1 2976
0 2978 7 1 2 2973 2977
0 2979 5 2 1 2978
0 2980 7 2 2 75813 84222
0 2981 7 4 2 65716 66824
0 2982 7 8 2 63850 64020
0 2983 7 2 2 84226 84230
0 2984 7 1 2 84224 84238
0 2985 5 1 1 2984
0 2986 7 1 2 633 2985
0 2987 5 1 1 2986
0 2988 7 1 2 72524 2987
0 2989 5 1 1 2988
0 2990 7 7 2 72899 74590
0 2991 5 16 1 84240
0 2992 7 4 2 84241 81390
0 2993 5 1 1 84263
0 2994 7 3 2 76366 84231
0 2995 7 4 2 71262 72094
0 2996 7 3 2 69723 74052
0 2997 7 1 2 84270 84274
0 2998 7 1 2 84267 2997
0 2999 7 1 2 84264 2998
0 3000 5 1 1 2999
0 3001 7 1 2 2989 3000
0 3002 5 1 1 3001
0 3003 7 1 2 65282 3002
0 3004 5 1 1 3003
0 3005 7 31 2 67517 67890
0 3006 5 2 1 84277
0 3007 7 2 2 67037 84278
0 3008 7 2 2 74082 84310
0 3009 7 19 2 68930 64021
0 3010 7 2 2 71263 75715
0 3011 7 1 2 84314 84333
0 3012 7 1 2 84312 3011
0 3013 5 1 1 3012
0 3014 7 10 2 65283 70763
0 3015 5 1 1 84335
0 3016 7 3 2 64950 84336
0 3017 7 1 2 75661 84345
0 3018 7 14 2 69096 64570
0 3019 7 5 2 74141 84348
0 3020 5 1 1 84362
0 3021 7 7 2 71995 72525
0 3022 7 11 2 72095 72900
0 3023 7 2 2 84367 84374
0 3024 7 1 2 84363 84385
0 3025 7 1 2 3017 3024
0 3026 5 1 1 3025
0 3027 7 1 2 3013 3026
0 3028 5 1 1 3027
0 3029 7 1 2 64266 3028
0 3030 5 1 1 3029
0 3031 7 4 2 70965 75896
0 3032 5 2 1 84387
0 3033 7 3 2 65894 74935
0 3034 5 1 1 84393
0 3035 7 2 2 84391 3034
0 3036 5 4 1 84396
0 3037 7 11 2 64571 70966
0 3038 5 1 1 84402
0 3039 7 1 2 74990 84403
0 3040 5 2 1 3039
0 3041 7 1 2 84397 84413
0 3042 5 1 1 3041
0 3043 7 2 2 69381 3042
0 3044 5 1 1 84415
0 3045 7 9 2 66927 67518
0 3046 7 5 2 64022 82409
0 3047 7 1 2 84417 84426
0 3048 7 1 2 77634 3047
0 3049 7 1 2 84416 3048
0 3050 5 1 1 3049
0 3051 7 1 2 3030 3050
0 3052 5 1 1 3051
0 3053 7 1 2 73937 3052
0 3054 5 1 1 3053
0 3055 7 1 2 78737 79296
0 3056 5 3 1 3055
0 3057 7 1 2 83656 84431
0 3058 5 1 1 3057
0 3059 7 5 2 67519 74094
0 3060 7 7 2 65717 84315
0 3061 7 4 2 70343 71891
0 3062 7 1 2 80111 84446
0 3063 7 1 2 84439 3062
0 3064 7 1 2 84434 3063
0 3065 7 1 2 3058 3064
0 3066 5 1 1 3065
0 3067 7 1 2 3054 3066
0 3068 7 1 2 3004 3067
0 3069 5 1 1 3068
0 3070 7 1 2 74021 3069
0 3071 5 1 1 3070
0 3072 7 16 2 64267 64572
0 3073 5 1 1 84450
0 3074 7 2 2 74349 84451
0 3075 7 2 2 81188 84466
0 3076 7 5 2 65567 70764
0 3077 7 1 2 84470 74159
0 3078 7 1 2 84468 3077
0 3079 5 1 1 3078
0 3080 7 2 2 84247 83385
0 3081 7 18 2 71264 71892
0 3082 7 2 2 76951 84477
0 3083 7 6 2 64023 74053
0 3084 5 1 1 84497
0 3085 7 3 2 68756 76878
0 3086 7 1 2 84498 84503
0 3087 7 1 2 84495 3086
0 3088 7 1 2 84475 3087
0 3089 5 1 1 3088
0 3090 7 1 2 3079 3089
0 3091 5 1 1 3090
0 3092 7 1 2 72526 3091
0 3093 5 1 1 3092
0 3094 7 7 2 64951 71893
0 3095 7 1 2 70601 79021
0 3096 7 1 2 84506 3095
0 3097 7 6 2 67520 74723
0 3098 7 3 2 65718 76930
0 3099 7 12 2 64024 64268
0 3100 7 3 2 68757 84522
0 3101 7 1 2 84519 84534
0 3102 7 1 2 84513 3101
0 3103 7 1 2 3096 3102
0 3104 5 1 1 3103
0 3105 7 1 2 3093 3104
0 3106 5 1 1 3105
0 3107 7 1 2 76761 3106
0 3108 5 1 1 3107
0 3109 7 1 2 3071 3108
0 3110 5 1 1 3109
0 3111 7 1 2 80386 3110
0 3112 5 1 1 3111
0 3113 7 1 2 81367 78773
0 3114 5 24 1 3113
0 3115 7 5 2 67038 74022
0 3116 7 1 2 74086 84561
0 3117 7 1 2 78505 3116
0 3118 5 1 1 3117
0 3119 7 13 2 63729 64952
0 3120 7 3 2 84566 79082
0 3121 7 9 2 66825 67521
0 3122 7 13 2 66628 72096
0 3123 7 1 2 74924 84591
0 3124 7 1 2 84582 3123
0 3125 7 1 2 84579 3124
0 3126 5 1 1 3125
0 3127 7 1 2 3118 3126
0 3128 5 1 1 3127
0 3129 7 1 2 71265 3128
0 3130 5 1 1 3129
0 3131 7 2 2 65568 66135
0 3132 7 7 2 66826 82753
0 3133 7 2 2 84604 84606
0 3134 7 10 2 72097 67522
0 3135 7 1 2 77399 84615
0 3136 7 1 2 84613 3135
0 3137 5 1 1 3136
0 3138 7 1 2 3130 3137
0 3139 5 1 1 3138
0 3140 7 1 2 70344 3139
0 3141 5 1 1 3140
0 3142 7 5 2 69724 75500
0 3143 7 2 2 84625 75778
0 3144 5 1 1 84630
0 3145 7 2 2 66136 77400
0 3146 5 1 1 84632
0 3147 7 1 2 3144 3146
0 3148 5 1 1 3147
0 3149 7 3 2 67523 77766
0 3150 7 15 2 63851 71738
0 3151 7 1 2 79624 84637
0 3152 7 1 2 84634 3151
0 3153 7 1 2 3148 3152
0 3154 5 1 1 3153
0 3155 7 1 2 3141 3154
0 3156 5 1 1 3155
0 3157 7 1 2 66928 3156
0 3158 5 1 1 3157
0 3159 7 2 2 81491 81543
0 3160 5 38 1 84652
0 3161 7 4 2 67039 84654
0 3162 7 4 2 69725 76701
0 3163 7 17 2 71266 66629
0 3164 5 2 1 84700
0 3165 7 1 2 84701 74295
0 3166 7 1 2 79128 3165
0 3167 7 1 2 84696 3166
0 3168 7 1 2 84692 3167
0 3169 5 1 1 3168
0 3170 7 1 2 3158 3169
0 3171 5 1 1 3170
0 3172 7 1 2 64025 3171
0 3173 5 1 1 3172
0 3174 7 3 2 81258 78425
0 3175 5 2 1 84719
0 3176 7 4 2 76445 78371
0 3177 5 1 1 84724
0 3178 7 3 2 72527 84725
0 3179 5 1 1 84728
0 3180 7 1 2 84722 3179
0 3181 5 3 1 3180
0 3182 7 15 2 66630 68573
0 3183 5 5 1 84734
0 3184 7 1 2 84749 83427
0 3185 5 6 1 3184
0 3186 7 4 2 65284 84754
0 3187 5 1 1 84760
0 3188 7 5 2 70345 82881
0 3189 5 4 1 84764
0 3190 7 1 2 3187 84769
0 3191 5 7 1 3190
0 3192 7 3 2 84567 77892
0 3193 7 3 2 84780 74261
0 3194 7 1 2 84773 84783
0 3195 7 1 2 84731 3194
0 3196 5 1 1 3195
0 3197 7 1 2 3173 3196
0 3198 5 1 1 3197
0 3199 7 1 2 65719 3198
0 3200 5 1 1 3199
0 3201 7 9 2 70346 66631
0 3202 5 4 1 84786
0 3203 7 6 2 1470 84795
0 3204 5 90 1 84799
0 3205 7 27 2 73655 84805
0 3206 5 4 1 84895
0 3207 7 2 2 64026 84732
0 3208 5 1 1 84926
0 3209 7 18 2 64269 72528
0 3210 5 2 1 84928
0 3211 7 1 2 84929 77849
0 3212 5 1 1 3211
0 3213 7 1 2 3208 3212
0 3214 5 2 1 3213
0 3215 7 1 2 84896 84948
0 3216 5 1 1 3215
0 3217 7 6 2 68574 74417
0 3218 5 1 1 84950
0 3219 7 2 2 72529 84951
0 3220 7 11 2 65895 66632
0 3221 7 12 2 65285 66137
0 3222 5 2 1 84969
0 3223 7 4 2 84958 84970
0 3224 7 1 2 84452 84983
0 3225 7 1 2 84956 3224
0 3226 5 1 1 3225
0 3227 7 1 2 3216 3226
0 3228 5 1 1 3227
0 3229 7 1 2 84784 3228
0 3230 5 1 1 3229
0 3231 7 1 2 3200 3230
0 3232 5 1 1 3231
0 3233 7 1 2 84537 3232
0 3234 5 1 1 3233
0 3235 7 55 2 72530 67891
0 3236 5 1 1 84987
0 3237 7 5 2 71267 84988
0 3238 5 7 1 85042
0 3239 7 4 2 79619 78145
0 3240 5 2 1 85054
0 3241 7 1 2 85047 85058
0 3242 5 5 1 3241
0 3243 7 1 2 70967 85060
0 3244 5 1 1 3243
0 3245 7 1 2 79462 84279
0 3246 5 6 1 3245
0 3247 7 1 2 3244 85065
0 3248 5 2 1 3247
0 3249 7 1 2 69382 85071
0 3250 5 1 1 3249
0 3251 7 17 2 71268 67524
0 3252 7 5 2 67892 85073
0 3253 7 1 2 85090 78372
0 3254 5 2 1 3253
0 3255 7 1 2 3250 85095
0 3256 5 1 1 3255
0 3257 7 14 2 68758 71894
0 3258 7 70 2 66929 85097
0 3259 7 3 2 74371 85111
0 3260 7 2 2 67040 82946
0 3261 7 3 2 65569 75997
0 3262 7 1 2 85184 85186
0 3263 5 1 1 3262
0 3264 7 1 2 63852 79759
0 3265 7 4 2 70602 71739
0 3266 7 1 2 74213 85189
0 3267 7 1 2 3264 3266
0 3268 5 1 1 3267
0 3269 7 1 2 3263 3268
0 3270 5 1 1 3269
0 3271 7 1 2 85181 3270
0 3272 5 1 1 3271
0 3273 7 160 2 63730 66930
0 3274 5 13 1 85193
0 3275 7 1 2 85194 83002
0 3276 7 5 2 67041 76795
0 3277 7 1 2 84440 85366
0 3278 7 1 2 3275 3277
0 3279 5 1 1 3278
0 3280 7 1 2 3272 3279
0 3281 5 1 1 3280
0 3282 7 1 2 3256 3281
0 3283 5 1 1 3282
0 3284 7 4 2 63731 77893
0 3285 7 5 2 71740 80208
0 3286 7 4 2 67525 76144
0 3287 7 2 2 74054 85380
0 3288 7 1 2 85375 85384
0 3289 5 1 1 3288
0 3290 7 4 2 69097 75897
0 3291 5 1 1 85386
0 3292 7 3 2 77983 83718
0 3293 7 2 2 85387 85390
0 3294 5 1 1 85393
0 3295 7 1 2 65286 85394
0 3296 5 1 1 3295
0 3297 7 1 2 3289 3296
0 3298 5 1 1 3297
0 3299 7 1 2 76762 3298
0 3300 5 1 1 3299
0 3301 7 3 2 74372 77401
0 3302 5 1 1 85395
0 3303 7 2 2 81817 85396
0 3304 7 1 2 84280 85398
0 3305 5 1 1 3304
0 3306 7 1 2 3294 3305
0 3307 5 1 1 3306
0 3308 7 1 2 75207 3307
0 3309 5 1 1 3308
0 3310 7 1 2 3300 3309
0 3311 5 1 1 3310
0 3312 7 1 2 64573 3311
0 3313 5 1 1 3312
0 3314 7 1 2 75208 82257
0 3315 5 1 1 3314
0 3316 7 7 2 68931 70968
0 3317 7 2 2 79159 85400
0 3318 5 1 1 85407
0 3319 7 1 2 80569 85408
0 3320 5 1 1 3319
0 3321 7 1 2 3315 3320
0 3322 5 1 1 3321
0 3323 7 5 2 67526 76066
0 3324 5 1 1 85409
0 3325 7 1 2 74373 85410
0 3326 7 1 2 3322 3325
0 3327 5 1 1 3326
0 3328 7 1 2 3313 3327
0 3329 5 1 1 3328
0 3330 7 1 2 64953 3329
0 3331 5 1 1 3330
0 3332 7 8 2 64027 64574
0 3333 7 3 2 68932 85414
0 3334 7 5 2 66138 71996
0 3335 7 1 2 71741 85425
0 3336 7 1 2 85422 3335
0 3337 7 1 2 84313 3336
0 3338 5 1 1 3337
0 3339 7 1 2 3331 3338
0 3340 5 1 1 3339
0 3341 7 1 2 85371 3340
0 3342 5 1 1 3341
0 3343 7 1 2 3283 3342
0 3344 5 1 1 3343
0 3345 7 1 2 73938 3344
0 3346 5 1 1 3345
0 3347 7 1 2 3234 3346
0 3348 7 1 2 3112 3347
0 3349 7 1 2 2959 3348
0 3350 7 1 2 2215 3349
0 3351 7 1 2 1403 3350
0 3352 5 1 1 3351
0 3353 7 1 2 73835 3352
0 3354 5 1 1 3353
0 3355 7 16 2 69098 65720
0 3356 5 1 1 85430
0 3357 7 28 2 64028 70765
0 3358 5 1 1 85446
0 3359 7 6 2 3356 3358
0 3360 5 87 1 85474
0 3361 7 9 2 70603 75716
0 3362 7 1 2 82882 79194
0 3363 5 10 1 3362
0 3364 7 3 2 67893 78587
0 3365 5 2 1 85586
0 3366 7 1 2 80570 85589
0 3367 5 1 1 3366
0 3368 7 1 2 85576 3367
0 3369 5 1 1 3368
0 3370 7 1 2 74591 3369
0 3371 5 1 1 3370
0 3372 7 4 2 65287 80334
0 3373 5 5 1 85591
0 3374 7 1 2 72901 85592
0 3375 5 1 1 3374
0 3376 7 2 2 3371 3375
0 3377 7 2 2 66633 79713
0 3378 5 2 1 85602
0 3379 7 1 2 75247 83575
0 3380 5 1 1 3379
0 3381 7 2 2 85604 3380
0 3382 5 1 1 85606
0 3383 7 1 2 70347 3382
0 3384 5 1 1 3383
0 3385 7 1 2 85600 3384
0 3386 5 1 1 3385
0 3387 7 1 2 66139 3386
0 3388 5 1 1 3387
0 3389 7 11 2 73349 80669
0 3390 5 26 1 85608
0 3391 7 14 2 68282 81818
0 3392 5 60 1 85645
0 3393 7 4 2 85659 74592
0 3394 5 2 1 85719
0 3395 7 2 2 85619 85720
0 3396 5 2 1 85725
0 3397 7 1 2 76984 85726
0 3398 5 1 1 3397
0 3399 7 2 2 3388 3398
0 3400 5 1 1 85729
0 3401 7 1 2 85567 3400
0 3402 5 1 1 3401
0 3403 7 22 2 73350 81674
0 3404 5 5 1 85731
0 3405 7 1 2 85732 76145
0 3406 5 4 1 3405
0 3407 7 7 2 70348 72902
0 3408 5 3 1 85762
0 3409 7 3 2 74869 85763
0 3410 5 1 1 85772
0 3411 7 1 2 71742 85773
0 3412 5 1 1 3411
0 3413 7 1 2 85758 3412
0 3414 5 3 1 3413
0 3415 7 1 2 85568 85775
0 3416 5 1 1 3415
0 3417 7 3 2 85660 76367
0 3418 7 1 2 65570 85778
0 3419 5 2 1 3418
0 3420 7 1 2 3416 85781
0 3421 5 2 1 3420
0 3422 7 1 2 79498 85783
0 3423 5 1 1 3422
0 3424 7 6 2 65571 76368
0 3425 5 3 1 85785
0 3426 7 2 2 71269 85646
0 3427 5 2 1 85794
0 3428 7 1 2 72903 85796
0 3429 5 1 1 3428
0 3430 7 1 2 74508 3429
0 3431 5 1 1 3430
0 3432 7 3 2 71270 82643
0 3433 5 2 1 85798
0 3434 7 1 2 67894 85799
0 3435 5 1 1 3434
0 3436 7 2 2 3431 3435
0 3437 7 1 2 85786 85803
0 3438 5 1 1 3437
0 3439 7 1 2 3423 3438
0 3440 7 1 2 3402 3439
0 3441 5 1 1 3440
0 3442 7 1 2 68759 3441
0 3443 5 1 1 3442
0 3444 7 1 2 74462 85804
0 3445 5 1 1 3444
0 3446 7 5 2 67895 82644
0 3447 5 4 1 85805
0 3448 7 1 2 85806 85723
0 3449 5 2 1 3448
0 3450 7 1 2 85814 82811
0 3451 5 1 1 3450
0 3452 7 1 2 85661 74463
0 3453 5 1 1 3452
0 3454 7 1 2 82833 3453
0 3455 5 2 1 3454
0 3456 7 1 2 79499 85816
0 3457 5 1 1 3456
0 3458 7 1 2 3451 3457
0 3459 7 1 2 3445 3458
0 3460 5 1 1 3459
0 3461 7 1 2 78155 3460
0 3462 5 1 1 3461
0 3463 7 1 2 3443 3462
0 3464 5 1 1 3463
0 3465 7 1 2 64575 3464
0 3466 5 1 1 3465
0 3467 7 7 2 72904 76670
0 3468 7 1 2 85818 85569
0 3469 5 1 1 3468
0 3470 7 7 2 71997 73351
0 3471 7 1 2 85825 77894
0 3472 5 1 1 3471
0 3473 7 1 2 3469 3472
0 3474 5 1 1 3473
0 3475 7 1 2 81675 3474
0 3476 5 1 1 3475
0 3477 7 4 2 66931 78563
0 3478 7 1 2 84447 85190
0 3479 7 1 2 85832 3478
0 3480 5 1 1 3479
0 3481 7 1 2 85791 3480
0 3482 5 1 1 3481
0 3483 7 1 2 72905 3482
0 3484 5 1 1 3483
0 3485 7 1 2 3476 3484
0 3486 5 1 1 3485
0 3487 7 1 2 68760 3486
0 3488 5 1 1 3487
0 3489 7 3 2 70604 74205
0 3490 5 1 1 85836
0 3491 7 1 2 82834 2277
0 3492 5 1 1 3491
0 3493 7 1 2 81819 2384
0 3494 5 1 1 3493
0 3495 7 2 2 3492 3494
0 3496 5 1 1 85839
0 3497 7 1 2 3490 3496
0 3498 5 1 1 3497
0 3499 7 1 2 78156 3498
0 3500 5 1 1 3499
0 3501 7 1 2 3488 3500
0 3502 5 1 1 3501
0 3503 7 1 2 66140 3502
0 3504 5 1 1 3503
0 3505 7 8 2 66827 72906
0 3506 7 1 2 63732 85840
0 3507 5 1 1 3506
0 3508 7 121 2 68761 71998
0 3509 5 1 1 85849
0 3510 7 1 2 65572 85850
0 3511 7 1 2 82629 3510
0 3512 5 1 1 3511
0 3513 7 1 2 3507 3512
0 3514 5 1 1 3513
0 3515 7 1 2 85841 3514
0 3516 5 1 1 3515
0 3517 7 1 2 3504 3516
0 3518 5 1 1 3517
0 3519 7 1 2 74593 3518
0 3520 5 1 1 3519
0 3521 7 1 2 74991 85817
0 3522 5 1 1 3521
0 3523 7 3 2 81676 82812
0 3524 5 1 1 85970
0 3525 7 1 2 73352 85971
0 3526 5 1 1 3525
0 3527 7 1 2 3522 3526
0 3528 5 1 1 3527
0 3529 7 1 2 78157 3528
0 3530 5 1 1 3529
0 3531 7 1 2 66141 85784
0 3532 5 1 1 3531
0 3533 7 2 2 66634 84478
0 3534 7 1 2 76879 85833
0 3535 7 1 2 85973 3534
0 3536 5 1 1 3535
0 3537 7 1 2 85782 3536
0 3538 5 1 1 3537
0 3539 7 1 2 72907 3538
0 3540 5 1 1 3539
0 3541 7 1 2 3532 3540
0 3542 5 1 1 3541
0 3543 7 1 2 68762 3542
0 3544 5 1 1 3543
0 3545 7 1 2 3530 3544
0 3546 5 1 1 3545
0 3547 7 1 2 75248 3546
0 3548 5 1 1 3547
0 3549 7 8 2 66932 79625
0 3550 5 1 1 85975
0 3551 7 8 2 71999 74023
0 3552 7 2 2 85662 85983
0 3553 5 1 1 85991
0 3554 7 1 2 3550 3553
0 3555 5 1 1 3554
0 3556 7 1 2 75898 3555
0 3557 5 1 1 3556
0 3558 7 3 2 65288 74992
0 3559 5 2 1 85993
0 3560 7 10 2 73353 85195
0 3561 5 1 1 85998
0 3562 7 4 2 65573 66635
0 3563 7 1 2 85999 86008
0 3564 7 1 2 85994 3563
0 3565 5 1 1 3564
0 3566 7 1 2 3557 3565
0 3567 5 1 1 3566
0 3568 7 1 2 66828 3567
0 3569 5 1 1 3568
0 3570 7 1 2 3548 3569
0 3571 7 1 2 3520 3570
0 3572 7 1 2 3466 3571
0 3573 5 1 1 3572
0 3574 7 1 2 65896 3573
0 3575 5 1 1 3574
0 3576 7 1 2 67527 3575
0 3577 5 1 1 3576
0 3578 7 1 2 81820 85787
0 3579 5 1 1 3578
0 3580 7 2 2 75324 84806
0 3581 7 1 2 85570 86012
0 3582 5 1 1 3581
0 3583 7 1 2 3579 3582
0 3584 5 1 1 3583
0 3585 7 1 2 68575 3584
0 3586 5 1 1 3585
0 3587 7 2 2 70081 76880
0 3588 7 2 2 71558 75717
0 3589 7 1 2 86014 86016
0 3590 5 1 1 3589
0 3591 7 1 2 80571 85788
0 3592 5 1 1 3591
0 3593 7 1 2 3590 3592
0 3594 7 1 2 3586 3593
0 3595 5 1 1 3594
0 3596 7 1 2 68763 3595
0 3597 5 1 1 3596
0 3598 7 2 2 70349 82947
0 3599 5 9 1 86018
0 3600 7 9 2 80387 86020
0 3601 5 42 1 86029
0 3602 7 3 2 76369 74004
0 3603 5 1 1 86080
0 3604 7 1 2 86038 86081
0 3605 5 1 1 3604
0 3606 7 1 2 3597 3605
0 3607 5 1 1 3606
0 3608 7 1 2 68283 3607
0 3609 5 1 1 3608
0 3610 7 3 2 66933 79817
0 3611 7 7 2 70082 70605
0 3612 7 1 2 86083 86086
0 3613 7 5 2 71743 71895
0 3614 7 5 2 68764 86093
0 3615 7 5 2 71559 75116
0 3616 7 1 2 86098 86103
0 3617 7 1 2 3612 3616
0 3618 5 1 1 3617
0 3619 7 1 2 3609 3618
0 3620 5 1 1 3619
0 3621 7 1 2 83238 3620
0 3622 5 1 1 3621
0 3623 7 4 2 71271 85663
0 3624 5 3 1 86108
0 3625 7 5 2 76446 74509
0 3626 5 2 1 86115
0 3627 7 2 2 64576 85664
0 3628 5 3 1 86122
0 3629 7 1 2 86120 86124
0 3630 5 1 1 3629
0 3631 7 1 2 86112 3630
0 3632 5 1 1 3631
0 3633 7 1 2 85984 3632
0 3634 5 1 1 3633
0 3635 7 1 2 81677 77959
0 3636 5 2 1 3635
0 3637 7 1 2 85976 86127
0 3638 5 1 1 3637
0 3639 7 1 2 3634 3638
0 3640 5 1 1 3639
0 3641 7 1 2 66829 3640
0 3642 5 1 1 3641
0 3643 7 14 2 66446 71744
0 3644 5 3 1 86129
0 3645 7 4 2 86130 79760
0 3646 5 2 1 86146
0 3647 7 2 2 86150 85727
0 3648 5 3 1 86152
0 3649 7 1 2 73656 86154
0 3650 5 2 1 3649
0 3651 7 4 2 71745 79832
0 3652 7 1 2 80478 86159
0 3653 5 1 1 3652
0 3654 7 2 2 86157 3653
0 3655 5 1 1 86163
0 3656 7 1 2 71272 86164
0 3657 5 1 1 3656
0 3658 7 2 2 66934 79129
0 3659 7 4 2 71560 74895
0 3660 5 1 1 86167
0 3661 7 4 2 69726 71746
0 3662 5 4 1 86171
0 3663 7 1 2 86019 86175
0 3664 5 1 1 3663
0 3665 7 2 2 85595 3664
0 3666 5 2 1 86179
0 3667 7 1 2 3660 86180
0 3668 5 1 1 3667
0 3669 7 1 2 80224 3668
0 3670 5 1 1 3669
0 3671 7 3 2 71747 74510
0 3672 5 2 1 86183
0 3673 7 3 2 80483 79708
0 3674 5 3 1 86188
0 3675 7 1 2 86184 86191
0 3676 5 1 1 3675
0 3677 7 1 2 66142 3676
0 3678 7 1 2 3670 3677
0 3679 5 1 1 3678
0 3680 7 1 2 86165 3679
0 3681 7 1 2 3657 3680
0 3682 5 1 1 3681
0 3683 7 1 2 3642 3682
0 3684 5 1 1 3683
0 3685 7 1 2 67896 3684
0 3686 5 1 1 3685
0 3687 7 8 2 71273 66830
0 3688 7 1 2 82645 86194
0 3689 7 1 2 85977 3688
0 3690 5 1 1 3689
0 3691 7 1 2 72531 3690
0 3692 7 1 2 3686 3691
0 3693 7 1 2 3622 3692
0 3694 5 1 1 3693
0 3695 7 1 2 65897 3694
0 3696 5 1 1 3695
0 3697 7 3 2 76370 74024
0 3698 7 21 2 66636 72908
0 3699 5 6 1 86205
0 3700 7 2 2 70969 86206
0 3701 5 2 1 86232
0 3702 7 4 2 66143 82339
0 3703 5 1 1 86236
0 3704 7 1 2 76146 86237
0 3705 5 1 1 3704
0 3706 7 1 2 86234 3705
0 3707 5 1 1 3706
0 3708 7 1 2 65289 3707
0 3709 5 1 1 3708
0 3710 7 1 2 75697 82560
0 3711 5 1 1 3710
0 3712 7 2 2 82883 75055
0 3713 7 1 2 81429 86240
0 3714 5 1 1 3713
0 3715 7 1 2 3711 3714
0 3716 7 1 2 3709 3715
0 3717 5 1 1 3716
0 3718 7 1 2 64577 3717
0 3719 5 1 1 3718
0 3720 7 5 2 72909 85665
0 3721 5 1 1 86242
0 3722 7 1 2 76868 86243
0 3723 5 1 1 3722
0 3724 7 1 2 3719 3723
0 3725 5 1 1 3724
0 3726 7 1 2 86202 3725
0 3727 5 1 1 3726
0 3728 7 12 2 64954 78611
0 3729 5 21 1 86247
0 3730 7 1 2 80572 86248
0 3731 5 2 1 3730
0 3732 7 1 2 86158 86280
0 3733 5 1 1 3732
0 3734 7 1 2 72910 3733
0 3735 5 1 1 3734
0 3736 7 2 2 81678 77297
0 3737 5 3 1 86282
0 3738 7 1 2 74724 86283
0 3739 5 2 1 3738
0 3740 7 1 2 3735 86287
0 3741 5 2 1 3740
0 3742 7 1 2 76541 86289
0 3743 5 1 1 3742
0 3744 7 4 2 73657 76179
0 3745 5 1 1 86291
0 3746 7 3 2 65290 83390
0 3747 5 8 1 86295
0 3748 7 4 2 70350 86131
0 3749 5 2 1 86306
0 3750 7 1 2 86298 86310
0 3751 5 1 1 3750
0 3752 7 1 2 64955 3751
0 3753 5 2 1 3752
0 3754 7 2 2 81679 79219
0 3755 5 2 1 86314
0 3756 7 1 2 86312 86316
0 3757 5 1 1 3756
0 3758 7 1 2 86292 3757
0 3759 5 1 1 3758
0 3760 7 6 2 64578 71748
0 3761 7 6 2 79062 86318
0 3762 5 2 1 86324
0 3763 7 25 2 64956 73658
0 3764 5 16 1 86332
0 3765 7 3 2 67897 86357
0 3766 5 1 1 86373
0 3767 7 1 2 80957 86374
0 3768 5 1 1 3767
0 3769 7 1 2 86325 3768
0 3770 5 1 1 3769
0 3771 7 6 2 64957 81680
0 3772 7 3 2 75779 77861
0 3773 5 1 1 86382
0 3774 7 1 2 86376 86383
0 3775 5 1 1 3774
0 3776 7 1 2 3770 3775
0 3777 5 1 1 3776
0 3778 7 1 2 73354 3777
0 3779 5 1 1 3778
0 3780 7 1 2 3759 3779
0 3781 7 1 2 3743 3780
0 3782 5 2 1 3781
0 3783 7 5 2 70970 66935
0 3784 7 1 2 86387 79130
0 3785 7 1 2 86385 3784
0 3786 5 1 1 3785
0 3787 7 1 2 3727 3786
0 3788 7 1 2 3696 3787
0 3789 5 1 1 3788
0 3790 7 1 2 3577 3789
0 3791 5 1 1 3790
0 3792 7 20 2 66637 71896
0 3793 7 10 2 66447 66936
0 3794 7 6 2 86392 86412
0 3795 7 5 2 76985 81391
0 3796 7 2 2 86422 86428
0 3797 7 1 2 76895 78333
0 3798 7 1 2 86433 3797
0 3799 5 1 1 3798
0 3800 7 1 2 3791 3799
0 3801 5 1 1 3800
0 3802 7 1 2 75872 3801
0 3803 5 1 1 3802
0 3804 7 3 2 85733 77862
0 3805 7 2 2 78793 86435
0 3806 5 2 1 86438
0 3807 7 5 2 73355 81821
0 3808 5 5 1 86442
0 3809 7 1 2 86447 86299
0 3810 5 2 1 3809
0 3811 7 1 2 74594 86452
0 3812 5 2 1 3811
0 3813 7 5 2 64958 81822
0 3814 5 3 1 86456
0 3815 7 3 2 66448 86457
0 3816 5 2 1 86464
0 3817 7 1 2 86454 86467
0 3818 5 2 1 3817
0 3819 7 1 2 72911 86469
0 3820 5 2 1 3819
0 3821 7 7 2 66638 81580
0 3822 5 1 1 86473
0 3823 7 2 2 83117 86474
0 3824 5 1 1 86480
0 3825 7 1 2 73659 86481
0 3826 5 2 1 3825
0 3827 7 1 2 86471 86482
0 3828 5 2 1 3827
0 3829 7 1 2 64579 86484
0 3830 5 1 1 3829
0 3831 7 1 2 86440 3830
0 3832 5 1 1 3831
0 3833 7 1 2 83197 3832
0 3834 5 1 1 3833
0 3835 7 8 2 68765 64580
0 3836 7 2 2 86486 84807
0 3837 7 15 2 64959 70606
0 3838 7 1 2 75522 86496
0 3839 7 1 2 85819 3838
0 3840 7 1 2 86494 3839
0 3841 5 1 1 3840
0 3842 7 1 2 3834 3841
0 3843 5 1 1 3842
0 3844 7 1 2 78399 3843
0 3845 5 1 1 3844
0 3846 7 2 2 83539 80462
0 3847 5 3 1 86511
0 3848 7 2 2 80239 82034
0 3849 5 1 1 86516
0 3850 7 1 2 82884 84248
0 3851 7 1 2 3849 3850
0 3852 5 1 1 3851
0 3853 7 1 2 86513 3852
0 3854 5 1 1 3853
0 3855 7 1 2 82813 3854
0 3856 5 1 1 3855
0 3857 7 3 2 76351 79714
0 3858 7 4 2 70607 71561
0 3859 7 10 2 70083 66639
0 3860 5 1 1 86525
0 3861 7 1 2 86521 86526
0 3862 7 1 2 86518 3861
0 3863 5 1 1 3862
0 3864 7 1 2 3856 3863
0 3865 5 1 1 3864
0 3866 7 1 2 69727 3865
0 3867 5 1 1 3866
0 3868 7 1 2 75036 82814
0 3869 5 1 1 3868
0 3870 7 15 2 64960 66640
0 3871 5 2 1 86535
0 3872 7 2 2 79220 74464
0 3873 5 1 1 86552
0 3874 7 1 2 86536 86553
0 3875 5 1 1 3874
0 3876 7 1 2 3869 3875
0 3877 5 1 1 3876
0 3878 7 1 2 68576 3877
0 3879 5 1 1 3878
0 3880 7 6 2 66641 66937
0 3881 7 2 2 74925 86554
0 3882 7 1 2 75325 86560
0 3883 5 1 1 3882
0 3884 7 1 2 3879 3883
0 3885 5 1 1 3884
0 3886 7 1 2 67898 3885
0 3887 5 1 1 3886
0 3888 7 1 2 86512 82815
0 3889 5 1 1 3888
0 3890 7 11 2 66938 73660
0 3891 7 3 2 65574 86562
0 3892 5 2 1 86573
0 3893 7 1 2 79833 81315
0 3894 5 1 1 3893
0 3895 7 1 2 86574 3894
0 3896 5 1 1 3895
0 3897 7 3 2 72000 74837
0 3898 7 1 2 76637 75863
0 3899 7 1 2 86578 3898
0 3900 5 1 1 3899
0 3901 7 1 2 3896 3900
0 3902 5 1 1 3901
0 3903 7 1 2 66642 3902
0 3904 5 1 1 3903
0 3905 7 1 2 3889 3904
0 3906 7 1 2 3887 3905
0 3907 5 1 1 3906
0 3908 7 1 2 71274 3907
0 3909 5 1 1 3908
0 3910 7 1 2 3867 3909
0 3911 5 1 1 3910
0 3912 7 1 2 65291 3911
0 3913 5 1 1 3912
0 3914 7 3 2 70084 76273
0 3915 5 2 1 86581
0 3916 7 4 2 72912 82816
0 3917 7 1 2 86582 86586
0 3918 5 1 1 3917
0 3919 7 3 2 79568 86333
0 3920 5 1 1 86590
0 3921 7 1 2 86591 83084
0 3922 5 1 1 3921
0 3923 7 1 2 3918 3922
0 3924 5 1 1 3923
0 3925 7 1 2 81823 3924
0 3926 5 1 1 3925
0 3927 7 4 2 71749 83889
0 3928 7 6 2 66449 79761
0 3929 7 1 2 86593 86597
0 3930 5 1 1 3929
0 3931 7 1 2 83239 86104
0 3932 5 1 1 3931
0 3933 7 1 2 3930 3932
0 3934 5 1 1 3933
0 3935 7 1 2 82817 3934
0 3936 5 1 1 3935
0 3937 7 1 2 3926 3936
0 3938 5 1 1 3937
0 3939 7 1 2 68284 3938
0 3940 5 1 1 3939
0 3941 7 14 2 70351 65575
0 3942 7 2 2 66939 86603
0 3943 7 2 2 70085 82712
0 3944 5 3 1 86619
0 3945 7 2 2 74870 86621
0 3946 5 1 1 86624
0 3947 7 1 2 67899 3946
0 3948 5 1 1 3947
0 3949 7 2 2 71275 84249
0 3950 7 1 2 3948 86626
0 3951 5 1 1 3950
0 3952 7 1 2 83354 3951
0 3953 5 1 1 3952
0 3954 7 1 2 86617 3953
0 3955 5 1 1 3954
0 3956 7 1 2 3940 3955
0 3957 7 1 2 3913 3956
0 3958 5 1 1 3957
0 3959 7 1 2 68766 3958
0 3960 5 1 1 3959
0 3961 7 1 2 74770 86105
0 3962 5 2 1 3961
0 3963 7 2 2 72913 85647
0 3964 5 4 1 86630
0 3965 7 2 2 66643 76671
0 3966 5 4 1 86636
0 3967 7 2 2 83442 86638
0 3968 5 1 1 86642
0 3969 7 1 2 65292 86643
0 3970 5 1 1 3969
0 3971 7 1 2 71562 1756
0 3972 7 1 2 3970 3971
0 3973 5 1 1 3972
0 3974 7 1 2 86632 3973
0 3975 5 1 1 3974
0 3976 7 1 2 70086 3975
0 3977 5 1 1 3976
0 3978 7 1 2 86628 3977
0 3979 5 1 1 3978
0 3980 7 1 2 76274 3979
0 3981 5 1 1 3980
0 3982 7 2 2 73661 75326
0 3983 5 2 1 86644
0 3984 7 9 2 69728 66644
0 3985 7 1 2 76405 86648
0 3986 7 1 2 86645 3985
0 3987 5 1 1 3986
0 3988 7 2 2 3981 3987
0 3989 7 1 2 82885 79864
0 3990 5 2 1 3989
0 3991 7 3 2 68577 75037
0 3992 7 1 2 71276 86661
0 3993 5 1 1 3992
0 3994 7 1 2 86659 3993
0 3995 5 1 1 3994
0 3996 7 1 2 65293 3995
0 3997 5 1 1 3996
0 3998 7 21 2 68578 80573
0 3999 5 4 1 86664
0 4000 7 1 2 86665 83091
0 4001 5 3 1 4000
0 4002 7 11 2 70352 71277
0 4003 7 1 2 86692 86625
0 4004 5 1 1 4003
0 4005 7 1 2 86689 4004
0 4006 7 1 2 3997 4005
0 4007 5 1 1 4006
0 4008 7 1 2 67900 4007
0 4009 5 1 1 4008
0 4010 7 1 2 86657 4009
0 4011 5 1 1 4010
0 4012 7 1 2 83104 4011
0 4013 5 1 1 4012
0 4014 7 1 2 3960 4013
0 4015 5 1 1 4014
0 4016 7 1 2 72532 4015
0 4017 5 1 1 4016
0 4018 7 3 2 64581 82035
0 4019 5 1 1 86703
0 4020 7 1 2 4019 83365
0 4021 5 1 1 4020
0 4022 7 1 2 81392 4021
0 4023 5 1 1 4022
0 4024 7 5 2 67528 74595
0 4025 7 1 2 75597 86706
0 4026 5 2 1 4025
0 4027 7 4 2 67901 81958
0 4028 5 2 1 86713
0 4029 7 1 2 74596 86714
0 4030 5 1 1 4029
0 4031 7 1 2 86711 4030
0 4032 7 1 2 4023 4031
0 4033 5 1 1 4032
0 4034 7 1 2 83198 4033
0 4035 5 1 1 4034
0 4036 7 4 2 64961 82131
0 4037 5 1 1 86719
0 4038 7 1 2 78981 75523
0 4039 7 1 2 85820 4038
0 4040 7 1 2 86720 4039
0 4041 5 1 1 4040
0 4042 7 1 2 4035 4041
0 4043 5 1 1 4042
0 4044 7 1 2 84808 4043
0 4045 5 1 1 4044
0 4046 7 5 2 82586 76147
0 4047 5 6 1 86723
0 4048 7 1 2 79744 86728
0 4049 5 2 1 4048
0 4050 7 1 2 65294 86734
0 4051 5 1 1 4050
0 4052 7 1 2 3410 4051
0 4053 5 1 1 4052
0 4054 7 1 2 64582 4053
0 4055 5 1 1 4054
0 4056 7 2 2 82587 75780
0 4057 5 4 1 86736
0 4058 7 2 2 72914 86737
0 4059 5 1 1 86742
0 4060 7 1 2 65295 86743
0 4061 5 1 1 4060
0 4062 7 1 2 4055 4061
0 4063 5 1 1 4062
0 4064 7 1 2 74597 4063
0 4065 5 1 1 4064
0 4066 7 1 2 81172 83710
0 4067 5 1 1 4066
0 4068 7 1 2 72915 83962
0 4069 5 1 1 4068
0 4070 7 3 2 70353 78564
0 4071 5 1 1 86744
0 4072 7 6 2 65296 78588
0 4073 5 3 1 86747
0 4074 7 1 2 4071 86753
0 4075 5 1 1 4074
0 4076 7 3 2 68285 83003
0 4077 5 2 1 86756
0 4078 7 1 2 82730 86759
0 4079 7 1 2 4075 4078
0 4080 5 1 1 4079
0 4081 7 1 2 4069 4080
0 4082 5 1 1 4081
0 4083 7 1 2 75249 4082
0 4084 5 1 1 4083
0 4085 7 1 2 4067 4084
0 4086 7 1 2 4065 4085
0 4087 5 1 1 4086
0 4088 7 1 2 67529 83199
0 4089 7 1 2 4087 4088
0 4090 5 1 1 4089
0 4091 7 1 2 4045 4090
0 4092 7 1 2 4017 4091
0 4093 5 1 1 4092
0 4094 7 1 2 65898 4093
0 4095 5 1 1 4094
0 4096 7 1 2 3845 4095
0 4097 5 1 1 4096
0 4098 7 1 2 71897 4097
0 4099 5 1 1 4098
0 4100 7 11 2 65297 82886
0 4101 5 10 1 86761
0 4102 7 5 2 67902 86772
0 4103 5 8 1 86782
0 4104 7 1 2 64583 86787
0 4105 5 4 1 4104
0 4106 7 2 2 72916 86762
0 4107 5 1 1 86799
0 4108 7 1 2 86795 4107
0 4109 5 2 1 4108
0 4110 7 1 2 75038 86801
0 4111 5 1 1 4110
0 4112 7 5 2 66450 78565
0 4113 5 6 1 86803
0 4114 7 1 2 83773 83825
0 4115 5 3 1 4114
0 4116 7 2 2 86808 86814
0 4117 5 2 1 86817
0 4118 7 1 2 82731 86819
0 4119 5 1 1 4118
0 4120 7 4 2 78612 86377
0 4121 5 6 1 86821
0 4122 7 1 2 75616 86825
0 4123 5 1 1 4122
0 4124 7 1 2 73662 4123
0 4125 5 1 1 4124
0 4126 7 1 2 4119 4125
0 4127 7 1 2 4111 4126
0 4128 5 1 1 4127
0 4129 7 1 2 67530 4128
0 4130 5 1 1 4129
0 4131 7 8 2 72533 80574
0 4132 7 7 2 69729 74511
0 4133 5 5 1 86839
0 4134 7 2 2 67903 86846
0 4135 5 1 1 86851
0 4136 7 2 2 4135 83250
0 4137 5 1 1 86853
0 4138 7 1 2 345 74751
0 4139 7 1 2 86854 4138
0 4140 5 1 1 4139
0 4141 7 1 2 86831 4140
0 4142 5 1 1 4141
0 4143 7 1 2 4130 4142
0 4144 5 1 1 4143
0 4145 7 5 2 72001 74309
0 4146 7 2 2 79626 86855
0 4147 7 1 2 4144 86860
0 4148 5 1 1 4147
0 4149 7 2 2 84800 83690
0 4150 5 6 1 86862
0 4151 7 1 2 80484 86863
0 4152 5 1 1 4151
0 4153 7 1 2 82732 4152
0 4154 5 1 1 4153
0 4155 7 1 2 85759 4154
0 4156 5 1 1 4155
0 4157 7 1 2 74598 4156
0 4158 5 1 1 4157
0 4159 7 1 2 83009 79343
0 4160 5 3 1 4159
0 4161 7 3 2 73356 86870
0 4162 5 1 1 86873
0 4163 7 2 2 66645 83054
0 4164 5 1 1 86876
0 4165 7 1 2 83165 86877
0 4166 5 1 1 4165
0 4167 7 2 2 4162 4166
0 4168 7 1 2 83980 86878
0 4169 5 1 1 4168
0 4170 7 1 2 82036 4169
0 4171 5 1 1 4170
0 4172 7 1 2 75327 86773
0 4173 5 2 1 4172
0 4174 7 1 2 72917 81589
0 4175 7 1 2 86880 4174
0 4176 5 1 1 4175
0 4177 7 4 2 73357 86864
0 4178 5 2 1 86882
0 4179 7 2 2 72918 82948
0 4180 5 3 1 86888
0 4181 7 10 2 66646 67904
0 4182 5 2 1 86893
0 4183 7 3 2 75094 86894
0 4184 5 3 1 86905
0 4185 7 1 2 86890 86908
0 4186 7 1 2 86886 4185
0 4187 5 1 1 4186
0 4188 7 1 2 64584 4187
0 4189 5 2 1 4188
0 4190 7 1 2 4176 86911
0 4191 7 1 2 4171 4190
0 4192 7 1 2 4158 4191
0 4193 5 1 1 4192
0 4194 7 1 2 65899 4193
0 4195 5 1 1 4194
0 4196 7 3 2 82588 76986
0 4197 5 2 1 86913
0 4198 7 1 2 76702 77947
0 4199 7 1 2 86914 4198
0 4200 5 1 1 4199
0 4201 7 1 2 4195 4200
0 4202 5 1 1 4201
0 4203 7 1 2 83200 4202
0 4204 5 1 1 4203
0 4205 7 1 2 84115 86639
0 4206 5 4 1 4205
0 4207 7 2 2 70354 86918
0 4208 5 3 1 86922
0 4209 7 3 2 86924 83572
0 4210 5 1 1 86927
0 4211 7 3 2 71750 76672
0 4212 5 5 1 86930
0 4213 7 2 2 70087 78589
0 4214 5 7 1 86938
0 4215 7 1 2 71563 78590
0 4216 5 5 1 4215
0 4217 7 3 2 86940 86947
0 4218 5 1 1 86952
0 4219 7 2 2 74871 86953
0 4220 5 1 1 86955
0 4221 7 1 2 74599 86956
0 4222 5 3 1 4221
0 4223 7 2 2 66647 86957
0 4224 5 1 1 86960
0 4225 7 1 2 86933 4224
0 4226 5 2 1 4225
0 4227 7 1 2 65298 86962
0 4228 5 1 1 4227
0 4229 7 1 2 86928 4228
0 4230 5 2 1 4229
0 4231 7 1 2 72919 86964
0 4232 5 1 1 4231
0 4233 7 3 2 82589 75642
0 4234 5 7 1 86966
0 4235 7 13 2 68286 84809
0 4236 5 1 1 86976
0 4237 7 5 2 73663 86977
0 4238 5 5 1 86989
0 4239 7 2 2 67905 85666
0 4240 5 2 1 86999
0 4241 7 1 2 86994 87001
0 4242 5 1 1 4241
0 4243 7 1 2 66451 4242
0 4244 5 1 1 4243
0 4245 7 1 2 86969 4244
0 4246 5 1 1 4245
0 4247 7 1 2 64962 4246
0 4248 5 1 1 4247
0 4249 7 3 2 66648 74725
0 4250 7 1 2 81581 87003
0 4251 5 1 1 4250
0 4252 7 1 2 4248 4251
0 4253 7 1 2 4232 4252
0 4254 5 1 1 4253
0 4255 7 1 2 64585 4254
0 4256 5 1 1 4255
0 4257 7 13 2 64963 72920
0 4258 5 3 1 87006
0 4259 7 2 2 87007 79221
0 4260 5 1 1 87022
0 4261 7 1 2 84897 87023
0 4262 5 1 1 4261
0 4263 7 1 2 4256 4262
0 4264 5 1 1 4263
0 4265 7 1 2 65900 83879
0 4266 7 1 2 4264 4265
0 4267 5 1 1 4266
0 4268 7 1 2 4204 4267
0 4269 5 1 1 4268
0 4270 7 1 2 71898 4269
0 4271 5 1 1 4270
0 4272 7 1 2 69730 86783
0 4273 5 1 1 4272
0 4274 7 1 2 75039 4273
0 4275 5 1 1 4274
0 4276 7 5 2 67906 78681
0 4277 5 14 1 87024
0 4278 7 1 2 73664 87029
0 4279 5 1 1 4278
0 4280 7 2 2 86815 4279
0 4281 7 1 2 64586 83917
0 4282 5 1 1 4281
0 4283 7 1 2 87043 4282
0 4284 7 1 2 4275 4283
0 4285 5 1 1 4284
0 4286 7 1 2 86861 4285
0 4287 5 1 1 4286
0 4288 7 1 2 67531 4287
0 4289 7 1 2 4271 4288
0 4290 5 1 1 4289
0 4291 7 10 2 65901 67907
0 4292 5 3 1 87045
0 4293 7 1 2 86186 2225
0 4294 5 6 1 4293
0 4295 7 1 2 64587 87058
0 4296 5 2 1 4295
0 4297 7 8 2 70088 81681
0 4298 5 3 1 87066
0 4299 7 1 2 77081 87067
0 4300 5 2 1 4299
0 4301 7 1 2 87064 87077
0 4302 5 2 1 4301
0 4303 7 1 2 87046 87079
0 4304 5 1 1 4303
0 4305 7 7 2 66452 80112
0 4306 7 2 2 71751 76987
0 4307 5 2 1 87088
0 4308 7 1 2 64588 84735
0 4309 5 1 1 4308
0 4310 7 1 2 87090 4309
0 4311 5 1 1 4310
0 4312 7 1 2 65299 4311
0 4313 5 1 1 4312
0 4314 7 3 2 64589 81824
0 4315 5 4 1 87092
0 4316 7 1 2 72921 84787
0 4317 5 1 1 4316
0 4318 7 1 2 87095 4317
0 4319 5 1 1 4318
0 4320 7 1 2 73665 4319
0 4321 5 1 1 4320
0 4322 7 1 2 4313 4321
0 4323 5 1 1 4322
0 4324 7 1 2 87081 4323
0 4325 5 1 1 4324
0 4326 7 1 2 4304 4325
0 4327 5 1 1 4326
0 4328 7 1 2 68287 4327
0 4329 5 1 1 4328
0 4330 7 1 2 82395 83611
0 4331 5 1 1 4330
0 4332 7 1 2 4329 4331
0 4333 5 1 1 4332
0 4334 7 1 2 79131 4333
0 4335 5 1 1 4334
0 4336 7 10 2 71752 66831
0 4337 7 4 2 63733 87099
0 4338 7 1 2 77650 86604
0 4339 7 1 2 87109 4338
0 4340 5 1 1 4339
0 4341 7 2 2 66649 74838
0 4342 5 2 1 87113
0 4343 7 1 2 87114 75643
0 4344 7 1 2 79525 4343
0 4345 5 1 1 4344
0 4346 7 1 2 4340 4345
0 4347 5 1 1 4346
0 4348 7 1 2 69731 4347
0 4349 5 1 1 4348
0 4350 7 1 2 64590 82561
0 4351 5 2 1 4350
0 4352 7 17 2 70355 65902
0 4353 7 3 2 87119 83596
0 4354 5 1 1 87136
0 4355 7 1 2 87117 4354
0 4356 5 1 1 4355
0 4357 7 1 2 78852 4356
0 4358 5 1 1 4357
0 4359 7 1 2 4349 4358
0 4360 7 1 2 4335 4359
0 4361 5 1 1 4360
0 4362 7 1 2 72002 4361
0 4363 5 1 1 4362
0 4364 7 1 2 66453 82362
0 4365 5 2 1 4364
0 4366 7 3 2 87139 82614
0 4367 5 1 1 87141
0 4368 7 1 2 86358 87142
0 4369 5 1 1 4368
0 4370 7 1 2 64591 4369
0 4371 5 1 1 4370
0 4372 7 1 2 77704 4371
0 4373 5 1 1 4372
0 4374 7 1 2 70356 4373
0 4375 5 1 1 4374
0 4376 7 1 2 81825 77596
0 4377 5 2 1 4376
0 4378 7 3 2 67908 77290
0 4379 5 4 1 87146
0 4380 7 1 2 81682 77685
0 4381 7 1 2 87149 4380
0 4382 5 1 1 4381
0 4383 7 1 2 87144 4382
0 4384 5 1 1 4383
0 4385 7 1 2 64964 4384
0 4386 5 3 1 4385
0 4387 7 4 2 66454 83435
0 4388 5 1 1 87156
0 4389 7 1 2 72922 87157
0 4390 5 1 1 4389
0 4391 7 1 2 87153 4390
0 4392 7 1 2 4375 4391
0 4393 5 1 1 4392
0 4394 7 1 2 70971 4393
0 4395 5 1 1 4394
0 4396 7 3 2 75546 82376
0 4397 5 1 1 87160
0 4398 7 1 2 82290 76703
0 4399 5 1 1 4398
0 4400 7 1 2 4397 4399
0 4401 5 1 1 4400
0 4402 7 1 2 82949 4401
0 4403 5 1 1 4402
0 4404 7 7 2 71753 87120
0 4405 7 1 2 87163 76750
0 4406 5 3 1 4405
0 4407 7 3 2 83037 86233
0 4408 5 1 1 87173
0 4409 7 1 2 75845 87121
0 4410 5 1 1 4409
0 4411 7 1 2 4408 4410
0 4412 5 1 1 4411
0 4413 7 1 2 70089 4412
0 4414 5 1 1 4413
0 4415 7 1 2 87170 4414
0 4416 7 1 2 4403 4415
0 4417 7 1 2 4395 4416
0 4418 5 1 1 4417
0 4419 7 1 2 75718 74025
0 4420 7 1 2 4418 4419
0 4421 5 1 1 4420
0 4422 7 1 2 72534 4421
0 4423 7 1 2 4363 4422
0 4424 5 1 1 4423
0 4425 7 1 2 66144 4424
0 4426 7 1 2 4290 4425
0 4427 5 1 1 4426
0 4428 7 1 2 4148 4427
0 4429 7 1 2 4099 4428
0 4430 5 1 1 4429
0 4431 7 1 2 74450 4430
0 4432 5 1 1 4431
0 4433 7 1 2 3803 4432
0 4434 5 1 1 4433
0 4435 7 1 2 64270 4434
0 4436 5 1 1 4435
0 4437 7 1 2 2103 86455
0 4438 5 1 1 4437
0 4439 7 1 2 72923 4438
0 4440 5 1 1 4439
0 4441 7 4 2 80920 83826
0 4442 7 1 2 70357 87176
0 4443 5 1 1 4442
0 4444 7 1 2 84796 83010
0 4445 5 16 1 4444
0 4446 7 1 2 73939 87180
0 4447 5 2 1 4446
0 4448 7 1 2 87196 85577
0 4449 7 1 2 4443 4448
0 4450 5 1 1 4449
0 4451 7 1 2 66145 4450
0 4452 5 1 1 4451
0 4453 7 1 2 4440 4452
0 4454 5 1 1 4453
0 4455 7 1 2 64592 4454
0 4456 5 1 1 4455
0 4457 7 12 2 86584 77928
0 4458 5 3 1 87198
0 4459 7 5 2 72924 81826
0 4460 5 2 1 87213
0 4461 7 1 2 87218 86909
0 4462 5 1 1 4461
0 4463 7 1 2 87199 4462
0 4464 5 1 1 4463
0 4465 7 1 2 81683 83558
0 4466 5 3 1 4465
0 4467 7 16 2 73358 74600
0 4468 5 14 1 87223
0 4469 7 1 2 81827 87224
0 4470 5 1 1 4469
0 4471 7 1 2 87220 4470
0 4472 5 1 1 4471
0 4473 7 1 2 66146 4472
0 4474 5 1 1 4473
0 4475 7 8 2 66650 78613
0 4476 7 1 2 64965 76406
0 4477 7 2 2 87253 4476
0 4478 5 2 1 87261
0 4479 7 1 2 4474 87263
0 4480 5 1 1 4479
0 4481 7 1 2 72925 4480
0 4482 5 1 1 4481
0 4483 7 1 2 4464 4482
0 4484 7 1 2 4456 4483
0 4485 5 1 1 4484
0 4486 7 1 2 65903 4485
0 4487 5 1 1 4486
0 4488 7 1 2 81298 87174
0 4489 5 1 1 4488
0 4490 7 1 2 4487 4489
0 4491 5 1 1 4490
0 4492 7 5 2 68933 84562
0 4493 7 1 2 4491 87265
0 4494 5 1 1 4493
0 4495 7 4 2 68767 72098
0 4496 7 3 2 87270 75152
0 4497 7 1 2 79500 85776
0 4498 5 1 1 4497
0 4499 7 1 2 85730 4498
0 4500 5 1 1 4499
0 4501 7 1 2 64593 4500
0 4502 5 1 1 4501
0 4503 7 5 2 65300 86537
0 4504 5 13 1 87277
0 4505 7 3 2 76988 79297
0 4506 5 1 1 87295
0 4507 7 1 2 87278 87296
0 4508 5 1 1 4507
0 4509 7 1 2 66147 86290
0 4510 5 1 1 4509
0 4511 7 1 2 4508 4510
0 4512 7 1 2 4502 4511
0 4513 5 2 1 4512
0 4514 7 1 2 65904 87298
0 4515 5 1 1 4514
0 4516 7 4 2 66651 76989
0 4517 5 2 1 87300
0 4518 7 3 2 78614 87301
0 4519 5 1 1 87306
0 4520 7 6 2 64966 76704
0 4521 7 1 2 76180 87309
0 4522 7 1 2 87307 4521
0 4523 5 1 1 4522
0 4524 7 1 2 4515 4523
0 4525 5 1 1 4524
0 4526 7 1 2 87274 4525
0 4527 5 1 1 4526
0 4528 7 1 2 4494 4527
0 4529 5 1 1 4528
0 4530 7 1 2 66940 4529
0 4531 5 1 1 4530
0 4532 7 6 2 64967 84898
0 4533 5 1 1 87315
0 4534 7 2 2 87316 79222
0 4535 5 1 1 87321
0 4536 7 1 2 78816 87322
0 4537 5 2 1 4536
0 4538 7 1 2 72926 83019
0 4539 5 1 1 4538
0 4540 7 2 2 86334 79223
0 4541 5 1 1 87325
0 4542 7 1 2 4539 4541
0 4543 5 1 1 4542
0 4544 7 1 2 81828 4543
0 4545 5 1 1 4544
0 4546 7 17 2 71564 66652
0 4547 5 2 1 87327
0 4548 7 4 2 87328 74896
0 4549 5 5 1 87346
0 4550 7 1 2 83453 86300
0 4551 5 11 1 4550
0 4552 7 1 2 75328 87355
0 4553 5 1 1 4552
0 4554 7 1 2 87350 4553
0 4555 5 2 1 4554
0 4556 7 1 2 72927 87366
0 4557 5 1 1 4556
0 4558 7 2 2 78615 83118
0 4559 5 2 1 87368
0 4560 7 15 2 67909 74601
0 4561 5 2 1 87372
0 4562 7 1 2 74872 87373
0 4563 5 1 1 4562
0 4564 7 4 2 64968 79224
0 4565 7 2 2 68579 87389
0 4566 5 1 1 87393
0 4567 7 1 2 4563 4566
0 4568 5 1 1 4567
0 4569 7 1 2 81684 4568
0 4570 5 1 1 4569
0 4571 7 1 2 87370 4570
0 4572 7 1 2 4557 4571
0 4573 7 1 2 4545 4572
0 4574 5 1 1 4573
0 4575 7 1 2 76181 4574
0 4576 5 1 1 4575
0 4577 7 1 2 87323 4576
0 4578 5 1 1 4577
0 4579 7 30 2 68768 68934
0 4580 7 6 2 70608 87395
0 4581 7 2 2 65905 76834
0 4582 7 1 2 87425 87431
0 4583 7 1 2 4578 4582
0 4584 5 1 1 4583
0 4585 7 1 2 71899 4584
0 4586 7 1 2 4531 4585
0 4587 5 1 1 4586
0 4588 7 1 2 65906 85992
0 4589 5 1 1 4588
0 4590 7 10 2 64969 65576
0 4591 7 2 2 79593 87433
0 4592 7 1 2 66941 87254
0 4593 7 1 2 87443 4592
0 4594 5 1 1 4593
0 4595 7 1 2 4589 4594
0 4596 5 1 1 4595
0 4597 7 1 2 79950 4596
0 4598 5 1 1 4597
0 4599 7 2 2 71565 81829
0 4600 5 16 1 87445
0 4601 7 2 2 85667 87447
0 4602 5 2 1 87463
0 4603 7 13 2 73940 87464
0 4604 5 6 1 87467
0 4605 7 1 2 83778 82281
0 4606 7 1 2 87480 4605
0 4607 5 5 1 4606
0 4608 7 1 2 85978 87486
0 4609 5 1 1 4608
0 4610 7 1 2 65907 85985
0 4611 5 1 1 4610
0 4612 7 1 2 4609 4611
0 4613 5 1 1 4612
0 4614 7 1 2 77557 4613
0 4615 5 1 1 4614
0 4616 7 1 2 4598 4615
0 4617 5 1 1 4616
0 4618 7 1 2 75873 4617
0 4619 5 1 1 4618
0 4620 7 5 2 72003 78717
0 4621 7 1 2 87491 79387
0 4622 7 1 2 82534 4621
0 4623 5 1 1 4622
0 4624 7 1 2 66832 4623
0 4625 7 1 2 4619 4624
0 4626 5 1 1 4625
0 4627 7 1 2 69383 4626
0 4628 7 1 2 4587 4627
0 4629 5 1 1 4628
0 4630 7 2 2 80821 87432
0 4631 7 1 2 68935 87496
0 4632 5 1 1 4631
0 4633 7 2 2 73359 74305
0 4634 7 17 2 66455 66653
0 4635 5 1 1 87500
0 4636 7 2 2 80113 87501
0 4637 7 1 2 87498 87517
0 4638 5 1 1 4637
0 4639 7 1 2 4632 4638
0 4640 5 1 1 4639
0 4641 7 1 2 65301 4640
0 4642 5 1 1 4641
0 4643 7 3 2 87329 74839
0 4644 5 1 1 87519
0 4645 7 1 2 70090 82363
0 4646 7 1 2 83835 4645
0 4647 5 1 1 4646
0 4648 7 1 2 4644 4647
0 4649 5 1 1 4648
0 4650 7 2 2 67042 4649
0 4651 7 5 2 65908 72004
0 4652 7 1 2 87524 75707
0 4653 7 1 2 87522 4652
0 4654 5 1 1 4653
0 4655 7 1 2 4642 4654
0 4656 5 1 1 4655
0 4657 7 1 2 72928 4656
0 4658 5 1 1 4657
0 4659 7 1 2 81685 87030
0 4660 5 1 1 4659
0 4661 7 1 2 77603 4660
0 4662 5 2 1 4661
0 4663 7 2 2 64970 87529
0 4664 5 1 1 87531
0 4665 7 1 2 72929 87468
0 4666 5 1 1 4665
0 4667 7 2 2 4664 4666
0 4668 5 3 1 87533
0 4669 7 1 2 70972 74262
0 4670 5 1 1 4669
0 4671 7 1 2 3318 4670
0 4672 5 1 1 4671
0 4673 7 1 2 87535 4672
0 4674 5 1 1 4673
0 4675 7 4 2 67910 84810
0 4676 7 2 2 68580 87538
0 4677 5 1 1 87542
0 4678 7 9 2 72930 75329
0 4679 5 2 1 87544
0 4680 7 1 2 87545 83679
0 4681 5 2 1 4680
0 4682 7 1 2 4677 87555
0 4683 5 1 1 4682
0 4684 7 1 2 65909 4683
0 4685 5 1 1 4684
0 4686 7 2 2 70973 78616
0 4687 7 1 2 87532 87557
0 4688 5 1 1 4687
0 4689 7 1 2 4685 4688
0 4690 5 1 1 4689
0 4691 7 1 2 78548 4690
0 4692 5 1 1 4691
0 4693 7 1 2 4674 4692
0 4694 5 1 1 4693
0 4695 7 1 2 64594 4694
0 4696 5 1 1 4695
0 4697 7 1 2 4658 4696
0 4698 5 1 1 4697
0 4699 7 1 2 78853 4698
0 4700 5 1 1 4699
0 4701 7 2 2 75330 82950
0 4702 5 3 1 87559
0 4703 7 5 2 65302 80388
0 4704 5 6 1 87564
0 4705 7 2 2 87560 87569
0 4706 7 1 2 87575 76723
0 4707 5 1 1 4706
0 4708 7 2 2 68936 75529
0 4709 7 5 2 71754 75719
0 4710 7 1 2 84141 87579
0 4711 7 1 2 87577 4710
0 4712 5 1 1 4711
0 4713 7 1 2 4707 4712
0 4714 5 1 1 4713
0 4715 7 1 2 87047 4714
0 4716 5 1 1 4715
0 4717 7 2 2 75720 79310
0 4718 7 4 2 67043 84811
0 4719 7 2 2 73666 87586
0 4720 7 1 2 87584 87590
0 4721 5 1 1 4720
0 4722 7 1 2 87448 76724
0 4723 5 1 1 4722
0 4724 7 1 2 4721 4723
0 4725 5 1 1 4724
0 4726 7 1 2 64971 4725
0 4727 5 1 1 4726
0 4728 7 2 2 87502 78108
0 4729 7 1 2 77737 87592
0 4730 5 1 1 4729
0 4731 7 1 2 4727 4730
0 4732 5 1 1 4731
0 4733 7 1 2 82562 4732
0 4734 5 1 1 4733
0 4735 7 1 2 4716 4734
0 4736 5 1 1 4735
0 4737 7 1 2 73360 4736
0 4738 5 1 1 4737
0 4739 7 6 2 68937 70091
0 4740 7 3 2 70358 87594
0 4741 7 1 2 77838 81978
0 4742 7 1 2 87600 4741
0 4743 5 1 1 4742
0 4744 7 4 2 70974 72005
0 4745 7 3 2 75662 87603
0 4746 7 4 2 64972 72099
0 4747 7 1 2 83662 87610
0 4748 7 1 2 87607 4747
0 4749 5 1 1 4748
0 4750 7 1 2 4743 4749
0 4751 5 1 1 4750
0 4752 7 1 2 66456 4751
0 4753 5 1 1 4752
0 4754 7 4 2 77302 87239
0 4755 7 2 2 67911 87614
0 4756 5 1 1 87618
0 4757 7 3 2 63853 75814
0 4758 7 1 2 74323 87620
0 4759 7 1 2 87619 4758
0 4760 5 1 1 4759
0 4761 7 1 2 4753 4760
0 4762 5 1 1 4761
0 4763 7 1 2 66654 4762
0 4764 5 1 1 4763
0 4765 7 9 2 68288 82951
0 4766 5 12 1 87623
0 4767 7 11 2 87624 87570
0 4768 5 4 1 87644
0 4769 7 3 2 72931 87645
0 4770 5 1 1 87659
0 4771 7 12 2 70092 82377
0 4772 5 1 1 87662
0 4773 7 1 2 87663 76725
0 4774 7 1 2 87660 4773
0 4775 5 1 1 4774
0 4776 7 1 2 4764 4775
0 4777 7 1 2 4738 4776
0 4778 5 1 1 4777
0 4779 7 1 2 64595 74026
0 4780 7 1 2 4778 4779
0 4781 5 1 1 4780
0 4782 7 1 2 4700 4781
0 4783 5 1 1 4782
0 4784 7 1 2 66148 4783
0 4785 5 1 1 4784
0 4786 7 2 2 81686 87434
0 4787 7 2 2 63734 84404
0 4788 7 1 2 66833 77863
0 4789 7 1 2 87676 4788
0 4790 7 1 2 87674 4789
0 4791 7 1 2 87499 4790
0 4792 5 1 1 4791
0 4793 7 1 2 4785 4792
0 4794 7 1 2 4629 4793
0 4795 5 1 1 4794
0 4796 7 1 2 72535 4795
0 4797 5 1 1 4796
0 4798 7 1 2 72536 83307
0 4799 5 2 1 4798
0 4800 7 1 2 75250 85061
0 4801 5 2 1 4800
0 4802 7 1 2 87678 87680
0 4803 5 1 1 4802
0 4804 7 1 2 68289 4803
0 4805 5 1 1 4804
0 4806 7 1 2 87553 74760
0 4807 5 3 1 4806
0 4808 7 1 2 83937 87682
0 4809 5 1 1 4808
0 4810 7 1 2 4805 4809
0 4811 5 2 1 4810
0 4812 7 1 2 64271 87685
0 4813 5 1 1 4812
0 4814 7 1 2 75899 87390
0 4815 5 3 1 4814
0 4816 7 23 2 74602 80240
0 4817 7 2 2 87690 77686
0 4818 5 1 1 87713
0 4819 7 1 2 87554 4818
0 4820 5 2 1 4819
0 4821 7 1 2 66149 87715
0 4822 5 1 1 4821
0 4823 7 1 2 4260 4822
0 4824 5 1 1 4823
0 4825 7 1 2 64596 4824
0 4826 5 1 1 4825
0 4827 7 1 2 87687 4826
0 4828 5 1 1 4827
0 4829 7 1 2 81454 4828
0 4830 5 1 1 4829
0 4831 7 1 2 4813 4830
0 4832 5 2 1 4831
0 4833 7 40 2 68769 63854
0 4834 7 5 2 72100 87719
0 4835 7 3 2 85571 87759
0 4836 7 1 2 87717 87764
0 4837 5 1 1 4836
0 4838 7 3 2 68770 76912
0 4839 7 3 2 87767 74214
0 4840 5 1 1 87770
0 4841 7 4 2 69732 81959
0 4842 5 4 1 87773
0 4843 7 33 2 67532 72932
0 4844 5 4 1 87781
0 4845 7 1 2 87691 87782
0 4846 5 2 1 4845
0 4847 7 1 2 87777 87818
0 4848 5 1 1 4847
0 4849 7 1 2 64272 4848
0 4850 5 1 1 4849
0 4851 7 3 2 74512 84989
0 4852 5 3 1 87820
0 4853 7 1 2 81544 87823
0 4854 5 1 1 4853
0 4855 7 1 2 76182 4854
0 4856 5 1 1 4855
0 4857 7 3 2 72933 81455
0 4858 5 1 1 87826
0 4859 7 1 2 81545 4858
0 4860 5 1 1 4859
0 4861 7 6 2 87025 83779
0 4862 5 3 1 87829
0 4863 7 1 2 76542 87835
0 4864 7 1 2 4860 4863
0 4865 5 1 1 4864
0 4866 7 1 2 4856 4865
0 4867 7 1 2 4850 4866
0 4868 5 1 1 4867
0 4869 7 1 2 87771 4868
0 4870 5 1 1 4869
0 4871 7 2 2 73667 75174
0 4872 5 1 1 87838
0 4873 7 5 2 70093 75846
0 4874 5 2 1 87840
0 4875 7 1 2 64597 87841
0 4876 5 1 1 4875
0 4877 7 1 2 81247 4876
0 4878 5 2 1 4877
0 4879 7 1 2 87839 87847
0 4880 5 1 1 4879
0 4881 7 2 2 64273 78034
0 4882 5 2 1 87849
0 4883 7 1 2 82037 87850
0 4884 5 1 1 4883
0 4885 7 2 2 82733 4884
0 4886 7 2 2 67044 87853
0 4887 7 1 2 78069 87855
0 4888 5 1 1 4887
0 4889 7 1 2 4880 4888
0 4890 5 1 1 4889
0 4891 7 1 2 72537 4890
0 4892 5 1 1 4891
0 4893 7 1 2 78103 4872
0 4894 5 3 1 4893
0 4895 7 1 2 82721 83785
0 4896 5 3 1 4895
0 4897 7 1 2 87860 81517
0 4898 7 1 2 87857 4897
0 4899 5 1 1 4898
0 4900 7 1 2 4892 4899
0 4901 5 1 1 4900
0 4902 7 1 2 66150 4901
0 4903 5 1 1 4902
0 4904 7 1 2 79614 78087
0 4905 5 1 1 4904
0 4906 7 8 2 69733 70609
0 4907 7 3 2 87863 75874
0 4908 5 1 1 87871
0 4909 7 1 2 75781 87872
0 4910 5 1 1 4909
0 4911 7 1 2 4905 4910
0 4912 5 1 1 4911
0 4913 7 1 2 84930 4912
0 4914 5 1 1 4913
0 4915 7 2 2 87692 82734
0 4916 5 1 1 87874
0 4917 7 1 2 75617 4916
0 4918 5 2 1 4917
0 4919 7 1 2 81518 87876
0 4920 5 1 1 4919
0 4921 7 11 2 64598 72538
0 4922 7 2 2 81229 87878
0 4923 5 1 1 87889
0 4924 7 1 2 4920 4923
0 4925 5 2 1 4924
0 4926 7 1 2 87858 87891
0 4927 5 1 1 4926
0 4928 7 1 2 4914 4927
0 4929 7 1 2 4903 4928
0 4930 5 1 1 4929
0 4931 7 1 2 63735 4930
0 4932 5 1 1 4931
0 4933 7 1 2 4870 4932
0 4934 5 1 1 4933
0 4935 7 1 2 66834 4934
0 4936 5 1 1 4935
0 4937 7 1 2 74757 84655
0 4938 5 1 1 4937
0 4939 7 5 2 71566 72539
0 4940 5 1 1 87893
0 4941 7 4 2 72934 87894
0 4942 7 1 2 83179 87898
0 4943 5 2 1 4942
0 4944 7 1 2 4938 87902
0 4945 5 1 1 4944
0 4946 7 2 2 74279 4945
0 4947 7 9 2 68938 64599
0 4948 7 17 2 66151 71900
0 4949 7 3 2 87906 87915
0 4950 7 1 2 78982 87932
0 4951 7 1 2 87904 4950
0 4952 5 1 1 4951
0 4953 7 1 2 4936 4952
0 4954 5 1 1 4953
0 4955 7 1 2 72006 4954
0 4956 5 1 1 4955
0 4957 7 1 2 4837 4956
0 4958 5 1 1 4957
0 4959 7 1 2 65910 4958
0 4960 5 1 1 4959
0 4961 7 2 2 72935 79398
0 4962 7 2 2 66152 80930
0 4963 5 1 1 87937
0 4964 7 1 2 69384 4963
0 4965 5 2 1 4964
0 4966 7 1 2 87935 87939
0 4967 5 2 1 4966
0 4968 7 3 2 66835 74206
0 4969 7 2 2 74926 87943
0 4970 7 1 2 77624 87946
0 4971 5 1 1 4970
0 4972 7 2 2 79184 75721
0 4973 7 17 2 64274 70610
0 4974 7 2 2 66457 87950
0 4975 7 1 2 87948 87967
0 4976 5 1 1 4975
0 4977 7 1 2 4971 4976
0 4978 5 1 1 4977
0 4979 7 1 2 64973 4978
0 4980 5 1 1 4979
0 4981 7 1 2 79877 87947
0 4982 5 1 1 4981
0 4983 7 1 2 4980 4982
0 4984 5 1 1 4983
0 4985 7 1 2 68771 4984
0 4986 5 1 1 4985
0 4987 7 1 2 76990 86082
0 4988 7 1 2 87940 4987
0 4989 5 1 1 4988
0 4990 7 1 2 4986 4989
0 4991 5 1 1 4990
0 4992 7 1 2 75875 4991
0 4993 5 1 1 4992
0 4994 7 1 2 87941 4993
0 4995 5 1 1 4994
0 4996 7 1 2 64600 4995
0 4997 5 1 1 4996
0 4998 7 2 2 87720 86497
0 4999 7 4 2 71901 74230
0 5000 7 4 2 79225 87971
0 5001 7 2 2 87969 87975
0 5002 5 1 1 87979
0 5003 7 1 2 63736 87859
0 5004 5 1 1 5003
0 5005 7 1 2 4840 5004
0 5006 5 2 1 5005
0 5007 7 1 2 76371 87981
0 5008 5 1 1 5007
0 5009 7 1 2 5002 5008
0 5010 5 1 1 5009
0 5011 7 1 2 64275 75900
0 5012 7 1 2 5010 5011
0 5013 5 1 1 5012
0 5014 7 1 2 4997 5013
0 5015 5 1 1 5014
0 5016 7 1 2 78400 5015
0 5017 5 1 1 5016
0 5018 7 1 2 4960 5017
0 5019 5 1 1 5018
0 5020 7 1 2 80670 5019
0 5021 5 1 1 5020
0 5022 7 7 2 64276 64974
0 5023 5 3 1 87983
0 5024 7 1 2 87990 87266
0 5025 5 1 1 5024
0 5026 7 13 2 69385 64975
0 5027 7 2 2 87993 75876
0 5028 7 1 2 78983 88006
0 5029 5 1 1 5028
0 5030 7 1 2 5025 5029
0 5031 5 1 1 5030
0 5032 7 3 2 84971 82524
0 5033 7 1 2 88008 86434
0 5034 7 1 2 5031 5033
0 5035 5 1 1 5034
0 5036 7 1 2 5021 5035
0 5037 7 1 2 4797 5036
0 5038 7 1 2 4436 5037
0 5039 5 1 1 5038
0 5040 7 1 2 73836 5039
0 5041 5 1 1 5040
0 5042 7 27 2 70611 70651
0 5043 7 8 2 69041 88011
0 5044 7 10 2 70702 71902
0 5045 7 32 2 88038 88046
0 5046 7 195 2 63855 67045
0 5047 5 12 1 88088
0 5048 7 1 2 66153 86847
0 5049 5 2 1 5048
0 5050 7 4 2 76638 88295
0 5051 7 3 2 64277 68581
0 5052 7 1 2 88297 88301
0 5053 5 1 1 5052
0 5054 7 1 2 1580 5053
0 5055 5 1 1 5054
0 5056 7 1 2 66655 5055
0 5057 5 1 1 5056
0 5058 7 7 2 73668 76543
0 5059 5 3 1 88304
0 5060 7 1 2 86132 87994
0 5061 7 1 2 88305 5060
0 5062 5 1 1 5061
0 5063 7 1 2 5057 5062
0 5064 5 1 1 5063
0 5065 7 1 2 65303 5064
0 5066 5 1 1 5065
0 5067 7 3 2 76275 82952
0 5068 5 1 1 88314
0 5069 7 2 2 77929 5068
0 5070 7 1 2 70359 88317
0 5071 5 1 1 5070
0 5072 7 1 2 84091 5071
0 5073 5 1 1 5072
0 5074 7 1 2 64976 5073
0 5075 5 1 1 5074
0 5076 7 6 2 64601 77040
0 5077 5 1 1 88319
0 5078 7 1 2 81830 88320
0 5079 5 1 1 5078
0 5080 7 1 2 5075 5079
0 5081 5 1 1 5080
0 5082 7 1 2 69386 5081
0 5083 5 1 1 5082
0 5084 7 1 2 5066 5083
0 5085 5 1 1 5084
0 5086 7 1 2 72936 5085
0 5087 5 1 1 5086
0 5088 7 1 2 81266 83233
0 5089 5 2 1 5088
0 5090 7 1 2 75251 88325
0 5091 5 1 1 5090
0 5092 7 5 2 66154 76639
0 5093 7 1 2 81202 88327
0 5094 5 1 1 5093
0 5095 7 1 2 5091 5094
0 5096 5 1 1 5095
0 5097 7 1 2 81687 5096
0 5098 5 1 1 5097
0 5099 7 6 2 64602 75331
0 5100 5 2 1 88332
0 5101 7 5 2 66155 88333
0 5102 5 1 1 88340
0 5103 7 13 2 64278 70360
0 5104 5 2 1 88345
0 5105 7 3 2 83597 88346
0 5106 5 1 1 88360
0 5107 7 1 2 88341 88361
0 5108 5 1 1 5107
0 5109 7 1 2 5098 5108
0 5110 5 1 1 5109
0 5111 7 1 2 68582 5110
0 5112 5 1 1 5111
0 5113 7 1 2 3920 82020
0 5114 5 1 1 5113
0 5115 7 1 2 81203 5114
0 5116 5 1 1 5115
0 5117 7 1 2 77298 81259
0 5118 5 1 1 5117
0 5119 7 1 2 5116 5118
0 5120 5 1 1 5119
0 5121 7 1 2 81831 5120
0 5122 5 1 1 5121
0 5123 7 1 2 5112 5122
0 5124 7 1 2 5087 5123
0 5125 5 1 1 5124
0 5126 7 1 2 68290 5125
0 5127 5 1 1 5126
0 5128 7 11 2 73669 80671
0 5129 5 8 1 88363
0 5130 7 5 2 81832 88374
0 5131 5 25 1 88382
0 5132 7 3 2 74603 88387
0 5133 5 1 1 88412
0 5134 7 2 2 5133 75332
0 5135 5 4 1 88415
0 5136 7 2 2 67912 88417
0 5137 5 1 1 88421
0 5138 7 1 2 87546 86039
0 5139 5 2 1 5138
0 5140 7 1 2 5137 88423
0 5141 5 1 1 5140
0 5142 7 1 2 73361 5141
0 5143 5 1 1 5142
0 5144 7 1 2 82887 87374
0 5145 5 2 1 5144
0 5146 7 5 2 70094 80389
0 5147 7 1 2 74486 88427
0 5148 5 1 1 5147
0 5149 7 1 2 88425 5148
0 5150 5 1 1 5149
0 5151 7 1 2 65304 5150
0 5152 5 1 1 5151
0 5153 7 4 2 71567 82888
0 5154 5 2 1 88432
0 5155 7 1 2 83342 88433
0 5156 5 2 1 5155
0 5157 7 1 2 5152 88438
0 5158 7 1 2 5143 5157
0 5159 5 1 1 5158
0 5160 7 1 2 80010 5159
0 5161 5 1 1 5160
0 5162 7 1 2 74513 88347
0 5163 7 1 2 83612 5162
0 5164 5 1 1 5163
0 5165 7 1 2 5161 5164
0 5166 5 1 1 5165
0 5167 7 1 2 66156 5166
0 5168 5 1 1 5167
0 5169 7 1 2 5127 5168
0 5170 5 1 1 5169
0 5171 7 1 2 72540 5170
0 5172 5 1 1 5171
0 5173 7 2 2 67913 73941
0 5174 7 4 2 80921 88440
0 5175 5 3 1 88442
0 5176 7 5 2 87547 74825
0 5177 5 1 1 88449
0 5178 7 1 2 88446 5177
0 5179 5 1 1 5178
0 5180 7 1 2 66656 5179
0 5181 5 1 1 5180
0 5182 7 9 2 67914 78566
0 5183 7 2 2 74604 88454
0 5184 5 1 1 88463
0 5185 7 1 2 77303 86207
0 5186 5 1 1 5185
0 5187 7 1 2 83416 82038
0 5188 5 1 1 5187
0 5189 7 1 2 5186 5188
0 5190 5 1 1 5189
0 5191 7 1 2 68291 5190
0 5192 5 1 1 5191
0 5193 7 1 2 5184 5192
0 5194 7 1 2 5181 5193
0 5195 5 1 1 5194
0 5196 7 1 2 65305 5195
0 5197 5 1 1 5196
0 5198 7 1 2 72937 4210
0 5199 5 1 1 5198
0 5200 7 4 2 66657 76148
0 5201 5 1 1 88465
0 5202 7 1 2 78617 88466
0 5203 5 1 1 5202
0 5204 7 1 2 71568 82953
0 5205 5 6 1 5204
0 5206 7 1 2 74726 88469
0 5207 5 1 1 5206
0 5208 7 2 2 82889 79226
0 5209 5 2 1 88475
0 5210 7 1 2 70361 88476
0 5211 5 1 1 5210
0 5212 7 1 2 5207 5211
0 5213 5 1 1 5212
0 5214 7 1 2 64977 5213
0 5215 5 1 1 5214
0 5216 7 1 2 5203 5215
0 5217 7 1 2 5199 5216
0 5218 7 1 2 5197 5217
0 5219 5 1 1 5218
0 5220 7 1 2 76183 5219
0 5221 5 1 1 5220
0 5222 7 1 2 87324 5221
0 5223 5 1 1 5222
0 5224 7 1 2 81519 5223
0 5225 5 1 1 5224
0 5226 7 1 2 5172 5225
0 5227 5 1 1 5226
0 5228 7 1 2 88089 5227
0 5229 5 1 1 5228
0 5230 7 160 2 68939 72101
0 5231 5 1 1 88479
0 5232 7 4 2 76184 88480
0 5233 5 1 1 88639
0 5234 7 5 2 72541 83890
0 5235 7 2 2 80575 88643
0 5236 5 1 1 88648
0 5237 7 5 2 67533 76991
0 5238 7 2 2 81688 88650
0 5239 5 2 1 88655
0 5240 7 1 2 5236 88657
0 5241 5 3 1 5240
0 5242 7 1 2 70095 88659
0 5243 5 1 1 5242
0 5244 7 2 2 64978 86865
0 5245 5 2 1 88662
0 5246 7 1 2 88663 87783
0 5247 5 1 1 5246
0 5248 7 1 2 5243 5247
0 5249 5 1 1 5248
0 5250 7 1 2 64279 5249
0 5251 5 1 1 5250
0 5252 7 2 2 75095 86527
0 5253 5 2 1 88666
0 5254 7 1 2 88664 88668
0 5255 5 2 1 5254
0 5256 7 1 2 88670 87827
0 5257 5 1 1 5256
0 5258 7 1 2 5251 5257
0 5259 5 1 1 5258
0 5260 7 1 2 73893 5259
0 5261 5 1 1 5260
0 5262 7 2 2 86249 84656
0 5263 5 1 1 88672
0 5264 7 11 2 70362 80335
0 5265 5 12 1 88674
0 5266 7 3 2 88685 86784
0 5267 7 1 2 88673 88697
0 5268 5 1 1 5267
0 5269 7 1 2 5261 5268
0 5270 5 1 1 5269
0 5271 7 1 2 88640 5270
0 5272 5 1 1 5271
0 5273 7 1 2 5229 5272
0 5274 5 1 1 5273
0 5275 7 1 2 65911 5274
0 5276 5 1 1 5275
0 5277 7 12 2 66157 66658
0 5278 5 2 1 88700
0 5279 7 2 2 68583 88701
0 5280 5 1 1 88714
0 5281 7 1 2 5280 87091
0 5282 5 1 1 5281
0 5283 7 1 2 65306 5282
0 5284 5 1 1 5283
0 5285 7 1 2 71278 86226
0 5286 5 3 1 5285
0 5287 7 1 2 83100 88716
0 5288 5 1 1 5287
0 5289 7 1 2 5284 5288
0 5290 5 1 1 5289
0 5291 7 1 2 64603 5290
0 5292 5 1 1 5291
0 5293 7 5 2 66158 73670
0 5294 5 2 1 88719
0 5295 7 6 2 72938 84812
0 5296 5 1 1 88726
0 5297 7 1 2 88720 88727
0 5298 5 1 1 5297
0 5299 7 1 2 5292 5298
0 5300 5 1 1 5299
0 5301 7 2 2 75252 84931
0 5302 7 1 2 77790 79322
0 5303 7 1 2 88732 5302
0 5304 7 1 2 5300 5303
0 5305 5 1 1 5304
0 5306 7 1 2 5276 5305
0 5307 5 1 1 5306
0 5308 7 1 2 85851 5307
0 5309 5 1 1 5308
0 5310 7 1 2 72542 86386
0 5311 5 1 1 5310
0 5312 7 3 2 67534 82590
0 5313 7 2 2 76992 88734
0 5314 5 1 1 88737
0 5315 7 2 2 81582 88738
0 5316 7 2 2 81664 88739
0 5317 5 1 1 88741
0 5318 7 1 2 5311 5317
0 5319 5 1 1 5318
0 5320 7 1 2 64280 5319
0 5321 5 1 1 5320
0 5322 7 2 2 72543 87308
0 5323 7 3 2 66159 78307
0 5324 5 1 1 88745
0 5325 7 1 2 79979 88746
0 5326 7 1 2 88743 5325
0 5327 5 1 1 5326
0 5328 7 1 2 5321 5327
0 5329 5 1 1 5328
0 5330 7 1 2 70975 5329
0 5331 5 1 1 5330
0 5332 7 1 2 65912 87718
0 5333 5 1 1 5332
0 5334 7 5 2 64281 75253
0 5335 7 2 2 78401 88748
0 5336 5 1 1 88753
0 5337 7 1 2 79189 88754
0 5338 5 1 1 5337
0 5339 7 1 2 5333 5338
0 5340 5 1 1 5339
0 5341 7 1 2 80672 5340
0 5342 5 1 1 5341
0 5343 7 1 2 84657 87299
0 5344 5 1 1 5343
0 5345 7 1 2 69387 88742
0 5346 5 1 1 5345
0 5347 7 13 2 68584 84813
0 5348 5 6 1 88755
0 5349 7 1 2 88756 83254
0 5350 5 1 1 5349
0 5351 7 2 2 66160 83598
0 5352 5 3 1 88774
0 5353 7 1 2 83963 88775
0 5354 5 1 1 5353
0 5355 7 1 2 5350 5354
0 5356 5 1 1 5355
0 5357 7 1 2 75333 5356
0 5358 5 1 1 5357
0 5359 7 1 2 1978 88426
0 5360 5 1 1 5359
0 5361 7 1 2 71279 5360
0 5362 5 1 1 5361
0 5363 7 1 2 78768 5362
0 5364 5 1 1 5363
0 5365 7 1 2 65307 5364
0 5366 5 1 1 5365
0 5367 7 1 2 5358 5366
0 5368 5 1 1 5367
0 5369 7 1 2 68292 5368
0 5370 5 1 1 5369
0 5371 7 1 2 86192 83266
0 5372 5 1 1 5371
0 5373 7 1 2 86816 2671
0 5374 5 2 1 5373
0 5375 7 2 2 71280 88779
0 5376 5 1 1 88781
0 5377 7 1 2 81430 88782
0 5378 5 1 1 5377
0 5379 7 1 2 5372 5378
0 5380 5 1 1 5379
0 5381 7 1 2 71755 5380
0 5382 5 1 1 5381
0 5383 7 1 2 5370 5382
0 5384 5 1 1 5383
0 5385 7 1 2 84932 5384
0 5386 5 1 1 5385
0 5387 7 1 2 5346 5386
0 5388 7 1 2 5344 5387
0 5389 5 1 1 5388
0 5390 7 1 2 65913 5389
0 5391 5 1 1 5390
0 5392 7 1 2 5342 5391
0 5393 7 1 2 5331 5392
0 5394 5 1 1 5393
0 5395 7 1 2 88481 5394
0 5396 5 1 1 5395
0 5397 7 2 2 70096 87503
0 5398 7 1 2 88783 86429
0 5399 5 1 1 5398
0 5400 7 3 2 71569 87625
0 5401 5 4 1 88785
0 5402 7 2 2 88788 86916
0 5403 7 1 2 72544 88792
0 5404 5 1 1 5403
0 5405 7 1 2 87255 88651
0 5406 5 1 1 5405
0 5407 7 1 2 5404 5406
0 5408 5 1 1 5407
0 5409 7 1 2 69388 5408
0 5410 5 1 1 5409
0 5411 7 1 2 5399 5410
0 5412 5 1 1 5411
0 5413 7 1 2 65308 5412
0 5414 5 1 1 5413
0 5415 7 1 2 69389 82364
0 5416 5 1 1 5415
0 5417 7 2 2 84116 83402
0 5418 5 4 1 88794
0 5419 7 1 2 88796 83134
0 5420 5 1 1 5419
0 5421 7 1 2 5416 5420
0 5422 5 1 1 5421
0 5423 7 1 2 66458 5422
0 5424 5 2 1 5423
0 5425 7 2 2 86359 82615
0 5426 5 1 1 88802
0 5427 7 1 2 67915 88803
0 5428 5 1 1 5427
0 5429 7 1 2 69390 5428
0 5430 5 1 1 5429
0 5431 7 1 2 88800 5430
0 5432 5 1 1 5431
0 5433 7 1 2 70363 5432
0 5434 5 1 1 5433
0 5435 7 1 2 69391 86889
0 5436 5 1 1 5435
0 5437 7 1 2 5434 5436
0 5438 5 1 1 5437
0 5439 7 1 2 72545 5438
0 5440 5 1 1 5439
0 5441 7 1 2 5414 5440
0 5442 5 1 1 5441
0 5443 7 1 2 66161 5442
0 5444 5 1 1 5443
0 5445 7 1 2 81456 86485
0 5446 5 1 1 5445
0 5447 7 1 2 5444 5446
0 5448 5 1 1 5447
0 5449 7 1 2 64604 5448
0 5450 5 1 1 5449
0 5451 7 1 2 85769 85578
0 5452 5 2 1 5451
0 5453 7 1 2 64605 88804
0 5454 5 1 1 5453
0 5455 7 1 2 79074 86879
0 5456 5 1 1 5455
0 5457 7 1 2 72939 5456
0 5458 5 1 1 5457
0 5459 7 1 2 5454 5458
0 5460 5 1 1 5459
0 5461 7 1 2 75254 5460
0 5462 5 1 1 5461
0 5463 7 1 2 74487 83059
0 5464 5 1 1 5463
0 5465 7 1 2 86912 5464
0 5466 5 1 1 5465
0 5467 7 1 2 66162 5466
0 5468 5 1 1 5467
0 5469 7 1 2 2308 86189
0 5470 5 1 1 5469
0 5471 7 1 2 79951 5470
0 5472 5 1 1 5471
0 5473 7 2 2 76149 83038
0 5474 5 3 1 88806
0 5475 7 1 2 85770 88808
0 5476 5 1 1 5475
0 5477 7 1 2 76544 5476
0 5478 5 1 1 5477
0 5479 7 5 2 66163 83964
0 5480 5 1 1 88811
0 5481 7 3 2 72940 78567
0 5482 7 1 2 76407 88816
0 5483 5 1 1 5482
0 5484 7 1 2 5480 5483
0 5485 7 1 2 5478 5484
0 5486 5 1 1 5485
0 5487 7 1 2 66659 5486
0 5488 5 1 1 5487
0 5489 7 1 2 5472 5488
0 5490 5 1 1 5489
0 5491 7 1 2 74605 5490
0 5492 5 1 1 5491
0 5493 7 1 2 83981 85579
0 5494 5 1 1 5493
0 5495 7 1 2 66164 5494
0 5496 5 1 1 5495
0 5497 7 1 2 76545 86883
0 5498 5 1 1 5497
0 5499 7 1 2 5496 5498
0 5500 5 1 1 5499
0 5501 7 1 2 82039 5500
0 5502 5 1 1 5501
0 5503 7 1 2 67535 5502
0 5504 7 1 2 5492 5503
0 5505 7 1 2 5468 5504
0 5506 7 1 2 5462 5505
0 5507 5 1 1 5506
0 5508 7 10 2 71756 74840
0 5509 5 4 1 88819
0 5510 7 2 2 74606 88829
0 5511 5 3 1 88833
0 5512 7 1 2 66165 88834
0 5513 5 1 1 5512
0 5514 7 2 2 75334 82616
0 5515 5 2 1 88838
0 5516 7 1 2 88835 88839
0 5517 5 1 1 5516
0 5518 7 1 2 70364 5517
0 5519 7 1 2 5513 5518
0 5520 5 1 1 5519
0 5521 7 1 2 70365 88836
0 5522 5 2 1 5521
0 5523 7 3 2 88842 88789
0 5524 5 1 1 88844
0 5525 7 1 2 66166 5524
0 5526 5 1 1 5525
0 5527 7 1 2 74514 82127
0 5528 5 1 1 5527
0 5529 7 1 2 71281 82954
0 5530 7 1 2 5528 5529
0 5531 5 1 1 5530
0 5532 7 1 2 86660 5531
0 5533 5 1 1 5532
0 5534 7 1 2 65309 5533
0 5535 5 1 1 5534
0 5536 7 1 2 5526 5535
0 5537 7 1 2 5520 5536
0 5538 5 1 1 5537
0 5539 7 1 2 67916 5538
0 5540 5 1 1 5539
0 5541 7 1 2 72546 5540
0 5542 7 1 2 86658 5541
0 5543 5 1 1 5542
0 5544 7 1 2 64282 5543
0 5545 7 1 2 5507 5544
0 5546 5 1 1 5545
0 5547 7 5 2 73362 87449
0 5548 7 2 2 88847 87282
0 5549 7 1 2 72941 88852
0 5550 5 2 1 5549
0 5551 7 1 2 87154 88854
0 5552 5 1 1 5551
0 5553 7 1 2 66167 5552
0 5554 5 1 1 5553
0 5555 7 1 2 86441 5554
0 5556 5 1 1 5555
0 5557 7 1 2 81457 5556
0 5558 5 1 1 5557
0 5559 7 1 2 65914 5558
0 5560 7 1 2 5546 5559
0 5561 7 1 2 5450 5560
0 5562 5 1 1 5561
0 5563 7 2 2 70366 78618
0 5564 5 3 1 88856
0 5565 7 1 2 88858 87197
0 5566 5 2 1 5565
0 5567 7 1 2 66168 88861
0 5568 5 1 1 5567
0 5569 7 9 2 68293 81689
0 5570 5 1 1 88863
0 5571 7 1 2 77864 88864
0 5572 5 1 1 5571
0 5573 7 1 2 5568 5572
0 5574 5 1 1 5573
0 5575 7 1 2 64606 5574
0 5576 5 1 1 5575
0 5577 7 1 2 77865 86443
0 5578 5 1 1 5577
0 5579 7 1 2 87155 5578
0 5580 5 1 1 5579
0 5581 7 1 2 76546 5580
0 5582 5 1 1 5581
0 5583 7 2 2 82630 83343
0 5584 5 1 1 88872
0 5585 7 1 2 66169 88873
0 5586 5 2 1 5585
0 5587 7 1 2 71282 86436
0 5588 5 1 1 5587
0 5589 7 1 2 73671 88812
0 5590 5 1 1 5589
0 5591 7 1 2 5588 5590
0 5592 5 1 1 5591
0 5593 7 1 2 64979 5592
0 5594 5 1 1 5593
0 5595 7 1 2 88874 5594
0 5596 7 1 2 5582 5595
0 5597 7 1 2 5576 5596
0 5598 5 1 1 5597
0 5599 7 1 2 64283 5598
0 5600 5 1 1 5599
0 5601 7 6 2 69392 66660
0 5602 5 1 1 88876
0 5603 7 1 2 84801 5602
0 5604 5 1 1 5603
0 5605 7 1 2 83806 81665
0 5606 7 1 2 77696 5605
0 5607 7 1 2 5604 5606
0 5608 5 1 1 5607
0 5609 7 1 2 5600 5608
0 5610 5 1 1 5609
0 5611 7 1 2 72547 5610
0 5612 5 1 1 5611
0 5613 7 6 2 66170 84453
0 5614 5 1 1 88882
0 5615 7 1 2 88883 88740
0 5616 5 1 1 5615
0 5617 7 1 2 70976 5616
0 5618 7 1 2 5612 5617
0 5619 5 1 1 5618
0 5620 7 1 2 88090 5619
0 5621 7 1 2 5562 5620
0 5622 5 1 1 5621
0 5623 7 1 2 5396 5622
0 5624 5 1 1 5623
0 5625 7 1 2 85196 5624
0 5626 5 1 1 5625
0 5627 7 1 2 5309 5626
0 5628 5 1 1 5627
0 5629 7 1 2 88056 5628
0 5630 5 1 1 5629
0 5631 7 14 2 65619 66836
0 5632 7 5 2 65577 88888
0 5633 7 26 2 63952 65671
0 5634 5 3 1 88907
0 5635 7 73 2 88902 88908
0 5636 5 7 1 88936
0 5637 7 2 2 85197 77402
0 5638 7 1 2 87487 89016
0 5639 5 1 1 5638
0 5640 7 3 2 71570 85648
0 5641 5 1 1 89018
0 5642 7 5 2 88375 89019
0 5643 7 4 2 70097 89021
0 5644 5 1 1 89026
0 5645 7 2 2 65915 89027
0 5646 5 2 1 89030
0 5647 7 1 2 87504 83039
0 5648 5 4 1 5647
0 5649 7 1 2 64980 87469
0 5650 5 1 1 5649
0 5651 7 3 2 89034 5650
0 5652 5 11 1 89038
0 5653 7 1 2 70977 89041
0 5654 5 1 1 5653
0 5655 7 2 2 89032 5654
0 5656 5 1 1 89052
0 5657 7 1 2 80998 89053
0 5658 5 1 1 5657
0 5659 7 1 2 85852 5658
0 5660 5 1 1 5659
0 5661 7 1 2 5639 5660
0 5662 5 1 1 5661
0 5663 7 1 2 88482 5662
0 5664 5 1 1 5663
0 5665 7 5 2 73672 82312
0 5666 5 2 1 89054
0 5667 7 1 2 73894 87283
0 5668 5 3 1 5667
0 5669 7 1 2 89055 89061
0 5670 5 1 1 5669
0 5671 7 3 2 73363 80863
0 5672 5 2 1 89064
0 5673 7 1 2 66459 89065
0 5674 5 1 1 5673
0 5675 7 1 2 5670 5674
0 5676 5 1 1 5675
0 5677 7 1 2 70978 5676
0 5678 5 1 1 5677
0 5679 7 3 2 75335 79800
0 5680 7 2 2 82664 89069
0 5681 5 3 1 89072
0 5682 7 1 2 80999 89074
0 5683 7 1 2 5678 5682
0 5684 5 1 1 5683
0 5685 7 1 2 85853 5684
0 5686 5 1 1 5685
0 5687 7 1 2 78619 89017
0 5688 5 1 1 5687
0 5689 7 1 2 5686 5688
0 5690 5 1 1 5689
0 5691 7 1 2 88091 5690
0 5692 5 1 1 5691
0 5693 7 1 2 5664 5692
0 5694 5 1 1 5693
0 5695 7 1 2 64607 5694
0 5696 5 1 1 5695
0 5697 7 16 2 68772 69393
0 5698 7 2 2 87525 89077
0 5699 5 1 1 89093
0 5700 7 2 2 86000 75255
0 5701 5 1 1 89095
0 5702 7 2 2 77403 89096
0 5703 5 1 1 89097
0 5704 7 1 2 5699 5703
0 5705 5 1 1 5704
0 5706 7 1 2 88483 5705
0 5707 5 1 1 5706
0 5708 7 4 2 73673 88092
0 5709 5 2 1 89099
0 5710 7 6 2 73364 85854
0 5711 7 1 2 89105 87082
0 5712 7 1 2 89100 5711
0 5713 5 1 1 5712
0 5714 7 1 2 5707 5713
0 5715 5 1 1 5714
0 5716 7 1 2 66661 5715
0 5717 5 1 1 5716
0 5718 7 1 2 87721 87497
0 5719 5 1 1 5718
0 5720 7 1 2 5717 5719
0 5721 5 1 1 5720
0 5722 7 1 2 65310 5721
0 5723 5 1 1 5722
0 5724 7 4 2 72007 79608
0 5725 7 19 2 68940 69394
0 5726 7 1 2 77012 89115
0 5727 5 2 1 5726
0 5728 7 9 2 63856 70367
0 5729 7 1 2 89136 87523
0 5730 5 1 1 5729
0 5731 7 1 2 89134 5730
0 5732 5 1 1 5731
0 5733 7 1 2 89111 5732
0 5734 5 1 1 5733
0 5735 7 1 2 5723 5734
0 5736 7 1 2 5696 5735
0 5737 5 1 1 5736
0 5738 7 1 2 66171 5737
0 5739 5 1 1 5738
0 5740 7 1 2 85668 89094
0 5741 5 1 1 5740
0 5742 7 1 2 81690 89098
0 5743 5 2 1 5742
0 5744 7 1 2 5741 89145
0 5745 5 1 1 5744
0 5746 7 1 2 88484 5745
0 5747 5 1 1 5746
0 5748 7 11 2 66662 72008
0 5749 7 2 2 89147 87722
0 5750 7 2 2 78620 74280
0 5751 7 1 2 87310 89160
0 5752 7 1 2 89158 5751
0 5753 5 1 1 5752
0 5754 7 1 2 5747 5753
0 5755 5 1 1 5754
0 5756 7 1 2 64608 5755
0 5757 5 1 1 5756
0 5758 7 1 2 5739 5757
0 5759 5 1 1 5758
0 5760 7 1 2 72942 5759
0 5761 5 1 1 5760
0 5762 7 11 2 82955 87571
0 5763 5 3 1 89162
0 5764 7 6 2 67917 89163
0 5765 7 1 2 75336 89176
0 5766 5 1 1 5765
0 5767 7 1 2 64284 5766
0 5768 5 1 1 5767
0 5769 7 1 2 73365 5768
0 5770 5 1 1 5769
0 5771 7 1 2 64285 4756
0 5772 5 1 1 5771
0 5773 7 1 2 81691 5772
0 5774 5 1 1 5773
0 5775 7 1 2 5770 5774
0 5776 5 1 1 5775
0 5777 7 1 2 89112 5776
0 5778 5 1 1 5777
0 5779 7 1 2 89146 5778
0 5780 5 1 1 5779
0 5781 7 1 2 88485 5780
0 5782 5 1 1 5781
0 5783 7 10 2 85855 88093
0 5784 7 2 2 82665 83891
0 5785 5 1 1 89192
0 5786 7 2 2 86538 78621
0 5787 7 1 2 70979 89194
0 5788 5 1 1 5787
0 5789 7 1 2 5785 5788
0 5790 5 1 1 5789
0 5791 7 1 2 65311 5790
0 5792 5 1 1 5791
0 5793 7 2 2 70368 84959
0 5794 7 1 2 83892 89196
0 5795 5 1 1 5794
0 5796 7 1 2 5792 5795
0 5797 5 1 1 5796
0 5798 7 1 2 89182 5797
0 5799 5 1 1 5798
0 5800 7 1 2 5782 5799
0 5801 5 1 1 5800
0 5802 7 1 2 76185 5801
0 5803 5 1 1 5802
0 5804 7 1 2 5761 5803
0 5805 5 1 1 5804
0 5806 7 1 2 72548 5805
0 5807 5 1 1 5806
0 5808 7 1 2 84899 76186
0 5809 5 2 1 5808
0 5810 7 5 2 66460 81833
0 5811 5 3 1 89200
0 5812 7 7 2 86461 89205
0 5813 5 3 1 89208
0 5814 7 1 2 65916 89215
0 5815 5 1 1 5814
0 5816 7 1 2 89198 5815
0 5817 5 1 1 5816
0 5818 7 1 2 67918 5817
0 5819 5 1 1 5818
0 5820 7 4 2 72943 89164
0 5821 7 1 2 81271 89218
0 5822 5 1 1 5821
0 5823 7 1 2 5819 5822
0 5824 5 1 1 5823
0 5825 7 1 2 68294 5824
0 5826 5 1 1 5825
0 5827 7 3 2 85669 76276
0 5828 5 1 1 89222
0 5829 7 1 2 87048 89223
0 5830 5 1 1 5829
0 5831 7 1 2 5826 5830
0 5832 5 1 1 5831
0 5833 7 1 2 72549 5832
0 5834 5 1 1 5833
0 5835 7 1 2 76277 81191
0 5836 5 2 1 5835
0 5837 7 1 2 81692 78426
0 5838 7 1 2 89225 5837
0 5839 5 1 1 5838
0 5840 7 1 2 5834 5839
0 5841 5 1 1 5840
0 5842 7 1 2 88486 5841
0 5843 5 1 1 5842
0 5844 7 2 2 73674 87488
0 5845 5 1 1 89227
0 5846 7 1 2 78427 89228
0 5847 5 1 1 5846
0 5848 7 1 2 70980 654
0 5849 5 1 1 5848
0 5850 7 8 2 72550 76278
0 5851 5 1 1 89229
0 5852 7 1 2 80576 89230
0 5853 7 1 2 5849 5852
0 5854 5 1 1 5853
0 5855 7 1 2 5847 5854
0 5856 5 1 1 5855
0 5857 7 1 2 72944 5856
0 5858 5 1 1 5857
0 5859 7 3 2 80577 84990
0 5860 5 4 1 89237
0 5861 7 6 2 66461 81393
0 5862 7 1 2 86763 89244
0 5863 5 1 1 5862
0 5864 7 1 2 89240 5863
0 5865 5 1 1 5864
0 5866 7 1 2 64981 5865
0 5867 5 1 1 5866
0 5868 7 3 2 68585 73895
0 5869 5 1 1 89250
0 5870 7 7 2 64609 73675
0 5871 5 1 1 89253
0 5872 7 1 2 89254 82186
0 5873 5 2 1 5872
0 5874 7 1 2 89241 89260
0 5875 5 1 1 5874
0 5876 7 1 2 5869 5875
0 5877 5 1 1 5876
0 5878 7 1 2 5867 5877
0 5879 5 1 1 5878
0 5880 7 1 2 65917 5879
0 5881 5 1 1 5880
0 5882 7 1 2 5858 5881
0 5883 5 1 1 5882
0 5884 7 1 2 88094 5883
0 5885 5 1 1 5884
0 5886 7 4 2 75901 87879
0 5887 7 3 2 70981 89262
0 5888 5 2 1 89266
0 5889 7 7 2 71571 75547
0 5890 5 4 1 89271
0 5891 7 1 2 76187 89278
0 5892 5 1 1 5891
0 5893 7 1 2 70098 5892
0 5894 5 1 1 5893
0 5895 7 2 2 76279 77705
0 5896 5 2 1 89282
0 5897 7 1 2 78428 89284
0 5898 7 1 2 5894 5897
0 5899 5 1 1 5898
0 5900 7 1 2 89269 5899
0 5901 7 1 2 5885 5900
0 5902 7 1 2 5843 5901
0 5903 5 1 1 5902
0 5904 7 1 2 88283 5231
0 5905 5 12 1 5904
0 5906 7 1 2 85856 89286
0 5907 7 1 2 5903 5906
0 5908 5 1 1 5907
0 5909 7 20 2 79359 74231
0 5910 5 8 1 89298
0 5911 7 1 2 87723 79160
0 5912 5 1 1 5911
0 5913 7 1 2 89318 5912
0 5914 5 3 1 5913
0 5915 7 1 2 74607 89326
0 5916 5 1 1 5915
0 5917 7 8 2 85857 88487
0 5918 7 1 2 82040 89329
0 5919 5 1 1 5918
0 5920 7 1 2 5916 5919
0 5921 5 1 1 5920
0 5922 7 1 2 78429 5921
0 5923 5 1 1 5922
0 5924 7 2 2 70982 87396
0 5925 7 1 2 89337 84386
0 5926 5 1 1 5925
0 5927 7 1 2 5923 5926
0 5928 5 1 1 5927
0 5929 7 1 2 85670 5928
0 5930 5 1 1 5929
0 5931 7 4 2 63857 78718
0 5932 5 1 1 89339
0 5933 7 1 2 85810 88488
0 5934 5 1 1 5933
0 5935 7 1 2 5932 5934
0 5936 5 1 1 5935
0 5937 7 1 2 74608 5936
0 5938 5 1 1 5937
0 5939 7 17 2 67046 73366
0 5940 7 7 2 63858 89343
0 5941 5 2 1 89360
0 5942 7 1 2 82041 89361
0 5943 5 1 1 5942
0 5944 7 1 2 5938 5943
0 5945 5 1 1 5944
0 5946 7 1 2 85858 5945
0 5947 5 1 1 5946
0 5948 7 1 2 85198 89362
0 5949 5 1 1 5948
0 5950 7 4 2 82313 87450
0 5951 5 2 1 89369
0 5952 7 2 2 80241 89370
0 5953 5 2 1 89375
0 5954 7 1 2 67919 89377
0 5955 5 1 1 5954
0 5956 7 1 2 89327 5955
0 5957 5 1 1 5956
0 5958 7 1 2 5949 5957
0 5959 7 1 2 5947 5958
0 5960 5 1 1 5959
0 5961 7 1 2 67536 5960
0 5962 5 1 1 5961
0 5963 7 1 2 89238 89183
0 5964 5 1 1 5963
0 5965 7 7 2 72009 87397
0 5966 7 14 2 72102 67920
0 5967 7 3 2 89379 89386
0 5968 7 1 2 72551 89400
0 5969 5 1 1 5968
0 5970 7 9 2 82754 74095
0 5971 5 1 1 89403
0 5972 7 1 2 79715 89404
0 5973 5 1 1 5972
0 5974 7 1 2 5969 5973
0 5975 5 1 1 5974
0 5976 7 1 2 81834 5975
0 5977 5 1 1 5976
0 5978 7 7 2 72945 85199
0 5979 5 1 1 89412
0 5980 7 3 2 70369 67047
0 5981 7 4 2 89419 84638
0 5982 5 1 1 89422
0 5983 7 1 2 89413 89423
0 5984 5 1 1 5983
0 5985 7 1 2 5977 5984
0 5986 5 1 1 5985
0 5987 7 1 2 68295 5986
0 5988 5 1 1 5987
0 5989 7 1 2 5964 5988
0 5990 7 1 2 5962 5989
0 5991 5 1 1 5990
0 5992 7 1 2 65918 5991
0 5993 5 1 1 5992
0 5994 7 1 2 5930 5993
0 5995 5 1 1 5994
0 5996 7 1 2 76547 5995
0 5997 5 1 1 5996
0 5998 7 6 2 63737 65919
0 5999 7 4 2 66942 89426
0 6000 7 1 2 76280 87534
0 6001 5 1 1 6000
0 6002 7 1 2 67537 6001
0 6003 5 1 1 6002
0 6004 7 6 2 72552 75955
0 6005 5 1 1 89436
0 6006 7 1 2 82631 74993
0 6007 5 1 1 6006
0 6008 7 1 2 89437 6007
0 6009 5 1 1 6008
0 6010 7 1 2 6003 6009
0 6011 5 1 1 6010
0 6012 7 1 2 88489 6011
0 6013 5 1 1 6012
0 6014 7 2 2 64610 81693
0 6015 5 2 1 89442
0 6016 7 1 2 89444 3721
0 6017 5 1 1 6016
0 6018 7 1 2 67538 6017
0 6019 5 1 1 6018
0 6020 7 1 2 68296 82071
0 6021 7 1 2 86040 6020
0 6022 5 1 1 6021
0 6023 7 1 2 1925 6022
0 6024 7 1 2 6019 6023
0 6025 5 1 1 6024
0 6026 7 1 2 88095 6025
0 6027 5 1 1 6026
0 6028 7 1 2 6013 6027
0 6029 5 1 1 6028
0 6030 7 1 2 89432 6029
0 6031 5 1 1 6030
0 6032 7 1 2 5997 6031
0 6033 7 1 2 5908 6032
0 6034 5 1 1 6033
0 6035 7 1 2 64286 6034
0 6036 5 1 1 6035
0 6037 7 2 2 73942 77404
0 6038 7 1 2 89446 89263
0 6039 5 1 1 6038
0 6040 7 2 2 65920 74994
0 6041 5 3 1 89448
0 6042 7 2 2 73676 81520
0 6043 5 1 1 89453
0 6044 7 1 2 89449 89454
0 6045 5 1 1 6044
0 6046 7 1 2 6039 6045
0 6047 5 1 1 6046
0 6048 7 1 2 89405 6047
0 6049 5 1 1 6048
0 6050 7 6 2 68941 74215
0 6051 5 1 1 89455
0 6052 7 1 2 87848 89456
0 6053 5 1 1 6052
0 6054 7 1 2 63859 87856
0 6055 5 1 1 6054
0 6056 7 1 2 6053 6055
0 6057 5 1 1 6056
0 6058 7 1 2 72553 6057
0 6059 5 1 1 6058
0 6060 7 1 2 88284 6051
0 6061 5 14 1 6060
0 6062 7 1 2 81521 89461
0 6063 7 1 2 87861 6062
0 6064 5 1 1 6063
0 6065 7 1 2 6059 6064
0 6066 5 1 1 6065
0 6067 7 1 2 66172 6066
0 6068 5 1 1 6067
0 6069 7 1 2 87892 89462
0 6070 5 1 1 6069
0 6071 7 2 2 76447 89457
0 6072 5 1 1 89475
0 6073 7 6 2 67921 88096
0 6074 7 1 2 76281 89477
0 6075 5 1 1 6074
0 6076 7 1 2 6072 6075
0 6077 5 1 1 6076
0 6078 7 2 2 72554 6077
0 6079 5 1 1 89483
0 6080 7 1 2 64287 89484
0 6081 5 1 1 6080
0 6082 7 1 2 6070 6081
0 6083 7 1 2 6068 6082
0 6084 5 1 1 6083
0 6085 7 1 2 65921 6084
0 6086 5 1 1 6085
0 6087 7 3 2 64611 87938
0 6088 5 2 1 89485
0 6089 7 1 2 80264 89488
0 6090 5 1 1 6089
0 6091 7 3 2 70983 82236
0 6092 5 1 1 89490
0 6093 7 1 2 89491 89463
0 6094 7 1 2 6090 6093
0 6095 5 1 1 6094
0 6096 7 1 2 6086 6095
0 6097 5 1 1 6096
0 6098 7 1 2 85859 6097
0 6099 5 1 1 6098
0 6100 7 1 2 6049 6099
0 6101 5 1 1 6100
0 6102 7 1 2 80673 6101
0 6103 5 1 1 6102
0 6104 7 1 2 6036 6103
0 6105 7 1 2 5807 6104
0 6106 5 1 1 6105
0 6107 7 1 2 88937 6106
0 6108 5 1 1 6107
0 6109 7 8 2 65578 70652
0 6110 5 1 1 89493
0 6111 7 27 2 69042 70703
0 6112 7 3 2 89494 89501
0 6113 5 1 1 89528
0 6114 7 22 2 65620 65672
0 6115 7 5 2 63953 70612
0 6116 7 2 2 89531 89553
0 6117 5 1 1 89558
0 6118 7 1 2 6113 6117
0 6119 5 32 1 6118
0 6120 7 3 2 89427 76372
0 6121 7 1 2 68586 80225
0 6122 7 1 2 89592 6121
0 6123 5 1 1 6122
0 6124 7 3 2 80114 78338
0 6125 7 1 2 86487 85834
0 6126 7 1 2 89595 6125
0 6127 5 1 1 6126
0 6128 7 1 2 6123 6127
0 6129 5 1 1 6128
0 6130 7 1 2 84814 6129
0 6131 5 1 1 6130
0 6132 7 1 2 86259 5845
0 6133 5 1 1 6132
0 6134 7 1 2 70984 6133
0 6135 5 1 1 6134
0 6136 7 1 2 89075 6135
0 6137 5 1 1 6136
0 6138 7 1 2 64612 6137
0 6139 5 1 1 6138
0 6140 7 2 2 65312 80511
0 6141 5 1 1 89598
0 6142 7 1 2 83454 6141
0 6143 5 2 1 6142
0 6144 7 1 2 87664 89600
0 6145 5 1 1 6144
0 6146 7 7 2 82890 78622
0 6147 5 2 1 89602
0 6148 7 1 2 89603 87311
0 6149 5 1 1 6148
0 6150 7 1 2 6145 6149
0 6151 7 1 2 6139 6150
0 6152 5 1 1 6151
0 6153 7 1 2 78191 6152
0 6154 5 1 1 6153
0 6155 7 1 2 6131 6154
0 6156 5 1 1 6155
0 6157 7 1 2 88097 6156
0 6158 5 1 1 6157
0 6159 7 3 2 76373 79444
0 6160 7 2 2 89611 88490
0 6161 5 1 1 89614
0 6162 7 1 2 5656 89615
0 6163 5 1 1 6162
0 6164 7 1 2 6158 6163
0 6165 5 1 1 6164
0 6166 7 1 2 66173 6165
0 6167 5 1 1 6166
0 6168 7 3 2 66462 82891
0 6169 5 2 1 89616
0 6170 7 3 2 79600 76835
0 6171 7 2 2 89617 89621
0 6172 7 10 2 63860 64613
0 6173 7 8 2 63738 89626
0 6174 7 1 2 89636 87312
0 6175 7 1 2 89624 6174
0 6176 5 1 1 6175
0 6177 7 4 2 66174 67048
0 6178 7 2 2 89627 89644
0 6179 5 1 1 89648
0 6180 7 1 2 85671 76548
0 6181 5 1 1 6180
0 6182 7 1 2 76282 6181
0 6183 5 2 1 6182
0 6184 7 1 2 88491 89650
0 6185 5 1 1 6184
0 6186 7 1 2 6179 6185
0 6187 5 2 1 6186
0 6188 7 1 2 89652 89593
0 6189 5 1 1 6188
0 6190 7 3 2 77280 88492
0 6191 7 1 2 68297 89654
0 6192 5 1 1 6191
0 6193 7 1 2 70099 89363
0 6194 5 1 1 6193
0 6195 7 1 2 6192 6194
0 6196 5 1 1 6195
0 6197 7 1 2 66175 6196
0 6198 5 2 1 6197
0 6199 7 1 2 64982 79307
0 6200 5 1 1 6199
0 6201 7 1 2 74609 82165
0 6202 5 2 1 6201
0 6203 7 1 2 6200 89659
0 6204 5 1 1 6203
0 6205 7 1 2 89464 6204
0 6206 5 1 1 6205
0 6207 7 1 2 89657 6206
0 6208 5 1 1 6207
0 6209 7 1 2 65922 6208
0 6210 5 1 1 6209
0 6211 7 3 2 64614 77960
0 6212 5 2 1 89661
0 6213 7 2 2 80115 89662
0 6214 5 1 1 89666
0 6215 7 1 2 66463 89667
0 6216 7 1 2 89465 6215
0 6217 5 1 1 6216
0 6218 7 1 2 6210 6217
0 6219 5 1 1 6218
0 6220 7 1 2 66663 6219
0 6221 5 1 1 6220
0 6222 7 11 2 72103 68587
0 6223 7 6 2 68942 89668
0 6224 5 1 1 89679
0 6225 7 1 2 76188 82666
0 6226 7 1 2 89680 6225
0 6227 5 1 1 6226
0 6228 7 1 2 6221 6227
0 6229 5 1 1 6228
0 6230 7 1 2 65313 6229
0 6231 5 1 1 6230
0 6232 7 11 2 68943 71757
0 6233 5 1 1 89685
0 6234 7 1 2 68588 321
0 6235 7 1 2 6233 6234
0 6236 7 1 2 89287 6235
0 6237 5 1 1 6236
0 6238 7 2 2 81835 88098
0 6239 5 6 1 89696
0 6240 7 1 2 77082 80089
0 6241 5 5 1 6240
0 6242 7 3 2 89686 76121
0 6243 5 1 1 89709
0 6244 7 1 2 89704 89710
0 6245 5 1 1 6244
0 6246 7 1 2 89698 6245
0 6247 7 1 2 6237 6246
0 6248 5 1 1 6247
0 6249 7 1 2 76189 6248
0 6250 5 1 1 6249
0 6251 7 2 2 76549 87693
0 6252 5 1 1 89712
0 6253 7 6 2 72104 89687
0 6254 7 1 2 79337 89714
0 6255 5 1 1 6254
0 6256 7 1 2 89699 6255
0 6257 5 1 1 6256
0 6258 7 1 2 89713 6257
0 6259 5 2 1 6258
0 6260 7 7 2 71758 72105
0 6261 7 5 2 68944 89722
0 6262 5 2 1 89729
0 6263 7 3 2 78623 89730
0 6264 7 5 2 64983 76550
0 6265 5 1 1 89739
0 6266 7 2 2 70370 89740
0 6267 7 1 2 89736 89744
0 6268 5 1 1 6267
0 6269 7 1 2 89720 6268
0 6270 7 1 2 6250 6269
0 6271 5 1 1 6270
0 6272 7 1 2 65923 6271
0 6273 5 1 1 6272
0 6274 7 1 2 6231 6273
0 6275 5 1 1 6274
0 6276 7 1 2 85112 6275
0 6277 5 1 1 6276
0 6278 7 1 2 6189 6277
0 6279 5 1 1 6278
0 6280 7 1 2 69395 6279
0 6281 5 1 1 6280
0 6282 7 1 2 6176 6281
0 6283 7 1 2 6167 6282
0 6284 5 1 1 6283
0 6285 7 1 2 72946 6284
0 6286 5 1 1 6285
0 6287 7 4 2 66176 78192
0 6288 7 2 2 80479 78738
0 6289 7 7 2 71759 67049
0 6290 7 5 2 63861 89752
0 6291 5 3 1 89759
0 6292 7 1 2 89750 89760
0 6293 5 1 1 6292
0 6294 7 5 2 72106 87907
0 6295 5 1 1 89767
0 6296 7 1 2 76673 89768
0 6297 7 1 2 87539 6296
0 6298 5 1 1 6297
0 6299 7 1 2 6293 6298
0 6300 5 1 1 6299
0 6301 7 1 2 89746 6300
0 6302 5 1 1 6301
0 6303 7 7 2 72947 78193
0 6304 5 1 1 89772
0 6305 7 1 2 89773 89653
0 6306 5 1 1 6305
0 6307 7 2 2 64984 74727
0 6308 5 1 1 89779
0 6309 7 1 2 75066 6308
0 6310 5 1 1 6309
0 6311 7 1 2 88493 6310
0 6312 5 1 1 6311
0 6313 7 1 2 64985 89478
0 6314 5 1 1 6313
0 6315 7 1 2 6312 6314
0 6316 5 1 1 6315
0 6317 7 1 2 82892 6316
0 6318 5 1 1 6317
0 6319 7 3 2 63862 82956
0 6320 7 1 2 89645 89781
0 6321 5 1 1 6320
0 6322 7 1 2 6318 6321
0 6323 5 1 1 6322
0 6324 7 1 2 65314 6323
0 6325 5 1 1 6324
0 6326 7 2 2 82365 88099
0 6327 5 1 1 89784
0 6328 7 1 2 86941 88494
0 6329 7 1 2 83576 6328
0 6330 5 1 1 6329
0 6331 7 1 2 6327 6330
0 6332 5 1 1 6331
0 6333 7 1 2 79063 6332
0 6334 5 1 1 6333
0 6335 7 1 2 6325 6334
0 6336 5 1 1 6335
0 6337 7 1 2 66464 6336
0 6338 5 1 1 6337
0 6339 7 5 2 85609 83076
0 6340 7 1 2 89786 88100
0 6341 5 1 1 6340
0 6342 7 4 2 67050 89137
0 6343 5 3 1 89791
0 6344 7 1 2 87356 88495
0 6345 5 1 1 6344
0 6346 7 1 2 89795 6345
0 6347 5 1 1 6346
0 6348 7 2 2 73677 6347
0 6349 5 1 1 89798
0 6350 7 1 2 64986 89799
0 6351 5 1 1 6350
0 6352 7 1 2 6341 6351
0 6353 5 1 1 6352
0 6354 7 1 2 66177 6353
0 6355 5 1 1 6354
0 6356 7 1 2 6338 6355
0 6357 5 1 1 6356
0 6358 7 1 2 64615 6357
0 6359 5 1 1 6358
0 6360 7 1 2 78624 78794
0 6361 5 4 1 6360
0 6362 7 1 2 68298 78964
0 6363 5 2 1 6362
0 6364 7 1 2 89800 89804
0 6365 5 1 1 6364
0 6366 7 1 2 89466 6365
0 6367 5 1 1 6366
0 6368 7 1 2 89658 6367
0 6369 5 1 1 6368
0 6370 7 1 2 81694 6369
0 6371 5 1 1 6370
0 6372 7 5 2 68945 76122
0 6373 5 1 1 89806
0 6374 7 1 2 83436 89807
0 6375 7 1 2 87200 6374
0 6376 5 1 1 6375
0 6377 7 1 2 89721 6376
0 6378 7 1 2 6371 6377
0 6379 5 1 1 6378
0 6380 7 1 2 72948 6379
0 6381 5 1 1 6380
0 6382 7 8 2 64987 77041
0 6383 5 2 1 89811
0 6384 7 2 2 81695 89812
0 6385 7 5 2 68946 77013
0 6386 5 3 1 89823
0 6387 7 1 2 88285 89828
0 6388 5 2 1 6387
0 6389 7 2 2 67922 89831
0 6390 5 1 1 89833
0 6391 7 2 2 73678 89834
0 6392 7 1 2 89821 89835
0 6393 5 1 1 6392
0 6394 7 1 2 6381 6393
0 6395 7 1 2 6359 6394
0 6396 5 1 1 6395
0 6397 7 1 2 85113 6396
0 6398 5 1 1 6397
0 6399 7 1 2 6306 6398
0 6400 5 1 1 6399
0 6401 7 1 2 70985 6400
0 6402 5 1 1 6401
0 6403 7 1 2 6302 6402
0 6404 5 1 1 6403
0 6405 7 1 2 64288 6404
0 6406 5 1 1 6405
0 6407 7 1 2 69396 5426
0 6408 5 1 1 6407
0 6409 7 1 2 88801 6408
0 6410 5 1 1 6409
0 6411 7 1 2 70371 6410
0 6412 5 1 1 6411
0 6413 7 1 2 79980 88793
0 6414 5 1 1 6413
0 6415 7 1 2 6412 6414
0 6416 5 1 1 6415
0 6417 7 1 2 88101 6416
0 6418 5 1 1 6417
0 6419 7 3 2 72107 89116
0 6420 7 1 2 86970 86153
0 6421 5 1 1 6420
0 6422 7 1 2 73679 6421
0 6423 5 1 1 6422
0 6424 7 1 2 86281 6423
0 6425 5 1 1 6424
0 6426 7 1 2 89837 6425
0 6427 5 1 1 6426
0 6428 7 1 2 6418 6427
0 6429 5 1 1 6428
0 6430 7 1 2 85114 6429
0 6431 5 1 1 6430
0 6432 7 6 2 63863 87587
0 6433 5 4 1 89840
0 6434 7 1 2 81836 81497
0 6435 5 2 1 6434
0 6436 7 1 2 86301 89850
0 6437 5 1 1 6436
0 6438 7 1 2 88496 6437
0 6439 5 1 1 6438
0 6440 7 1 2 89846 6439
0 6441 5 1 1 6440
0 6442 7 1 2 68589 6441
0 6443 5 1 1 6442
0 6444 7 1 2 88497 87367
0 6445 5 1 1 6444
0 6446 7 1 2 6443 6445
0 6447 5 1 1 6446
0 6448 7 1 2 67923 6447
0 6449 5 1 1 6448
0 6450 7 2 2 69397 85672
0 6451 5 3 1 89852
0 6452 7 1 2 89853 88498
0 6453 5 1 1 6452
0 6454 7 1 2 6449 6453
0 6455 5 1 1 6454
0 6456 7 1 2 78194 6455
0 6457 5 1 1 6456
0 6458 7 1 2 6431 6457
0 6459 5 1 1 6458
0 6460 7 1 2 76190 6459
0 6461 5 1 1 6460
0 6462 7 3 2 76551 75501
0 6463 7 1 2 89078 86423
0 6464 7 1 2 89857 6463
0 6465 7 1 2 89836 6464
0 6466 5 1 1 6465
0 6467 7 1 2 6461 6466
0 6468 5 1 1 6467
0 6469 7 1 2 65924 6468
0 6470 5 1 1 6469
0 6471 7 14 2 63864 69398
0 6472 7 7 2 67051 89860
0 6473 5 1 1 89874
0 6474 7 5 2 75337 88102
0 6475 5 2 1 89881
0 6476 7 1 2 74216 83875
0 6477 5 1 1 6476
0 6478 7 1 2 89886 6477
0 6479 5 1 1 6478
0 6480 7 1 2 67924 6479
0 6481 5 1 1 6480
0 6482 7 1 2 6473 6481
0 6483 5 1 1 6482
0 6484 7 1 2 65925 6483
0 6485 5 1 1 6484
0 6486 7 2 2 87694 89467
0 6487 7 1 2 82563 89888
0 6488 5 1 1 6487
0 6489 7 1 2 6485 6488
0 6490 5 1 1 6489
0 6491 7 1 2 78195 6490
0 6492 5 1 1 6491
0 6493 7 13 2 72108 75722
0 6494 7 7 2 87398 89890
0 6495 7 1 2 80980 89903
0 6496 7 1 2 87716 6495
0 6497 5 1 1 6496
0 6498 7 1 2 6492 6497
0 6499 5 1 1 6498
0 6500 7 1 2 64616 6499
0 6501 5 1 1 6500
0 6502 7 9 2 65926 72949
0 6503 7 1 2 88103 87851
0 6504 5 1 1 6503
0 6505 7 1 2 74217 89117
0 6506 5 1 1 6505
0 6507 7 1 2 6504 6506
0 6508 5 1 1 6507
0 6509 7 1 2 78196 6508
0 6510 5 1 1 6509
0 6511 7 1 2 87995 87399
0 6512 7 1 2 87976 6511
0 6513 5 1 1 6512
0 6514 7 1 2 6510 6513
0 6515 5 1 1 6514
0 6516 7 1 2 89910 6515
0 6517 5 1 1 6516
0 6518 7 1 2 6501 6517
0 6519 5 1 1 6518
0 6520 7 1 2 66178 6519
0 6521 5 1 1 6520
0 6522 7 3 2 75723 77720
0 6523 7 11 2 68773 64988
0 6524 5 1 1 89922
0 6525 7 2 2 89923 79311
0 6526 7 1 2 89919 89933
0 6527 5 1 1 6526
0 6528 7 1 2 78197 89468
0 6529 5 1 1 6528
0 6530 7 1 2 6527 6529
0 6531 5 2 1 6530
0 6532 7 1 2 75598 80981
0 6533 7 1 2 89935 6532
0 6534 5 1 1 6533
0 6535 7 1 2 6521 6534
0 6536 5 1 1 6535
0 6537 7 1 2 80674 6536
0 6538 5 1 1 6537
0 6539 7 4 2 66179 87505
0 6540 7 2 2 89937 89637
0 6541 7 1 2 87313 89622
0 6542 7 1 2 89941 6541
0 6543 5 1 1 6542
0 6544 7 1 2 6538 6543
0 6545 7 1 2 6470 6544
0 6546 7 1 2 6406 6545
0 6547 7 1 2 6286 6546
0 6548 5 1 1 6547
0 6549 7 1 2 72555 6548
0 6550 5 1 1 6549
0 6551 7 3 2 66180 82735
0 6552 5 3 1 89943
0 6553 7 1 2 86764 74995
0 6554 5 2 1 6553
0 6555 7 1 2 89946 89949
0 6556 7 1 2 86796 6555
0 6557 5 1 1 6556
0 6558 7 1 2 75040 6557
0 6559 5 1 1 6558
0 6560 7 1 2 66181 83918
0 6561 5 1 1 6560
0 6562 7 1 2 87044 6561
0 6563 5 1 1 6562
0 6564 7 1 2 64617 6563
0 6565 5 1 1 6564
0 6566 7 1 2 74996 86820
0 6567 5 1 1 6566
0 6568 7 1 2 75956 86826
0 6569 5 1 1 6568
0 6570 7 1 2 73680 6569
0 6571 5 1 1 6570
0 6572 7 1 2 6567 6571
0 6573 7 1 2 6565 6572
0 6574 7 1 2 6559 6573
0 6575 5 1 1 6574
0 6576 7 1 2 67539 6575
0 6577 5 1 1 6576
0 6578 7 6 2 80090 83317
0 6579 5 1 1 89951
0 6580 7 1 2 89952 83865
0 6581 5 1 1 6580
0 6582 7 2 2 67925 6581
0 6583 5 1 1 89957
0 6584 7 1 2 83251 6583
0 6585 5 1 1 6584
0 6586 7 1 2 86832 6585
0 6587 5 1 1 6586
0 6588 7 1 2 6577 6587
0 6589 5 1 1 6588
0 6590 7 1 2 88104 6589
0 6591 5 1 1 6590
0 6592 7 1 2 67926 86121
0 6593 5 1 1 6592
0 6594 7 1 2 68590 83240
0 6595 5 1 1 6594
0 6596 7 1 2 6593 6595
0 6597 5 1 1 6596
0 6598 7 1 2 81837 6597
0 6599 5 1 1 6598
0 6600 7 3 2 70372 76283
0 6601 7 2 2 71760 89959
0 6602 5 1 1 89962
0 6603 7 1 2 72950 89963
0 6604 5 1 1 6603
0 6605 7 1 2 6599 6604
0 6606 5 1 1 6605
0 6607 7 1 2 68299 6606
0 6608 5 1 1 6607
0 6609 7 1 2 76284 87000
0 6610 5 2 1 6609
0 6611 7 1 2 72556 89964
0 6612 7 1 2 6608 6611
0 6613 5 1 1 6612
0 6614 7 1 2 75957 82282
0 6615 5 1 1 6614
0 6616 7 3 2 74997 6615
0 6617 5 1 1 89966
0 6618 7 1 2 74936 87284
0 6619 5 2 1 6618
0 6620 7 1 2 64618 89969
0 6621 5 1 1 6620
0 6622 7 1 2 6617 6621
0 6623 5 1 1 6622
0 6624 7 1 2 73943 6623
0 6625 5 1 1 6624
0 6626 7 3 2 67540 77565
0 6627 5 1 1 89971
0 6628 7 2 2 76552 87031
0 6629 5 1 1 89974
0 6630 7 1 2 89283 6629
0 6631 5 1 1 6630
0 6632 7 1 2 82314 6631
0 6633 5 1 1 6632
0 6634 7 1 2 89972 6633
0 6635 7 1 2 6625 6634
0 6636 5 1 1 6635
0 6637 7 1 2 88499 6636
0 6638 7 1 2 6613 6637
0 6639 5 1 1 6638
0 6640 7 1 2 6591 6639
0 6641 5 1 1 6640
0 6642 7 1 2 78198 6641
0 6643 5 1 1 6642
0 6644 7 1 2 88500 89601
0 6645 5 1 1 6644
0 6646 7 1 2 89796 6645
0 6647 5 2 1 6646
0 6648 7 1 2 72951 89976
0 6649 5 1 1 6648
0 6650 7 13 2 67052 77496
0 6651 5 5 1 89978
0 6652 7 1 2 89979 3968
0 6653 5 1 1 6652
0 6654 7 1 2 6649 6653
0 6655 5 1 1 6654
0 6656 7 1 2 70100 6655
0 6657 5 1 1 6656
0 6658 7 3 2 74841 88105
0 6659 5 1 1 89996
0 6660 7 1 2 72952 89997
0 6661 5 1 1 6660
0 6662 7 1 2 6657 6661
0 6663 5 1 1 6662
0 6664 7 1 2 76285 6663
0 6665 5 1 1 6664
0 6666 7 1 2 70101 89977
0 6667 5 1 1 6666
0 6668 7 2 2 79323 89782
0 6669 5 1 1 89999
0 6670 7 1 2 6667 6669
0 6671 5 1 1 6670
0 6672 7 1 2 76021 6671
0 6673 5 1 1 6672
0 6674 7 1 2 6665 6673
0 6675 5 1 1 6674
0 6676 7 1 2 71572 6675
0 6677 5 1 1 6676
0 6678 7 2 2 75117 74937
0 6679 7 4 2 80336 79801
0 6680 5 4 1 90003
0 6681 7 1 2 74610 90007
0 6682 5 1 1 6681
0 6683 7 1 2 85620 6682
0 6684 5 1 1 6683
0 6685 7 1 2 90001 6684
0 6686 5 1 1 6685
0 6687 7 1 2 74842 84126
0 6688 5 2 1 6687
0 6689 7 1 2 372 90011
0 6690 5 1 1 6689
0 6691 7 1 2 64989 6690
0 6692 5 1 1 6691
0 6693 7 4 2 65315 79569
0 6694 5 3 1 90013
0 6695 7 1 2 79064 74843
0 6696 5 2 1 6695
0 6697 7 1 2 90017 90020
0 6698 7 1 2 6692 6697
0 6699 5 1 1 6698
0 6700 7 1 2 67927 6699
0 6701 5 1 1 6700
0 6702 7 1 2 76286 74812
0 6703 5 1 1 6702
0 6704 7 1 2 6701 6703
0 6705 5 1 1 6704
0 6706 7 1 2 71761 6705
0 6707 5 1 1 6706
0 6708 7 1 2 6686 6707
0 6709 5 1 1 6708
0 6710 7 1 2 88106 6709
0 6711 5 1 1 6710
0 6712 7 1 2 84815 89681
0 6713 5 2 1 6712
0 6714 7 1 2 89797 90022
0 6715 5 1 1 6714
0 6716 7 1 2 83241 6715
0 6717 5 1 1 6716
0 6718 7 10 2 68947 66182
0 6719 7 1 2 89387 90024
0 6720 7 1 2 86181 6719
0 6721 5 1 1 6720
0 6722 7 1 2 6717 6721
0 6723 5 1 1 6722
0 6724 7 1 2 68300 6723
0 6725 5 1 1 6724
0 6726 7 4 2 74998 79179
0 6727 5 12 1 90034
0 6728 7 5 2 63865 81696
0 6729 7 3 2 74281 90050
0 6730 5 1 1 90055
0 6731 7 1 2 90038 90056
0 6732 5 1 1 6731
0 6733 7 1 2 6725 6732
0 6734 5 1 1 6733
0 6735 7 1 2 75338 6734
0 6736 5 1 1 6735
0 6737 7 3 2 74938 88501
0 6738 5 1 1 90058
0 6739 7 1 2 3655 90059
0 6740 5 1 1 6739
0 6741 7 1 2 72557 6740
0 6742 7 1 2 6736 6741
0 6743 7 1 2 6711 6742
0 6744 7 1 2 6677 6743
0 6745 5 1 1 6744
0 6746 7 27 2 68774 75724
0 6747 7 5 2 73681 78682
0 6748 7 2 2 86208 89980
0 6749 7 1 2 90088 90093
0 6750 5 1 1 6749
0 6751 7 5 2 72953 80390
0 6752 5 2 1 90095
0 6753 7 6 2 66664 78568
0 6754 5 9 1 90102
0 6755 7 1 2 67928 90108
0 6756 5 4 1 6755
0 6757 7 4 2 90100 90117
0 6758 5 1 1 90121
0 6759 7 1 2 90122 88502
0 6760 5 1 1 6759
0 6761 7 1 2 83175 5201
0 6762 5 1 1 6761
0 6763 7 1 2 88107 6762
0 6764 5 1 1 6763
0 6765 7 1 2 65316 6764
0 6766 7 1 2 6760 6765
0 6767 5 1 1 6766
0 6768 7 6 2 72954 88503
0 6769 7 1 2 68591 90125
0 6770 5 1 1 6769
0 6771 7 1 2 89367 6770
0 6772 5 1 1 6771
0 6773 7 1 2 66665 6772
0 6774 5 1 1 6773
0 6775 7 1 2 75339 85587
0 6776 5 1 1 6775
0 6777 7 1 2 88108 6776
0 6778 5 1 1 6777
0 6779 7 2 2 71762 82042
0 6780 7 2 2 74873 88504
0 6781 5 1 1 90133
0 6782 7 1 2 90131 90134
0 6783 5 1 1 6782
0 6784 7 1 2 70373 6783
0 6785 7 1 2 6778 6784
0 6786 7 1 2 6774 6785
0 6787 5 1 1 6786
0 6788 7 1 2 6767 6787
0 6789 5 1 1 6788
0 6790 7 1 2 82957 89340
0 6791 5 1 1 6790
0 6792 7 1 2 6789 6791
0 6793 5 1 1 6792
0 6794 7 1 2 64619 6793
0 6795 5 1 1 6794
0 6796 7 1 2 6750 6795
0 6797 5 1 1 6796
0 6798 7 1 2 66183 6797
0 6799 5 1 1 6798
0 6800 7 1 2 84802 86190
0 6801 5 1 1 6800
0 6802 7 2 2 67053 6801
0 6803 7 1 2 63866 90135
0 6804 5 1 1 6803
0 6805 7 1 2 6349 6804
0 6806 5 1 1 6805
0 6807 7 1 2 79952 6806
0 6808 5 1 1 6807
0 6809 7 1 2 81697 78569
0 6810 7 3 2 88109 6809
0 6811 5 1 1 90137
0 6812 7 1 2 78903 90138
0 6813 5 1 1 6812
0 6814 7 4 2 82893 76408
0 6815 5 1 1 90140
0 6816 7 1 2 90141 89364
0 6817 5 1 1 6816
0 6818 7 1 2 88813 89715
0 6819 5 1 1 6818
0 6820 7 1 2 6817 6819
0 6821 5 1 1 6820
0 6822 7 1 2 72955 6821
0 6823 5 1 1 6822
0 6824 7 1 2 6813 6823
0 6825 7 1 2 6808 6824
0 6826 5 1 1 6825
0 6827 7 1 2 74611 6826
0 6828 5 1 1 6827
0 6829 7 1 2 75256 88805
0 6830 5 1 1 6829
0 6831 7 1 2 82043 86884
0 6832 5 1 1 6831
0 6833 7 1 2 6830 6832
0 6834 5 1 1 6833
0 6835 7 1 2 88110 6834
0 6836 5 1 1 6835
0 6837 7 5 2 66465 72109
0 6838 7 3 2 77818 90144
0 6839 5 1 1 90149
0 6840 7 1 2 85777 90150
0 6841 5 1 1 6840
0 6842 7 1 2 6836 6841
0 6843 5 1 1 6842
0 6844 7 1 2 76553 6843
0 6845 5 1 1 6844
0 6846 7 1 2 85580 86887
0 6847 5 2 1 6846
0 6848 7 1 2 90152 88111
0 6849 5 1 1 6848
0 6850 7 2 2 73367 84702
0 6851 7 2 2 74218 75998
0 6852 7 1 2 90154 90156
0 6853 5 1 1 6852
0 6854 7 1 2 6849 6853
0 6855 5 1 1 6854
0 6856 7 1 2 83359 6855
0 6857 5 1 1 6856
0 6858 7 1 2 67541 6857
0 6859 7 1 2 6845 6858
0 6860 7 1 2 6828 6859
0 6861 7 1 2 6799 6860
0 6862 5 1 1 6861
0 6863 7 1 2 90061 6862
0 6864 7 1 2 6745 6863
0 6865 5 1 1 6864
0 6866 7 1 2 6643 6865
0 6867 5 1 1 6866
0 6868 7 1 2 65927 6867
0 6869 5 1 1 6868
0 6870 7 1 2 89904 87686
0 6871 5 1 1 6870
0 6872 7 2 2 87695 80157
0 6873 5 2 1 90158
0 6874 7 1 2 80172 90160
0 6875 5 2 1 6874
0 6876 7 1 2 67542 89469
0 6877 7 1 2 90162 6876
0 6878 5 1 1 6877
0 6879 7 1 2 6079 6878
0 6880 5 1 1 6879
0 6881 7 1 2 78199 6880
0 6882 5 1 1 6881
0 6883 7 1 2 6871 6882
0 6884 5 1 1 6883
0 6885 7 1 2 65928 6884
0 6886 5 1 1 6885
0 6887 7 1 2 78817 89936
0 6888 5 1 1 6887
0 6889 7 3 2 87400 81666
0 6890 7 1 2 90164 87977
0 6891 5 1 1 6890
0 6892 7 1 2 6888 6891
0 6893 5 1 1 6892
0 6894 7 1 2 78402 6893
0 6895 5 1 1 6894
0 6896 7 1 2 6886 6895
0 6897 5 1 1 6896
0 6898 7 1 2 80675 6897
0 6899 5 1 1 6898
0 6900 7 10 2 72110 77819
0 6901 5 3 1 90167
0 6902 7 1 2 88286 90177
0 6903 5 4 1 6902
0 6904 7 11 2 73682 77651
0 6905 7 1 2 66943 90184
0 6906 7 3 2 90180 6905
0 6907 7 2 2 67543 86393
0 6908 7 2 2 90195 90198
0 6909 7 3 2 68775 76705
0 6910 7 1 2 88321 90202
0 6911 7 1 2 90200 6910
0 6912 5 1 1 6911
0 6913 7 1 2 6899 6912
0 6914 7 1 2 6869 6913
0 6915 5 1 1 6914
0 6916 7 1 2 64289 6915
0 6917 5 1 1 6916
0 6918 7 2 2 68776 66466
0 6919 7 1 2 90205 87991
0 6920 7 1 2 88009 6919
0 6921 7 1 2 90201 6920
0 6922 5 1 1 6921
0 6923 7 1 2 6917 6922
0 6924 7 1 2 6550 6923
0 6925 5 1 1 6924
0 6926 7 1 2 89560 6925
0 6927 5 1 1 6926
0 6928 7 1 2 6108 6927
0 6929 7 1 2 5630 6928
0 6930 7 1 2 5041 6929
0 6931 5 1 1 6930
0 6932 7 1 2 85480 6931
0 6933 5 1 1 6932
0 6934 7 8 2 85200 88938
0 6935 7 6 2 69399 77652
0 6936 5 2 1 90215
0 6937 7 2 2 83893 82786
0 6938 5 1 1 90223
0 6939 7 1 2 90221 6938
0 6940 5 1 1 6939
0 6941 7 1 2 71763 6940
0 6942 5 1 1 6941
0 6943 7 3 2 69400 79716
0 6944 5 1 1 90225
0 6945 7 1 2 73368 90226
0 6946 5 1 1 6945
0 6947 7 1 2 75548 83630
0 6948 5 1 1 6947
0 6949 7 1 2 6946 6948
0 6950 7 1 2 6942 6949
0 6951 5 1 1 6950
0 6952 7 1 2 88112 6951
0 6953 5 1 1 6952
0 6954 7 1 2 89716 82688
0 6955 5 1 1 6954
0 6956 7 1 2 6953 6955
0 6957 5 1 1 6956
0 6958 7 1 2 70102 6957
0 6959 5 1 1 6958
0 6960 7 7 2 64290 71764
0 6961 7 1 2 76820 90228
0 6962 5 1 1 6961
0 6963 7 1 2 81230 83170
0 6964 5 1 1 6963
0 6965 7 1 2 6962 6964
0 6966 5 1 1 6965
0 6967 7 1 2 71573 6966
0 6968 5 1 1 6967
0 6969 7 1 2 69401 74612
0 6970 7 1 2 74771 6969
0 6971 5 1 1 6970
0 6972 7 1 2 6968 6971
0 6973 5 1 1 6972
0 6974 7 1 2 88113 6973
0 6975 5 1 1 6974
0 6976 7 1 2 6959 6975
0 6977 5 1 1 6976
0 6978 7 1 2 67544 6977
0 6979 5 1 1 6978
0 6980 7 3 2 74515 81458
0 6981 5 1 1 90235
0 6982 7 1 2 90236 88114
0 6983 7 1 2 76751 6982
0 6984 5 1 1 6983
0 6985 7 1 2 6979 6984
0 6986 5 1 1 6985
0 6987 7 1 2 64620 6986
0 6988 5 1 1 6987
0 6989 7 2 2 74728 84181
0 6990 7 2 2 67054 90238
0 6991 7 3 2 64291 74516
0 6992 5 1 1 90242
0 6993 7 1 2 90243 84639
0 6994 7 1 2 90240 6993
0 6995 5 1 1 6994
0 6996 7 1 2 6988 6995
0 6997 5 1 1 6996
0 6998 7 1 2 74142 6997
0 6999 5 1 1 6998
0 7000 7 2 2 74282 84640
0 7001 5 1 1 90245
0 7002 7 1 2 87008 78373
0 7003 7 1 2 82086 7002
0 7004 7 1 2 90246 7003
0 7005 5 1 1 7004
0 7006 7 1 2 6999 7005
0 7007 5 1 1 7006
0 7008 7 1 2 90207 7007
0 7009 5 1 1 7008
0 7010 7 8 2 70653 89502
0 7011 7 2 2 66944 76975
0 7012 5 1 1 90255
0 7013 7 1 2 78795 74465
0 7014 5 1 1 7013
0 7015 7 1 2 7012 7014
0 7016 5 1 1 7015
0 7017 7 1 2 88115 7016
0 7018 5 1 1 7017
0 7019 7 3 2 71574 77820
0 7020 7 4 2 73683 75815
0 7021 7 1 2 75590 90260
0 7022 7 1 2 90257 7021
0 7023 5 1 1 7022
0 7024 7 1 2 7018 7023
0 7025 5 1 1 7024
0 7026 7 1 2 69734 7025
0 7027 5 1 1 7026
0 7028 7 9 2 63867 71283
0 7029 7 2 2 83951 90264
0 7030 7 1 2 82818 90273
0 7031 5 1 1 7030
0 7032 7 1 2 7027 7031
0 7033 5 1 1 7032
0 7034 7 1 2 72956 7033
0 7035 5 1 1 7034
0 7036 7 2 2 82819 88116
0 7037 7 1 2 83628 90275
0 7038 5 1 1 7037
0 7039 7 1 2 7035 7038
0 7040 5 1 1 7039
0 7041 7 1 2 90247 7040
0 7042 5 1 1 7041
0 7043 7 2 2 72957 77916
0 7044 5 1 1 90277
0 7045 7 1 2 2584 7044
0 7046 5 1 1 7045
0 7047 7 2 2 74096 7046
0 7048 7 12 2 63868 63954
0 7049 7 4 2 65673 90281
0 7050 7 2 2 70613 90293
0 7051 5 1 1 90297
0 7052 7 1 2 65621 90298
0 7053 7 1 2 90279 7052
0 7054 5 1 1 7053
0 7055 7 1 2 7042 7054
0 7056 5 1 1 7055
0 7057 7 1 2 68777 7056
0 7058 5 1 1 7057
0 7059 7 2 2 82755 88039
0 7060 7 5 2 70704 90299
0 7061 7 1 2 90301 90280
0 7062 5 1 1 7061
0 7063 7 1 2 7058 7062
0 7064 5 1 1 7063
0 7065 7 1 2 71903 7064
0 7066 5 1 1 7065
0 7067 7 4 2 63955 65622
0 7068 5 1 1 90306
0 7069 7 14 2 65674 90307
0 7070 7 7 2 73998 90310
0 7071 5 1 1 90324
0 7072 7 1 2 63739 89561
0 7073 5 1 1 7072
0 7074 7 1 2 7071 7073
0 7075 5 12 1 7074
0 7076 7 13 2 66837 90331
0 7077 7 1 2 76554 89388
0 7078 7 1 2 74296 7077
0 7079 7 1 2 90343 7078
0 7080 5 1 1 7079
0 7081 7 1 2 7066 7080
0 7082 5 1 1 7081
0 7083 7 1 2 70986 7082
0 7084 5 1 1 7083
0 7085 7 3 2 79463 82722
0 7086 5 3 1 90356
0 7087 7 7 2 63740 70654
0 7088 7 7 2 69043 70614
0 7089 7 3 2 70705 90369
0 7090 7 6 2 90362 90376
0 7091 5 1 1 90379
0 7092 7 2 2 68778 89562
0 7093 5 1 1 90385
0 7094 7 1 2 7091 7093
0 7095 5 13 1 7094
0 7096 7 2 2 68592 75725
0 7097 7 8 2 72111 87595
0 7098 5 2 1 90402
0 7099 7 1 2 90410 89764
0 7100 5 2 1 7099
0 7101 7 1 2 90400 90412
0 7102 7 1 2 90387 7101
0 7103 5 1 1 7102
0 7104 7 8 2 65579 89532
0 7105 7 7 2 68948 63956
0 7106 7 3 2 68779 90422
0 7107 7 4 2 90414 90429
0 7108 5 1 1 90432
0 7109 7 4 2 75830 90433
0 7110 5 2 1 90436
0 7111 7 8 2 72010 89563
0 7112 7 2 2 79360 77767
0 7113 7 1 2 90442 90450
0 7114 5 1 1 7113
0 7115 7 1 2 90440 7114
0 7116 7 1 2 7103 7115
0 7117 5 1 1 7116
0 7118 7 1 2 90357 7117
0 7119 5 1 1 7118
0 7120 7 1 2 7084 7119
0 7121 5 1 1 7120
0 7122 7 1 2 84658 7121
0 7123 5 1 1 7122
0 7124 7 3 2 70103 81459
0 7125 5 1 1 90452
0 7126 7 4 2 64621 86335
0 7127 5 1 1 90455
0 7128 7 1 2 82212 90456
0 7129 5 1 1 7128
0 7130 7 1 2 7125 7129
0 7131 5 1 1 7130
0 7132 7 1 2 66184 7131
0 7133 5 1 1 7132
0 7134 7 2 2 71765 83985
0 7135 5 1 1 90459
0 7136 7 1 2 83856 90460
0 7137 5 1 1 7136
0 7138 7 1 2 7133 7137
0 7139 5 1 1 7138
0 7140 7 1 2 88117 7139
0 7141 5 1 1 7140
0 7142 7 6 2 70104 82958
0 7143 5 18 1 90461
0 7144 7 1 2 80471 90467
0 7145 5 1 1 7144
0 7146 7 11 2 72112 83616
0 7147 7 1 2 87774 90485
0 7148 7 1 2 7145 7147
0 7149 5 1 1 7148
0 7150 7 1 2 7141 7149
0 7151 5 1 1 7150
0 7152 7 1 2 67929 7151
0 7153 5 1 1 7152
0 7154 7 1 2 83344 89231
0 7155 7 1 2 89875 7154
0 7156 5 1 1 7155
0 7157 7 1 2 7153 7156
0 7158 5 2 1 7157
0 7159 7 1 2 66945 89564
0 7160 7 1 2 90496 7159
0 7161 5 1 1 7160
0 7162 7 3 2 75340 82801
0 7163 7 4 2 67930 79271
0 7164 7 1 2 90498 90501
0 7165 5 1 1 7164
0 7166 7 1 2 79165 75618
0 7167 7 1 2 3766 7166
0 7168 5 1 1 7167
0 7169 7 1 2 7165 7168
0 7170 5 1 1 7169
0 7171 7 1 2 88118 7170
0 7172 5 1 1 7171
0 7173 7 1 2 86840 86594
0 7174 7 1 2 90486 7173
0 7175 5 1 1 7174
0 7176 7 1 2 7172 7175
0 7177 5 1 1 7176
0 7178 7 3 2 71284 72011
0 7179 7 2 2 72558 90505
0 7180 7 9 2 70615 70706
0 7181 7 8 2 69044 70655
0 7182 7 10 2 90510 90519
0 7183 7 1 2 90508 90527
0 7184 7 1 2 7177 7183
0 7185 5 1 1 7184
0 7186 7 1 2 7161 7185
0 7187 5 1 1 7186
0 7188 7 1 2 71904 7187
0 7189 5 1 1 7188
0 7190 7 5 2 67055 84641
0 7191 7 1 2 75341 90537
0 7192 5 1 1 7191
0 7193 7 5 2 72113 82959
0 7194 5 1 1 90542
0 7195 7 1 2 68949 90543
0 7196 7 1 2 78782 7195
0 7197 5 1 1 7196
0 7198 7 1 2 7192 7197
0 7199 5 1 1 7198
0 7200 7 1 2 81231 7199
0 7201 5 1 1 7200
0 7202 7 8 2 67931 88505
0 7203 5 1 1 90547
0 7204 7 2 2 71575 83180
0 7205 5 1 1 90555
0 7206 7 1 2 76448 7205
0 7207 7 1 2 90548 7206
0 7208 5 1 1 7207
0 7209 7 1 2 7201 7208
0 7210 5 1 1 7209
0 7211 7 1 2 72559 7210
0 7212 5 1 1 7211
0 7213 7 1 2 67932 5324
0 7214 5 1 1 7213
0 7215 7 2 2 72958 78838
0 7216 5 1 1 90557
0 7217 7 3 2 67545 88506
0 7218 7 1 2 7216 90559
0 7219 7 1 2 7214 7218
0 7220 5 1 1 7219
0 7221 7 1 2 7212 7220
0 7222 5 2 1 7221
0 7223 7 2 2 90311 85789
0 7224 7 1 2 90562 90564
0 7225 5 1 1 7224
0 7226 7 1 2 68780 7225
0 7227 7 1 2 7189 7226
0 7228 5 1 1 7227
0 7229 7 1 2 90443 90563
0 7230 5 1 1 7229
0 7231 7 4 2 75342 88507
0 7232 5 1 1 90566
0 7233 7 1 2 89765 7232
0 7234 5 1 1 7233
0 7235 7 25 2 65580 65623
0 7236 7 6 2 63957 69402
0 7237 7 2 2 90570 90595
0 7238 7 6 2 65675 66946
0 7239 7 2 2 72560 90603
0 7240 7 1 2 90601 90609
0 7241 7 1 2 7234 7240
0 7242 5 1 1 7241
0 7243 7 1 2 7230 7242
0 7244 5 1 1 7243
0 7245 7 1 2 66838 7244
0 7246 5 1 1 7245
0 7247 7 2 2 66947 88057
0 7248 7 1 2 90611 90497
0 7249 5 1 1 7248
0 7250 7 1 2 63741 7249
0 7251 7 1 2 7246 7250
0 7252 5 1 1 7251
0 7253 7 1 2 70987 7252
0 7254 7 1 2 7228 7253
0 7255 5 1 1 7254
0 7256 7 4 2 63869 75530
0 7257 5 2 1 90613
0 7258 7 1 2 75343 89769
0 7259 5 1 1 7258
0 7260 7 1 2 90617 7259
0 7261 5 1 1 7260
0 7262 7 2 2 68781 66185
0 7263 7 1 2 90619 87580
0 7264 7 1 2 7261 7263
0 7265 5 1 1 7264
0 7266 7 1 2 6161 7265
0 7267 5 1 1 7266
0 7268 7 1 2 67933 7267
0 7269 5 1 1 7268
0 7270 7 5 2 79361 76374
0 7271 7 5 2 72114 90621
0 7272 5 2 1 90626
0 7273 7 3 2 63870 71576
0 7274 7 6 2 67056 90633
0 7275 5 1 1 90636
0 7276 7 1 2 90062 90637
0 7277 5 1 1 7276
0 7278 7 1 2 90631 7277
0 7279 5 1 1 7278
0 7280 7 1 2 83255 7279
0 7281 5 1 1 7280
0 7282 7 1 2 7269 7281
0 7283 5 1 1 7282
0 7284 7 1 2 65929 7283
0 7285 5 1 1 7284
0 7286 7 2 2 77508 84375
0 7287 7 8 2 63742 70105
0 7288 7 4 2 76375 90644
0 7289 7 1 2 76191 90652
0 7290 7 1 2 90642 7289
0 7291 5 1 1 7290
0 7292 7 1 2 7285 7291
0 7293 5 1 1 7292
0 7294 7 1 2 69403 7293
0 7295 5 1 1 7294
0 7296 7 4 2 66467 66839
0 7297 7 6 2 72012 90656
0 7298 7 1 2 79362 89389
0 7299 7 1 2 83857 7298
0 7300 7 1 2 90660 7299
0 7301 5 1 1 7300
0 7302 7 1 2 7295 7301
0 7303 5 1 1 7302
0 7304 7 1 2 89565 7303
0 7305 5 1 1 7304
0 7306 7 2 2 87401 80982
0 7307 7 1 2 75816 90666
0 7308 5 1 1 7307
0 7309 7 4 2 63743 84044
0 7310 7 3 2 67057 74613
0 7311 7 4 2 63871 90672
0 7312 5 1 1 90675
0 7313 7 1 2 90668 90676
0 7314 5 1 1 7313
0 7315 7 1 2 7308 7314
0 7316 5 1 1 7315
0 7317 7 1 2 69735 7316
0 7318 5 1 1 7317
0 7319 7 1 2 79483 82021
0 7320 5 2 1 7319
0 7321 7 4 2 68782 89118
0 7322 7 1 2 75817 90681
0 7323 7 1 2 90679 7322
0 7324 5 1 1 7323
0 7325 7 1 2 7318 7324
0 7326 5 1 1 7325
0 7327 7 1 2 72959 7326
0 7328 5 1 1 7327
0 7329 7 1 2 64292 80134
0 7330 5 1 1 7329
0 7331 7 1 2 81980 7330
0 7332 5 1 1 7331
0 7333 7 1 2 89401 7332
0 7334 5 1 1 7333
0 7335 7 1 2 7328 7334
0 7336 5 1 1 7335
0 7337 7 1 2 88939 7336
0 7338 5 1 1 7337
0 7339 7 2 2 80983 88058
0 7340 7 10 2 72013 86488
0 7341 7 8 2 71577 80337
0 7342 5 1 1 90697
0 7343 7 1 2 90687 90698
0 7344 5 1 1 7343
0 7345 7 1 2 85353 3509
0 7346 5 7 1 7345
0 7347 7 12 2 68783 69736
0 7348 5 1 1 90712
0 7349 7 1 2 7348 6524
0 7350 7 1 2 80497 7349
0 7351 7 1 2 90705 7350
0 7352 5 1 1 7351
0 7353 7 1 2 7344 7352
0 7354 5 1 1 7353
0 7355 7 1 2 76022 7354
0 7356 5 1 1 7355
0 7357 7 1 2 77917 89414
0 7358 5 1 1 7357
0 7359 7 1 2 7356 7358
0 7360 5 1 1 7359
0 7361 7 1 2 88119 7360
0 7362 5 1 1 7361
0 7363 7 2 2 85201 75344
0 7364 5 2 1 90724
0 7365 7 5 2 68784 79048
0 7366 7 1 2 74517 90728
0 7367 5 1 1 7366
0 7368 7 1 2 90726 7367
0 7369 5 4 1 7368
0 7370 7 4 2 68950 89390
0 7371 7 1 2 84089 90737
0 7372 7 1 2 90733 7371
0 7373 5 1 1 7372
0 7374 7 1 2 7362 7373
0 7375 5 1 1 7374
0 7376 7 1 2 90685 7375
0 7377 5 1 1 7376
0 7378 7 1 2 7338 7377
0 7379 7 1 2 7305 7378
0 7380 5 1 1 7379
0 7381 7 1 2 67546 7380
0 7382 5 1 1 7381
0 7383 7 8 2 63958 90571
0 7384 7 8 2 90741 90604
0 7385 7 4 2 71766 76449
0 7386 5 1 1 90757
0 7387 7 1 2 67934 88315
0 7388 5 1 1 7387
0 7389 7 1 2 7386 7388
0 7390 5 1 1 7389
0 7391 7 1 2 72561 7390
0 7392 5 1 1 7391
0 7393 7 1 2 85059 7392
0 7394 5 1 1 7393
0 7395 7 1 2 88120 7394
0 7396 5 1 1 7395
0 7397 7 6 2 66186 87784
0 7398 5 9 1 90761
0 7399 7 1 2 72562 80173
0 7400 5 1 1 7399
0 7401 7 1 2 90767 7400
0 7402 5 3 1 7401
0 7403 7 1 2 90567 90776
0 7404 5 1 1 7403
0 7405 7 1 2 7396 7404
0 7406 5 1 1 7405
0 7407 7 1 2 90749 7406
0 7408 5 1 1 7407
0 7409 7 2 2 72115 83876
0 7410 5 1 1 90779
0 7411 7 1 2 89887 7410
0 7412 5 1 1 7411
0 7413 7 1 2 71767 7412
0 7414 5 1 1 7413
0 7415 7 1 2 89669 83877
0 7416 5 1 1 7415
0 7417 7 1 2 7414 7416
0 7418 5 1 1 7417
0 7419 7 1 2 81960 74207
0 7420 7 2 2 7418 7419
0 7421 7 1 2 69737 89566
0 7422 7 1 2 90781 7421
0 7423 5 1 1 7422
0 7424 7 1 2 7408 7423
0 7425 5 1 1 7424
0 7426 7 1 2 63744 7425
0 7427 5 1 1 7426
0 7428 7 10 2 90572 88909
0 7429 7 2 2 90713 90783
0 7430 7 1 2 90782 90793
0 7431 5 1 1 7430
0 7432 7 1 2 7427 7431
0 7433 5 1 1 7432
0 7434 7 1 2 66840 7433
0 7435 5 1 1 7434
0 7436 7 2 2 78339 74097
0 7437 7 3 2 76450 75798
0 7438 7 2 2 73684 84991
0 7439 7 1 2 90797 90800
0 7440 7 1 2 90795 7439
0 7441 7 1 2 90388 7440
0 7442 5 1 1 7441
0 7443 7 1 2 7435 7442
0 7444 5 1 1 7443
0 7445 7 1 2 77405 7444
0 7446 5 1 1 7445
0 7447 7 1 2 7382 7446
0 7448 7 1 2 7255 7447
0 7449 7 1 2 7123 7448
0 7450 5 1 1 7449
0 7451 7 1 2 68301 7450
0 7452 5 1 1 7451
0 7453 7 2 2 78455 88508
0 7454 7 1 2 80071 90802
0 7455 5 1 1 7454
0 7456 7 1 2 84108 83945
0 7457 5 18 1 7456
0 7458 7 7 2 66468 68593
0 7459 5 1 1 90822
0 7460 7 1 2 90823 88121
0 7461 7 1 2 90804 7460
0 7462 5 1 1 7461
0 7463 7 1 2 7455 7462
0 7464 5 1 1 7463
0 7465 7 1 2 67935 7464
0 7466 5 1 1 7465
0 7467 7 1 2 90803 90278
0 7468 5 1 1 7467
0 7469 7 1 2 7466 7468
0 7470 5 1 1 7469
0 7471 7 1 2 85202 7470
0 7472 5 1 1 7471
0 7473 7 4 2 76451 78403
0 7474 5 2 1 90829
0 7475 7 3 2 65930 84182
0 7476 5 2 1 90835
0 7477 7 1 2 71578 90836
0 7478 5 1 1 7477
0 7479 7 1 2 90833 7478
0 7480 5 1 1 7479
0 7481 7 1 2 83242 7480
0 7482 5 1 1 7481
0 7483 7 3 2 80072 83894
0 7484 5 1 1 90840
0 7485 7 1 2 83742 90841
0 7486 5 1 1 7485
0 7487 7 1 2 7482 7486
0 7488 5 1 1 7487
0 7489 7 1 2 89184 7488
0 7490 5 1 1 7489
0 7491 7 1 2 7472 7490
0 7492 5 1 1 7491
0 7493 7 1 2 69404 7492
0 7494 5 1 1 7493
0 7495 7 4 2 83895 88122
0 7496 5 1 1 90843
0 7497 7 5 2 72563 85203
0 7498 7 1 2 90847 80135
0 7499 7 1 2 90844 7498
0 7500 5 1 1 7499
0 7501 7 1 2 68594 89185
0 7502 5 1 1 7501
0 7503 7 1 2 89319 7502
0 7504 5 1 1 7503
0 7505 7 1 2 64293 82213
0 7506 7 1 2 83256 7505
0 7507 7 1 2 7504 7506
0 7508 5 1 1 7507
0 7509 7 1 2 7500 7508
0 7510 5 1 1 7509
0 7511 7 1 2 70988 7510
0 7512 5 1 1 7511
0 7513 7 1 2 7494 7512
0 7514 5 1 1 7513
0 7515 7 1 2 70106 7514
0 7516 5 1 1 7515
0 7517 7 2 2 86360 80962
0 7518 5 2 1 90852
0 7519 7 2 2 67936 89299
0 7520 7 1 2 84659 90856
0 7521 7 1 2 90854 7520
0 7522 5 1 1 7521
0 7523 7 12 2 69405 67547
0 7524 5 1 1 90858
0 7525 7 1 2 7524 87492
0 7526 7 2 2 69738 87724
0 7527 7 1 2 80886 2945
0 7528 5 1 1 7527
0 7529 7 1 2 90870 7528
0 7530 7 1 2 7525 7529
0 7531 5 1 1 7530
0 7532 7 1 2 7522 7531
0 7533 5 1 1 7532
0 7534 7 1 2 71285 7533
0 7535 5 1 1 7534
0 7536 7 6 2 64622 75902
0 7537 5 5 1 90872
0 7538 7 2 2 74614 79953
0 7539 7 1 2 75478 90883
0 7540 5 1 1 7539
0 7541 7 1 2 90878 7540
0 7542 5 1 1 7541
0 7543 7 3 2 68951 67548
0 7544 7 12 2 63745 69406
0 7545 7 1 2 90888 74232
0 7546 7 2 2 90885 7545
0 7547 7 1 2 7542 90900
0 7548 5 1 1 7547
0 7549 7 1 2 7535 7548
0 7550 5 1 1 7549
0 7551 7 1 2 70989 7550
0 7552 5 1 1 7551
0 7553 7 1 2 84394 90901
0 7554 7 1 2 90855 7553
0 7555 5 1 1 7554
0 7556 7 1 2 7552 7555
0 7557 7 1 2 7516 7556
0 7558 5 1 1 7557
0 7559 7 1 2 88059 7558
0 7560 5 1 1 7559
0 7561 7 13 2 76376 90325
0 7562 5 2 1 90902
0 7563 7 3 2 64623 76067
0 7564 5 7 1 90917
0 7565 7 1 2 90920 219
0 7566 5 1 1 7565
0 7567 7 2 2 81568 7566
0 7568 7 1 2 67549 90927
0 7569 5 1 1 7568
0 7570 7 7 2 72564 74518
0 7571 7 5 2 64294 74999
0 7572 5 3 1 90936
0 7573 7 2 2 79180 90937
0 7574 5 1 1 90944
0 7575 7 1 2 90929 7574
0 7576 5 1 1 7575
0 7577 7 1 2 7569 7576
0 7578 5 1 1 7577
0 7579 7 1 2 88123 7578
0 7580 5 1 1 7579
0 7581 7 1 2 88509 81561
0 7582 5 1 1 7581
0 7583 7 1 2 7580 7582
0 7584 5 1 1 7583
0 7585 7 1 2 70990 7584
0 7586 5 1 1 7585
0 7587 7 1 2 82052 89682
0 7588 5 1 1 7587
0 7589 7 1 2 83858 88124
0 7590 5 1 1 7589
0 7591 7 1 2 7588 7590
0 7592 5 1 1 7591
0 7593 7 1 2 67550 7592
0 7594 5 1 1 7593
0 7595 7 2 2 77918 88125
0 7596 5 1 1 90946
0 7597 7 6 2 68952 69739
0 7598 7 4 2 72116 90948
0 7599 7 1 2 71286 90954
0 7600 5 1 1 7599
0 7601 7 1 2 7596 7600
0 7602 5 1 1 7601
0 7603 7 1 2 70107 7602
0 7604 5 1 1 7603
0 7605 7 3 2 71579 72117
0 7606 7 6 2 68953 90958
0 7607 5 2 1 90961
0 7608 7 1 2 76452 90962
0 7609 5 1 1 7608
0 7610 7 1 2 7604 7609
0 7611 5 1 1 7610
0 7612 7 1 2 81460 7611
0 7613 5 1 1 7612
0 7614 7 1 2 7594 7613
0 7615 5 1 1 7614
0 7616 7 1 2 67937 7615
0 7617 5 1 1 7616
0 7618 7 1 2 81461 83952
0 7619 7 1 2 90798 7618
0 7620 5 1 1 7619
0 7621 7 1 2 7617 7620
0 7622 7 1 2 7586 7621
0 7623 5 1 1 7622
0 7624 7 1 2 90903 7623
0 7625 5 1 1 7624
0 7626 7 1 2 7560 7625
0 7627 5 1 1 7626
0 7628 7 1 2 73369 7627
0 7629 5 1 1 7628
0 7630 7 2 2 80846 90805
0 7631 5 1 1 90969
0 7632 7 1 2 89479 90970
0 7633 5 1 1 7632
0 7634 7 1 2 79954 78470
0 7635 5 1 1 7634
0 7636 7 1 2 74939 83743
0 7637 5 1 1 7636
0 7638 7 1 2 7635 7637
0 7639 5 1 1 7638
0 7640 7 1 2 80864 88510
0 7641 7 1 2 7639 7640
0 7642 5 1 1 7641
0 7643 7 1 2 7633 7642
0 7644 5 1 1 7643
0 7645 7 1 2 66469 7644
0 7646 5 1 1 7645
0 7647 7 1 2 86336 79955
0 7648 5 1 1 7647
0 7649 7 1 2 90879 7648
0 7650 5 1 1 7649
0 7651 7 1 2 78471 7650
0 7652 5 1 1 7651
0 7653 7 1 2 69740 86361
0 7654 5 2 1 7653
0 7655 7 1 2 74940 90971
0 7656 5 1 1 7655
0 7657 7 1 2 2404 7656
0 7658 5 1 1 7657
0 7659 7 1 2 83744 7658
0 7660 5 1 1 7659
0 7661 7 1 2 7652 7660
0 7662 5 1 1 7661
0 7663 7 1 2 88511 7662
0 7664 5 1 1 7663
0 7665 7 1 2 7646 7664
0 7666 5 1 1 7665
0 7667 7 1 2 85115 7666
0 7668 5 1 1 7667
0 7669 7 3 2 69741 83953
0 7670 7 1 2 75799 90973
0 7671 5 2 1 7670
0 7672 7 6 2 72118 75345
0 7673 7 1 2 85401 90978
0 7674 5 1 1 7673
0 7675 7 1 2 90976 7674
0 7676 5 1 1 7675
0 7677 7 1 2 75958 7676
0 7678 5 1 1 7677
0 7679 7 2 2 75800 83954
0 7680 5 1 1 90984
0 7681 7 1 2 75346 90955
0 7682 5 1 1 7681
0 7683 7 1 2 7680 7682
0 7684 5 1 1 7683
0 7685 7 1 2 89450 7684
0 7686 5 1 1 7685
0 7687 7 1 2 7678 7686
0 7688 5 1 1 7687
0 7689 7 1 2 72565 7688
0 7690 5 1 1 7689
0 7691 7 7 2 67551 83896
0 7692 7 1 2 90986 88641
0 7693 5 1 1 7692
0 7694 7 1 2 7690 7693
0 7695 5 1 1 7694
0 7696 7 1 2 78200 7695
0 7697 5 1 1 7696
0 7698 7 1 2 7668 7697
0 7699 5 1 1 7698
0 7700 7 1 2 69407 7699
0 7701 5 1 1 7700
0 7702 7 1 2 67938 90853
0 7703 5 1 1 7702
0 7704 7 1 2 86627 7703
0 7705 5 1 1 7704
0 7706 7 1 2 78769 7705
0 7707 5 1 1 7706
0 7708 7 1 2 84151 89891
0 7709 7 1 2 7707 7708
0 7710 5 1 1 7709
0 7711 7 33 2 63746 76377
0 7712 5 6 1 90993
0 7713 7 10 2 90994 88126
0 7714 5 2 1 91032
0 7715 7 1 2 91033 90928
0 7716 5 1 1 7715
0 7717 7 1 2 67552 7716
0 7718 7 1 2 7710 7717
0 7719 5 1 1 7718
0 7720 7 5 2 74519 75959
0 7721 5 1 1 91044
0 7722 7 1 2 88127 91045
0 7723 5 1 1 7722
0 7724 7 1 2 6738 7723
0 7725 5 1 1 7724
0 7726 7 1 2 79824 7725
0 7727 5 1 1 7726
0 7728 7 1 2 81607 89480
0 7729 5 1 1 7728
0 7730 7 1 2 7727 7729
0 7731 5 1 1 7730
0 7732 7 1 2 78201 7731
0 7733 5 1 1 7732
0 7734 7 5 2 86413 85098
0 7735 7 1 2 77813 91049
0 7736 7 1 2 90845 7735
0 7737 5 1 1 7736
0 7738 7 1 2 72566 7737
0 7739 7 1 2 7733 7738
0 7740 5 1 1 7739
0 7741 7 1 2 70991 7740
0 7742 7 1 2 7719 7741
0 7743 5 1 1 7742
0 7744 7 2 2 79272 85091
0 7745 5 1 1 91054
0 7746 7 1 2 91034 91055
0 7747 5 1 1 7746
0 7748 7 1 2 7743 7747
0 7749 7 1 2 7701 7748
0 7750 5 1 1 7749
0 7751 7 1 2 73370 7750
0 7752 5 1 1 7751
0 7753 7 2 2 67939 80984
0 7754 5 1 1 91056
0 7755 7 4 2 74520 85116
0 7756 5 1 1 91058
0 7757 7 1 2 91059 88512
0 7758 5 1 1 7757
0 7759 7 1 2 91042 7758
0 7760 5 1 1 7759
0 7761 7 1 2 91057 7760
0 7762 5 1 1 7761
0 7763 7 16 2 66948 72960
0 7764 7 2 2 91062 85099
0 7765 7 1 2 91078 89838
0 7766 5 1 1 7765
0 7767 7 3 2 72014 77744
0 7768 7 3 2 84607 91080
0 7769 5 1 1 91083
0 7770 7 1 2 7766 7769
0 7771 5 1 1 7770
0 7772 7 1 2 70992 77117
0 7773 7 1 2 7771 7772
0 7774 5 1 1 7773
0 7775 7 1 2 7762 7774
0 7776 5 1 1 7775
0 7777 7 1 2 72567 7776
0 7778 5 1 1 7777
0 7779 7 3 2 72961 77118
0 7780 5 1 1 91086
0 7781 7 2 2 75726 84616
0 7782 7 1 2 79098 85402
0 7783 7 1 2 91089 7782
0 7784 7 1 2 91087 7783
0 7785 5 1 1 7784
0 7786 7 1 2 7778 7785
0 7787 5 1 1 7786
0 7788 7 1 2 69742 7787
0 7789 5 1 1 7788
0 7790 7 3 2 69408 77304
0 7791 5 1 1 91091
0 7792 7 2 2 84608 87493
0 7793 5 1 1 91094
0 7794 7 1 2 7791 91095
0 7795 5 1 1 7794
0 7796 7 2 2 75257 90063
0 7797 5 1 1 91096
0 7798 7 1 2 76150 90487
0 7799 7 1 2 91097 7798
0 7800 5 1 1 7799
0 7801 7 1 2 7795 7800
0 7802 5 1 1 7801
0 7803 7 1 2 78472 7802
0 7804 5 1 1 7803
0 7805 7 1 2 7789 7804
0 7806 5 1 1 7805
0 7807 7 1 2 71287 7806
0 7808 5 1 1 7807
0 7809 7 1 2 71288 77291
0 7810 5 3 1 7809
0 7811 7 1 2 91098 91084
0 7812 5 1 1 7811
0 7813 7 10 2 89079 75727
0 7814 5 1 1 91101
0 7815 7 1 2 75000 91102
0 7816 7 1 2 89655 7815
0 7817 5 1 1 7816
0 7818 7 1 2 7812 7817
0 7819 5 1 1 7818
0 7820 7 1 2 64990 7819
0 7821 5 1 1 7820
0 7822 7 1 2 66187 77093
0 7823 5 2 1 7822
0 7824 7 1 2 69409 91111
0 7825 5 1 1 7824
0 7826 7 1 2 91085 7825
0 7827 5 1 1 7826
0 7828 7 1 2 7821 7827
0 7829 5 1 1 7828
0 7830 7 1 2 64624 7829
0 7831 5 1 1 7830
0 7832 7 2 2 86337 75903
0 7833 7 3 2 75728 90145
0 7834 7 2 2 69410 87402
0 7835 7 2 2 91115 91118
0 7836 7 1 2 91113 91120
0 7837 5 1 1 7836
0 7838 7 1 2 75001 81169
0 7839 5 1 1 7838
0 7840 7 1 2 78950 79752
0 7841 5 1 1 7840
0 7842 7 1 2 7839 7841
0 7843 5 1 1 7842
0 7844 7 1 2 91035 7843
0 7845 5 1 1 7844
0 7846 7 1 2 7837 7845
0 7847 7 1 2 7831 7846
0 7848 5 1 1 7847
0 7849 7 1 2 78473 7848
0 7850 5 1 1 7849
0 7851 7 20 2 64295 70108
0 7852 7 3 2 83318 91122
0 7853 5 1 1 91142
0 7854 7 1 2 69411 77299
0 7855 5 1 1 7854
0 7856 7 1 2 7853 7855
0 7857 5 1 1 7856
0 7858 7 1 2 89905 7857
0 7859 5 1 1 7858
0 7860 7 12 2 63872 64296
0 7861 7 1 2 84052 91145
0 7862 7 1 2 79347 7861
0 7863 5 1 1 7862
0 7864 7 1 2 7859 7863
0 7865 5 1 1 7864
0 7866 7 1 2 71289 7865
0 7867 5 1 1 7866
0 7868 7 1 2 78844 91036
0 7869 5 1 1 7868
0 7870 7 1 2 7867 7869
0 7871 5 1 1 7870
0 7872 7 1 2 67940 7871
0 7873 5 1 1 7872
0 7874 7 1 2 76287 81232
0 7875 7 1 2 91037 7874
0 7876 5 1 1 7875
0 7877 7 1 2 7873 7876
0 7878 5 1 1 7877
0 7879 7 1 2 83745 7878
0 7880 5 1 1 7879
0 7881 7 1 2 7850 7880
0 7882 7 1 2 7808 7881
0 7883 7 1 2 7752 7882
0 7884 5 1 1 7883
0 7885 7 1 2 89567 7884
0 7886 5 1 1 7885
0 7887 7 24 2 70656 70707
0 7888 7 3 2 69045 70109
0 7889 7 3 2 91157 91181
0 7890 7 4 2 86522 91184
0 7891 7 1 2 79363 89892
0 7892 7 2 2 91187 7891
0 7893 5 1 1 91191
0 7894 7 8 2 71905 68595
0 7895 7 2 2 91193 91188
0 7896 5 1 1 91201
0 7897 7 1 2 89009 7896
0 7898 5 1 1 7897
0 7899 7 1 2 89186 7898
0 7900 5 1 1 7899
0 7901 7 1 2 7893 7900
0 7902 5 1 1 7901
0 7903 7 1 2 90358 7902
0 7904 5 1 1 7903
0 7905 7 4 2 68785 90282
0 7906 7 5 2 90415 91203
0 7907 7 2 2 76836 91207
0 7908 7 9 2 66841 91212
0 7909 7 1 2 77551 75619
0 7910 7 2 2 91214 7909
0 7911 5 1 1 91223
0 7912 7 1 2 72962 91215
0 7913 5 3 1 7912
0 7914 7 1 2 77305 7780
0 7915 5 1 1 7914
0 7916 7 3 2 79364 90528
0 7917 5 1 1 91228
0 7918 7 4 2 89893 91229
0 7919 7 1 2 75620 91231
0 7920 7 1 2 7915 7919
0 7921 5 1 1 7920
0 7922 7 1 2 91225 7921
0 7923 5 1 1 7922
0 7924 7 1 2 71290 7923
0 7925 5 1 1 7924
0 7926 7 1 2 7911 7925
0 7927 5 1 1 7926
0 7928 7 1 2 70993 7927
0 7929 5 1 1 7928
0 7930 7 1 2 7904 7929
0 7931 5 1 1 7930
0 7932 7 1 2 84660 7931
0 7933 5 1 1 7932
0 7934 7 13 2 67058 72568
0 7935 7 2 2 91235 90283
0 7936 7 8 2 65676 66842
0 7937 7 5 2 90573 91250
0 7938 7 1 2 83319 91258
0 7939 7 1 2 91248 7938
0 7940 5 1 1 7939
0 7941 7 5 2 69046 64991
0 7942 7 7 2 68954 70657
0 7943 5 1 1 91268
0 7944 7 2 2 91269 90511
0 7945 7 2 2 91263 91275
0 7946 7 10 2 65931 72119
0 7947 7 1 2 78340 91279
0 7948 7 1 2 85381 7947
0 7949 7 1 2 91277 7948
0 7950 5 1 1 7949
0 7951 7 1 2 7940 7950
0 7952 5 1 1 7951
0 7953 7 1 2 85204 7952
0 7954 5 1 1 7953
0 7955 7 3 2 67059 87785
0 7956 7 1 2 86856 91289
0 7957 7 1 2 91208 7956
0 7958 5 1 1 7957
0 7959 7 1 2 7954 7958
0 7960 5 1 1 7959
0 7961 7 1 2 71291 7960
0 7962 5 1 1 7961
0 7963 7 1 2 78430 91224
0 7964 5 1 1 7963
0 7965 7 1 2 7962 7964
0 7966 5 1 1 7965
0 7967 7 1 2 69412 7966
0 7968 5 1 1 7967
0 7969 7 4 2 87435 89533
0 7970 7 1 2 86384 91292
0 7971 5 1 1 7970
0 7972 7 2 2 64992 91099
0 7973 5 1 1 91296
0 7974 7 1 2 7973 91112
0 7975 5 1 1 7974
0 7976 7 1 2 64625 7975
0 7977 5 1 1 7976
0 7978 7 3 2 73685 77042
0 7979 5 1 1 91298
0 7980 7 1 2 64993 91299
0 7981 5 1 1 7980
0 7982 7 1 2 7977 7981
0 7983 5 1 1 7982
0 7984 7 1 2 67941 90416
0 7985 7 1 2 7983 7984
0 7986 5 1 1 7985
0 7987 7 1 2 7971 7986
0 7988 5 1 1 7987
0 7989 7 2 2 79348 91204
0 7990 7 1 2 67553 91301
0 7991 7 1 2 7988 7990
0 7992 5 1 1 7991
0 7993 7 3 2 67060 91251
0 7994 7 6 2 65624 76913
0 7995 7 1 2 63959 91306
0 7996 7 5 2 91303 7995
0 7997 7 1 2 80265 87895
0 7998 7 1 2 91312 7997
0 7999 5 1 1 7998
0 8000 7 3 2 84061 90520
0 8001 7 1 2 77281 84507
0 8002 7 3 2 70708 72120
0 8003 7 1 2 90859 91320
0 8004 7 1 2 8001 8003
0 8005 7 1 2 91317 8004
0 8006 7 1 2 79956 8005
0 8007 5 1 1 8006
0 8008 7 1 2 7999 8007
0 8009 5 1 1 8008
0 8010 7 1 2 85205 8009
0 8011 5 1 1 8010
0 8012 7 5 2 76453 84992
0 8013 5 2 1 91323
0 8014 7 1 2 91216 80890
0 8015 5 1 1 8014
0 8016 7 1 2 64297 91192
0 8017 5 1 1 8016
0 8018 7 1 2 8015 8017
0 8019 5 1 1 8018
0 8020 7 1 2 91324 8019
0 8021 5 1 1 8020
0 8022 7 1 2 8011 8021
0 8023 7 1 2 7992 8022
0 8024 5 1 1 8023
0 8025 7 1 2 70994 8024
0 8026 5 1 1 8025
0 8027 7 1 2 7968 8026
0 8028 7 1 2 7933 8027
0 8029 7 1 2 7886 8028
0 8030 7 1 2 7629 8029
0 8031 5 1 1 8030
0 8032 7 1 2 71768 8031
0 8033 5 1 1 8032
0 8034 7 5 2 71906 72963
0 8035 7 2 2 67061 91158
0 8036 7 2 2 91330 91335
0 8037 7 6 2 69047 69413
0 8038 7 1 2 75153 91339
0 8039 7 1 2 91337 8038
0 8040 5 1 1 8039
0 8041 7 9 2 66843 90574
0 8042 7 4 2 65677 90423
0 8043 5 2 1 91354
0 8044 7 6 2 91345 91355
0 8045 5 1 1 91360
0 8046 7 16 2 72121 91361
0 8047 7 1 2 67942 91366
0 8048 5 1 1 8047
0 8049 7 1 2 8040 8048
0 8050 5 3 1 8049
0 8051 7 1 2 75470 91382
0 8052 5 1 1 8051
0 8053 7 6 2 64994 88012
0 8054 7 1 2 79753 91385
0 8055 7 3 2 72122 88047
0 8056 7 2 2 68955 91340
0 8057 7 1 2 91391 91394
0 8058 7 1 2 8054 8057
0 8059 5 1 1 8058
0 8060 7 1 2 8052 8059
0 8061 5 1 1 8060
0 8062 7 1 2 76454 8061
0 8063 5 1 1 8062
0 8064 7 4 2 68956 65678
0 8065 7 1 2 77768 91396
0 8066 7 1 2 75471 8065
0 8067 7 1 2 90602 8066
0 8068 5 1 1 8067
0 8069 7 1 2 8063 8068
0 8070 5 1 1 8069
0 8071 7 1 2 72569 8070
0 8072 5 1 1 8071
0 8073 7 1 2 79754 90168
0 8074 5 1 1 8073
0 8075 7 2 2 75801 78719
0 8076 5 1 1 91400
0 8077 7 1 2 8074 8076
0 8078 5 1 1 8077
0 8079 7 5 2 71907 91159
0 8080 7 4 2 69048 87951
0 8081 7 6 2 91402 91407
0 8082 7 1 2 78392 91411
0 8083 7 1 2 8078 8082
0 8084 5 1 1 8083
0 8085 7 1 2 8072 8084
0 8086 5 1 1 8085
0 8087 7 1 2 77574 8086
0 8088 5 1 1 8087
0 8089 7 1 2 83946 84007
0 8090 5 1 1 8089
0 8091 7 3 2 75347 8090
0 8092 7 4 2 66844 89391
0 8093 7 4 2 69414 90575
0 8094 7 1 2 91356 91424
0 8095 7 1 2 91420 8094
0 8096 7 1 2 91417 8095
0 8097 5 1 1 8096
0 8098 7 1 2 8088 8097
0 8099 5 1 1 8098
0 8100 7 1 2 89106 8099
0 8101 5 1 1 8100
0 8102 7 10 2 71580 81129
0 8103 5 1 1 91428
0 8104 7 1 2 72570 8103
0 8105 5 2 1 8104
0 8106 7 1 2 81204 91438
0 8107 5 1 1 8106
0 8108 7 15 2 69743 64995
0 8109 5 1 1 91440
0 8110 7 4 2 66470 87786
0 8111 7 1 2 91441 91455
0 8112 5 1 1 8111
0 8113 7 1 2 8107 8112
0 8114 5 1 1 8113
0 8115 7 1 2 75072 8114
0 8116 5 1 1 8115
0 8117 7 1 2 78796 84993
0 8118 5 4 1 8117
0 8119 7 1 2 73944 85055
0 8120 5 1 1 8119
0 8121 7 1 2 91459 8120
0 8122 5 1 1 8121
0 8123 7 1 2 69415 8122
0 8124 5 2 1 8123
0 8125 7 6 2 71292 84281
0 8126 5 1 1 91465
0 8127 7 1 2 82677 91466
0 8128 5 1 1 8127
0 8129 7 1 2 91463 8128
0 8130 7 1 2 8116 8129
0 8131 5 1 1 8130
0 8132 7 1 2 73686 8131
0 8133 5 1 1 8132
0 8134 7 1 2 75621 87032
0 8135 7 1 2 84661 8134
0 8136 5 1 1 8135
0 8137 7 1 2 87903 8136
0 8138 5 1 1 8137
0 8139 7 1 2 71293 8138
0 8140 5 1 1 8139
0 8141 7 1 2 78625 85056
0 8142 5 1 1 8141
0 8143 7 1 2 78761 90930
0 8144 5 1 1 8143
0 8145 7 1 2 8142 8144
0 8146 5 1 1 8145
0 8147 7 1 2 69416 8146
0 8148 5 1 1 8147
0 8149 7 1 2 8140 8148
0 8150 7 1 2 8133 8149
0 8151 5 1 1 8150
0 8152 7 6 2 90064 88128
0 8153 7 1 2 8151 91471
0 8154 5 1 1 8153
0 8155 7 3 2 75348 81550
0 8156 5 1 1 91477
0 8157 7 11 2 72123 72571
0 8158 7 2 2 91480 90622
0 8159 7 1 2 82100 91491
0 8160 7 1 2 91478 8159
0 8161 5 1 1 8160
0 8162 7 1 2 8154 8161
0 8163 5 1 1 8162
0 8164 7 1 2 70995 8163
0 8165 5 1 1 8164
0 8166 7 1 2 91418 90627
0 8167 5 1 1 8166
0 8168 7 2 2 79464 87725
0 8169 7 1 2 77094 75767
0 8170 7 1 2 91493 8169
0 8171 7 1 2 91439 8170
0 8172 5 1 1 8171
0 8173 7 1 2 8167 8172
0 8174 5 1 1 8173
0 8175 7 1 2 73371 8174
0 8176 5 1 1 8175
0 8177 7 12 2 67554 73687
0 8178 7 3 2 65932 79570
0 8179 7 1 2 91495 91507
0 8180 7 1 2 91472 8179
0 8181 5 1 1 8180
0 8182 7 1 2 8176 8181
0 8183 5 1 1 8182
0 8184 7 1 2 74128 8183
0 8185 5 1 1 8184
0 8186 7 1 2 8165 8185
0 8187 5 1 1 8186
0 8188 7 1 2 89568 8187
0 8189 5 1 1 8188
0 8190 7 3 2 67062 88048
0 8191 7 4 2 90521 75154
0 8192 7 4 2 91510 91513
0 8193 7 2 2 86338 78626
0 8194 5 2 1 91521
0 8195 7 1 2 69417 91523
0 8196 5 1 1 8195
0 8197 7 1 2 76455 8196
0 8198 5 1 1 8197
0 8199 7 2 2 78591 80145
0 8200 5 2 1 91525
0 8201 7 1 2 78845 91527
0 8202 5 1 1 8201
0 8203 7 1 2 8198 8202
0 8204 5 1 1 8203
0 8205 7 1 2 72964 8204
0 8206 5 1 1 8205
0 8207 7 1 2 91528 88326
0 8208 5 1 1 8207
0 8209 7 1 2 8206 8208
0 8210 5 1 1 8209
0 8211 7 1 2 91517 8210
0 8212 5 1 1 8211
0 8213 7 1 2 75960 90159
0 8214 5 1 1 8213
0 8215 7 1 2 84250 89944
0 8216 5 1 1 8215
0 8217 7 1 2 8214 8216
0 8218 5 1 1 8217
0 8219 7 1 2 91367 8218
0 8220 5 1 1 8219
0 8221 7 1 2 8212 8220
0 8222 5 1 1 8221
0 8223 7 1 2 70996 8222
0 8224 5 1 1 8223
0 8225 7 17 2 65625 88910
0 8226 7 2 2 77821 91529
0 8227 7 3 2 77895 84376
0 8228 7 1 2 91546 91548
0 8229 5 1 1 8228
0 8230 7 14 2 63873 69049
0 8231 7 11 2 91551 91160
0 8232 5 1 1 91565
0 8233 7 1 2 76151 79514
0 8234 7 1 2 84193 8233
0 8235 7 1 2 91566 8234
0 8236 5 1 1 8235
0 8237 7 1 2 8229 8236
0 8238 5 1 1 8237
0 8239 7 1 2 71294 8238
0 8240 5 1 1 8239
0 8241 7 2 2 88513 88940
0 8242 5 4 1 91576
0 8243 7 1 2 67943 89741
0 8244 7 1 2 91577 8243
0 8245 5 1 1 8244
0 8246 7 1 2 8240 8245
0 8247 5 1 1 8246
0 8248 7 1 2 73945 8247
0 8249 5 1 1 8248
0 8250 7 2 2 77924 77936
0 8251 5 1 1 91582
0 8252 7 1 2 78904 91583
0 8253 5 2 1 8252
0 8254 7 5 2 73372 79571
0 8255 5 1 1 91586
0 8256 7 1 2 1571 8255
0 8257 5 2 1 8256
0 8258 7 1 2 72965 91591
0 8259 5 1 1 8258
0 8260 7 1 2 91584 8259
0 8261 5 1 1 8260
0 8262 7 1 2 91368 8261
0 8263 5 1 1 8262
0 8264 7 4 2 71295 78341
0 8265 7 7 2 70709 65933
0 8266 5 1 1 91597
0 8267 7 3 2 91593 91598
0 8268 7 6 2 67063 74729
0 8269 7 1 2 91514 91607
0 8270 7 1 2 91604 8269
0 8271 5 1 1 8270
0 8272 7 1 2 8263 8271
0 8273 7 1 2 8249 8272
0 8274 5 1 1 8273
0 8275 7 1 2 69418 8274
0 8276 5 1 1 8275
0 8277 7 1 2 8224 8276
0 8278 5 1 1 8277
0 8279 7 1 2 67555 8278
0 8280 5 1 1 8279
0 8281 7 2 2 77204 82736
0 8282 5 1 1 91613
0 8283 7 3 2 77406 8282
0 8284 7 1 2 91615 91369
0 8285 5 1 1 8284
0 8286 7 3 2 76796 78720
0 8287 7 4 2 70997 91161
0 8288 7 1 2 76952 91552
0 8289 7 1 2 91621 8288
0 8290 7 1 2 91618 8289
0 8291 5 1 1 8290
0 8292 7 1 2 8285 8291
0 8293 5 1 1 8292
0 8294 7 1 2 81279 8293
0 8295 5 1 1 8294
0 8296 7 1 2 65934 81617
0 8297 5 4 1 8296
0 8298 7 1 2 77407 91625
0 8299 7 2 2 81624 8298
0 8300 7 1 2 75622 91370
0 8301 7 1 2 91629 8300
0 8302 5 1 1 8301
0 8303 7 1 2 74941 87177
0 8304 5 1 1 8303
0 8305 7 1 2 83304 8304
0 8306 5 1 1 8305
0 8307 7 6 2 70998 71908
0 8308 7 5 2 67064 91631
0 8309 7 6 2 70616 91162
0 8310 7 5 2 69419 91553
0 8311 7 3 2 91642 91648
0 8312 7 1 2 91637 91653
0 8313 7 1 2 8306 8312
0 8314 5 1 1 8313
0 8315 7 1 2 8302 8314
0 8316 7 1 2 8295 8315
0 8317 5 1 1 8316
0 8318 7 1 2 72572 8317
0 8319 5 1 1 8318
0 8320 7 2 2 75802 88040
0 8321 7 1 2 83407 81015
0 8322 7 4 2 70710 71581
0 8323 7 3 2 84479 91658
0 8324 7 1 2 91662 91608
0 8325 7 1 2 8321 8324
0 8326 7 1 2 91656 8325
0 8327 5 1 1 8326
0 8328 7 1 2 8319 8327
0 8329 7 1 2 8280 8328
0 8330 5 1 1 8329
0 8331 7 1 2 85206 8330
0 8332 5 1 1 8331
0 8333 7 1 2 8189 8332
0 8334 7 1 2 8101 8333
0 8335 7 1 2 8033 8334
0 8336 7 1 2 7452 8335
0 8337 5 1 1 8336
0 8338 7 1 2 64029 8337
0 8339 5 1 1 8338
0 8340 7 1 2 7009 8339
0 8341 5 1 1 8340
0 8342 7 1 2 70374 8341
0 8343 5 1 1 8342
0 8344 7 6 2 69050 69744
0 8345 7 2 2 88013 91665
0 8346 7 6 2 65935 68596
0 8347 7 3 2 70711 84480
0 8348 7 2 2 91673 91679
0 8349 7 1 2 91671 91682
0 8350 5 1 1 8349
0 8351 7 4 2 65317 88941
0 8352 7 1 2 76288 91684
0 8353 5 1 1 8352
0 8354 7 1 2 8350 8353
0 8355 5 1 1 8354
0 8356 7 1 2 72573 8355
0 8357 5 1 1 8356
0 8358 7 13 2 70712 88014
0 8359 7 1 2 71769 74143
0 8360 7 8 2 71909 67556
0 8361 7 6 2 69051 64626
0 8362 7 1 2 91701 91709
0 8363 7 1 2 8359 8362
0 8364 7 1 2 91688 8363
0 8365 5 1 1 8364
0 8366 7 1 2 8357 8365
0 8367 5 1 1 8366
0 8368 7 1 2 68302 8367
0 8369 5 1 1 8368
0 8370 7 4 2 65318 65626
0 8371 7 4 2 63960 65581
0 8372 7 2 2 91715 91719
0 8373 7 2 2 91252 91723
0 8374 5 1 1 91725
0 8375 7 1 2 80338 89232
0 8376 7 1 2 91726 8375
0 8377 5 1 1 8376
0 8378 7 1 2 8369 8377
0 8379 5 1 1 8378
0 8380 7 1 2 71582 8379
0 8381 5 1 1 8380
0 8382 7 1 2 90806 91685
0 8383 5 1 1 8382
0 8384 7 1 2 8381 8383
0 8385 5 1 1 8384
0 8386 7 1 2 70110 8385
0 8387 5 1 1 8386
0 8388 7 1 2 73373 80489
0 8389 5 3 1 8388
0 8390 7 1 2 90807 91727
0 8391 5 1 1 8390
0 8392 7 1 2 76289 78431
0 8393 5 2 1 8392
0 8394 7 1 2 8391 91730
0 8395 5 1 1 8394
0 8396 7 1 2 91686 8395
0 8397 5 1 1 8396
0 8398 7 1 2 8387 8397
0 8399 5 1 1 8398
0 8400 7 1 2 88129 8399
0 8401 5 1 1 8400
0 8402 7 1 2 731 87778
0 8403 5 1 1 8402
0 8404 7 1 2 79782 8403
0 8405 5 1 1 8404
0 8406 7 1 2 73374 91419
0 8407 5 1 1 8406
0 8408 7 1 2 8405 8407
0 8409 5 1 1 8408
0 8410 7 1 2 71770 8409
0 8411 5 1 1 8410
0 8412 7 1 2 1974 8411
0 8413 5 1 1 8412
0 8414 7 1 2 91371 8413
0 8415 5 1 1 8414
0 8416 7 1 2 8401 8415
0 8417 5 1 1 8416
0 8418 7 1 2 85860 8417
0 8419 5 1 1 8418
0 8420 7 1 2 64627 82617
0 8421 5 4 1 8420
0 8422 7 5 2 71771 73946
0 8423 7 1 2 64996 91736
0 8424 5 1 1 8423
0 8425 7 1 2 91732 8424
0 8426 5 1 1 8425
0 8427 7 1 2 88942 8426
0 8428 5 1 1 8427
0 8429 7 6 2 68303 76640
0 8430 5 4 1 91741
0 8431 7 2 2 74521 80339
0 8432 5 3 1 91751
0 8433 7 1 2 91747 91753
0 8434 5 2 1 8433
0 8435 7 1 2 77972 88060
0 8436 7 1 2 91756 8435
0 8437 5 1 1 8436
0 8438 7 1 2 8428 8437
0 8439 5 1 1 8438
0 8440 7 1 2 66188 8439
0 8441 5 1 1 8440
0 8442 7 4 2 65319 88015
0 8443 7 1 2 69052 83525
0 8444 7 1 2 91758 8443
0 8445 7 1 2 91605 8444
0 8446 5 1 1 8445
0 8447 7 2 2 80922 82291
0 8448 5 5 1 91762
0 8449 7 3 2 71772 88943
0 8450 5 1 1 91769
0 8451 7 1 2 91763 91770
0 8452 5 1 1 8451
0 8453 7 1 2 8446 8452
0 8454 7 1 2 8441 8453
0 8455 5 1 1 8454
0 8456 7 1 2 88514 8455
0 8457 5 1 1 8456
0 8458 7 1 2 76555 88944
0 8459 5 1 1 8458
0 8460 7 7 2 65320 70658
0 8461 7 2 2 91772 90370
0 8462 7 1 2 91779 91683
0 8463 5 1 1 8462
0 8464 7 1 2 8459 8463
0 8465 5 1 1 8464
0 8466 7 1 2 73375 8465
0 8467 5 1 1 8466
0 8468 7 3 2 66189 73896
0 8469 5 4 1 91781
0 8470 7 1 2 91784 90018
0 8471 5 1 1 8470
0 8472 7 3 2 88016 79515
0 8473 7 4 2 91788 89503
0 8474 7 1 2 68597 91791
0 8475 7 1 2 8471 8474
0 8476 5 1 1 8475
0 8477 7 1 2 8467 8476
0 8478 5 1 1 8477
0 8479 7 1 2 88130 8478
0 8480 5 1 1 8479
0 8481 7 1 2 67557 8480
0 8482 7 1 2 8457 8481
0 8483 5 1 1 8482
0 8484 7 1 2 82366 86622
0 8485 5 1 1 8484
0 8486 7 1 2 90568 8485
0 8487 5 1 1 8486
0 8488 7 1 2 88820 88131
0 8489 5 1 1 8488
0 8490 7 1 2 8487 8489
0 8491 5 1 1 8490
0 8492 7 1 2 76290 8491
0 8493 5 1 1 8492
0 8494 7 2 2 78627 77822
0 8495 5 1 1 91795
0 8496 7 1 2 66666 91796
0 8497 5 1 1 8496
0 8498 7 1 2 76456 89288
0 8499 7 1 2 8497 8498
0 8500 5 1 1 8499
0 8501 7 1 2 8493 8500
0 8502 5 1 1 8501
0 8503 7 1 2 88945 8502
0 8504 5 1 1 8503
0 8505 7 1 2 68304 90638
0 8506 5 1 1 8505
0 8507 7 1 2 89734 8506
0 8508 5 1 1 8507
0 8509 7 2 2 68598 91666
0 8510 7 3 2 88017 91599
0 8511 7 1 2 84481 91799
0 8512 7 1 2 91797 8511
0 8513 7 1 2 80934 8512
0 8514 7 1 2 8508 8513
0 8515 5 1 1 8514
0 8516 7 1 2 72574 8515
0 8517 7 1 2 8504 8516
0 8518 5 1 1 8517
0 8519 7 1 2 85207 8518
0 8520 7 1 2 8483 8519
0 8521 5 1 1 8520
0 8522 7 1 2 8419 8521
0 8523 5 1 1 8522
0 8524 7 1 2 69420 8523
0 8525 5 1 1 8524
0 8526 7 4 2 68786 65321
0 8527 7 3 2 65936 76352
0 8528 7 1 2 91802 91806
0 8529 5 1 1 8528
0 8530 7 1 2 5701 8529
0 8531 5 1 1 8530
0 8532 7 1 2 88132 8531
0 8533 5 1 1 8532
0 8534 7 2 2 68305 81989
0 8535 7 1 2 90229 89330
0 8536 7 1 2 91809 8535
0 8537 5 1 1 8536
0 8538 7 1 2 8533 8537
0 8539 5 1 1 8538
0 8540 7 1 2 88946 8539
0 8541 5 1 1 8540
0 8542 7 1 2 88287 89735
0 8543 5 3 1 8542
0 8544 7 2 2 85208 91811
0 8545 5 2 1 91814
0 8546 7 4 2 70111 72015
0 8547 7 5 2 68787 91818
0 8548 5 1 1 91822
0 8549 7 1 2 91823 88133
0 8550 5 1 1 8549
0 8551 7 1 2 91816 8550
0 8552 5 1 1 8551
0 8553 7 1 2 73897 8552
0 8554 5 1 1 8553
0 8555 7 1 2 83495 78683
0 8556 7 1 2 89300 8555
0 8557 5 1 1 8556
0 8558 7 1 2 8554 8557
0 8559 5 1 1 8558
0 8560 7 1 2 91674 91412
0 8561 7 1 2 8559 8560
0 8562 5 1 1 8561
0 8563 7 1 2 8541 8562
0 8564 5 1 1 8563
0 8565 7 1 2 71296 8564
0 8566 5 1 1 8565
0 8567 7 7 2 71583 66845
0 8568 7 3 2 80512 76837
0 8569 7 2 2 91827 91834
0 8570 7 1 2 84172 87726
0 8571 7 1 2 76130 8570
0 8572 7 1 2 91530 8571
0 8573 7 1 2 91837 8572
0 8574 5 1 1 8573
0 8575 7 1 2 8566 8574
0 8576 5 1 1 8575
0 8577 7 1 2 69745 8576
0 8578 5 1 1 8577
0 8579 7 5 2 76131 89534
0 8580 7 4 2 63961 70112
0 8581 7 1 2 91839 91844
0 8582 7 1 2 91494 8581
0 8583 7 1 2 91838 8582
0 8584 5 1 1 8583
0 8585 7 1 2 8578 8584
0 8586 5 1 1 8585
0 8587 7 1 2 67558 8586
0 8588 5 1 1 8587
0 8589 7 1 2 8525 8588
0 8590 5 1 1 8589
0 8591 7 1 2 67944 8590
0 8592 5 1 1 8591
0 8593 7 6 2 66846 67945
0 8594 7 3 2 82340 89301
0 8595 5 1 1 91854
0 8596 7 2 2 68788 77497
0 8597 7 1 2 91835 91857
0 8598 5 2 1 8597
0 8599 7 1 2 82618 89302
0 8600 5 1 1 8599
0 8601 7 1 2 91859 8600
0 8602 5 1 1 8601
0 8603 7 1 2 71584 8602
0 8604 5 1 1 8603
0 8605 7 1 2 8595 8604
0 8606 5 1 1 8605
0 8607 7 1 2 70113 8606
0 8608 5 1 1 8607
0 8609 7 1 2 90967 90618
0 8610 5 1 1 8609
0 8611 7 1 2 85209 82341
0 8612 7 1 2 8610 8611
0 8613 5 1 1 8612
0 8614 7 1 2 8608 8613
0 8615 5 1 1 8614
0 8616 7 2 2 91848 8615
0 8617 7 1 2 90784 91861
0 8618 5 1 1 8617
0 8619 7 1 2 84111 88515
0 8620 5 1 1 8619
0 8621 7 1 2 89991 8620
0 8622 5 1 1 8621
0 8623 7 1 2 85861 8622
0 8624 5 1 1 8623
0 8625 7 1 2 89320 8624
0 8626 5 1 1 8625
0 8627 7 1 2 75349 8626
0 8628 5 1 1 8627
0 8629 7 1 2 79049 89753
0 8630 7 1 2 91858 8629
0 8631 5 1 1 8630
0 8632 7 1 2 91817 8631
0 8633 7 1 2 8628 8632
0 8634 5 1 1 8633
0 8635 7 1 2 67946 8634
0 8636 5 1 1 8635
0 8637 7 1 2 70114 91855
0 8638 5 1 1 8637
0 8639 7 5 2 71773 72016
0 8640 7 6 2 68789 91863
0 8641 7 1 2 91868 76782
0 8642 5 1 1 8641
0 8643 7 1 2 85210 82619
0 8644 5 1 1 8643
0 8645 7 1 2 8642 8644
0 8646 5 1 1 8645
0 8647 7 1 2 88516 8646
0 8648 5 1 1 8647
0 8649 7 1 2 91860 8648
0 8650 5 1 1 8649
0 8651 7 1 2 70115 8650
0 8652 5 1 1 8651
0 8653 7 1 2 68306 91815
0 8654 5 1 1 8653
0 8655 7 1 2 8652 8654
0 8656 5 1 1 8655
0 8657 7 1 2 71585 8656
0 8658 5 1 1 8657
0 8659 7 1 2 8638 8658
0 8660 7 1 2 8636 8659
0 8661 5 1 1 8660
0 8662 7 1 2 88947 8661
0 8663 5 1 1 8662
0 8664 7 12 2 71586 71910
0 8665 7 3 2 70713 91874
0 8666 7 2 2 91886 91657
0 8667 7 1 2 75531 91889
0 8668 5 1 1 8667
0 8669 7 1 2 71774 91372
0 8670 5 1 1 8669
0 8671 7 1 2 8668 8670
0 8672 5 1 1 8671
0 8673 7 1 2 85862 8672
0 8674 5 1 1 8673
0 8675 7 1 2 89688 90979
0 8676 5 1 1 8675
0 8677 7 1 2 7275 8676
0 8678 5 1 1 8677
0 8679 7 10 2 63747 69053
0 8680 7 2 2 75729 91689
0 8681 7 10 2 91891 91901
0 8682 7 1 2 68599 91903
0 8683 7 1 2 8678 8682
0 8684 5 1 1 8683
0 8685 7 1 2 8674 8684
0 8686 5 1 1 8685
0 8687 7 1 2 64298 8686
0 8688 5 1 1 8687
0 8689 7 3 2 91253 75674
0 8690 7 2 2 90308 91913
0 8691 7 1 2 85863 89689
0 8692 7 1 2 91916 8691
0 8693 5 1 1 8692
0 8694 7 1 2 79704 74098
0 8695 7 1 2 91887 8694
0 8696 7 1 2 90300 8695
0 8697 5 1 1 8696
0 8698 7 1 2 8693 8697
0 8699 5 1 1 8698
0 8700 7 1 2 64997 8699
0 8701 5 1 1 8700
0 8702 7 2 2 86133 88517
0 8703 5 1 1 91918
0 8704 7 1 2 89992 8703
0 8705 5 1 1 8704
0 8706 7 1 2 85864 8705
0 8707 5 1 1 8706
0 8708 7 1 2 89321 8707
0 8709 5 1 1 8708
0 8710 7 1 2 88948 8709
0 8711 5 1 1 8710
0 8712 7 1 2 8701 8711
0 8713 7 1 2 8688 8712
0 8714 5 1 1 8713
0 8715 7 1 2 68307 8714
0 8716 5 1 1 8715
0 8717 7 3 2 69054 79365
0 8718 7 1 2 72124 91123
0 8719 7 1 2 83580 8718
0 8720 7 1 2 91920 8719
0 8721 7 1 2 91902 8720
0 8722 5 1 1 8721
0 8723 7 1 2 8716 8722
0 8724 5 1 1 8723
0 8725 7 1 2 67947 8724
0 8726 5 1 1 8725
0 8727 7 1 2 8663 8726
0 8728 5 1 1 8727
0 8729 7 1 2 71297 8728
0 8730 5 1 1 8729
0 8731 7 1 2 8618 8730
0 8732 5 1 1 8731
0 8733 7 1 2 69746 8732
0 8734 5 1 1 8733
0 8735 7 2 2 75961 80513
0 8736 5 1 1 91923
0 8737 7 1 2 76641 80514
0 8738 5 3 1 8737
0 8739 7 1 2 79957 91925
0 8740 7 1 2 8736 8739
0 8741 5 1 1 8740
0 8742 7 1 2 88949 8741
0 8743 5 1 1 8742
0 8744 7 4 2 91690 91667
0 8745 7 1 2 91594 88455
0 8746 7 1 2 91928 8745
0 8747 5 1 1 8746
0 8748 7 1 2 8743 8747
0 8749 5 1 1 8748
0 8750 7 1 2 65322 8749
0 8751 5 1 1 8750
0 8752 7 4 2 70714 71298
0 8753 7 3 2 76797 90522
0 8754 7 2 2 91932 91936
0 8755 7 1 2 72966 82367
0 8756 5 2 1 8755
0 8757 7 2 2 87033 91941
0 8758 7 1 2 69747 91943
0 8759 5 1 1 8758
0 8760 7 1 2 83417 81353
0 8761 5 1 1 8760
0 8762 7 1 2 8759 8761
0 8763 5 1 1 8762
0 8764 7 1 2 64998 8763
0 8765 5 1 1 8764
0 8766 7 7 2 69748 66471
0 8767 5 1 1 91945
0 8768 7 4 2 71775 74772
0 8769 7 1 2 91946 91952
0 8770 5 1 1 8769
0 8771 7 1 2 8765 8770
0 8772 5 1 1 8771
0 8773 7 1 2 91939 8772
0 8774 5 1 1 8773
0 8775 7 1 2 8751 8774
0 8776 5 1 1 8775
0 8777 7 1 2 85865 8776
0 8778 5 1 1 8777
0 8779 7 1 2 83540 83110
0 8780 7 1 2 77566 8779
0 8781 5 1 1 8780
0 8782 7 1 2 83287 8781
0 8783 5 1 1 8782
0 8784 7 1 2 82960 8783
0 8785 5 1 1 8784
0 8786 7 2 2 73947 83897
0 8787 7 1 2 76409 91956
0 8788 5 1 1 8787
0 8789 7 1 2 8785 8788
0 8790 5 1 1 8789
0 8791 7 1 2 88061 8790
0 8792 5 1 1 8791
0 8793 7 1 2 76192 77597
0 8794 5 1 1 8793
0 8795 7 1 2 88950 8794
0 8796 5 1 1 8795
0 8797 7 1 2 8792 8796
0 8798 5 1 1 8797
0 8799 7 1 2 85211 8798
0 8800 5 1 1 8799
0 8801 7 3 2 66847 85866
0 8802 7 3 2 63962 91958
0 8803 7 3 2 91961 91840
0 8804 5 2 1 91964
0 8805 7 3 2 66190 75730
0 8806 7 1 2 74844 91969
0 8807 7 1 2 90380 8806
0 8808 5 1 1 8807
0 8809 7 1 2 91967 8808
0 8810 5 1 1 8809
0 8811 7 1 2 67948 8810
0 8812 5 1 1 8811
0 8813 7 2 2 75731 76783
0 8814 7 1 2 91972 90381
0 8815 5 1 1 8814
0 8816 7 1 2 91968 8815
0 8817 5 1 1 8816
0 8818 7 1 2 76291 8817
0 8819 5 1 1 8818
0 8820 7 3 2 71299 86094
0 8821 7 2 2 91643 91974
0 8822 7 2 2 85867 77653
0 8823 7 1 2 91979 91798
0 8824 7 1 2 91977 8823
0 8825 5 1 1 8824
0 8826 7 1 2 8819 8825
0 8827 7 1 2 8812 8826
0 8828 5 1 1 8827
0 8829 7 1 2 75350 8828
0 8830 5 1 1 8829
0 8831 7 1 2 8800 8830
0 8832 7 1 2 8778 8831
0 8833 5 1 1 8832
0 8834 7 1 2 88134 8833
0 8835 5 1 1 8834
0 8836 7 5 2 88049 91780
0 8837 7 2 2 79834 91926
0 8838 5 1 1 91986
0 8839 7 1 2 72967 8838
0 8840 5 1 1 8839
0 8841 7 4 2 80923 79240
0 8842 5 1 1 91988
0 8843 7 1 2 67949 91989
0 8844 5 2 1 8843
0 8845 7 1 2 8840 91992
0 8846 5 2 1 8845
0 8847 7 1 2 91981 91994
0 8848 5 1 1 8847
0 8849 7 10 2 64999 77948
0 8850 5 2 1 91996
0 8851 7 4 2 66667 77654
0 8852 7 1 2 91997 92008
0 8853 5 1 1 8852
0 8854 7 1 2 88951 8853
0 8855 5 1 1 8854
0 8856 7 1 2 8848 8855
0 8857 5 1 1 8856
0 8858 7 1 2 71300 8857
0 8859 5 1 1 8858
0 8860 7 2 2 80515 78762
0 8861 7 1 2 91982 92012
0 8862 5 1 1 8861
0 8863 7 1 2 82620 88952
0 8864 5 1 1 8863
0 8865 7 1 2 8862 8864
0 8866 5 1 1 8865
0 8867 7 1 2 74522 8866
0 8868 5 1 1 8867
0 8869 7 2 2 82368 75599
0 8870 5 1 1 92014
0 8871 7 1 2 75351 8870
0 8872 5 1 1 8871
0 8873 7 1 2 82621 75623
0 8874 5 1 1 8873
0 8875 7 1 2 82737 8874
0 8876 7 1 2 8872 8875
0 8877 5 1 1 8876
0 8878 7 1 2 88953 8877
0 8879 5 1 1 8878
0 8880 7 2 2 70715 91759
0 8881 7 2 2 75549 91668
0 8882 7 1 2 87916 92018
0 8883 7 1 2 92016 8882
0 8884 5 1 1 8883
0 8885 7 1 2 8879 8884
0 8886 7 1 2 8868 8885
0 8887 7 1 2 8859 8886
0 8888 5 1 1 8887
0 8889 7 1 2 85212 8888
0 8890 5 1 1 8889
0 8891 7 1 2 73376 79944
0 8892 5 3 1 8891
0 8893 7 1 2 77567 81498
0 8894 5 2 1 8893
0 8895 7 1 2 72968 78788
0 8896 5 1 1 8895
0 8897 7 1 2 92023 8896
0 8898 5 1 1 8897
0 8899 7 1 2 68600 8898
0 8900 5 1 1 8899
0 8901 7 1 2 81655 8900
0 8902 5 1 1 8901
0 8903 7 1 2 71776 8902
0 8904 5 1 1 8903
0 8905 7 1 2 92020 8904
0 8906 5 1 1 8905
0 8907 7 1 2 90904 8906
0 8908 5 1 1 8907
0 8909 7 1 2 8890 8908
0 8910 5 1 1 8909
0 8911 7 1 2 88518 8910
0 8912 5 1 1 8911
0 8913 7 1 2 8835 8912
0 8914 5 1 1 8913
0 8915 7 1 2 69421 8914
0 8916 5 1 1 8915
0 8917 7 3 2 65679 71301
0 8918 7 5 2 90742 92025
0 8919 7 1 2 92028 91862
0 8920 5 1 1 8919
0 8921 7 1 2 72575 8920
0 8922 7 1 2 8916 8921
0 8923 7 1 2 8734 8922
0 8924 5 1 1 8923
0 8925 7 4 2 67065 79717
0 8926 7 3 2 63874 75258
0 8927 7 1 2 92033 92037
0 8928 5 1 1 8927
0 8929 7 2 2 74615 90738
0 8930 5 2 1 92040
0 8931 7 1 2 64299 92041
0 8932 5 1 1 8931
0 8933 7 1 2 8928 8932
0 8934 5 1 1 8933
0 8935 7 1 2 73377 8934
0 8936 5 1 1 8935
0 8937 7 2 2 83345 90488
0 8938 5 1 1 92044
0 8939 7 1 2 8936 8938
0 8940 5 1 1 8939
0 8941 7 1 2 69749 8940
0 8942 5 1 1 8941
0 8943 7 1 2 73948 90614
0 8944 5 1 1 8943
0 8945 7 3 2 68957 75259
0 8946 7 1 2 77721 92046
0 8947 5 1 1 8946
0 8948 7 1 2 8944 8947
0 8949 5 2 1 8948
0 8950 7 1 2 81205 92049
0 8951 5 1 1 8950
0 8952 7 1 2 8942 8951
0 8953 5 1 1 8952
0 8954 7 1 2 71302 8953
0 8955 5 1 1 8954
0 8956 7 3 2 68958 84377
0 8957 5 1 1 92051
0 8958 7 1 2 83271 92052
0 8959 5 1 1 8958
0 8960 7 2 2 83898 79324
0 8961 7 13 2 63875 65000
0 8962 7 1 2 76193 92056
0 8963 7 1 2 92054 8962
0 8964 5 1 1 8963
0 8965 7 1 2 8959 8964
0 8966 5 1 1 8965
0 8967 7 1 2 71587 8966
0 8968 5 1 1 8967
0 8969 7 1 2 83468 92050
0 8970 5 1 1 8969
0 8971 7 3 2 68959 79273
0 8972 7 7 2 66191 72125
0 8973 7 1 2 75550 92072
0 8974 7 1 2 92069 8973
0 8975 5 1 1 8974
0 8976 7 1 2 8970 8975
0 8977 7 1 2 8968 8976
0 8978 7 1 2 8955 8977
0 8979 5 1 1 8978
0 8980 7 1 2 85213 8979
0 8981 5 1 1 8980
0 8982 7 3 2 79083 76170
0 8983 7 2 2 75524 79099
0 8984 7 1 2 88456 92082
0 8985 7 1 2 92079 8984
0 8986 5 1 1 8985
0 8987 7 1 2 8981 8986
0 8988 5 1 1 8987
0 8989 7 1 2 88062 8988
0 8990 5 1 1 8989
0 8991 7 1 2 91217 1677
0 8992 5 1 1 8991
0 8993 7 3 2 80073 83346
0 8994 5 4 1 92084
0 8995 7 1 2 92085 91218
0 8996 5 1 1 8995
0 8997 7 2 2 79553 75847
0 8998 5 1 1 92091
0 8999 7 1 2 72969 88298
0 9000 5 1 1 8999
0 9001 7 1 2 8998 9000
0 9002 5 2 1 9001
0 9003 7 1 2 89303 91413
0 9004 7 1 2 92093 9003
0 9005 5 1 1 9004
0 9006 7 1 2 8996 9005
0 9007 5 1 1 9006
0 9008 7 1 2 80516 9007
0 9009 5 1 1 9008
0 9010 7 1 2 8992 9009
0 9011 7 1 2 8990 9010
0 9012 5 1 1 9011
0 9013 7 1 2 65323 9012
0 9014 5 1 1 9013
0 9015 7 1 2 67950 83774
0 9016 5 1 1 9015
0 9017 7 1 2 74816 9016
0 9018 5 1 1 9017
0 9019 7 1 2 71777 9018
0 9020 5 1 1 9019
0 9021 7 1 2 74497 79421
0 9022 5 2 1 9021
0 9023 7 1 2 82622 92095
0 9024 5 1 1 9023
0 9025 7 1 2 81248 9024
0 9026 7 1 2 9020 9025
0 9027 5 1 1 9026
0 9028 7 1 2 66192 9027
0 9029 5 1 1 9028
0 9030 7 1 2 71778 75962
0 9031 7 1 2 87875 9030
0 9032 5 1 1 9031
0 9033 7 1 2 9029 9032
0 9034 5 1 1 9033
0 9035 7 1 2 85214 9034
0 9036 5 1 1 9035
0 9037 7 2 2 76556 82342
0 9038 5 1 1 92097
0 9039 7 1 2 67951 92098
0 9040 5 1 1 9039
0 9041 7 1 2 92021 9040
0 9042 5 1 1 9041
0 9043 7 1 2 64300 9042
0 9044 5 1 1 9043
0 9045 7 2 2 78846 77937
0 9046 5 1 1 92099
0 9047 7 1 2 82343 78832
0 9048 5 1 1 9047
0 9049 7 1 2 9046 9048
0 9050 5 1 1 9049
0 9051 7 1 2 72970 9050
0 9052 5 1 1 9051
0 9053 7 1 2 79408 86238
0 9054 5 1 1 9053
0 9055 7 1 2 84432 9054
0 9056 5 1 1 9055
0 9057 7 1 2 65001 9056
0 9058 5 1 1 9057
0 9059 7 1 2 9052 9058
0 9060 7 1 2 9044 9059
0 9061 5 1 1 9060
0 9062 7 1 2 85868 9061
0 9063 5 1 1 9062
0 9064 7 1 2 9036 9063
0 9065 5 1 1 9064
0 9066 7 1 2 88519 9065
0 9067 5 1 1 9066
0 9068 7 2 2 63748 83213
0 9069 5 1 1 92101
0 9070 7 2 2 86489 85426
0 9071 5 1 1 92103
0 9072 7 1 2 9069 9071
0 9073 5 1 1 9072
0 9074 7 1 2 69422 9073
0 9075 5 1 1 9074
0 9076 7 2 2 73378 76292
0 9077 5 1 1 92105
0 9078 7 1 2 9077 9038
0 9079 5 1 1 9078
0 9080 7 1 2 85215 9079
0 9081 5 1 1 9080
0 9082 7 1 2 9075 9081
0 9083 5 1 1 9082
0 9084 7 1 2 72971 9083
0 9085 5 1 1 9084
0 9086 7 1 2 84078 82166
0 9087 5 1 1 9086
0 9088 7 7 2 73379 76557
0 9089 5 1 1 92107
0 9090 7 1 2 67952 92108
0 9091 5 1 1 9090
0 9092 7 1 2 9087 9091
0 9093 5 1 1 9092
0 9094 7 1 2 85216 9093
0 9095 5 1 1 9094
0 9096 7 1 2 9085 9095
0 9097 5 1 1 9096
0 9098 7 1 2 88135 9097
0 9099 5 1 1 9098
0 9100 7 1 2 9067 9099
0 9101 5 1 1 9100
0 9102 7 1 2 88954 9101
0 9103 5 1 1 9102
0 9104 7 1 2 91869 83559
0 9105 5 1 1 9104
0 9106 7 1 2 85217 82961
0 9107 5 1 1 9106
0 9108 7 1 2 72972 9107
0 9109 7 1 2 9105 9108
0 9110 5 1 1 9109
0 9111 7 1 2 85869 86250
0 9112 5 2 1 9111
0 9113 7 1 2 67953 92114
0 9114 5 1 1 9113
0 9115 7 1 2 76457 9114
0 9116 7 1 2 9110 9115
0 9117 5 1 1 9116
0 9118 7 1 2 85218 74886
0 9119 7 1 2 83257 9118
0 9120 5 1 1 9119
0 9121 7 1 2 9117 9120
0 9122 5 1 1 9121
0 9123 7 29 2 71911 67066
0 9124 7 6 2 70659 87952
0 9125 7 3 2 63876 89504
0 9126 5 1 1 92151
0 9127 7 3 2 92145 92152
0 9128 7 1 2 92116 92154
0 9129 7 1 2 9122 9128
0 9130 5 1 1 9129
0 9131 7 1 2 67559 9130
0 9132 7 1 2 9103 9131
0 9133 7 1 2 9014 9132
0 9134 5 1 1 9133
0 9135 7 1 2 70999 9134
0 9136 7 1 2 8924 9135
0 9137 5 1 1 9136
0 9138 7 1 2 67560 90680
0 9139 5 1 1 9138
0 9140 7 1 2 77109 81961
0 9141 5 1 1 9140
0 9142 7 1 2 78443 9141
0 9143 5 1 1 9142
0 9144 7 1 2 69750 9143
0 9145 5 1 1 9144
0 9146 7 1 2 9139 9145
0 9147 5 1 1 9146
0 9148 7 1 2 85870 9147
0 9149 5 1 1 9148
0 9150 7 5 2 66949 90645
0 9151 7 1 2 92157 82187
0 9152 5 1 1 9151
0 9153 7 1 2 9149 9152
0 9154 5 1 1 9153
0 9155 7 1 2 68308 9154
0 9156 5 1 1 9155
0 9157 7 5 2 70116 80074
0 9158 5 5 1 92162
0 9159 7 3 2 71303 87696
0 9160 5 2 1 92172
0 9161 7 1 2 92167 92175
0 9162 5 2 1 9161
0 9163 7 4 2 67561 85219
0 9164 7 1 2 92177 92179
0 9165 5 1 1 9164
0 9166 7 1 2 9156 9165
0 9167 5 1 1 9166
0 9168 7 1 2 72973 9167
0 9169 5 1 1 9168
0 9170 7 2 2 87240 81554
0 9171 7 2 2 69751 92183
0 9172 5 1 1 92185
0 9173 7 1 2 90669 92186
0 9174 5 1 1 9173
0 9175 7 1 2 9169 9174
0 9176 5 1 1 9175
0 9177 7 1 2 88520 9176
0 9178 5 1 1 9177
0 9179 7 1 2 79190 92180
0 9180 5 1 1 9179
0 9181 7 8 2 72974 82188
0 9182 5 3 1 92187
0 9183 7 1 2 84109 92195
0 9184 5 4 1 9183
0 9185 7 4 2 70117 83111
0 9186 7 1 2 90729 92202
0 9187 7 1 2 92198 9186
0 9188 5 1 1 9187
0 9189 7 1 2 9180 9188
0 9190 5 1 1 9189
0 9191 7 1 2 88136 9190
0 9192 5 1 1 9191
0 9193 7 1 2 9178 9192
0 9194 5 1 1 9193
0 9195 7 1 2 71779 9194
0 9196 5 1 1 9195
0 9197 7 2 2 63749 79084
0 9198 7 1 2 84045 91236
0 9199 7 1 2 92206 9198
0 9200 5 1 1 9199
0 9201 7 3 2 65324 89187
0 9202 5 1 1 92208
0 9203 7 1 2 89322 9202
0 9204 5 1 1 9203
0 9205 7 1 2 70118 92199
0 9206 7 1 2 9204 9205
0 9207 5 1 1 9206
0 9208 7 1 2 9200 9207
0 9209 5 1 1 9208
0 9210 7 1 2 73898 9209
0 9211 5 1 1 9210
0 9212 7 3 2 84418 78721
0 9213 7 1 2 82756 92211
0 9214 7 1 2 92106 9213
0 9215 5 1 1 9214
0 9216 7 1 2 9211 9215
0 9217 7 1 2 9196 9216
0 9218 5 1 1 9217
0 9219 7 1 2 88955 9218
0 9220 5 1 1 9219
0 9221 7 1 2 90403 89599
0 9222 5 1 1 9221
0 9223 7 1 2 6659 9222
0 9224 5 1 1 9223
0 9225 7 1 2 77919 9224
0 9226 5 1 1 9225
0 9227 7 1 2 71304 77722
0 9228 7 1 2 79042 9227
0 9229 5 1 1 9228
0 9230 7 1 2 9226 9229
0 9231 5 1 1 9230
0 9232 7 3 2 91892 91800
0 9233 7 1 2 87787 75732
0 9234 7 1 2 92214 9233
0 9235 7 1 2 9231 9234
0 9236 5 1 1 9235
0 9237 7 1 2 9220 9236
0 9238 5 1 1 9237
0 9239 7 1 2 69423 9238
0 9240 5 1 1 9239
0 9241 7 1 2 89415 78892
0 9242 5 1 1 9241
0 9243 7 2 2 68790 74897
0 9244 7 1 2 82378 79050
0 9245 7 1 2 92217 9244
0 9246 5 1 1 9245
0 9247 7 1 2 9242 9246
0 9248 5 1 1 9247
0 9249 7 1 2 71780 9248
0 9250 5 1 1 9249
0 9251 7 7 2 68309 85871
0 9252 7 1 2 65325 87665
0 9253 7 1 2 92219 9252
0 9254 5 1 1 9253
0 9255 7 1 2 9250 9254
0 9256 5 1 1 9255
0 9257 7 7 2 65680 90576
0 9258 7 9 2 66848 67067
0 9259 7 1 2 92233 90284
0 9260 7 4 2 92226 9259
0 9261 5 1 1 92242
0 9262 7 1 2 78393 92243
0 9263 7 1 2 9256 9262
0 9264 5 1 1 9263
0 9265 7 1 2 9240 9264
0 9266 7 1 2 9137 9265
0 9267 7 1 2 8592 9266
0 9268 5 1 1 9267
0 9269 7 1 2 64030 9268
0 9270 5 1 1 9269
0 9271 7 1 2 78684 83672
0 9272 5 1 1 9271
0 9273 7 3 2 77604 9272
0 9274 7 1 2 92246 84729
0 9275 5 1 1 9274
0 9276 7 1 2 84720 91944
0 9277 5 1 1 9276
0 9278 7 1 2 9275 9277
0 9279 5 1 1 9278
0 9280 7 1 2 65002 9279
0 9281 5 1 1 9280
0 9282 7 1 2 73899 84994
0 9283 5 3 1 9282
0 9284 7 9 2 73380 87788
0 9285 5 1 1 92252
0 9286 7 1 2 92249 9285
0 9287 5 2 1 9286
0 9288 7 1 2 70119 92261
0 9289 5 1 1 9288
0 9290 7 1 2 2800 9289
0 9291 5 1 1 9290
0 9292 7 1 2 68601 9291
0 9293 5 1 1 9292
0 9294 7 1 2 68310 91456
0 9295 5 1 1 9294
0 9296 7 1 2 9293 9295
0 9297 5 1 1 9296
0 9298 7 1 2 71781 9297
0 9299 5 1 1 9298
0 9300 7 6 2 66472 67562
0 9301 7 1 2 92263 88807
0 9302 5 1 1 9301
0 9303 7 1 2 9299 9302
0 9304 5 1 1 9303
0 9305 7 1 2 69424 9304
0 9306 5 1 1 9305
0 9307 7 2 2 89272 91124
0 9308 5 1 1 92269
0 9309 7 2 2 67563 92270
0 9310 5 1 1 92271
0 9311 7 1 2 71782 92272
0 9312 5 1 1 9311
0 9313 7 1 2 9306 9312
0 9314 5 1 1 9313
0 9315 7 1 2 82535 9314
0 9316 5 1 1 9315
0 9317 7 1 2 9281 9316
0 9318 5 1 1 9317
0 9319 7 9 2 63750 63963
0 9320 7 2 2 76914 92273
0 9321 7 4 2 66849 89535
0 9322 7 1 2 74099 92284
0 9323 7 1 2 92282 9322
0 9324 7 1 2 9318 9323
0 9325 5 1 1 9324
0 9326 7 1 2 9270 9325
0 9327 7 1 2 8343 9326
0 9328 5 1 1 9327
0 9329 7 1 2 65721 9328
0 9330 5 1 1 9329
0 9331 7 2 2 64301 78404
0 9332 5 3 1 92288
0 9333 7 1 2 82555 92290
0 9334 5 2 1 9333
0 9335 7 2 2 79652 91531
0 9336 7 3 2 86563 92295
0 9337 7 1 2 92293 92297
0 9338 5 1 1 9337
0 9339 7 11 2 71912 72017
0 9340 7 7 2 68791 69055
0 9341 7 1 2 92300 92311
0 9342 7 2 2 84662 9341
0 9343 7 1 2 74055 91691
0 9344 7 1 2 92318 9343
0 9345 5 1 1 9344
0 9346 7 1 2 9338 9345
0 9347 5 1 1 9346
0 9348 7 1 2 76458 9347
0 9349 5 1 1 9348
0 9350 7 2 2 66950 89536
0 9351 7 2 2 79445 91720
0 9352 7 1 2 82189 74310
0 9353 7 1 2 92322 9352
0 9354 7 2 2 92320 9353
0 9355 5 1 1 92324
0 9356 7 2 2 69425 92325
0 9357 5 1 1 92326
0 9358 7 1 2 73688 92327
0 9359 5 1 1 9358
0 9360 7 1 2 9349 9359
0 9361 5 1 1 9360
0 9362 7 1 2 64031 9361
0 9363 5 1 1 9362
0 9364 7 2 2 76459 74056
0 9365 5 2 1 92328
0 9366 7 1 2 92330 77853
0 9367 5 3 1 9366
0 9368 7 1 2 84933 92332
0 9369 5 1 1 9368
0 9370 7 9 2 64628 65722
0 9371 7 1 2 92335 82190
0 9372 7 1 2 80985 9371
0 9373 5 1 1 9372
0 9374 7 1 2 9369 9373
0 9375 5 1 1 9374
0 9376 7 1 2 92298 9375
0 9377 5 1 1 9376
0 9378 7 1 2 9363 9377
0 9379 5 1 1 9378
0 9380 7 1 2 84538 9379
0 9381 5 1 1 9380
0 9382 7 14 2 67564 68311
0 9383 7 4 2 73689 92344
0 9384 7 7 2 71000 66473
0 9385 7 1 2 92362 78527
0 9386 7 1 2 92358 9385
0 9387 7 1 2 78911 9386
0 9388 7 1 2 90332 9387
0 9389 5 1 1 9388
0 9390 7 1 2 9381 9389
0 9391 5 1 1 9390
0 9392 7 1 2 88521 9391
0 9393 5 1 1 9392
0 9394 7 1 2 64302 92274
0 9395 7 2 2 90417 9394
0 9396 7 3 2 66850 68312
0 9397 7 3 2 88306 92371
0 9398 7 1 2 92369 92374
0 9399 5 1 1 9398
0 9400 7 10 2 69752 65723
0 9401 7 1 2 73381 84482
0 9402 7 1 2 92377 9401
0 9403 7 1 2 90389 9402
0 9404 5 1 1 9403
0 9405 7 1 2 9399 9404
0 9406 5 1 1 9405
0 9407 7 1 2 71001 9406
0 9408 5 1 1 9407
0 9409 7 1 2 65937 79627
0 9410 7 1 2 89537 90596
0 9411 7 1 2 9409 9410
0 9412 7 1 2 92375 9411
0 9413 5 1 1 9412
0 9414 7 1 2 9408 9413
0 9415 5 1 1 9414
0 9416 7 1 2 72975 9415
0 9417 5 1 1 9416
0 9418 7 3 2 65724 74942
0 9419 5 1 1 92387
0 9420 7 3 2 74144 80011
0 9421 5 2 1 92390
0 9422 7 1 2 64303 77585
0 9423 7 1 2 89451 9422
0 9424 5 1 1 9423
0 9425 7 2 2 92393 9424
0 9426 5 1 1 92395
0 9427 7 1 2 9419 92396
0 9428 5 1 1 9427
0 9429 7 1 2 76674 92296
0 9430 7 1 2 9428 9429
0 9431 5 1 1 9430
0 9432 7 1 2 9417 9431
0 9433 5 1 1 9432
0 9434 7 1 2 66474 9433
0 9435 5 1 1 9434
0 9436 7 2 2 75551 90390
0 9437 7 7 2 64629 71588
0 9438 5 1 1 92399
0 9439 7 10 2 65725 66193
0 9440 7 1 2 92400 92406
0 9441 7 1 2 91632 9440
0 9442 7 1 2 92397 9441
0 9443 5 1 1 9442
0 9444 7 1 2 9435 9443
0 9445 5 1 1 9444
0 9446 7 1 2 67565 9445
0 9447 5 1 1 9446
0 9448 7 8 2 65726 71589
0 9449 7 1 2 92416 91633
0 9450 7 1 2 84098 9449
0 9451 7 1 2 92398 9450
0 9452 5 1 1 9451
0 9453 7 1 2 9447 9452
0 9454 5 1 1 9453
0 9455 7 1 2 64032 9454
0 9456 5 1 1 9455
0 9457 7 2 2 79465 81206
0 9458 5 2 1 92424
0 9459 7 3 2 75002 81016
0 9460 7 1 2 79181 92428
0 9461 5 2 1 9460
0 9462 7 1 2 92426 92431
0 9463 5 1 1 9462
0 9464 7 4 2 90577 90657
0 9465 7 10 2 65681 65727
0 9466 7 1 2 92275 92437
0 9467 7 1 2 92433 9466
0 9468 7 1 2 92359 9467
0 9469 7 1 2 9463 9468
0 9470 5 1 1 9469
0 9471 7 1 2 9456 9470
0 9472 5 1 1 9471
0 9473 7 1 2 66951 9472
0 9474 5 1 1 9473
0 9475 7 1 2 71002 79257
0 9476 5 1 1 9475
0 9477 7 1 2 3044 9476
0 9478 5 1 1 9477
0 9479 7 8 2 69056 64033
0 9480 7 3 2 68792 92447
0 9481 7 2 2 92301 91644
0 9482 7 2 2 92455 92458
0 9483 7 5 2 65728 66475
0 9484 7 1 2 92462 92360
0 9485 7 1 2 92460 9484
0 9486 7 1 2 9478 9485
0 9487 5 1 1 9486
0 9488 7 1 2 9474 9487
0 9489 5 1 1 9488
0 9490 7 1 2 88137 9489
0 9491 5 1 1 9490
0 9492 7 1 2 9393 9491
0 9493 5 1 1 9492
0 9494 7 1 2 65003 9493
0 9495 5 1 1 9494
0 9496 7 3 2 78158 90743
0 9497 7 4 2 90605 92467
0 9498 5 2 1 92470
0 9499 7 5 2 68793 87953
0 9500 7 2 2 92476 90248
0 9501 7 3 2 92302 92481
0 9502 7 1 2 71003 92483
0 9503 5 1 1 9502
0 9504 7 1 2 92474 9503
0 9505 5 1 1 9504
0 9506 7 1 2 83408 74773
0 9507 7 1 2 9505 9506
0 9508 5 1 1 9507
0 9509 7 3 2 75733 81017
0 9510 7 1 2 88441 92486
0 9511 7 1 2 90391 9510
0 9512 5 1 1 9511
0 9513 7 1 2 9508 9512
0 9514 5 1 1 9513
0 9515 7 1 2 71305 9514
0 9516 5 1 1 9515
0 9517 7 2 2 73949 90392
0 9518 7 5 2 69426 71913
0 9519 7 2 2 86388 92491
0 9520 7 1 2 79958 92496
0 9521 7 1 2 92489 9520
0 9522 5 1 1 9521
0 9523 7 1 2 9516 9522
0 9524 5 1 1 9523
0 9525 7 1 2 67566 9524
0 9526 5 1 1 9525
0 9527 7 4 2 67954 84483
0 9528 7 1 2 77138 78359
0 9529 7 1 2 92498 9528
0 9530 7 1 2 92490 9529
0 9531 5 1 1 9530
0 9532 7 1 2 9526 9531
0 9533 5 1 1 9532
0 9534 7 1 2 65729 9533
0 9535 5 1 1 9534
0 9536 7 2 2 71306 77408
0 9537 5 2 1 92502
0 9538 7 1 2 92323 92361
0 9539 7 1 2 92504 9538
0 9540 7 1 2 75003 81003
0 9541 5 1 1 9540
0 9542 7 7 2 66851 66952
0 9543 7 2 2 92506 89538
0 9544 7 1 2 2145 92513
0 9545 7 1 2 9541 9544
0 9546 7 1 2 9539 9545
0 9547 5 1 1 9546
0 9548 7 1 2 9535 9547
0 9549 5 1 1 9548
0 9550 7 1 2 88138 9549
0 9551 5 1 1 9550
0 9552 7 3 2 68313 90333
0 9553 7 3 2 68960 76194
0 9554 7 1 2 76898 92518
0 9555 7 1 2 85385 9554
0 9556 7 1 2 92515 9555
0 9557 5 1 1 9556
0 9558 7 1 2 9551 9557
0 9559 5 1 1 9558
0 9560 7 1 2 64034 9559
0 9561 5 1 1 9560
0 9562 7 6 2 76195 77316
0 9563 7 2 2 92521 88911
0 9564 7 3 2 73382 74418
0 9565 5 1 1 92529
0 9566 7 1 2 90578 91063
0 9567 7 1 2 92530 9566
0 9568 7 1 2 92527 9567
0 9569 5 1 1 9568
0 9570 7 2 2 64035 89569
0 9571 7 1 2 77205 79959
0 9572 5 2 1 9571
0 9573 7 5 2 65730 77409
0 9574 5 1 1 92536
0 9575 7 1 2 76353 92537
0 9576 7 1 2 92534 9575
0 9577 7 1 2 92532 9576
0 9578 5 1 1 9577
0 9579 7 1 2 9569 9578
0 9580 5 1 1 9579
0 9581 7 1 2 72576 9580
0 9582 5 1 1 9581
0 9583 7 2 2 89570 80954
0 9584 7 1 2 76354 78534
0 9585 7 1 2 92541 9584
0 9586 5 1 1 9585
0 9587 7 1 2 9582 9586
0 9588 5 1 1 9587
0 9589 7 1 2 63751 9588
0 9590 5 1 1 9589
0 9591 7 1 2 77410 90777
0 9592 5 1 1 9591
0 9593 7 8 2 72577 77139
0 9594 5 4 1 92543
0 9595 7 1 2 78432 80174
0 9596 5 1 1 9595
0 9597 7 1 2 92551 9596
0 9598 7 1 2 9592 9597
0 9599 5 1 1 9598
0 9600 7 4 2 64036 65582
0 9601 7 4 2 68794 92555
0 9602 7 4 2 90312 92559
0 9603 7 5 2 65731 68314
0 9604 7 1 2 72018 92567
0 9605 7 1 2 92563 9604
0 9606 7 1 2 9599 9605
0 9607 5 1 1 9606
0 9608 7 1 2 9590 9607
0 9609 5 1 1 9608
0 9610 7 1 2 67068 75663
0 9611 7 1 2 9609 9610
0 9612 5 1 1 9611
0 9613 7 2 2 83258 78506
0 9614 5 1 1 92572
0 9615 7 1 2 84441 89920
0 9616 7 1 2 90393 9615
0 9617 7 1 2 92573 9616
0 9618 5 1 1 9617
0 9619 7 1 2 9612 9618
0 9620 5 1 1 9619
0 9621 7 1 2 75352 9620
0 9622 5 1 1 9621
0 9623 7 11 2 72578 73383
0 9624 7 2 2 92574 91064
0 9625 7 2 2 67069 92585
0 9626 7 1 2 65732 91146
0 9627 7 1 2 92276 9626
0 9628 7 2 2 81130 86195
0 9629 7 3 2 65682 71004
0 9630 7 3 2 90579 92591
0 9631 7 1 2 92589 92594
0 9632 7 1 2 9627 9631
0 9633 7 1 2 92587 9632
0 9634 5 1 1 9633
0 9635 7 1 2 9622 9634
0 9636 5 1 1 9635
0 9637 7 1 2 68602 9636
0 9638 5 1 1 9637
0 9639 7 5 2 67955 76675
0 9640 7 1 2 82525 76008
0 9641 7 1 2 92597 9640
0 9642 7 2 2 84419 86196
0 9643 7 2 2 91147 92277
0 9644 7 4 2 65627 92438
0 9645 7 1 2 92604 92606
0 9646 7 1 2 92602 9645
0 9647 7 1 2 9641 9646
0 9648 5 1 1 9647
0 9649 7 1 2 9638 9648
0 9650 7 1 2 9561 9649
0 9651 7 1 2 9495 9650
0 9652 5 1 1 9651
0 9653 7 1 2 84816 9652
0 9654 5 1 1 9653
0 9655 7 10 2 72126 75999
0 9656 5 1 1 92610
0 9657 7 1 2 88288 9656
0 9658 5 6 1 9657
0 9659 7 1 2 92620 78531
0 9660 5 1 1 9659
0 9661 7 1 2 78893 85062
0 9662 5 1 1 9661
0 9663 7 9 2 65004 67567
0 9664 7 3 2 77866 92626
0 9665 5 3 1 92635
0 9666 7 1 2 69753 84995
0 9667 5 3 1 9666
0 9668 7 1 2 92638 92641
0 9669 5 1 1 9668
0 9670 7 1 2 71307 9669
0 9671 5 1 1 9670
0 9672 7 7 2 67956 75260
0 9673 7 1 2 78146 92644
0 9674 5 1 1 9673
0 9675 7 1 2 9671 9674
0 9676 5 1 1 9675
0 9677 7 1 2 73384 9676
0 9678 5 1 1 9677
0 9679 7 1 2 9662 9678
0 9680 5 1 1 9679
0 9681 7 1 2 88522 9680
0 9682 5 1 1 9681
0 9683 7 2 2 72579 87210
0 9684 5 1 1 92651
0 9685 7 1 2 76558 89245
0 9686 5 1 1 9685
0 9687 7 1 2 9684 9686
0 9688 5 1 1 9687
0 9689 7 1 2 67957 9688
0 9690 5 1 1 9689
0 9691 7 1 2 86260 92200
0 9692 5 1 1 9691
0 9693 7 1 2 79572 92253
0 9694 5 1 1 9693
0 9695 7 4 2 74523 76293
0 9696 7 1 2 81410 92653
0 9697 5 1 1 9696
0 9698 7 1 2 9694 9697
0 9699 7 1 2 9692 9698
0 9700 7 1 2 9690 9699
0 9701 5 1 1 9700
0 9702 7 1 2 88139 9701
0 9703 5 1 1 9702
0 9704 7 1 2 9682 9703
0 9705 5 1 1 9704
0 9706 7 1 2 75096 9705
0 9707 5 1 1 9706
0 9708 7 2 2 79227 85063
0 9709 5 1 1 92657
0 9710 7 1 2 82162 9709
0 9711 5 1 1 9710
0 9712 7 1 2 65005 9711
0 9713 5 1 1 9712
0 9714 7 1 2 67958 79304
0 9715 5 1 1 9714
0 9716 7 2 2 72976 79501
0 9717 5 2 1 92659
0 9718 7 16 2 69754 72580
0 9719 5 1 1 92663
0 9720 7 1 2 92661 92664
0 9721 7 1 2 9715 9720
0 9722 5 1 1 9721
0 9723 7 1 2 9713 9722
0 9724 5 2 1 9723
0 9725 7 1 2 88523 92679
0 9726 5 1 1 9725
0 9727 7 1 2 9707 9726
0 9728 5 1 1 9727
0 9729 7 1 2 69427 9728
0 9730 5 1 1 9729
0 9731 7 2 2 63877 74898
0 9732 7 1 2 89161 92681
0 9733 5 1 1 9732
0 9734 7 1 2 83617 90980
0 9735 5 1 1 9734
0 9736 7 1 2 9733 9735
0 9737 5 1 1 9736
0 9738 7 1 2 72977 9737
0 9739 5 1 1 9738
0 9740 7 3 2 78685 88140
0 9741 5 1 1 92683
0 9742 7 1 2 6390 9741
0 9743 5 1 1 9742
0 9744 7 1 2 75097 9743
0 9745 5 1 1 9744
0 9746 7 10 2 73385 88524
0 9747 7 1 2 87375 92686
0 9748 5 1 1 9747
0 9749 7 1 2 9745 9748
0 9750 5 1 1 9749
0 9751 7 1 2 64304 9750
0 9752 5 1 1 9751
0 9753 7 1 2 9739 9752
0 9754 5 1 1 9753
0 9755 7 1 2 69755 9754
0 9756 5 1 1 9755
0 9757 7 7 2 68315 88525
0 9758 5 1 1 92696
0 9759 7 1 2 92697 75493
0 9760 5 1 1 9759
0 9761 7 2 2 75098 90639
0 9762 5 2 1 92703
0 9763 7 1 2 9760 92705
0 9764 5 1 1 9763
0 9765 7 1 2 81207 9764
0 9766 5 1 1 9765
0 9767 7 1 2 9756 9766
0 9768 5 1 1 9767
0 9769 7 1 2 71308 9768
0 9770 5 1 1 9769
0 9771 7 2 2 77723 90025
0 9772 5 1 1 92707
0 9773 7 1 2 9772 92706
0 9774 5 1 1 9773
0 9775 7 2 2 82723 9774
0 9776 5 1 1 92709
0 9777 7 1 2 64305 92710
0 9778 5 1 1 9777
0 9779 7 1 2 9770 9778
0 9780 5 1 1 9779
0 9781 7 1 2 67568 9780
0 9782 5 1 1 9781
0 9783 7 1 2 9730 9782
0 9784 5 1 1 9783
0 9785 7 1 2 71005 9784
0 9786 5 1 1 9785
0 9787 7 1 2 65326 89101
0 9788 5 1 1 9787
0 9789 7 1 2 8957 9788
0 9790 5 1 1 9789
0 9791 7 1 2 69756 9790
0 9792 5 1 1 9791
0 9793 7 1 2 90549 75494
0 9794 5 1 1 9793
0 9795 7 1 2 9792 9794
0 9796 5 1 1 9795
0 9797 7 1 2 68316 9796
0 9798 5 1 1 9797
0 9799 7 1 2 75624 92704
0 9800 5 1 1 9799
0 9801 7 1 2 9798 9800
0 9802 5 1 1 9801
0 9803 7 1 2 71309 9802
0 9804 5 1 1 9803
0 9805 7 1 2 9776 9804
0 9806 5 1 1 9805
0 9807 7 1 2 65938 9806
0 9808 5 1 1 9807
0 9809 7 3 2 71310 74899
0 9810 7 1 2 66476 92711
0 9811 7 3 2 67070 79085
0 9812 5 1 1 92714
0 9813 7 1 2 90185 92715
0 9814 7 1 2 9810 9813
0 9815 5 1 1 9814
0 9816 7 1 2 9808 9815
0 9817 5 1 1 9816
0 9818 7 1 2 90860 9817
0 9819 5 1 1 9818
0 9820 7 1 2 9786 9819
0 9821 5 1 1 9820
0 9822 7 1 2 85182 9821
0 9823 5 1 1 9822
0 9824 7 1 2 9660 9823
0 9825 5 1 1 9824
0 9826 7 1 2 66668 9825
0 9827 5 1 1 9826
0 9828 7 1 2 83282 89824
0 9829 5 1 1 9828
0 9830 7 1 2 68317 89981
0 9831 7 1 2 78912 9830
0 9832 5 1 1 9831
0 9833 7 1 2 9829 9832
0 9834 5 1 1 9833
0 9835 7 1 2 74616 9834
0 9836 5 1 1 9835
0 9837 7 1 2 89982 78945
0 9838 5 1 1 9837
0 9839 7 1 2 9836 9838
0 9840 5 1 1 9839
0 9841 7 1 2 67569 9840
0 9842 5 1 1 9841
0 9843 7 1 2 71590 81551
0 9844 5 1 1 9843
0 9845 7 1 2 69428 77931
0 9846 5 1 1 9845
0 9847 7 1 2 9844 9846
0 9848 5 1 1 9847
0 9849 7 1 2 70120 9848
0 9850 5 1 1 9849
0 9851 7 1 2 69429 84213
0 9852 5 1 1 9851
0 9853 7 1 2 9850 9852
0 9854 5 1 1 9853
0 9855 7 1 2 68961 91481
0 9856 7 1 2 9854 9855
0 9857 5 1 1 9856
0 9858 7 1 2 9842 9857
0 9859 5 1 1 9858
0 9860 7 1 2 71006 9859
0 9861 5 1 1 9860
0 9862 7 1 2 72581 90739
0 9863 7 1 2 81635 9862
0 9864 5 1 1 9863
0 9865 7 1 2 9861 9864
0 9866 5 1 1 9865
0 9867 7 1 2 73690 9866
0 9868 5 1 1 9867
0 9869 7 5 2 64630 82191
0 9870 5 2 1 92717
0 9871 7 1 2 92722 87779
0 9872 5 2 1 9871
0 9873 7 2 2 69430 92724
0 9874 5 2 1 92726
0 9875 7 1 2 78444 81492
0 9876 5 2 1 9875
0 9877 7 1 2 77131 92730
0 9878 5 1 1 9877
0 9879 7 1 2 92728 9878
0 9880 5 1 1 9879
0 9881 7 1 2 67959 77306
0 9882 7 1 2 9880 9881
0 9883 5 1 1 9882
0 9884 7 1 2 74524 84183
0 9885 7 1 2 81337 9884
0 9886 5 1 1 9885
0 9887 7 1 2 9883 9886
0 9888 5 1 1 9887
0 9889 7 1 2 68318 9888
0 9890 5 1 1 9889
0 9891 7 2 2 70121 77292
0 9892 5 2 1 92732
0 9893 7 2 2 77095 92734
0 9894 5 4 1 92736
0 9895 7 2 2 84282 92738
0 9896 7 1 2 82053 92742
0 9897 5 1 1 9896
0 9898 7 1 2 79573 91442
0 9899 5 3 1 9898
0 9900 7 2 2 77083 75056
0 9901 5 1 1 92747
0 9902 7 1 2 70122 92748
0 9903 5 1 1 9902
0 9904 7 1 2 92744 9903
0 9905 5 2 1 9904
0 9906 7 1 2 87789 92749
0 9907 5 1 1 9906
0 9908 7 10 2 72582 75552
0 9909 5 1 1 92751
0 9910 7 1 2 77307 80266
0 9911 5 1 1 9910
0 9912 7 1 2 77133 9911
0 9913 5 1 1 9912
0 9914 7 1 2 92752 9913
0 9915 5 1 1 9914
0 9916 7 1 2 9907 9915
0 9917 5 1 1 9916
0 9918 7 1 2 71007 9917
0 9919 5 1 1 9918
0 9920 7 1 2 9897 9919
0 9921 7 1 2 9890 9920
0 9922 5 1 1 9921
0 9923 7 1 2 92611 9922
0 9924 5 1 1 9923
0 9925 7 16 2 69757 65939
0 9926 7 6 2 71311 92761
0 9927 5 1 1 92777
0 9928 7 1 2 92345 92778
0 9929 5 2 1 9928
0 9930 7 1 2 90808 78059
0 9931 5 1 1 9930
0 9932 7 1 2 92783 9931
0 9933 5 1 1 9932
0 9934 7 1 2 67960 9933
0 9935 5 1 1 9934
0 9936 7 1 2 67570 79442
0 9937 5 1 1 9936
0 9938 7 4 2 71312 76953
0 9939 5 2 1 92785
0 9940 7 1 2 72583 92789
0 9941 7 1 2 8156 9940
0 9942 5 1 1 9941
0 9943 7 1 2 71008 9942
0 9944 7 1 2 9937 9943
0 9945 5 1 1 9944
0 9946 7 1 2 9935 9945
0 9947 5 1 1 9946
0 9948 7 1 2 88141 9947
0 9949 5 1 1 9948
0 9950 7 1 2 9924 9949
0 9951 7 1 2 9868 9950
0 9952 5 1 1 9951
0 9953 7 1 2 74374 9952
0 9954 5 1 1 9953
0 9955 7 1 2 74341 83642
0 9956 7 2 2 65940 91237
0 9957 7 1 2 74203 92791
0 9958 7 1 2 9955 9957
0 9959 5 1 1 9958
0 9960 7 6 2 74617 88526
0 9961 7 1 2 80242 92793
0 9962 5 1 1 9961
0 9963 7 1 2 75041 89983
0 9964 5 1 1 9963
0 9965 7 1 2 9962 9964
0 9966 5 1 1 9965
0 9967 7 1 2 76196 9966
0 9968 5 1 1 9967
0 9969 7 2 2 63878 75502
0 9970 7 3 2 67071 76559
0 9971 7 1 2 78628 92801
0 9972 7 1 2 92799 9971
0 9973 5 1 1 9972
0 9974 7 1 2 9968 9973
0 9975 5 1 1 9974
0 9976 7 1 2 82237 78299
0 9977 7 1 2 9975 9976
0 9978 5 1 1 9977
0 9979 7 1 2 9959 9978
0 9980 7 1 2 9954 9979
0 9981 5 1 1 9980
0 9982 7 1 2 66669 9981
0 9983 5 1 1 9982
0 9984 7 7 2 64037 67571
0 9985 5 2 1 92804
0 9986 7 4 2 69431 74057
0 9987 5 1 1 92813
0 9988 7 1 2 92805 92814
0 9989 5 2 1 9988
0 9990 7 13 2 69099 65006
0 9991 5 1 1 92819
0 9992 7 2 2 92820 85391
0 9993 7 1 2 78629 92832
0 9994 5 1 1 9993
0 9995 7 1 2 92817 9994
0 9996 5 1 1 9995
0 9997 7 1 2 89289 9996
0 9998 5 1 1 9997
0 9999 7 2 2 82344 82214
0 10000 7 11 2 70123 65733
0 10001 7 3 2 69432 92836
0 10002 7 7 2 72127 84316
0 10003 7 1 2 92847 92850
0 10004 7 1 2 92834 10003
0 10005 5 1 1 10004
0 10006 7 1 2 9998 10005
0 10007 5 1 1 10006
0 10008 7 1 2 66194 10007
0 10009 5 1 1 10008
0 10010 7 1 2 79922 82542
0 10011 7 8 2 64038 72128
0 10012 7 1 2 92857 85403
0 10013 7 1 2 10010 10012
0 10014 5 1 1 10013
0 10015 7 1 2 10009 10014
0 10016 5 1 1 10015
0 10017 7 1 2 75600 10016
0 10018 5 1 1 10017
0 10019 7 7 2 71009 73386
0 10020 7 2 2 79274 85074
0 10021 5 1 1 92872
0 10022 7 1 2 80340 75353
0 10023 5 1 1 10022
0 10024 7 1 2 76560 10023
0 10025 5 1 1 10024
0 10026 7 1 2 69433 89233
0 10027 7 1 2 10025 10026
0 10028 5 1 1 10027
0 10029 7 1 2 10021 10028
0 10030 5 1 1 10029
0 10031 7 1 2 92865 10030
0 10032 5 1 1 10031
0 10033 7 2 2 80012 82192
0 10034 5 2 1 92874
0 10035 7 3 2 72584 80277
0 10036 5 2 1 92878
0 10037 7 2 2 68603 92879
0 10038 5 1 1 92883
0 10039 7 1 2 92876 10038
0 10040 5 1 1 10039
0 10041 7 1 2 81499 10040
0 10042 5 1 1 10041
0 10043 7 1 2 65007 92725
0 10044 5 1 1 10043
0 10045 7 1 2 76561 84663
0 10046 5 1 1 10045
0 10047 7 1 2 80887 84099
0 10048 5 1 1 10047
0 10049 7 1 2 10046 10048
0 10050 7 1 2 10044 10049
0 10051 5 1 1 10050
0 10052 7 1 2 71010 10051
0 10053 5 1 1 10052
0 10054 7 1 2 84100 80986
0 10055 5 4 1 10054
0 10056 7 1 2 67572 81997
0 10057 5 1 1 10056
0 10058 7 1 2 92885 10057
0 10059 7 1 2 10053 10058
0 10060 5 1 1 10059
0 10061 7 1 2 68319 10060
0 10062 5 1 1 10061
0 10063 7 1 2 10042 10062
0 10064 5 1 1 10063
0 10065 7 1 2 71783 10064
0 10066 5 1 1 10065
0 10067 7 3 2 73387 78507
0 10068 7 1 2 76294 92889
0 10069 5 1 1 10068
0 10070 7 1 2 67961 10069
0 10071 7 1 2 10066 10070
0 10072 5 1 1 10071
0 10073 7 9 2 67573 81018
0 10074 5 2 1 92892
0 10075 7 1 2 68604 92544
0 10076 5 1 1 10075
0 10077 7 1 2 92901 10076
0 10078 5 1 1 10077
0 10079 7 1 2 76295 10078
0 10080 5 1 1 10079
0 10081 7 1 2 74525 92884
0 10082 5 1 1 10081
0 10083 7 1 2 10080 10082
0 10084 5 1 1 10083
0 10085 7 1 2 82345 10084
0 10086 5 1 1 10085
0 10087 7 2 2 73388 78474
0 10088 7 1 2 92745 83852
0 10089 5 1 1 10088
0 10090 7 1 2 92903 10089
0 10091 5 1 1 10090
0 10092 7 1 2 72978 10091
0 10093 7 1 2 10086 10092
0 10094 5 1 1 10093
0 10095 7 1 2 10072 10094
0 10096 5 1 1 10095
0 10097 7 1 2 10032 10096
0 10098 5 1 1 10097
0 10099 7 1 2 65734 92851
0 10100 7 1 2 10098 10099
0 10101 5 1 1 10100
0 10102 7 1 2 10018 10101
0 10103 7 1 2 9983 10102
0 10104 5 1 1 10103
0 10105 7 1 2 78202 10104
0 10106 5 1 1 10105
0 10107 7 1 2 66477 80436
0 10108 5 9 1 10107
0 10109 7 2 2 72979 92905
0 10110 5 2 1 92914
0 10111 7 1 2 66195 91754
0 10112 5 1 1 10111
0 10113 7 1 2 92915 10112
0 10114 5 1 1 10113
0 10115 7 3 2 71313 74618
0 10116 7 1 2 74730 92918
0 10117 5 1 1 10116
0 10118 7 1 2 10114 10117
0 10119 5 1 1 10118
0 10120 7 1 2 69758 10119
0 10121 5 1 1 10120
0 10122 7 1 2 90699 78968
0 10123 5 1 1 10122
0 10124 7 1 2 83357 10123
0 10125 7 1 2 10121 10124
0 10126 5 1 1 10125
0 10127 7 1 2 72585 10126
0 10128 5 1 1 10127
0 10129 7 1 2 65008 92658
0 10130 5 1 1 10129
0 10131 7 1 2 10128 10130
0 10132 5 1 1 10131
0 10133 7 1 2 69434 10132
0 10134 5 1 1 10133
0 10135 7 1 2 71314 91995
0 10136 5 1 1 10135
0 10137 7 9 2 69759 66196
0 10138 5 4 1 92921
0 10139 7 1 2 92922 75553
0 10140 5 2 1 10139
0 10141 7 1 2 74526 92013
0 10142 5 1 1 10141
0 10143 7 1 2 92934 10142
0 10144 7 1 2 10136 10143
0 10145 5 1 1 10144
0 10146 7 1 2 81522 10145
0 10147 5 1 1 10146
0 10148 7 1 2 10134 10147
0 10149 5 1 1 10148
0 10150 7 1 2 71011 10149
0 10151 5 1 1 10150
0 10152 7 5 2 67574 80987
0 10153 5 1 1 92936
0 10154 7 3 2 78797 78921
0 10155 5 4 1 92941
0 10156 7 1 2 83310 92944
0 10157 5 1 1 10156
0 10158 7 2 2 68320 10157
0 10159 5 1 1 92948
0 10160 7 1 2 80517 83267
0 10161 5 1 1 10160
0 10162 7 1 2 10159 10161
0 10163 5 1 1 10162
0 10164 7 1 2 92937 10163
0 10165 5 1 1 10164
0 10166 7 1 2 10151 10165
0 10167 5 1 1 10166
0 10168 7 1 2 89906 10167
0 10169 5 1 1 10168
0 10170 7 1 2 83181 83171
0 10171 5 1 1 10170
0 10172 7 3 2 67962 78798
0 10173 5 1 1 92950
0 10174 7 1 2 74845 92951
0 10175 5 1 1 10174
0 10176 7 1 2 10171 10175
0 10177 5 1 1 10176
0 10178 7 1 2 87896 10177
0 10179 5 1 1 10178
0 10180 7 1 2 78812 84094
0 10181 5 1 1 10180
0 10182 7 1 2 10179 10181
0 10183 5 1 1 10182
0 10184 7 1 2 69760 10183
0 10185 5 1 1 10184
0 10186 7 5 2 83899 92346
0 10187 7 2 2 76197 82869
0 10188 7 1 2 92953 92958
0 10189 5 1 1 10188
0 10190 7 1 2 10185 10189
0 10191 5 1 1 10190
0 10192 7 1 2 85117 10191
0 10193 5 1 1 10192
0 10194 7 1 2 71315 91990
0 10195 5 3 1 10194
0 10196 7 1 2 66197 91757
0 10197 5 1 1 10196
0 10198 7 1 2 92960 10197
0 10199 5 1 1 10198
0 10200 7 1 2 72980 10199
0 10201 5 1 1 10200
0 10202 7 1 2 81254 83234
0 10203 7 1 2 10201 10202
0 10204 5 1 1 10203
0 10205 7 1 2 67575 10204
0 10206 5 1 1 10205
0 10207 7 1 2 2074 91987
0 10208 5 1 1 10207
0 10209 7 1 2 72586 90941
0 10210 7 1 2 10208 10209
0 10211 5 1 1 10210
0 10212 7 1 2 10206 10211
0 10213 5 1 1 10212
0 10214 7 1 2 90995 10213
0 10215 5 1 1 10214
0 10216 7 1 2 10193 10215
0 10217 5 1 1 10216
0 10218 7 1 2 71012 10217
0 10219 5 1 1 10218
0 10220 7 9 2 72587 77411
0 10221 5 1 1 92963
0 10222 7 3 2 69761 80518
0 10223 5 1 1 92972
0 10224 7 3 2 74527 90996
0 10225 7 1 2 92973 92975
0 10226 5 1 1 10225
0 10227 7 5 2 68795 71591
0 10228 7 3 2 92978 75734
0 10229 7 1 2 83172 92983
0 10230 5 1 1 10229
0 10231 7 1 2 91026 10230
0 10232 5 1 1 10231
0 10233 7 1 2 70124 10232
0 10234 5 1 1 10233
0 10235 7 5 2 64631 78630
0 10236 5 2 1 92986
0 10237 7 1 2 80391 92987
0 10238 5 1 1 10237
0 10239 7 1 2 78203 10238
0 10240 5 1 1 10239
0 10241 7 1 2 10234 10240
0 10242 5 1 1 10241
0 10243 7 1 2 77140 10242
0 10244 5 1 1 10243
0 10245 7 1 2 10226 10244
0 10246 5 1 1 10245
0 10247 7 1 2 92964 10246
0 10248 5 1 1 10247
0 10249 7 4 2 69762 67576
0 10250 5 1 1 92993
0 10251 7 2 2 78204 92994
0 10252 7 1 2 87666 80519
0 10253 5 1 1 10252
0 10254 7 1 2 78389 10253
0 10255 5 1 1 10254
0 10256 7 1 2 92997 10255
0 10257 5 1 1 10256
0 10258 7 1 2 10248 10257
0 10259 5 1 1 10258
0 10260 7 1 2 75963 10259
0 10261 5 1 1 10260
0 10262 7 1 2 90809 80452
0 10263 5 1 1 10262
0 10264 7 1 2 91731 10263
0 10265 5 1 1 10264
0 10266 7 1 2 69435 10265
0 10267 5 1 1 10266
0 10268 7 1 2 10267 92784
0 10269 5 1 1 10268
0 10270 7 1 2 67963 10269
0 10271 5 1 1 10270
0 10272 7 1 2 86717 92196
0 10273 5 28 1 10272
0 10274 7 2 2 69436 92999
0 10275 5 2 1 93027
0 10276 7 1 2 85066 93029
0 10277 5 1 1 10276
0 10278 7 3 2 70125 80520
0 10279 7 1 2 71592 93031
0 10280 7 1 2 10277 10279
0 10281 5 1 1 10280
0 10282 7 1 2 10271 10281
0 10283 5 1 1 10282
0 10284 7 1 2 78205 10283
0 10285 5 1 1 10284
0 10286 7 1 2 10261 10285
0 10287 7 1 2 10219 10286
0 10288 5 1 1 10287
0 10289 7 1 2 88142 10288
0 10290 5 1 1 10289
0 10291 7 1 2 10169 10290
0 10292 5 1 1 10291
0 10293 7 1 2 74375 10292
0 10294 5 1 1 10293
0 10295 7 2 2 74350 84368
0 10296 7 1 2 72981 93034
0 10297 7 1 2 74179 10296
0 10298 5 1 1 10297
0 10299 7 12 2 68796 64039
0 10300 7 2 2 93036 75735
0 10301 7 1 2 90987 93048
0 10302 7 1 2 84520 10301
0 10303 5 1 1 10302
0 10304 7 1 2 10298 10303
0 10305 5 1 1 10304
0 10306 7 1 2 64306 10305
0 10307 5 1 1 10306
0 10308 7 15 2 69437 65735
0 10309 7 2 2 93037 93050
0 10310 7 1 2 90401 93065
0 10311 7 1 2 85072 10310
0 10312 5 1 1 10311
0 10313 7 1 2 10307 10312
0 10314 5 1 1 10313
0 10315 7 1 2 73950 10314
0 10316 5 1 1 10315
0 10317 7 5 2 66198 66852
0 10318 7 1 2 75601 78631
0 10319 7 1 2 93067 10318
0 10320 7 3 2 65941 77984
0 10321 5 1 1 93072
0 10322 7 1 2 93073 93035
0 10323 7 1 2 10319 10322
0 10324 5 1 1 10323
0 10325 7 1 2 10316 10324
0 10326 5 1 1 10325
0 10327 7 1 2 88143 10326
0 10328 5 1 1 10327
0 10329 7 1 2 10294 10328
0 10330 5 1 1 10329
0 10331 7 1 2 65327 10330
0 10332 5 1 1 10331
0 10333 7 4 2 67577 76931
0 10334 7 5 2 64040 92378
0 10335 7 1 2 93075 93079
0 10336 5 1 1 10335
0 10337 7 12 2 66199 72588
0 10338 7 2 2 78287 93084
0 10339 5 1 1 93096
0 10340 7 1 2 74328 93097
0 10341 5 1 1 10340
0 10342 7 1 2 10336 10341
0 10343 5 2 1 10342
0 10344 7 1 2 92612 93098
0 10345 5 1 1 10344
0 10346 7 10 2 63879 69100
0 10347 7 6 2 70766 93100
0 10348 7 1 2 93110 88884
0 10349 7 1 2 92792 10348
0 10350 5 1 1 10349
0 10351 7 1 2 10345 10350
0 10352 5 1 1 10351
0 10353 7 1 2 87225 10352
0 10354 5 1 1 10353
0 10355 7 7 2 66478 72589
0 10356 7 2 2 66200 93116
0 10357 7 5 2 69101 78308
0 10358 7 1 2 70767 93125
0 10359 7 2 2 93123 10358
0 10360 5 1 1 93130
0 10361 7 2 2 77317 93131
0 10362 5 1 1 93132
0 10363 7 1 2 92621 93133
0 10364 5 1 1 10363
0 10365 7 1 2 10354 10364
0 10366 5 1 1 10365
0 10367 7 1 2 72982 10366
0 10368 5 1 1 10367
0 10369 7 2 2 72590 84223
0 10370 7 9 2 65328 65736
0 10371 7 1 2 93136 92852
0 10372 7 1 2 93134 10371
0 10373 5 1 1 10372
0 10374 7 1 2 10368 10373
0 10375 5 1 1 10374
0 10376 7 1 2 78206 10375
0 10377 5 1 1 10376
0 10378 7 4 2 68797 75503
0 10379 7 1 2 89628 93145
0 10380 7 2 2 80313 87917
0 10381 7 1 2 78001 93149
0 10382 7 1 2 10379 10381
0 10383 7 1 2 92588 10382
0 10384 5 1 1 10383
0 10385 7 1 2 10377 10384
0 10386 5 1 1 10385
0 10387 7 1 2 80392 10386
0 10388 5 1 1 10387
0 10389 7 1 2 87814 85048
0 10390 5 9 1 10389
0 10391 7 1 2 93151 88144
0 10392 5 1 1 10391
0 10393 7 5 2 71784 84996
0 10394 7 3 2 71316 88527
0 10395 7 1 2 93160 93165
0 10396 5 1 1 10395
0 10397 7 1 2 10392 10396
0 10398 5 1 1 10397
0 10399 7 1 2 68321 10398
0 10400 5 1 1 10399
0 10401 7 2 2 77801 84997
0 10402 7 1 2 93168 89717
0 10403 5 1 1 10402
0 10404 7 1 2 10400 10403
0 10405 5 1 1 10404
0 10406 7 1 2 71593 10405
0 10407 5 1 1 10406
0 10408 7 2 2 81411 89392
0 10409 7 1 2 84157 87596
0 10410 7 1 2 93170 10409
0 10411 5 1 1 10410
0 10412 7 1 2 10407 10411
0 10413 5 1 1 10412
0 10414 7 1 2 69763 10413
0 10415 5 1 1 10414
0 10416 7 5 2 67072 67578
0 10417 7 1 2 93172 90634
0 10418 7 1 2 76116 10417
0 10419 5 1 1 10418
0 10420 7 1 2 10415 10419
0 10421 5 1 1 10420
0 10422 7 1 2 81019 10421
0 10423 5 1 1 10422
0 10424 7 3 2 82564 81462
0 10425 5 1 1 93177
0 10426 7 1 2 88145 93178
0 10427 5 1 1 10426
0 10428 7 1 2 82667 81523
0 10429 7 1 2 90060 10428
0 10430 5 1 1 10429
0 10431 7 1 2 10427 10430
0 10432 5 1 1 10431
0 10433 7 1 2 69764 10432
0 10434 5 1 1 10433
0 10435 7 4 2 72591 76068
0 10436 5 1 1 93180
0 10437 7 3 2 77141 88146
0 10438 7 1 2 93181 93184
0 10439 5 1 1 10438
0 10440 7 1 2 10434 10439
0 10441 5 1 1 10440
0 10442 7 1 2 75354 10441
0 10443 5 1 1 10442
0 10444 7 6 2 67073 91148
0 10445 7 4 2 79466 83320
0 10446 7 1 2 84283 93193
0 10447 7 1 2 93187 10446
0 10448 5 1 1 10447
0 10449 7 1 2 10443 10448
0 10450 5 1 1 10449
0 10451 7 1 2 68322 10450
0 10452 5 1 1 10451
0 10453 7 2 2 72983 77791
0 10454 7 1 2 93197 84693
0 10455 5 1 1 10454
0 10456 7 3 2 65942 84284
0 10457 5 2 1 93199
0 10458 7 1 2 86185 93200
0 10459 7 1 2 90489 10458
0 10460 5 1 1 10459
0 10461 7 1 2 10455 10460
0 10462 5 1 1 10461
0 10463 7 1 2 76460 10462
0 10464 5 1 1 10463
0 10465 7 1 2 10452 10464
0 10466 7 1 2 10423 10465
0 10467 5 1 1 10466
0 10468 7 1 2 68605 10467
0 10469 5 1 1 10468
0 10470 7 2 2 71013 84158
0 10471 7 1 2 72984 79086
0 10472 7 1 2 93204 10471
0 10473 7 1 2 84694 10472
0 10474 5 1 1 10473
0 10475 7 1 2 10469 10474
0 10476 5 1 1 10475
0 10477 7 1 2 85183 10476
0 10478 5 1 1 10477
0 10479 7 1 2 10388 10478
0 10480 7 1 2 10332 10479
0 10481 7 1 2 10106 10480
0 10482 7 1 2 9827 10481
0 10483 5 1 1 10482
0 10484 7 1 2 89571 10483
0 10485 5 1 1 10484
0 10486 7 2 2 64307 74145
0 10487 7 1 2 74846 93206
0 10488 5 1 1 10487
0 10489 7 16 2 65737 71317
0 10490 7 1 2 93208 75261
0 10491 5 1 1 10490
0 10492 7 1 2 10488 10491
0 10493 5 1 1 10492
0 10494 7 1 2 69765 10493
0 10495 5 1 1 10494
0 10496 7 1 2 75262 92391
0 10497 5 1 1 10496
0 10498 7 1 2 76562 92538
0 10499 5 1 1 10498
0 10500 7 1 2 10497 10499
0 10501 7 1 2 10495 10500
0 10502 5 1 1 10501
0 10503 7 1 2 67964 10502
0 10504 5 1 1 10503
0 10505 7 3 2 69438 76296
0 10506 5 4 1 93224
0 10507 7 2 2 93227 77586
0 10508 5 1 1 93231
0 10509 7 3 2 77206 93232
0 10510 5 1 1 93233
0 10511 7 9 2 65738 72985
0 10512 7 1 2 10510 93236
0 10513 5 1 1 10512
0 10514 7 1 2 10504 10513
0 10515 5 1 1 10514
0 10516 7 1 2 64041 10515
0 10517 5 1 1 10516
0 10518 7 22 2 65739 65943
0 10519 5 1 1 93245
0 10520 7 3 2 71594 83900
0 10521 5 1 1 93267
0 10522 7 1 2 91125 93268
0 10523 5 1 1 10522
0 10524 7 1 2 64632 86362
0 10525 7 1 2 81233 10524
0 10526 5 1 1 10525
0 10527 7 1 2 10523 10526
0 10528 5 1 1 10527
0 10529 7 1 2 68323 10528
0 10530 5 1 1 10529
0 10531 7 1 2 80013 78928
0 10532 5 1 1 10531
0 10533 7 1 2 10530 10532
0 10534 5 1 1 10533
0 10535 7 1 2 66201 10534
0 10536 5 1 1 10535
0 10537 7 1 2 81356 91126
0 10538 7 1 2 83930 10537
0 10539 5 1 1 10538
0 10540 7 1 2 10536 10539
0 10541 5 1 1 10540
0 10542 7 1 2 93246 10541
0 10543 5 1 1 10542
0 10544 7 1 2 10517 10543
0 10545 5 1 1 10544
0 10546 7 1 2 67579 10545
0 10547 5 1 1 10546
0 10548 7 2 2 82484 80828
0 10549 7 1 2 71318 93270
0 10550 5 1 1 10549
0 10551 7 1 2 77854 10550
0 10552 5 1 1 10551
0 10553 7 2 2 76676 82238
0 10554 7 1 2 93272 83631
0 10555 7 1 2 10552 10554
0 10556 5 1 1 10555
0 10557 7 1 2 10547 10556
0 10558 5 1 1 10557
0 10559 7 1 2 88147 10558
0 10560 5 1 1 10559
0 10561 7 1 2 73389 79590
0 10562 5 1 1 10561
0 10563 7 1 2 89805 10562
0 10564 5 1 1 10563
0 10565 7 1 2 67965 10564
0 10566 5 1 1 10565
0 10567 7 2 2 87009 75689
0 10568 5 2 1 93274
0 10569 7 1 2 73390 79548
0 10570 5 1 1 10569
0 10571 7 1 2 93276 10570
0 10572 7 1 2 10566 10571
0 10573 5 1 1 10572
0 10574 7 1 2 77412 10573
0 10575 5 1 1 10574
0 10576 7 3 2 73391 77142
0 10577 5 1 1 93278
0 10578 7 1 2 75004 93279
0 10579 5 1 1 10578
0 10580 7 1 2 10575 10579
0 10581 5 1 1 10580
0 10582 7 1 2 78535 10581
0 10583 5 1 1 10582
0 10584 7 3 2 78632 75904
0 10585 5 1 1 93281
0 10586 7 3 2 66202 87034
0 10587 5 3 1 93284
0 10588 7 2 2 93287 77706
0 10589 5 2 1 93290
0 10590 7 1 2 64633 93292
0 10591 5 1 1 10590
0 10592 7 1 2 10585 10591
0 10593 5 4 1 10592
0 10594 7 1 2 92833 93294
0 10595 5 1 1 10594
0 10596 7 1 2 10583 10595
0 10597 5 1 1 10596
0 10598 7 1 2 88528 10597
0 10599 5 1 1 10598
0 10600 7 1 2 10560 10599
0 10601 5 1 1 10600
0 10602 7 1 2 88956 10601
0 10603 5 1 1 10602
0 10604 7 2 2 71319 77879
0 10605 5 1 1 93298
0 10606 7 1 2 75855 10605
0 10607 5 3 1 10606
0 10608 7 1 2 64308 93300
0 10609 5 1 1 10608
0 10610 7 1 2 77802 77697
0 10611 5 1 1 10610
0 10612 7 1 2 10609 10611
0 10613 5 1 1 10612
0 10614 7 1 2 88148 10613
0 10615 5 1 1 10614
0 10616 7 1 2 89825 83231
0 10617 5 1 1 10616
0 10618 7 1 2 10615 10617
0 10619 5 1 1 10618
0 10620 7 1 2 69766 10619
0 10621 5 1 1 10620
0 10622 7 1 2 77709 89481
0 10623 5 1 1 10622
0 10624 7 1 2 64309 10623
0 10625 5 1 1 10624
0 10626 7 1 2 78633 81569
0 10627 7 1 2 90181 10626
0 10628 5 1 1 10627
0 10629 7 1 2 75905 89882
0 10630 5 1 1 10629
0 10631 7 1 2 90861 10630
0 10632 7 1 2 10628 10631
0 10633 5 1 1 10632
0 10634 7 1 2 10625 10633
0 10635 5 1 1 10634
0 10636 7 1 2 10621 10635
0 10637 5 1 1 10636
0 10638 7 1 2 88149 80185
0 10639 5 1 1 10638
0 10640 7 1 2 77532 89826
0 10641 5 1 1 10640
0 10642 7 1 2 10639 10641
0 10643 5 1 1 10642
0 10644 7 1 2 69439 10643
0 10645 5 1 1 10644
0 10646 7 1 2 72592 10645
0 10647 5 1 1 10646
0 10648 7 1 2 71014 10647
0 10649 7 1 2 10637 10648
0 10650 5 1 1 10649
0 10651 7 2 2 76642 88150
0 10652 5 1 1 93303
0 10653 7 1 2 92042 10652
0 10654 5 1 1 10653
0 10655 7 1 2 71320 10654
0 10656 5 1 1 10655
0 10657 7 1 2 72593 90977
0 10658 7 1 2 10656 10657
0 10659 5 1 1 10658
0 10660 7 1 2 79960 92794
0 10661 5 1 1 10660
0 10662 7 1 2 66203 89341
0 10663 5 1 1 10662
0 10664 7 1 2 67580 10663
0 10665 7 1 2 10661 10664
0 10666 5 1 1 10665
0 10667 7 1 2 69440 10666
0 10668 7 1 2 10659 10667
0 10669 5 1 1 10668
0 10670 7 1 2 81004 10669
0 10671 5 1 1 10670
0 10672 7 1 2 92043 9812
0 10673 5 1 1 10672
0 10674 7 1 2 85075 10673
0 10675 5 1 1 10674
0 10676 7 1 2 77207 10675
0 10677 5 1 1 10676
0 10678 7 1 2 68324 10677
0 10679 7 1 2 10671 10678
0 10680 5 1 1 10679
0 10681 7 1 2 82379 80175
0 10682 5 1 1 10681
0 10683 7 1 2 79975 10682
0 10684 5 1 1 10683
0 10685 7 1 2 67581 89876
0 10686 7 1 2 10684 10685
0 10687 5 1 1 10686
0 10688 7 1 2 10680 10687
0 10689 7 1 2 10650 10688
0 10690 5 1 1 10689
0 10691 7 8 2 64042 70617
0 10692 7 4 2 93305 90523
0 10693 7 5 2 71914 73691
0 10694 7 8 2 70716 65740
0 10695 5 1 1 93322
0 10696 7 1 2 93317 93323
0 10697 7 1 2 93313 10696
0 10698 7 1 2 10690 10697
0 10699 5 1 1 10698
0 10700 7 1 2 10603 10699
0 10701 5 1 1 10700
0 10702 7 1 2 85220 10701
0 10703 5 1 1 10702
0 10704 7 1 2 72986 74874
0 10705 5 3 1 10704
0 10706 7 1 2 69441 93330
0 10707 7 1 2 89945 10706
0 10708 5 1 1 10707
0 10709 7 1 2 80005 80055
0 10710 7 1 2 10708 10709
0 10711 5 1 1 10710
0 10712 7 1 2 80057 10711
0 10713 5 1 1 10712
0 10714 7 1 2 80147 10713
0 10715 5 1 1 10714
0 10716 7 1 2 88529 10715
0 10717 5 1 1 10716
0 10718 7 1 2 88530 92750
0 10719 5 1 1 10718
0 10720 7 1 2 73692 81181
0 10721 7 2 2 81316 10720
0 10722 7 2 2 67074 90265
0 10723 7 1 2 93333 93335
0 10724 5 1 1 10723
0 10725 7 1 2 10719 10724
0 10726 5 1 1 10725
0 10727 7 1 2 72987 10726
0 10728 5 1 1 10727
0 10729 7 1 2 76563 78894
0 10730 5 1 1 10729
0 10731 7 1 2 89801 10730
0 10732 5 1 1 10731
0 10733 7 1 2 76152 88151
0 10734 7 1 2 10732 10733
0 10735 5 1 1 10734
0 10736 7 1 2 10728 10735
0 10737 5 1 1 10736
0 10738 7 1 2 71015 10737
0 10739 5 1 1 10738
0 10740 7 1 2 10717 10739
0 10741 5 1 1 10740
0 10742 7 1 2 67582 10741
0 10743 5 1 1 10742
0 10744 7 1 2 84998 92698
0 10745 7 1 2 77494 10744
0 10746 5 1 1 10745
0 10747 7 1 2 10743 10746
0 10748 5 1 1 10747
0 10749 7 1 2 74376 10748
0 10750 5 1 1 10749
0 10751 7 3 2 87035 83827
0 10752 7 1 2 65009 93337
0 10753 5 1 1 10752
0 10754 7 1 2 73951 76993
0 10755 5 1 1 10754
0 10756 7 1 2 10753 10755
0 10757 5 1 1 10756
0 10758 7 1 2 76198 10757
0 10759 5 1 1 10758
0 10760 7 6 2 76564 75263
0 10761 7 1 2 90186 93340
0 10762 5 1 1 10761
0 10763 7 1 2 10759 10762
0 10764 5 1 1 10763
0 10765 7 9 2 69102 72594
0 10766 5 1 1 93346
0 10767 7 5 2 77058 93347
0 10768 5 1 1 93355
0 10769 7 1 2 93188 93356
0 10770 7 1 2 10764 10769
0 10771 5 1 1 10770
0 10772 7 1 2 10750 10771
0 10773 5 1 1 10772
0 10774 7 1 2 88957 10773
0 10775 5 1 1 10774
0 10776 7 4 2 88018 93324
0 10777 7 2 2 71915 93360
0 10778 7 3 2 92448 93364
0 10779 7 1 2 72988 88311
0 10780 7 1 2 644 10779
0 10781 5 1 1 10780
0 10782 7 1 2 7484 10781
0 10783 5 1 1 10782
0 10784 7 1 2 88152 10783
0 10785 5 1 1 10784
0 10786 7 1 2 74488 89476
0 10787 5 1 1 10786
0 10788 7 1 2 10785 10787
0 10789 5 1 1 10788
0 10790 7 1 2 70126 10789
0 10791 5 1 1 10790
0 10792 7 1 2 79718 92080
0 10793 5 1 1 10792
0 10794 7 1 2 10791 10793
0 10795 5 1 1 10794
0 10796 7 1 2 84664 10795
0 10797 5 1 1 10796
0 10798 7 1 2 76297 79502
0 10799 7 1 2 89877 88644
0 10800 7 1 2 10798 10799
0 10801 5 1 1 10800
0 10802 7 1 2 10797 10801
0 10803 5 1 1 10802
0 10804 7 1 2 68325 10803
0 10805 5 1 1 10804
0 10806 7 1 2 74821 81463
0 10807 5 1 1 10806
0 10808 7 1 2 67583 88749
0 10809 5 1 1 10808
0 10810 7 1 2 10807 10809
0 10811 5 1 1 10810
0 10812 7 1 2 67966 10811
0 10813 5 1 1 10812
0 10814 7 1 2 81524 88450
0 10815 5 1 1 10814
0 10816 7 1 2 10813 10815
0 10817 5 1 1 10816
0 10818 7 1 2 92081 10817
0 10819 5 1 1 10818
0 10820 7 1 2 10805 10819
0 10821 5 1 1 10820
0 10822 7 1 2 71016 10821
0 10823 5 1 1 10822
0 10824 7 3 2 67584 84173
0 10825 7 1 2 89861 83955
0 10826 7 1 2 93369 10825
0 10827 7 1 2 83640 10826
0 10828 5 1 1 10827
0 10829 7 1 2 10823 10828
0 10830 5 1 1 10829
0 10831 7 1 2 93366 10830
0 10832 5 1 1 10831
0 10833 7 1 2 10775 10832
0 10834 5 1 1 10833
0 10835 7 1 2 85872 10834
0 10836 5 1 1 10835
0 10837 7 1 2 10703 10836
0 10838 5 1 1 10837
0 10839 7 1 2 65329 10838
0 10840 5 1 1 10839
0 10841 7 1 2 74377 87403
0 10842 7 1 2 84225 10841
0 10843 5 1 1 10842
0 10844 7 2 2 82768 77745
0 10845 5 1 1 93372
0 10846 7 6 2 69103 72989
0 10847 5 1 1 93374
0 10848 7 2 2 93375 89331
0 10849 5 1 1 93380
0 10850 7 1 2 10845 10849
0 10851 5 1 1 10850
0 10852 7 1 2 77850 10851
0 10853 5 1 1 10852
0 10854 7 1 2 82757 84048
0 10855 7 1 2 93271 10854
0 10856 5 1 1 10855
0 10857 7 1 2 10853 10856
0 10858 5 1 1 10857
0 10859 7 1 2 64310 87697
0 10860 7 1 2 10858 10859
0 10861 5 1 1 10860
0 10862 7 1 2 10843 10861
0 10863 5 1 1 10862
0 10864 7 1 2 73693 10863
0 10865 5 1 1 10864
0 10866 7 3 2 72019 75355
0 10867 7 1 2 93382 93066
0 10868 5 1 1 10867
0 10869 7 1 2 64311 83143
0 10870 5 1 1 10869
0 10871 7 3 2 85873 74378
0 10872 7 1 2 10870 93385
0 10873 5 1 1 10872
0 10874 7 1 2 67967 93386
0 10875 5 1 1 10874
0 10876 7 3 2 64312 82485
0 10877 7 7 2 66953 84568
0 10878 5 1 1 93391
0 10879 7 1 2 74774 93392
0 10880 7 1 2 93388 10879
0 10881 5 1 1 10880
0 10882 7 1 2 10875 10881
0 10883 5 1 1 10882
0 10884 7 1 2 71595 10883
0 10885 5 1 1 10884
0 10886 7 1 2 10873 10885
0 10887 5 1 1 10886
0 10888 7 1 2 76461 10887
0 10889 5 1 1 10888
0 10890 7 1 2 10868 10889
0 10891 5 1 1 10890
0 10892 7 1 2 77575 10891
0 10893 5 1 1 10892
0 10894 7 5 2 66954 79446
0 10895 7 2 2 66204 93398
0 10896 7 2 2 77318 74164
0 10897 7 1 2 81357 93405
0 10898 7 1 2 93403 10897
0 10899 5 1 1 10898
0 10900 7 2 2 72020 82024
0 10901 7 5 2 69767 93209
0 10902 5 1 1 93409
0 10903 7 1 2 69442 93038
0 10904 7 1 2 93410 10903
0 10905 7 1 2 93407 10904
0 10906 5 1 1 10905
0 10907 7 1 2 10899 10906
0 10908 7 1 2 10893 10907
0 10909 5 1 1 10908
0 10910 7 1 2 88153 10909
0 10911 5 1 1 10910
0 10912 7 1 2 72595 10911
0 10913 7 1 2 10865 10912
0 10914 5 1 1 10913
0 10915 7 6 2 68798 74208
0 10916 5 1 1 93414
0 10917 7 1 2 93415 92329
0 10918 5 1 1 10917
0 10919 7 1 2 10902 92394
0 10920 5 2 1 10919
0 10921 7 1 2 85221 76153
0 10922 7 1 2 93420 10921
0 10923 5 1 1 10922
0 10924 7 1 2 10918 10923
0 10925 5 1 1 10924
0 10926 7 1 2 88154 10925
0 10927 5 1 1 10926
0 10928 7 1 2 76045 74219
0 10929 7 1 2 89380 10928
0 10930 7 1 2 84275 10929
0 10931 5 1 1 10930
0 10932 7 1 2 10927 10931
0 10933 5 1 1 10932
0 10934 7 1 2 64043 10933
0 10935 5 1 1 10934
0 10936 7 6 2 65741 74146
0 10937 7 2 2 80014 93422
0 10938 5 1 1 93428
0 10939 7 1 2 76154 89406
0 10940 7 1 2 93429 10939
0 10941 5 1 1 10940
0 10942 7 1 2 10935 10941
0 10943 5 1 1 10942
0 10944 7 1 2 87226 10943
0 10945 5 1 1 10944
0 10946 7 2 2 65742 88155
0 10947 7 4 2 66205 81999
0 10948 7 4 2 66955 90889
0 10949 7 4 2 65944 73694
0 10950 7 1 2 74489 93440
0 10951 7 1 2 93436 10950
0 10952 7 1 2 93432 10951
0 10953 5 1 1 10952
0 10954 7 7 2 65010 92363
0 10955 5 1 1 93444
0 10956 7 1 2 76565 93445
0 10957 5 1 1 10956
0 10958 7 1 2 81327 10957
0 10959 5 1 1 10958
0 10960 7 1 2 67968 10959
0 10961 5 1 1 10960
0 10962 7 1 2 77583 92660
0 10963 5 1 1 10962
0 10964 7 1 2 82065 10963
0 10965 7 1 2 10961 10964
0 10966 5 1 1 10965
0 10967 7 10 2 72021 93039
0 10968 7 1 2 93451 82067
0 10969 7 1 2 10966 10968
0 10970 5 1 1 10969
0 10971 7 1 2 10953 10970
0 10972 5 1 1 10971
0 10973 7 1 2 93430 10972
0 10974 5 1 1 10973
0 10975 7 1 2 67585 10974
0 10976 7 1 2 10945 10975
0 10977 5 1 1 10976
0 10978 7 1 2 88958 10977
0 10979 7 1 2 10914 10978
0 10980 5 1 1 10979
0 10981 7 1 2 69443 92680
0 10982 5 1 1 10981
0 10983 7 1 2 72990 79825
0 10984 5 2 1 10983
0 10985 7 1 2 91993 93461
0 10986 5 1 1 10985
0 10987 7 1 2 71321 10986
0 10988 5 1 1 10987
0 10989 7 1 2 92935 10988
0 10990 5 1 1 10989
0 10991 7 1 2 81525 10990
0 10992 5 1 1 10991
0 10993 7 1 2 10982 10992
0 10994 5 1 1 10993
0 10995 7 1 2 89304 10994
0 10996 5 1 1 10995
0 10997 7 2 2 71322 85874
0 10998 7 1 2 93463 79087
0 10999 7 1 2 87905 10998
0 11000 5 1 1 10999
0 11001 7 1 2 10996 11000
0 11002 5 1 1 11001
0 11003 7 1 2 71017 11002
0 11004 5 1 1 11003
0 11005 7 1 2 92938 89305
0 11006 7 1 2 92949 11005
0 11007 5 1 1 11006
0 11008 7 1 2 11004 11007
0 11009 5 1 1 11008
0 11010 7 1 2 93367 11009
0 11011 5 1 1 11010
0 11012 7 1 2 85875 79993
0 11013 7 4 2 67586 75964
0 11014 5 2 1 93465
0 11015 7 1 2 93466 84499
0 11016 7 1 2 11012 11015
0 11017 5 1 1 11016
0 11018 7 1 2 73952 93376
0 11019 7 1 2 90848 11018
0 11020 7 1 2 77851 11019
0 11021 5 1 1 11020
0 11022 7 1 2 11017 11021
0 11023 5 1 1 11022
0 11024 7 1 2 88959 11023
0 11025 5 1 1 11024
0 11026 7 1 2 84349 78360
0 11027 7 1 2 90187 11026
0 11028 7 7 2 70717 70768
0 11029 7 4 2 70660 93471
0 11030 7 2 2 86498 91893
0 11031 7 1 2 93482 93150
0 11032 7 1 2 93478 11031
0 11033 7 1 2 11027 11032
0 11034 5 1 1 11033
0 11035 7 1 2 11025 11034
0 11036 5 1 1 11035
0 11037 7 1 2 64313 11036
0 11038 5 1 1 11037
0 11039 7 1 2 78818 78475
0 11040 5 1 1 11039
0 11041 7 1 2 79615 83746
0 11042 5 1 1 11041
0 11043 7 1 2 11040 11042
0 11044 5 1 1 11043
0 11045 7 2 2 93051 88912
0 11046 7 1 2 93452 88903
0 11047 7 1 2 93484 11046
0 11048 7 1 2 11044 11047
0 11049 5 1 1 11048
0 11050 7 1 2 11038 11049
0 11051 5 1 1 11050
0 11052 7 1 2 92622 11051
0 11053 5 1 1 11052
0 11054 7 1 2 11011 11053
0 11055 7 1 2 10980 11054
0 11056 7 1 2 10840 11055
0 11057 5 1 1 11056
0 11058 7 1 2 66670 11057
0 11059 5 1 1 11058
0 11060 7 1 2 88289 6224
0 11061 5 1 1 11060
0 11062 7 4 2 64044 71596
0 11063 7 1 2 93486 84014
0 11064 7 1 2 92542 11063
0 11065 5 1 1 11064
0 11066 7 1 2 79574 78405
0 11067 7 1 2 91065 11066
0 11068 7 2 2 63964 79275
0 11069 7 1 2 92227 93490
0 11070 7 1 2 11067 11069
0 11071 5 1 1 11070
0 11072 7 1 2 11065 11071
0 11073 5 1 1 11072
0 11074 7 1 2 65743 11073
0 11075 5 1 1 11074
0 11076 7 2 2 64634 90580
0 11077 7 1 2 86414 88913
0 11078 7 1 2 93492 11077
0 11079 7 5 2 75906 83719
0 11080 7 2 2 64314 74419
0 11081 7 1 2 93494 93499
0 11082 7 1 2 11078 11081
0 11083 5 1 1 11082
0 11084 7 1 2 11075 11083
0 11085 5 1 1 11084
0 11086 7 1 2 63752 11085
0 11087 5 1 1 11086
0 11088 7 1 2 92417 84015
0 11089 7 1 2 92564 11088
0 11090 7 1 2 80955 11089
0 11091 5 1 1 11090
0 11092 7 1 2 11087 11091
0 11093 5 1 1 11092
0 11094 7 1 2 73392 11093
0 11095 5 1 1 11094
0 11096 7 4 2 72022 87790
0 11097 7 1 2 92565 93501
0 11098 5 1 1 11097
0 11099 7 1 2 92533 93502
0 11100 5 1 1 11099
0 11101 7 2 2 67969 82380
0 11102 7 1 2 72596 93505
0 11103 7 1 2 90750 11102
0 11104 5 1 1 11103
0 11105 7 1 2 11100 11104
0 11106 5 1 1 11105
0 11107 7 1 2 63753 11106
0 11108 5 1 1 11107
0 11109 7 1 2 11098 11108
0 11110 5 1 1 11109
0 11111 7 1 2 82054 92568
0 11112 7 1 2 11110 11111
0 11113 5 1 1 11112
0 11114 7 1 2 11095 11113
0 11115 5 1 1 11114
0 11116 7 1 2 70127 11115
0 11117 5 1 1 11116
0 11118 7 3 2 64635 80075
0 11119 7 2 2 64045 93052
0 11120 7 1 2 93507 93510
0 11121 7 1 2 93503 11120
0 11122 7 1 2 92516 11121
0 11123 5 1 1 11122
0 11124 7 1 2 11117 11123
0 11125 5 1 1 11124
0 11126 7 1 2 87100 11125
0 11127 5 1 1 11126
0 11128 7 3 2 69444 83720
0 11129 5 1 1 93512
0 11130 7 5 2 64315 78433
0 11131 5 3 1 93515
0 11132 7 1 2 93520 92291
0 11133 7 1 2 11129 11132
0 11134 5 11 1 11133
0 11135 7 4 2 68326 91875
0 11136 7 1 2 74134 75143
0 11137 7 1 2 92379 11136
0 11138 7 1 2 93534 11137
0 11139 7 1 2 93523 11138
0 11140 7 1 2 90394 11139
0 11141 5 1 1 11140
0 11142 7 1 2 11127 11141
0 11143 5 1 1 11142
0 11144 7 1 2 11061 11143
0 11145 5 1 1 11144
0 11146 7 1 2 83428 84723
0 11147 5 1 1 11146
0 11148 7 1 2 84927 11147
0 11149 5 1 1 11148
0 11150 7 2 2 86319 79892
0 11151 7 3 2 70769 83721
0 11152 5 1 1 93540
0 11153 7 1 2 73695 93541
0 11154 7 1 2 93538 11153
0 11155 5 1 1 11154
0 11156 7 1 2 11149 11155
0 11157 5 1 1 11156
0 11158 7 1 2 65011 11157
0 11159 5 1 1 11158
0 11160 7 1 2 64046 92264
0 11161 7 1 2 92392 11160
0 11162 5 1 1 11161
0 11163 7 1 2 11159 11162
0 11164 5 1 1 11163
0 11165 7 2 2 82758 90785
0 11166 7 1 2 72991 92507
0 11167 7 1 2 79325 11166
0 11168 7 1 2 93543 11167
0 11169 7 1 2 11164 11168
0 11170 5 1 1 11169
0 11171 7 1 2 11145 11170
0 11172 5 1 1 11171
0 11173 7 1 2 70375 11172
0 11174 5 1 1 11173
0 11175 7 1 2 92811 92292
0 11176 5 1 1 11175
0 11177 7 1 2 87227 11176
0 11178 5 1 1 11177
0 11179 7 1 2 5336 11178
0 11180 5 1 1 11179
0 11181 7 1 2 90208 11180
0 11182 5 1 1 11181
0 11183 7 3 2 86499 91163
0 11184 7 2 2 92456 93545
0 11185 7 2 2 92303 81394
0 11186 7 1 2 78374 93550
0 11187 7 1 2 93548 11186
0 11188 5 1 1 11187
0 11189 7 1 2 11182 11188
0 11190 5 1 1 11189
0 11191 7 1 2 77533 11190
0 11192 5 1 1 11191
0 11193 7 2 2 93453 88063
0 11194 7 1 2 90830 93552
0 11195 5 1 1 11194
0 11196 7 1 2 9355 11195
0 11197 5 1 1 11196
0 11198 7 1 2 69445 84476
0 11199 7 1 2 11197 11198
0 11200 5 1 1 11199
0 11201 7 1 2 11192 11200
0 11202 5 1 1 11201
0 11203 7 1 2 65744 11202
0 11204 5 1 1 11203
0 11205 7 2 2 67970 88960
0 11206 7 1 2 87228 84949
0 11207 5 1 1 11206
0 11208 7 7 2 64047 71018
0 11209 7 2 2 76462 93556
0 11210 5 1 1 93563
0 11211 7 1 2 77855 11210
0 11212 5 2 1 11211
0 11213 7 1 2 88733 93565
0 11214 5 1 1 11213
0 11215 7 1 2 11207 11214
0 11216 5 1 1 11215
0 11217 7 1 2 93554 11216
0 11218 5 1 1 11217
0 11219 7 1 2 77655 84454
0 11220 7 5 2 71916 72597
0 11221 7 6 2 69057 69104
0 11222 5 1 1 93572
0 11223 7 1 2 93567 93573
0 11224 7 1 2 11219 11223
0 11225 7 1 2 77077 93546
0 11226 7 1 2 11224 11225
0 11227 5 1 1 11226
0 11228 7 1 2 11218 11227
0 11229 5 1 1 11228
0 11230 7 1 2 85222 11229
0 11231 5 1 1 11230
0 11232 7 1 2 11204 11231
0 11233 5 1 1 11232
0 11234 7 1 2 88156 11233
0 11235 5 1 1 11234
0 11236 7 1 2 87229 93099
0 11237 5 1 1 11236
0 11238 7 1 2 10362 11237
0 11239 5 1 1 11238
0 11240 7 1 2 72992 11239
0 11241 5 1 1 11240
0 11242 7 1 2 74379 93135
0 11243 5 1 1 11242
0 11244 7 1 2 11241 11243
0 11245 5 1 1 11244
0 11246 7 1 2 90437 11245
0 11247 5 1 1 11246
0 11248 7 1 2 11235 11247
0 11249 5 1 1 11248
0 11250 7 1 2 65330 11249
0 11251 5 1 1 11250
0 11252 7 2 2 72598 81189
0 11253 7 11 2 63880 90581
0 11254 7 8 2 68799 70770
0 11255 7 3 2 69105 93591
0 11256 7 1 2 93580 93599
0 11257 7 1 2 79349 11256
0 11258 7 1 2 92528 11257
0 11259 7 1 2 93578 11258
0 11260 5 1 1 11259
0 11261 7 1 2 11251 11260
0 11262 5 1 1 11261
0 11263 7 1 2 80393 11262
0 11264 5 1 1 11263
0 11265 7 12 2 64048 69768
0 11266 7 9 2 71323 93602
0 11267 7 6 2 70718 71019
0 11268 7 4 2 88019 93623
0 11269 7 1 2 93614 93629
0 11270 7 1 2 92319 11269
0 11271 5 1 1 11270
0 11272 7 1 2 9357 11271
0 11273 5 1 1 11272
0 11274 7 1 2 88157 11273
0 11275 5 1 1 11274
0 11276 7 1 2 63965 65012
0 11277 7 1 2 68606 11276
0 11278 7 1 2 89306 11277
0 11279 7 1 2 91259 11278
0 11280 7 1 2 84733 11279
0 11281 5 1 1 11280
0 11282 7 1 2 11275 11281
0 11283 5 1 1 11282
0 11284 7 1 2 66671 11283
0 11285 5 1 1 11284
0 11286 7 3 2 68607 84665
0 11287 7 1 2 93603 84484
0 11288 7 1 2 91264 11287
0 11289 7 1 2 89332 93630
0 11290 7 1 2 11288 11289
0 11291 7 1 2 93633 11290
0 11292 5 1 1 11291
0 11293 7 1 2 11285 11292
0 11294 5 1 1 11293
0 11295 7 1 2 65331 11294
0 11296 5 1 1 11295
0 11297 7 5 2 65683 66206
0 11298 7 5 2 63754 71785
0 11299 7 1 2 93641 74233
0 11300 7 1 2 93636 11299
0 11301 7 7 2 63966 64049
0 11302 5 1 1 93646
0 11303 7 2 2 68962 93647
0 11304 7 10 2 67587 77413
0 11305 5 1 1 93655
0 11306 7 1 2 91346 93656
0 11307 7 1 2 93653 11306
0 11308 7 1 2 11300 11307
0 11309 5 1 1 11308
0 11310 7 1 2 11296 11309
0 11311 5 1 1 11310
0 11312 7 1 2 65745 11311
0 11313 5 1 1 11312
0 11314 7 8 2 66672 66853
0 11315 7 2 2 76132 93665
0 11316 7 2 2 63967 89539
0 11317 7 1 2 89307 93675
0 11318 7 1 2 93673 11317
0 11319 7 3 2 65013 65945
0 11320 5 1 1 93677
0 11321 7 1 2 88885 93678
0 11322 7 1 2 84957 11321
0 11323 7 1 2 11318 11322
0 11324 5 1 1 11323
0 11325 7 1 2 11313 11324
0 11326 5 1 1 11325
0 11327 7 1 2 84539 11326
0 11328 5 1 1 11327
0 11329 7 2 2 65332 73953
0 11330 5 6 1 93680
0 11331 7 1 2 93682 78686
0 11332 5 3 1 11331
0 11333 7 4 2 69106 77059
0 11334 5 1 1 93691
0 11335 7 1 2 77558 93692
0 11336 7 1 2 93688 11335
0 11337 5 1 1 11336
0 11338 7 1 2 65014 92247
0 11339 7 1 2 93566 11338
0 11340 5 1 1 11339
0 11341 7 1 2 11337 11340
0 11342 5 1 1 11341
0 11343 7 1 2 85223 11342
0 11344 5 1 1 11343
0 11345 7 23 2 68800 69107
0 11346 7 1 2 80307 93695
0 11347 7 1 2 74209 11346
0 11348 7 1 2 80924 77852
0 11349 7 1 2 11347 11348
0 11350 7 1 2 93689 11349
0 11351 5 1 1 11350
0 11352 7 1 2 11344 11351
0 11353 5 1 1 11352
0 11354 7 1 2 88158 11353
0 11355 5 1 1 11354
0 11356 7 6 2 85224 74619
0 11357 5 1 1 93718
0 11358 7 1 2 80243 93719
0 11359 5 1 1 11358
0 11360 7 1 2 92115 11359
0 11361 5 1 1 11360
0 11362 7 20 2 68963 69108
0 11363 7 2 2 93724 74329
0 11364 7 1 2 75907 91280
0 11365 7 1 2 93744 11364
0 11366 7 1 2 11361 11365
0 11367 5 1 1 11366
0 11368 7 1 2 11355 11367
0 11369 5 1 1 11368
0 11370 7 1 2 84934 11369
0 11371 5 1 1 11370
0 11372 7 8 2 73393 75264
0 11373 5 6 1 93746
0 11374 7 1 2 84251 93754
0 11375 5 2 1 11374
0 11376 7 8 2 63755 64050
0 11377 7 2 2 93762 89862
0 11378 7 1 2 93770 84435
0 11379 7 1 2 82536 91942
0 11380 7 1 2 11378 11379
0 11381 7 1 2 93760 11380
0 11382 5 1 1 11381
0 11383 7 1 2 11371 11382
0 11384 5 1 1 11383
0 11385 7 1 2 88961 11384
0 11386 5 1 1 11385
0 11387 7 1 2 11328 11386
0 11388 7 1 2 11264 11387
0 11389 7 1 2 11174 11388
0 11390 7 1 2 11059 11389
0 11391 7 1 2 10485 11390
0 11392 7 1 2 9654 11391
0 11393 7 1 2 9330 11392
0 11394 7 1 2 6933 11393
0 11395 7 1 2 3354 11394
0 11396 5 1 1 11395
0 11397 7 1 2 72297 11396
0 11398 5 1 1 11397
0 11399 7 3 2 81698 86363
0 11400 5 1 1 93772
0 11401 7 2 2 93773 80958
0 11402 5 3 1 93775
0 11403 7 2 2 81699 77308
0 11404 5 2 1 93780
0 11405 7 2 2 86462 93782
0 11406 5 3 1 93784
0 11407 7 1 2 84922 93785
0 11408 5 2 1 11407
0 11409 7 1 2 68327 93789
0 11410 5 1 1 11409
0 11411 7 2 2 93777 11410
0 11412 5 1 1 93791
0 11413 7 3 2 65015 78024
0 11414 5 5 1 93793
0 11415 7 1 2 93796 83437
0 11416 5 1 1 11415
0 11417 7 1 2 93792 11416
0 11418 5 1 1 11417
0 11419 7 1 2 88159 11418
0 11420 5 1 1 11419
0 11421 7 6 2 65016 80676
0 11422 5 10 1 93801
0 11423 7 1 2 86774 93807
0 11424 5 5 1 11423
0 11425 7 2 2 71597 93817
0 11426 5 1 1 93822
0 11427 7 5 2 65017 80578
0 11428 5 4 1 93824
0 11429 7 1 2 73696 93825
0 11430 5 1 1 11429
0 11431 7 1 2 11426 11430
0 11432 5 2 1 11431
0 11433 7 3 2 68328 93833
0 11434 5 3 1 93835
0 11435 7 1 2 73394 83496
0 11436 7 1 2 75118 83156
0 11437 7 1 2 11435 11436
0 11438 5 1 1 11437
0 11439 7 1 2 93838 11438
0 11440 5 1 1 11439
0 11441 7 1 2 88531 11440
0 11442 5 1 1 11441
0 11443 7 1 2 11420 11442
0 11444 5 1 1 11443
0 11445 7 1 2 72993 11444
0 11446 5 1 1 11445
0 11447 7 12 2 63881 66673
0 11448 7 4 2 67075 93841
0 11449 7 2 2 79228 79762
0 11450 5 2 1 93857
0 11451 7 1 2 93853 93858
0 11452 5 1 1 11451
0 11453 7 7 2 74620 87561
0 11454 5 1 1 93861
0 11455 7 2 2 73395 92623
0 11456 7 1 2 93862 93868
0 11457 5 1 1 11456
0 11458 7 2 2 65018 89290
0 11459 7 1 2 81583 7194
0 11460 7 1 2 93870 11459
0 11461 5 1 1 11460
0 11462 7 1 2 11457 11461
0 11463 5 1 1 11462
0 11464 7 1 2 67971 11463
0 11465 5 1 1 11464
0 11466 7 1 2 11452 11465
0 11467 7 1 2 11446 11466
0 11468 5 1 1 11467
0 11469 7 1 2 85876 11468
0 11470 5 1 1 11469
0 11471 7 1 2 65333 82369
0 11472 5 2 1 11471
0 11473 7 1 2 87842 93872
0 11474 5 1 1 11473
0 11475 7 1 2 88160 11474
0 11476 5 1 1 11475
0 11477 7 6 2 71786 75119
0 11478 5 1 1 93874
0 11479 7 1 2 87836 93875
0 11480 5 1 1 11479
0 11481 7 1 2 73396 78025
0 11482 5 8 1 11481
0 11483 7 2 2 74621 87632
0 11484 5 1 1 93888
0 11485 7 1 2 93880 93889
0 11486 5 1 1 11485
0 11487 7 2 2 90824 79763
0 11488 5 1 1 93890
0 11489 7 1 2 86729 11488
0 11490 7 1 2 11486 11489
0 11491 7 1 2 11480 11490
0 11492 5 1 1 11491
0 11493 7 1 2 88532 11492
0 11494 5 1 1 11493
0 11495 7 1 2 11476 11494
0 11496 5 1 1 11495
0 11497 7 1 2 85225 11496
0 11498 5 1 1 11497
0 11499 7 1 2 11470 11498
0 11500 5 1 1 11499
0 11501 7 1 2 66207 11500
0 11502 5 1 1 11501
0 11503 7 5 2 66956 79366
0 11504 7 3 2 87572 90544
0 11505 7 1 2 93892 93897
0 11506 5 1 1 11505
0 11507 7 1 2 68801 86995
0 11508 5 1 1 11507
0 11509 7 1 2 90706 88161
0 11510 7 1 2 11508 11509
0 11511 5 1 1 11510
0 11512 7 1 2 11506 11511
0 11513 5 1 1 11512
0 11514 7 1 2 66479 11513
0 11515 5 1 1 11514
0 11516 7 2 2 79818 88162
0 11517 5 2 1 93900
0 11518 7 4 2 73397 89165
0 11519 5 2 1 93904
0 11520 7 1 2 86640 93908
0 11521 5 1 1 11520
0 11522 7 1 2 88533 11521
0 11523 5 1 1 11522
0 11524 7 1 2 93902 11523
0 11525 5 2 1 11524
0 11526 7 1 2 85226 93910
0 11527 5 1 1 11526
0 11528 7 1 2 11515 11527
0 11529 5 1 1 11528
0 11530 7 1 2 65019 11529
0 11531 5 2 1 11530
0 11532 7 1 2 66480 93911
0 11533 5 1 1 11532
0 11534 7 3 2 87633 88163
0 11535 5 1 1 93914
0 11536 7 1 2 65334 93915
0 11537 5 1 1 11536
0 11538 7 1 2 11533 11537
0 11539 5 1 1 11538
0 11540 7 1 2 85227 11539
0 11541 5 1 1 11540
0 11542 7 1 2 93912 11541
0 11543 5 1 1 11542
0 11544 7 1 2 72994 11543
0 11545 5 1 1 11544
0 11546 7 2 2 66674 74622
0 11547 5 2 1 93917
0 11548 7 1 2 86954 93918
0 11549 5 1 1 11548
0 11550 7 1 2 86261 11549
0 11551 5 1 1 11550
0 11552 7 1 2 89984 11551
0 11553 5 1 1 11552
0 11554 7 1 2 77823 89393
0 11555 7 1 2 89604 11554
0 11556 5 1 1 11555
0 11557 7 1 2 11553 11556
0 11558 5 1 1 11557
0 11559 7 1 2 85228 11558
0 11560 5 1 1 11559
0 11561 7 1 2 11545 11560
0 11562 7 1 2 11502 11561
0 11563 5 1 1 11562
0 11564 7 1 2 11563 88064
0 11565 5 1 1 11564
0 11566 7 1 2 74875 88164
0 11567 5 2 1 11566
0 11568 7 4 2 65335 87634
0 11569 5 2 1 93923
0 11570 7 7 2 65336 74623
0 11571 5 3 1 93929
0 11572 7 1 2 74943 87241
0 11573 7 1 2 93936 11572
0 11574 7 1 2 93927 11573
0 11575 5 1 1 11574
0 11576 7 1 2 88534 11575
0 11577 5 1 1 11576
0 11578 7 1 2 93921 11577
0 11579 5 1 1 11578
0 11580 7 1 2 85229 11579
0 11581 5 1 1 11580
0 11582 7 4 2 66481 87635
0 11583 5 1 1 93939
0 11584 7 2 2 90109 11583
0 11585 5 3 1 93943
0 11586 7 1 2 65020 93945
0 11587 5 2 1 11586
0 11588 7 1 2 66208 75586
0 11589 5 3 1 11588
0 11590 7 1 2 67972 89619
0 11591 5 2 1 11590
0 11592 7 1 2 73398 93953
0 11593 5 1 1 11592
0 11594 7 1 2 93950 11593
0 11595 7 1 2 93948 11594
0 11596 5 1 1 11595
0 11597 7 1 2 88535 11596
0 11598 5 1 1 11597
0 11599 7 1 2 71598 90462
0 11600 5 4 1 11599
0 11601 7 2 2 77498 89344
0 11602 5 2 1 93959
0 11603 7 2 2 72129 75005
0 11604 7 1 2 68964 93963
0 11605 5 1 1 11604
0 11606 7 1 2 93961 11605
0 11607 5 1 1 11606
0 11608 7 1 2 93955 11607
0 11609 5 1 1 11608
0 11610 7 6 2 67973 82962
0 11611 5 2 1 93965
0 11612 7 2 2 74624 93971
0 11613 5 1 1 93973
0 11614 7 1 2 79494 81514
0 11615 7 1 2 11613 11614
0 11616 5 1 1 11615
0 11617 7 1 2 88165 11616
0 11618 5 1 1 11617
0 11619 7 1 2 11609 11618
0 11620 7 1 2 11598 11619
0 11621 5 1 1 11620
0 11622 7 1 2 85877 11621
0 11623 5 1 1 11622
0 11624 7 1 2 11581 11623
0 11625 5 1 1 11624
0 11626 7 1 2 11625 88962
0 11627 5 1 1 11626
0 11628 7 1 2 11565 11627
0 11629 5 1 1 11628
0 11630 7 1 2 64636 11629
0 11631 5 1 1 11630
0 11632 7 1 2 83157 88166
0 11633 5 1 1 11632
0 11634 7 2 2 70128 82894
0 11635 5 5 1 93975
0 11636 7 1 2 88376 89201
0 11637 5 4 1 11636
0 11638 7 1 2 93977 93982
0 11639 5 1 1 11638
0 11640 7 1 2 88536 11639
0 11641 5 1 1 11640
0 11642 7 1 2 11633 11641
0 11643 5 1 1 11642
0 11644 7 1 2 73399 11643
0 11645 5 1 1 11644
0 11646 7 2 2 67076 88470
0 11647 7 1 2 77499 93986
0 11648 5 1 1 11647
0 11649 7 1 2 11645 11648
0 11650 5 1 1 11649
0 11651 7 1 2 85230 11650
0 11652 5 1 1 11651
0 11653 7 1 2 93913 11652
0 11654 5 1 1 11653
0 11655 7 1 2 88065 11654
0 11656 5 1 1 11655
0 11657 7 1 2 75042 89291
0 11658 5 1 1 11657
0 11659 7 3 2 82895 88537
0 11660 5 2 1 93988
0 11661 7 1 2 89993 93991
0 11662 7 1 2 11658 11661
0 11663 5 1 1 11662
0 11664 7 1 2 85878 11663
0 11665 5 1 1 11664
0 11666 7 1 2 89323 11665
0 11667 5 1 1 11666
0 11668 7 1 2 88963 11667
0 11669 5 1 1 11668
0 11670 7 1 2 11656 11669
0 11671 5 1 1 11670
0 11672 7 1 2 66209 11671
0 11673 5 1 1 11672
0 11674 7 2 2 75265 91692
0 11675 7 1 2 92117 91554
0 11676 7 1 2 93993 11675
0 11677 5 1 1 11676
0 11678 7 1 2 91578 11677
0 11679 5 1 1 11678
0 11680 7 1 2 85231 11679
0 11681 5 1 1 11680
0 11682 7 2 2 74625 90905
0 11683 5 1 1 93995
0 11684 7 1 2 88167 93996
0 11685 5 1 1 11684
0 11686 7 1 2 11681 11685
0 11687 5 1 1 11686
0 11688 7 1 2 65337 11687
0 11689 5 1 1 11688
0 11690 7 4 2 68802 63968
0 11691 7 2 2 87436 93997
0 11692 7 3 2 65628 66482
0 11693 7 1 2 94003 91397
0 11694 7 1 2 76899 11693
0 11695 7 1 2 94001 11694
0 11696 5 1 1 11695
0 11697 7 1 2 11689 11696
0 11698 5 1 1 11697
0 11699 7 1 2 87636 11698
0 11700 5 1 1 11699
0 11701 7 1 2 79819 91373
0 11702 5 1 1 11701
0 11703 7 2 2 78570 89985
0 11704 7 1 2 86394 90529
0 11705 7 1 2 94006 11704
0 11706 5 1 1 11705
0 11707 7 1 2 11702 11706
0 11708 5 1 1 11707
0 11709 7 1 2 85232 11708
0 11710 5 1 1 11709
0 11711 7 5 2 73697 82591
0 11712 7 1 2 94008 76900
0 11713 7 1 2 90434 11712
0 11714 5 1 1 11713
0 11715 7 1 2 11710 11714
0 11716 5 1 1 11715
0 11717 7 1 2 74626 11716
0 11718 5 1 1 11717
0 11719 7 2 2 71324 87506
0 11720 5 1 1 94013
0 11721 7 3 2 71917 72130
0 11722 7 1 2 73698 94015
0 11723 7 1 2 94014 11722
0 11724 7 1 2 91278 11723
0 11725 5 1 1 11724
0 11726 7 1 2 9261 11725
0 11727 5 1 1 11726
0 11728 7 1 2 85233 11727
0 11729 5 1 1 11728
0 11730 7 1 2 86881 91219
0 11731 5 1 1 11730
0 11732 7 1 2 11729 11731
0 11733 5 1 1 11732
0 11734 7 1 2 73400 11733
0 11735 5 1 1 11734
0 11736 7 1 2 75525 89924
0 11737 5 3 1 11736
0 11738 7 1 2 63756 86555
0 11739 5 3 1 11738
0 11740 7 1 2 94018 94021
0 11741 5 1 1 11740
0 11742 7 1 2 65338 92244
0 11743 7 1 2 11741 11742
0 11744 5 1 1 11743
0 11745 7 1 2 11735 11744
0 11746 7 1 2 11718 11745
0 11747 7 1 2 11700 11746
0 11748 7 1 2 11673 11747
0 11749 5 1 1 11748
0 11750 7 1 2 72995 11749
0 11751 5 1 1 11750
0 11752 7 1 2 82896 89107
0 11753 5 1 1 11752
0 11754 7 2 2 63757 86084
0 11755 5 1 1 94024
0 11756 7 1 2 11753 11755
0 11757 5 1 1 11756
0 11758 7 1 2 88538 11757
0 11759 5 1 1 11758
0 11760 7 2 2 86021 93916
0 11761 5 1 1 94026
0 11762 7 1 2 85879 94027
0 11763 5 1 1 11762
0 11764 7 1 2 11759 11763
0 11765 5 1 1 11764
0 11766 7 1 2 66210 11765
0 11767 5 1 1 11766
0 11768 7 6 2 63758 66675
0 11769 7 3 2 94028 86564
0 11770 5 1 1 94034
0 11771 7 1 2 65339 92687
0 11772 5 1 1 11771
0 11773 7 1 2 93903 11772
0 11774 5 2 1 11773
0 11775 7 1 2 94035 94037
0 11776 5 1 1 11775
0 11777 7 1 2 11767 11776
0 11778 5 1 1 11777
0 11779 7 1 2 88964 11778
0 11780 5 1 1 11779
0 11781 7 2 2 83214 74283
0 11782 7 1 2 81700 87918
0 11783 7 1 2 94039 11782
0 11784 7 1 2 90302 11783
0 11785 5 1 1 11784
0 11786 7 1 2 11780 11785
0 11787 5 1 1 11786
0 11788 7 1 2 74627 11787
0 11789 5 1 1 11788
0 11790 7 2 2 82897 83040
0 11791 5 3 1 94041
0 11792 7 1 2 75356 94043
0 11793 5 1 1 11792
0 11794 7 1 2 88168 11793
0 11795 5 1 1 11794
0 11796 7 1 2 93940 90169
0 11797 5 1 1 11796
0 11798 7 1 2 11795 11797
0 11799 5 1 1 11798
0 11800 7 1 2 90906 11799
0 11801 5 1 1 11800
0 11802 7 1 2 93924 88539
0 11803 5 1 1 11802
0 11804 7 1 2 93922 11803
0 11805 5 1 1 11804
0 11806 7 1 2 88965 11805
0 11807 5 1 1 11806
0 11808 7 3 2 73401 93989
0 11809 5 1 1 94046
0 11810 7 1 2 67974 94047
0 11811 5 2 1 11810
0 11812 7 1 2 65340 89785
0 11813 5 1 1 11812
0 11814 7 1 2 94049 11813
0 11815 5 1 1 11814
0 11816 7 2 2 78342 90530
0 11817 7 1 2 65021 94051
0 11818 7 1 2 11815 11817
0 11819 5 1 1 11818
0 11820 7 1 2 11807 11819
0 11821 5 1 1 11820
0 11822 7 1 2 85234 11821
0 11823 5 1 1 11822
0 11824 7 1 2 11801 11823
0 11825 5 1 1 11824
0 11826 7 1 2 66211 11825
0 11827 5 1 1 11826
0 11828 7 1 2 85235 92624
0 11829 5 1 1 11828
0 11830 7 1 2 82898 92209
0 11831 5 1 1 11830
0 11832 7 1 2 11829 11831
0 11833 5 1 1 11832
0 11834 7 1 2 73402 11833
0 11835 5 1 1 11834
0 11836 7 5 2 66957 94029
0 11837 7 1 2 94053 90157
0 11838 5 1 1 11837
0 11839 7 1 2 11835 11838
0 11840 5 1 1 11839
0 11841 7 1 2 75266 88966
0 11842 7 1 2 11840 11841
0 11843 5 1 1 11842
0 11844 7 1 2 11827 11843
0 11845 7 1 2 11789 11844
0 11846 7 1 2 11751 11845
0 11847 7 1 2 11631 11846
0 11848 5 1 1 11847
0 11849 7 1 2 65946 11848
0 11850 5 1 1 11849
0 11851 7 1 2 74731 87919
0 11852 7 1 2 90531 11851
0 11853 5 1 1 11852
0 11854 7 1 2 8374 11853
0 11855 5 1 1 11854
0 11856 7 1 2 90688 11855
0 11857 5 1 1 11856
0 11858 7 1 2 76069 91983
0 11859 5 1 1 11858
0 11860 7 1 2 89010 11859
0 11861 5 1 1 11860
0 11862 7 1 2 86001 11861
0 11863 5 1 1 11862
0 11864 7 1 2 11857 11863
0 11865 5 1 1 11864
0 11866 7 1 2 66483 11865
0 11867 5 1 1 11866
0 11868 7 3 2 91894 92017
0 11869 7 5 2 66958 68329
0 11870 7 3 2 72996 87920
0 11871 7 1 2 94061 94066
0 11872 7 1 2 94058 11871
0 11873 5 1 1 11872
0 11874 7 1 2 11867 11873
0 11875 5 1 1 11874
0 11876 7 1 2 65022 11875
0 11877 5 1 1 11876
0 11878 7 7 2 64637 65583
0 11879 7 2 2 88889 94069
0 11880 7 1 2 88914 94076
0 11881 5 1 1 11880
0 11882 7 11 2 69058 91164
0 11883 7 1 2 94067 86015
0 11884 7 1 2 94078 11883
0 11885 5 1 1 11884
0 11886 7 1 2 11881 11885
0 11887 5 1 1 11886
0 11888 7 1 2 86002 11887
0 11889 5 1 1 11888
0 11890 7 2 2 72997 91962
0 11891 7 1 2 84972 92228
0 11892 7 1 2 94089 11891
0 11893 5 1 1 11892
0 11894 7 1 2 11889 11893
0 11895 7 1 2 11877 11894
0 11896 5 1 1 11895
0 11897 7 1 2 88540 11896
0 11898 5 1 1 11897
0 11899 7 3 2 91165 91710
0 11900 7 1 2 79689 76881
0 11901 7 1 2 94091 11900
0 11902 5 1 1 11901
0 11903 7 1 2 89011 11902
0 11904 5 1 1 11903
0 11905 7 1 2 85236 11904
0 11906 5 1 1 11905
0 11907 7 1 2 73403 91965
0 11908 5 1 1 11907
0 11909 7 1 2 11906 11908
0 11910 5 1 1 11909
0 11911 7 1 2 88541 11910
0 11912 5 1 1 11911
0 11913 7 1 2 79601 91213
0 11914 5 1 1 11913
0 11915 7 1 2 11912 11914
0 11916 5 1 1 11915
0 11917 7 1 2 74628 11916
0 11918 5 1 1 11917
0 11919 7 1 2 65341 90438
0 11920 5 1 1 11919
0 11921 7 4 2 75736 89345
0 11922 7 1 2 90303 94094
0 11923 5 1 1 11922
0 11924 7 1 2 11920 11923
0 11925 5 1 1 11924
0 11926 7 1 2 79835 11925
0 11927 5 1 1 11926
0 11928 7 3 2 63969 79367
0 11929 7 1 2 79077 94098
0 11930 7 1 2 91260 11929
0 11931 5 1 1 11930
0 11932 7 1 2 11927 11931
0 11933 7 1 2 11918 11932
0 11934 5 1 1 11933
0 11935 7 1 2 75006 11934
0 11936 5 1 1 11935
0 11937 7 1 2 93962 6295
0 11938 5 1 1 11937
0 11939 7 1 2 85237 11938
0 11940 5 1 1 11939
0 11941 7 1 2 64638 94038
0 11942 5 1 1 11941
0 11943 7 1 2 66212 89986
0 11944 5 1 1 11943
0 11945 7 1 2 11942 11944
0 11946 5 1 1 11945
0 11947 7 1 2 85880 11946
0 11948 5 1 1 11947
0 11949 7 1 2 11940 11948
0 11950 5 1 1 11949
0 11951 7 1 2 88967 11950
0 11952 5 1 1 11951
0 11953 7 1 2 85238 78819
0 11954 5 1 1 11953
0 11955 7 1 2 68803 75644
0 11956 7 1 2 77961 77027
0 11957 7 1 2 11955 11956
0 11958 5 1 1 11957
0 11959 7 1 2 11954 11958
0 11960 5 1 1 11959
0 11961 7 1 2 91518 11960
0 11962 5 1 1 11961
0 11963 7 1 2 11952 11962
0 11964 5 1 1 11963
0 11965 7 1 2 74629 11964
0 11966 5 1 1 11965
0 11967 7 2 2 79368 91403
0 11968 7 4 2 74732 74234
0 11969 7 2 2 64639 76882
0 11970 7 1 2 69059 94107
0 11971 7 1 2 94103 11970
0 11972 7 1 2 94101 11971
0 11973 5 1 1 11972
0 11974 7 1 2 91226 11973
0 11975 5 1 1 11974
0 11976 7 1 2 79503 11975
0 11977 5 1 1 11976
0 11978 7 3 2 94070 89540
0 11979 7 3 2 94090 94109
0 11980 5 1 1 94112
0 11981 7 1 2 75965 92006
0 11982 5 2 1 11981
0 11983 7 2 2 73404 94115
0 11984 5 1 1 94117
0 11985 7 1 2 94118 91904
0 11986 5 1 1 11985
0 11987 7 1 2 11980 11986
0 11988 5 1 1 11987
0 11989 7 1 2 88169 11988
0 11990 5 1 1 11989
0 11991 7 1 2 11977 11990
0 11992 7 1 2 11966 11991
0 11993 7 1 2 11936 11992
0 11994 7 1 2 11898 11993
0 11995 5 1 1 11994
0 11996 7 1 2 65947 11995
0 11997 5 1 1 11996
0 11998 7 2 2 77656 89894
0 11999 7 2 2 70618 94119
0 12000 7 1 2 70661 91895
0 12001 7 3 2 93624 12000
0 12002 7 3 2 78951 81584
0 12003 7 1 2 87908 94126
0 12004 7 1 2 94123 12003
0 12005 7 1 2 94121 12004
0 12006 5 1 1 12005
0 12007 7 1 2 11997 12006
0 12008 5 1 1 12007
0 12009 7 1 2 80394 12008
0 12010 5 1 1 12009
0 12011 7 2 2 90188 74235
0 12012 7 2 2 88702 78343
0 12013 7 9 2 64640 70619
0 12014 7 1 2 77824 94133
0 12015 7 1 2 94131 12014
0 12016 7 1 2 94124 12015
0 12017 7 1 2 94129 12016
0 12018 5 1 1 12017
0 12019 7 1 2 12010 12018
0 12020 7 1 2 11850 12019
0 12021 5 1 1 12020
0 12022 7 1 2 64316 12021
0 12023 5 1 1 12022
0 12024 7 3 2 78952 82526
0 12025 7 2 2 66484 94142
0 12026 7 1 2 86395 91693
0 12027 7 1 2 94145 12026
0 12028 7 1 2 94130 12027
0 12029 5 1 1 12028
0 12030 7 4 2 70662 91600
0 12031 7 1 2 87565 81299
0 12032 7 1 2 94147 12031
0 12033 7 1 2 94122 12032
0 12034 5 1 1 12033
0 12035 7 1 2 12029 12034
0 12036 5 1 1 12035
0 12037 7 1 2 91896 89119
0 12038 7 1 2 12036 12037
0 12039 5 1 1 12038
0 12040 7 1 2 12023 12039
0 12041 5 1 1 12040
0 12042 7 1 2 67588 12041
0 12043 5 1 1 12042
0 12044 7 2 2 73954 86866
0 12045 5 2 1 94151
0 12046 7 1 2 81701 90089
0 12047 5 1 1 12046
0 12048 7 1 2 94153 12047
0 12049 5 1 1 12048
0 12050 7 1 2 81020 12049
0 12051 5 1 1 12050
0 12052 7 3 2 86666 73900
0 12053 5 1 1 94155
0 12054 7 2 2 65948 94156
0 12055 5 2 1 94158
0 12056 7 2 2 69446 81585
0 12057 7 1 2 90103 94162
0 12058 5 1 1 12057
0 12059 7 1 2 94160 12058
0 12060 5 1 1 12059
0 12061 7 1 2 70129 12060
0 12062 5 1 1 12061
0 12063 7 1 2 86775 80988
0 12064 5 1 1 12063
0 12065 7 1 2 69447 86765
0 12066 5 1 1 12065
0 12067 7 1 2 88665 12066
0 12068 5 1 1 12067
0 12069 7 1 2 87558 12068
0 12070 5 1 1 12069
0 12071 7 1 2 12064 12070
0 12072 7 1 2 12062 12071
0 12073 5 1 1 12072
0 12074 7 1 2 64641 12073
0 12075 5 1 1 12074
0 12076 7 1 2 12051 12075
0 12077 5 1 1 12076
0 12078 7 1 2 88066 12077
0 12079 5 1 1 12078
0 12080 7 1 2 85673 77414
0 12081 5 1 1 12080
0 12082 7 1 2 84923 89209
0 12083 5 2 1 12082
0 12084 7 1 2 68330 94164
0 12085 5 1 1 12084
0 12086 7 1 2 12081 12085
0 12087 5 1 1 12086
0 12088 7 1 2 64642 12087
0 12089 5 1 1 12088
0 12090 7 1 2 12089 4535
0 12091 5 1 1 12090
0 12092 7 1 2 88968 12091
0 12093 5 1 1 12092
0 12094 7 1 2 12079 12093
0 12095 5 1 1 12094
0 12096 7 1 2 85239 12095
0 12097 5 1 1 12096
0 12098 7 4 2 66485 84817
0 12099 5 1 1 94166
0 12100 7 1 2 86339 94167
0 12101 5 1 1 12100
0 12102 7 1 2 69769 12101
0 12103 5 1 1 12102
0 12104 7 2 2 93790 12103
0 12105 7 1 2 94170 80989
0 12106 5 1 1 12105
0 12107 7 5 2 64317 84818
0 12108 7 2 2 73699 94172
0 12109 5 2 1 94177
0 12110 7 1 2 93446 94178
0 12111 5 1 1 12110
0 12112 7 1 2 12106 12111
0 12113 5 1 1 12112
0 12114 7 1 2 68331 12113
0 12115 5 1 1 12114
0 12116 7 2 2 82315 88686
0 12117 5 5 1 94181
0 12118 7 1 2 73405 94183
0 12119 5 3 1 12118
0 12120 7 2 2 94188 93778
0 12121 5 2 1 94191
0 12122 7 2 2 65949 94193
0 12123 5 1 1 94195
0 12124 7 1 2 80015 94196
0 12125 5 1 1 12124
0 12126 7 1 2 12115 12125
0 12127 5 1 1 12126
0 12128 7 1 2 88067 12127
0 12129 5 1 1 12128
0 12130 7 1 2 68608 82668
0 12131 7 1 2 83786 12130
0 12132 5 1 1 12131
0 12133 7 1 2 64643 88790
0 12134 5 2 1 12133
0 12135 7 1 2 89609 94197
0 12136 5 1 1 12135
0 12137 7 1 2 65023 12136
0 12138 5 1 1 12137
0 12139 7 1 2 64644 93946
0 12140 5 1 1 12139
0 12141 7 1 2 12138 12140
0 12142 5 1 1 12141
0 12143 7 1 2 71020 12142
0 12144 5 1 1 12143
0 12145 7 1 2 12132 12144
0 12146 5 1 1 12145
0 12147 7 1 2 65342 12146
0 12148 5 1 1 12147
0 12149 7 2 2 80395 87698
0 12150 5 2 1 94199
0 12151 7 1 2 86262 94201
0 12152 5 1 1 12151
0 12153 7 1 2 84405 12152
0 12154 5 1 1 12153
0 12155 7 2 2 68332 84960
0 12156 5 1 1 94203
0 12157 7 6 2 70376 90230
0 12158 7 1 2 73406 94205
0 12159 5 1 1 12158
0 12160 7 1 2 12156 12159
0 12161 5 1 1 12160
0 12162 7 1 2 69770 12161
0 12163 5 1 1 12162
0 12164 7 1 2 80912 81021
0 12165 5 1 1 12164
0 12166 7 1 2 82963 86176
0 12167 7 1 2 80226 12166
0 12168 5 1 1 12167
0 12169 7 1 2 86514 12168
0 12170 5 1 1 12169
0 12171 7 1 2 87122 12170
0 12172 5 1 1 12171
0 12173 7 1 2 12165 12172
0 12174 7 1 2 12163 12173
0 12175 7 1 2 12154 12174
0 12176 7 1 2 12148 12175
0 12177 5 1 1 12176
0 12178 7 1 2 88969 12177
0 12179 5 1 1 12178
0 12180 7 1 2 12129 12179
0 12181 5 1 1 12180
0 12182 7 1 2 85881 12181
0 12183 5 1 1 12182
0 12184 7 1 2 12097 12183
0 12185 5 1 1 12184
0 12186 7 1 2 88170 12185
0 12187 5 1 1 12186
0 12188 7 1 2 82305 80396
0 12189 5 1 1 12188
0 12190 7 1 2 88768 12189
0 12191 5 2 1 12190
0 12192 7 1 2 71599 94211
0 12193 5 1 1 12192
0 12194 7 2 2 80541 80847
0 12195 5 1 1 94213
0 12196 7 1 2 12193 12195
0 12197 5 1 1 12196
0 12198 7 1 2 89113 12197
0 12199 5 1 1 12198
0 12200 7 6 2 65343 87507
0 12201 5 1 1 94215
0 12202 7 2 2 76745 94216
0 12203 7 1 2 94221 93393
0 12204 5 1 1 12203
0 12205 7 1 2 12199 12204
0 12206 5 1 1 12205
0 12207 7 1 2 73407 12206
0 12208 5 1 1 12207
0 12209 7 5 2 72023 90206
0 12210 5 1 1 94223
0 12211 7 1 2 68333 94224
0 12212 5 1 1 12211
0 12213 7 1 2 85354 12212
0 12214 5 1 1 12213
0 12215 7 1 2 93876 12214
0 12216 5 1 1 12215
0 12217 7 3 2 81702 89067
0 12218 5 1 1 94228
0 12219 7 1 2 71600 94229
0 12220 5 1 1 12219
0 12221 7 1 2 90012 12220
0 12222 5 1 1 12221
0 12223 7 1 2 85882 12222
0 12224 5 1 1 12223
0 12225 7 1 2 12216 12224
0 12226 5 1 1 12225
0 12227 7 1 2 65950 12226
0 12228 5 1 1 12227
0 12229 7 1 2 12208 12228
0 12230 5 1 1 12229
0 12231 7 8 2 69448 70620
0 12232 7 5 2 88050 90524
0 12233 7 5 2 94231 94239
0 12234 7 1 2 12230 94244
0 12235 5 1 1 12234
0 12236 7 1 2 84797 79709
0 12237 5 3 1 12236
0 12238 7 1 2 65024 94249
0 12239 5 1 1 12238
0 12240 7 1 2 88669 12239
0 12241 5 1 1 12240
0 12242 7 1 2 71601 12241
0 12243 5 1 1 12242
0 12244 7 1 2 82866 12243
0 12245 5 2 1 12244
0 12246 7 2 2 68334 94252
0 12247 5 2 1 94254
0 12248 7 4 2 66486 80677
0 12249 5 10 1 94258
0 12250 7 4 2 85621 94262
0 12251 5 3 1 94272
0 12252 7 8 2 78687 94273
0 12253 5 7 1 94279
0 12254 7 1 2 86364 94280
0 12255 5 1 1 12254
0 12256 7 1 2 77415 12255
0 12257 5 1 1 12256
0 12258 7 1 2 94256 12257
0 12259 5 1 1 12258
0 12260 7 1 2 85240 12259
0 12261 5 1 1 12260
0 12262 7 1 2 80397 93925
0 12263 5 1 1 12262
0 12264 7 2 2 90110 12263
0 12265 5 3 1 94294
0 12266 7 1 2 66487 94296
0 12267 5 2 1 12266
0 12268 7 1 2 68609 85649
0 12269 5 1 1 12268
0 12270 7 1 2 66488 12269
0 12271 5 1 1 12270
0 12272 7 1 2 94295 12271
0 12273 5 2 1 12272
0 12274 7 1 2 65025 94301
0 12275 5 1 1 12274
0 12276 7 1 2 94299 12275
0 12277 5 2 1 12276
0 12278 7 1 2 69449 94303
0 12279 5 1 1 12278
0 12280 7 4 2 68335 87059
0 12281 7 1 2 64318 94305
0 12282 5 1 1 12281
0 12283 7 1 2 81005 12282
0 12284 7 1 2 12279 12283
0 12285 5 1 1 12284
0 12286 7 1 2 85883 12285
0 12287 5 1 1 12286
0 12288 7 1 2 12261 12287
0 12289 5 1 1 12288
0 12290 7 1 2 88970 12289
0 12291 5 1 1 12290
0 12292 7 1 2 12235 12291
0 12293 5 1 1 12292
0 12294 7 1 2 64645 12293
0 12295 5 1 1 12294
0 12296 7 1 2 75267 75120
0 12297 5 1 1 12296
0 12298 7 1 2 83695 87230
0 12299 5 1 1 12298
0 12300 7 1 2 12297 12299
0 12301 5 1 1 12300
0 12302 7 1 2 71787 12301
0 12303 5 1 1 12302
0 12304 7 1 2 65026 78013
0 12305 7 1 2 82715 12304
0 12306 5 1 1 12305
0 12307 7 1 2 12303 12306
0 12308 5 1 1 12307
0 12309 7 1 2 91905 12308
0 12310 5 1 1 12309
0 12311 7 1 2 85779 90326
0 12312 5 1 1 12311
0 12313 7 1 2 12310 12312
0 12314 5 1 1 12313
0 12315 7 1 2 81022 12314
0 12316 5 1 1 12315
0 12317 7 5 2 70130 87123
0 12318 7 1 2 89108 90700
0 12319 7 2 2 94309 12318
0 12320 5 1 1 94314
0 12321 7 4 2 85241 75268
0 12322 5 1 1 94316
0 12323 7 6 2 65344 77416
0 12324 7 5 2 82899 94320
0 12325 5 1 1 94326
0 12326 7 1 2 94317 94327
0 12327 5 1 1 12326
0 12328 7 1 2 12320 12327
0 12329 5 1 1 12328
0 12330 7 1 2 88971 12329
0 12331 5 1 1 12330
0 12332 7 1 2 12316 12331
0 12333 7 1 2 12295 12332
0 12334 5 1 1 12333
0 12335 7 1 2 88542 12334
0 12336 5 1 1 12335
0 12337 7 1 2 12187 12336
0 12338 5 1 1 12337
0 12339 7 1 2 72998 12338
0 12340 5 1 1 12339
0 12341 7 2 2 80244 74822
0 12342 7 1 2 94331 94245
0 12343 5 1 1 12342
0 12344 7 1 2 87615 88972
0 12345 5 1 1 12344
0 12346 7 1 2 12343 12345
0 12347 5 1 1 12346
0 12348 7 1 2 66676 12347
0 12349 5 1 1 12348
0 12350 7 2 2 86500 91341
0 12351 7 2 2 78634 88051
0 12352 7 1 2 70663 94335
0 12353 7 1 2 94333 12352
0 12354 5 1 1 12353
0 12355 7 1 2 12349 12354
0 12356 5 1 1 12355
0 12357 7 1 2 65345 12356
0 12358 5 1 1 12357
0 12359 7 4 2 92146 89505
0 12360 7 3 2 70131 71918
0 12361 7 2 2 73901 94341
0 12362 7 1 2 94337 94344
0 12363 5 1 1 12362
0 12364 7 1 2 82101 91254
0 12365 7 1 2 90744 12364
0 12366 5 1 1 12365
0 12367 7 1 2 12363 12366
0 12368 5 1 1 12367
0 12369 7 1 2 80579 12368
0 12370 5 1 1 12369
0 12371 7 2 2 78344 91166
0 12372 7 1 2 80503 94334
0 12373 7 1 2 94346 12372
0 12374 5 1 1 12373
0 12375 7 1 2 12370 12374
0 12376 7 1 2 12358 12375
0 12377 5 1 1 12376
0 12378 7 1 2 90689 12377
0 12379 5 1 1 12378
0 12380 7 2 2 87242 75486
0 12381 5 1 1 94348
0 12382 7 1 2 77119 12381
0 12383 5 1 1 12382
0 12384 7 1 2 90231 12383
0 12385 5 1 1 12384
0 12386 7 2 2 69450 86251
0 12387 5 1 1 94350
0 12388 7 1 2 86030 94351
0 12389 5 1 1 12388
0 12390 7 1 2 12385 12389
0 12391 5 1 1 12390
0 12392 7 1 2 91906 12391
0 12393 5 1 1 12392
0 12394 7 1 2 12379 12393
0 12395 5 1 1 12394
0 12396 7 1 2 88543 12395
0 12397 5 1 1 12396
0 12398 7 4 2 81703 75269
0 12399 5 3 1 94352
0 12400 7 4 2 73408 88418
0 12401 5 1 1 94359
0 12402 7 1 2 94356 12401
0 12403 5 2 1 12402
0 12404 7 1 2 94363 94246
0 12405 5 1 1 12404
0 12406 7 1 2 88757 88973
0 12407 5 1 1 12406
0 12408 7 1 2 93666 90786
0 12409 5 1 1 12408
0 12410 7 3 2 79802 90232
0 12411 5 1 1 94365
0 12412 7 2 2 68610 88068
0 12413 7 1 2 94366 94368
0 12414 5 1 1 12413
0 12415 7 1 2 12409 12414
0 12416 5 1 1 12415
0 12417 7 1 2 75357 12416
0 12418 5 1 1 12417
0 12419 7 1 2 12407 12418
0 12420 7 1 2 12405 12419
0 12421 5 1 1 12420
0 12422 7 1 2 64646 12421
0 12423 5 1 1 12422
0 12424 7 1 2 87357 91202
0 12425 5 1 1 12424
0 12426 7 5 2 86605 93676
0 12427 7 1 2 87101 94370
0 12428 5 1 1 12427
0 12429 7 1 2 12425 12428
0 12430 5 1 1 12429
0 12431 7 1 2 64319 12430
0 12432 5 1 1 12431
0 12433 7 1 2 12423 12432
0 12434 5 1 1 12433
0 12435 7 1 2 85884 12434
0 12436 5 1 1 12435
0 12437 7 1 2 83173 91728
0 12438 5 1 1 12437
0 12439 7 1 2 79237 12438
0 12440 5 2 1 12439
0 12441 7 1 2 82000 94375
0 12442 5 1 1 12441
0 12443 7 3 2 82900 79904
0 12444 5 1 1 94377
0 12445 7 1 2 69451 94378
0 12446 5 1 1 12445
0 12447 7 1 2 12442 12446
0 12448 5 1 1 12447
0 12449 7 1 2 65346 12448
0 12450 5 1 1 12449
0 12451 7 3 2 66489 83391
0 12452 5 3 1 94380
0 12453 7 3 2 75636 7459
0 12454 5 3 1 94386
0 12455 7 1 2 80480 94389
0 12456 5 1 1 12455
0 12457 7 1 2 94383 12456
0 12458 5 2 1 12457
0 12459 7 1 2 82001 94392
0 12460 5 1 1 12459
0 12461 7 1 2 12411 12460
0 12462 7 1 2 12450 12461
0 12463 5 1 1 12462
0 12464 7 1 2 91907 12463
0 12465 5 1 1 12464
0 12466 7 1 2 12436 12465
0 12467 5 1 1 12466
0 12468 7 1 2 88171 12467
0 12469 5 1 1 12468
0 12470 7 1 2 12397 12469
0 12471 5 1 1 12470
0 12472 7 1 2 67975 12471
0 12473 5 1 1 12472
0 12474 7 6 2 68804 82002
0 12475 7 1 2 94394 77764
0 12476 5 2 1 12475
0 12477 7 1 2 90727 94400
0 12478 5 1 1 12477
0 12479 7 1 2 94369 12478
0 12480 5 1 1 12479
0 12481 7 1 2 90915 12480
0 12482 5 1 1 12481
0 12483 7 1 2 82787 12482
0 12484 5 1 1 12483
0 12485 7 1 2 63970 89109
0 12486 7 2 2 65584 82003
0 12487 7 1 2 94402 92285
0 12488 7 1 2 12485 12487
0 12489 5 1 1 12488
0 12490 7 1 2 12484 12489
0 12491 5 1 1 12490
0 12492 7 1 2 67976 12491
0 12493 5 1 1 12492
0 12494 7 2 2 63759 80016
0 12495 7 2 2 68611 73955
0 12496 7 3 2 80925 94406
0 12497 7 1 2 94404 94408
0 12498 7 1 2 90612 12497
0 12499 5 1 1 12498
0 12500 7 1 2 12493 12499
0 12501 5 1 1 12500
0 12502 7 1 2 88544 12501
0 12503 5 1 1 12502
0 12504 7 3 2 68805 91555
0 12505 7 2 2 91888 94411
0 12506 7 2 2 75554 76838
0 12507 7 1 2 82004 92147
0 12508 7 1 2 94416 12507
0 12509 7 1 2 94414 12508
0 12510 5 1 1 12509
0 12511 7 1 2 12503 12510
0 12512 5 1 1 12511
0 12513 7 1 2 81838 12512
0 12514 5 1 1 12513
0 12515 7 1 2 75121 94025
0 12516 5 1 1 12515
0 12517 7 1 2 68806 83537
0 12518 5 1 1 12517
0 12519 7 2 2 90707 12518
0 12520 7 1 2 68612 85355
0 12521 5 2 1 12520
0 12522 7 1 2 84819 94420
0 12523 7 1 2 94418 12522
0 12524 5 1 1 12523
0 12525 7 1 2 12516 12524
0 12526 5 1 1 12525
0 12527 7 1 2 66490 12526
0 12528 5 1 1 12527
0 12529 7 1 2 85242 86874
0 12530 5 1 1 12529
0 12531 7 1 2 12528 12530
0 12532 5 2 1 12531
0 12533 7 1 2 88172 94422
0 12534 5 1 1 12533
0 12535 7 1 2 88388 83560
0 12536 5 2 1 12535
0 12537 7 2 2 74630 80580
0 12538 5 1 1 94426
0 12539 7 2 2 80245 94427
0 12540 5 4 1 94428
0 12541 7 1 2 94424 94430
0 12542 5 1 1 12541
0 12543 7 1 2 89308 12542
0 12544 5 1 1 12543
0 12545 7 1 2 12534 12544
0 12546 5 1 1 12545
0 12547 7 1 2 88069 12546
0 12548 5 1 1 12547
0 12549 7 5 2 67077 80678
0 12550 7 5 2 63882 94434
0 12551 5 5 1 94439
0 12552 7 2 2 72131 85674
0 12553 7 1 2 68965 94449
0 12554 5 1 1 12553
0 12555 7 1 2 94444 12554
0 12556 5 2 1 12555
0 12557 7 2 2 76378 94451
0 12558 7 1 2 90327 94453
0 12559 5 1 1 12558
0 12560 7 1 2 12548 12559
0 12561 5 1 1 12560
0 12562 7 1 2 80017 12561
0 12563 5 1 1 12562
0 12564 7 1 2 12514 12563
0 12565 7 1 2 12473 12564
0 12566 5 1 1 12565
0 12567 7 1 2 65951 12566
0 12568 5 1 1 12567
0 12569 7 3 2 85572 94125
0 12570 7 1 2 94409 94455
0 12571 5 1 1 12570
0 12572 7 1 2 75555 90661
0 12573 7 1 2 90328 12572
0 12574 5 1 1 12573
0 12575 7 1 2 12571 12574
0 12576 5 1 1 12575
0 12577 7 1 2 81839 12576
0 12578 5 1 1 12577
0 12579 7 1 2 88389 83526
0 12580 5 1 1 12579
0 12581 7 1 2 94431 12580
0 12582 5 1 1 12581
0 12583 7 1 2 94456 12582
0 12584 5 1 1 12583
0 12585 7 1 2 12578 12584
0 12586 5 1 1 12585
0 12587 7 1 2 88545 12586
0 12588 5 1 1 12587
0 12589 7 1 2 71021 94423
0 12590 5 1 1 12589
0 12591 7 2 2 87330 82102
0 12592 5 1 1 94458
0 12593 7 1 2 85243 81431
0 12594 7 1 2 94459 12593
0 12595 5 1 1 12594
0 12596 7 1 2 12590 12595
0 12597 5 1 1 12596
0 12598 7 1 2 91519 12597
0 12599 5 1 1 12598
0 12600 7 1 2 12588 12599
0 12601 5 1 1 12600
0 12602 7 1 2 64320 12601
0 12603 5 1 1 12602
0 12604 7 2 2 75708 87611
0 12605 5 1 1 94460
0 12606 7 1 2 89994 12605
0 12607 5 2 1 12606
0 12608 7 1 2 80398 94462
0 12609 5 1 1 12608
0 12610 7 1 2 90468 88173
0 12611 5 1 1 12610
0 12612 7 1 2 83004 90170
0 12613 5 1 1 12612
0 12614 7 1 2 12611 12613
0 12615 7 1 2 12609 12614
0 12616 5 1 1 12615
0 12617 7 1 2 67977 12616
0 12618 5 1 1 12617
0 12619 7 1 2 94328 88546
0 12620 5 1 1 12619
0 12621 7 1 2 12618 12620
0 12622 5 1 1 12621
0 12623 7 1 2 85244 12622
0 12624 5 1 1 12623
0 12625 7 3 2 75504 87727
0 12626 7 13 2 71022 66677
0 12627 7 1 2 94467 79161
0 12628 7 1 2 94464 12627
0 12629 5 1 1 12628
0 12630 7 1 2 12624 12629
0 12631 5 1 1 12630
0 12632 7 1 2 73409 12631
0 12633 5 1 1 12632
0 12634 7 8 2 67978 81704
0 12635 5 2 1 94480
0 12636 7 1 2 86996 94488
0 12637 5 1 1 12636
0 12638 7 2 2 65027 89407
0 12639 7 1 2 12637 94490
0 12640 5 1 1 12639
0 12641 7 1 2 12633 12640
0 12642 5 1 1 12641
0 12643 7 1 2 66491 12642
0 12644 5 1 1 12643
0 12645 7 2 2 88390 74733
0 12646 7 1 2 94492 94491
0 12647 5 1 1 12646
0 12648 7 1 2 12644 12647
0 12649 5 1 1 12648
0 12650 7 1 2 88974 12649
0 12651 5 1 1 12650
0 12652 7 1 2 12603 12651
0 12653 5 1 1 12652
0 12654 7 1 2 64647 12653
0 12655 5 1 1 12654
0 12656 7 5 2 72132 80679
0 12657 7 4 2 83807 94494
0 12658 7 1 2 77825 94499
0 12659 5 1 1 12658
0 12660 7 1 2 12659 6730
0 12661 5 1 1 12660
0 12662 7 1 2 73410 75144
0 12663 7 2 2 12661 12662
0 12664 7 2 2 78345 94503
0 12665 7 1 2 87954 91897
0 12666 7 1 2 91622 12665
0 12667 7 1 2 94505 12666
0 12668 5 1 1 12667
0 12669 7 1 2 12655 12668
0 12670 7 1 2 12568 12669
0 12671 7 1 2 12340 12670
0 12672 5 1 1 12671
0 12673 7 1 2 66213 12672
0 12674 5 1 1 12673
0 12675 7 7 2 66678 77417
0 12676 7 1 2 94507 92613
0 12677 5 1 1 12676
0 12678 7 1 2 86978 88174
0 12679 5 1 1 12678
0 12680 7 1 2 12677 12679
0 12681 5 1 1 12680
0 12682 7 1 2 85245 12681
0 12683 5 1 1 12682
0 12684 7 2 2 89148 89346
0 12685 7 1 2 87728 76706
0 12686 7 1 2 94514 12685
0 12687 5 1 1 12686
0 12688 7 1 2 12683 12687
0 12689 5 1 1 12688
0 12690 7 1 2 88975 12689
0 12691 5 1 1 12690
0 12692 7 2 2 68336 87729
0 12693 7 1 2 72024 94516
0 12694 7 1 2 87588 12693
0 12695 7 1 2 90686 12694
0 12696 5 1 1 12695
0 12697 7 1 2 12691 12696
0 12698 5 1 1 12697
0 12699 7 1 2 73700 12698
0 12700 5 1 1 12699
0 12701 7 2 2 89166 89895
0 12702 7 1 2 89120 92215
0 12703 7 1 2 94518 12702
0 12704 5 1 1 12703
0 12705 7 1 2 12700 12704
0 12706 5 1 1 12705
0 12707 7 1 2 65028 12706
0 12708 5 1 1 12707
0 12709 7 1 2 83691 89847
0 12710 5 1 1 12709
0 12711 7 1 2 71788 92688
0 12712 5 1 1 12711
0 12713 7 1 2 88290 12712
0 12714 5 1 1 12713
0 12715 7 2 2 80990 90382
0 12716 7 3 2 75737 94520
0 12717 5 1 1 94522
0 12718 7 1 2 12714 94523
0 12719 7 1 2 12710 12718
0 12720 5 1 1 12719
0 12721 7 1 2 12708 12720
0 12722 5 1 1 12721
0 12723 7 1 2 66492 12722
0 12724 5 1 1 12723
0 12725 7 5 2 84592 76000
0 12726 5 1 1 94525
0 12727 7 1 2 94445 12726
0 12728 5 1 1 12727
0 12729 7 1 2 90907 12728
0 12730 5 1 1 12729
0 12731 7 6 2 65029 68613
0 12732 5 1 1 94530
0 12733 7 1 2 72133 12732
0 12734 5 1 1 12733
0 12735 7 2 2 89292 12734
0 12736 7 1 2 84820 94536
0 12737 5 1 1 12736
0 12738 7 1 2 83696 88175
0 12739 5 1 1 12738
0 12740 7 1 2 83418 94461
0 12741 5 1 1 12740
0 12742 7 1 2 12739 12741
0 12743 7 1 2 12737 12742
0 12744 5 1 1 12743
0 12745 7 1 2 91908 12744
0 12746 5 1 1 12745
0 12747 7 1 2 90441 12746
0 12748 5 1 1 12747
0 12749 7 1 2 73411 12748
0 12750 5 1 1 12749
0 12751 7 1 2 12730 12750
0 12752 5 1 1 12751
0 12753 7 1 2 80991 12752
0 12754 5 1 1 12753
0 12755 7 1 2 12724 12754
0 12756 5 1 1 12755
0 12757 7 1 2 72999 12756
0 12758 5 1 1 12757
0 12759 7 1 2 94506 94521
0 12760 5 1 1 12759
0 12761 7 1 2 12758 12760
0 12762 5 1 1 12761
0 12763 7 1 2 64648 12762
0 12764 5 1 1 12763
0 12765 7 2 2 88391 81500
0 12766 7 2 2 69771 94538
0 12767 5 1 1 94540
0 12768 7 1 2 8109 83554
0 12769 5 1 1 12768
0 12770 7 1 2 89173 12769
0 12771 5 2 1 12770
0 12772 7 1 2 94542 94432
0 12773 5 1 1 12772
0 12774 7 1 2 71325 12773
0 12775 5 1 1 12774
0 12776 7 1 2 12767 12775
0 12777 5 1 1 12776
0 12778 7 1 2 88070 12777
0 12779 5 1 1 12778
0 12780 7 1 2 88724 88976
0 12781 5 1 1 12780
0 12782 7 1 2 12779 12781
0 12783 5 1 1 12782
0 12784 7 1 2 85246 12783
0 12785 5 1 1 12784
0 12786 7 1 2 86997 5828
0 12787 5 1 1 12786
0 12788 7 1 2 90908 12787
0 12789 5 1 1 12788
0 12790 7 1 2 12785 12789
0 12791 5 1 1 12790
0 12792 7 1 2 88547 12791
0 12793 5 1 1 12792
0 12794 7 5 2 69772 68614
0 12795 5 5 1 94544
0 12796 7 1 2 94549 90909
0 12797 5 1 1 12796
0 12798 7 2 2 68337 75481
0 12799 7 1 2 94554 91909
0 12800 5 1 1 12799
0 12801 7 1 2 12797 12800
0 12802 5 1 1 12801
0 12803 7 1 2 71789 12802
0 12804 5 1 1 12803
0 12805 7 1 2 77120 92102
0 12806 5 1 1 12805
0 12807 7 2 2 82901 87391
0 12808 5 1 1 94556
0 12809 7 1 2 85885 94557
0 12810 5 1 1 12809
0 12811 7 1 2 12806 12810
0 12812 5 1 1 12811
0 12813 7 1 2 91940 12812
0 12814 5 1 1 12813
0 12815 7 1 2 12804 12814
0 12816 5 1 1 12815
0 12817 7 1 2 70377 12816
0 12818 5 1 1 12817
0 12819 7 1 2 80581 90418
0 12820 7 1 2 91963 12819
0 12821 5 2 1 12820
0 12822 7 9 2 63760 71326
0 12823 7 5 2 66959 94560
0 12824 5 2 1 94569
0 12825 7 1 2 94570 87181
0 12826 7 1 2 88071 12825
0 12827 5 1 1 12826
0 12828 7 1 2 94558 12827
0 12829 5 1 1 12828
0 12830 7 1 2 75043 12829
0 12831 5 1 1 12830
0 12832 7 4 2 80680 76379
0 12833 7 1 2 94576 90329
0 12834 5 1 1 12833
0 12835 7 3 2 66960 86396
0 12836 7 1 2 75634 94580
0 12837 7 1 2 94059 12836
0 12838 5 1 1 12837
0 12839 7 1 2 12834 12838
0 12840 5 1 1 12839
0 12841 7 1 2 76298 12840
0 12842 5 1 1 12841
0 12843 7 14 2 70664 71919
0 12844 7 5 2 94583 90512
0 12845 7 2 2 91265 94597
0 12846 7 3 2 85886 79575
0 12847 5 1 1 94604
0 12848 7 2 2 82346 75099
0 12849 5 1 1 94607
0 12850 7 1 2 94605 94608
0 12851 7 1 2 94602 12850
0 12852 5 1 1 12851
0 12853 7 1 2 12852 92475
0 12854 7 1 2 12842 12853
0 12855 7 1 2 12831 12854
0 12856 7 1 2 12818 12855
0 12857 5 1 1 12856
0 12858 7 1 2 88176 12857
0 12859 5 1 1 12858
0 12860 7 1 2 12793 12859
0 12861 5 1 1 12860
0 12862 7 1 2 67979 12861
0 12863 5 1 1 12862
0 12864 7 1 2 85247 75122
0 12865 5 1 1 12864
0 12866 7 5 2 89149 91803
0 12867 5 1 1 94609
0 12868 7 2 2 68615 94610
0 12869 5 1 1 94614
0 12870 7 1 2 70132 94615
0 12871 5 1 1 12870
0 12872 7 1 2 12865 12871
0 12873 5 1 1 12872
0 12874 7 1 2 68338 12873
0 12875 5 1 1 12874
0 12876 7 4 2 80582 90730
0 12877 5 2 1 94616
0 12878 7 1 2 83541 94617
0 12879 5 1 1 12878
0 12880 7 1 2 12875 12879
0 12881 5 1 1 12880
0 12882 7 1 2 88177 12881
0 12883 5 1 1 12882
0 12884 7 1 2 79820 81601
0 12885 5 1 1 12884
0 12886 7 1 2 85248 89718
0 12887 7 1 2 12885 12886
0 12888 5 1 1 12887
0 12889 7 1 2 12883 12888
0 12890 5 1 1 12889
0 12891 7 1 2 71602 12890
0 12892 5 1 1 12891
0 12893 7 1 2 80290 91856
0 12894 5 1 1 12893
0 12895 7 1 2 12892 12894
0 12896 5 1 1 12895
0 12897 7 1 2 88072 12896
0 12898 5 1 1 12897
0 12899 7 4 2 68807 84642
0 12900 7 1 2 79350 94622
0 12901 7 1 2 94371 12900
0 12902 5 1 1 12901
0 12903 7 1 2 12898 12902
0 12904 5 1 1 12903
0 12905 7 1 2 83243 12904
0 12906 5 1 1 12905
0 12907 7 3 2 66854 75966
0 12908 7 4 2 94626 90787
0 12909 5 1 1 94629
0 12910 7 1 2 90532 92499
0 12911 7 1 2 94410 12910
0 12912 5 1 1 12911
0 12913 7 1 2 12909 12912
0 12914 5 1 1 12913
0 12915 7 1 2 85249 12914
0 12916 5 1 1 12915
0 12917 7 1 2 90910 4137
0 12918 5 1 1 12917
0 12919 7 2 2 73000 75738
0 12920 7 1 2 75358 83931
0 12921 7 1 2 94633 12920
0 12922 7 1 2 90383 12921
0 12923 5 1 1 12922
0 12924 7 1 2 12918 12923
0 12925 5 1 1 12924
0 12926 7 1 2 68339 12925
0 12927 5 1 1 12926
0 12928 7 1 2 12916 12927
0 12929 5 1 1 12928
0 12930 7 1 2 88548 12929
0 12931 5 1 1 12930
0 12932 7 3 2 82759 90745
0 12933 7 1 2 94062 91304
0 12934 7 1 2 94635 12933
0 12935 5 1 1 12934
0 12936 7 1 2 12931 12935
0 12937 5 1 1 12936
0 12938 7 1 2 81840 12937
0 12939 5 1 1 12938
0 12940 7 1 2 89103 89829
0 12941 5 1 1 12940
0 12942 7 1 2 66679 78688
0 12943 7 1 2 12941 12942
0 12944 5 1 1 12943
0 12945 7 1 2 78601 77509
0 12946 5 1 1 12945
0 12947 7 1 2 12944 12946
0 12948 5 1 1 12947
0 12949 7 1 2 65347 12948
0 12950 5 1 1 12949
0 12951 7 1 2 88434 92689
0 12952 5 1 1 12951
0 12953 7 1 2 12950 12952
0 12954 5 1 1 12953
0 12955 7 2 2 88052 91672
0 12956 7 1 2 12954 94638
0 12957 5 1 1 12956
0 12958 7 1 2 68616 91374
0 12959 5 1 1 12958
0 12960 7 1 2 12957 12959
0 12961 5 1 1 12960
0 12962 7 1 2 94571 12961
0 12963 5 1 1 12962
0 12964 7 1 2 65952 12963
0 12965 7 1 2 12939 12964
0 12966 7 1 2 12906 12965
0 12967 7 1 2 12863 12966
0 12968 5 1 1 12967
0 12969 7 3 2 63761 66493
0 12970 7 1 2 94640 94504
0 12971 5 1 1 12970
0 12972 7 1 2 94152 88178
0 12973 5 1 1 12972
0 12974 7 1 2 83697 89737
0 12975 5 1 1 12974
0 12976 7 1 2 83430 93983
0 12977 5 1 1 12976
0 12978 7 1 2 90171 12977
0 12979 5 1 1 12978
0 12980 7 1 2 12975 12979
0 12981 7 1 2 12973 12980
0 12982 5 1 1 12981
0 12983 7 1 2 85250 12982
0 12984 5 1 1 12983
0 12985 7 1 2 82103 89309
0 12986 5 1 1 12985
0 12987 7 2 2 72025 76677
0 12988 7 5 2 63883 66494
0 12989 7 1 2 68808 94645
0 12990 7 2 2 94643 12989
0 12991 7 1 2 67078 94650
0 12992 5 1 1 12991
0 12993 7 1 2 12986 12992
0 12994 5 1 1 12993
0 12995 7 1 2 65030 84821
0 12996 7 1 2 12994 12995
0 12997 5 1 1 12996
0 12998 7 1 2 12984 12997
0 12999 5 1 1 12998
0 13000 7 1 2 73001 12999
0 13001 5 1 1 13000
0 13002 7 1 2 12971 13001
0 13003 5 1 1 13002
0 13004 7 1 2 64649 13003
0 13005 5 1 1 13004
0 13006 7 2 2 94561 86475
0 13007 7 1 2 90196 94652
0 13008 5 1 1 13007
0 13009 7 1 2 13005 13008
0 13010 5 1 1 13009
0 13011 7 1 2 88073 13010
0 13012 5 1 1 13011
0 13013 7 1 2 94113 94452
0 13014 5 1 1 13013
0 13015 7 1 2 71023 13014
0 13016 7 1 2 13012 13015
0 13017 5 1 1 13016
0 13018 7 1 2 64321 13017
0 13019 7 1 2 12968 13018
0 13020 5 1 1 13019
0 13021 7 8 2 66680 79981
0 13022 5 1 1 94654
0 13023 7 1 2 94655 91595
0 13024 7 1 2 92216 13023
0 13025 7 1 2 90197 13024
0 13026 5 1 1 13025
0 13027 7 1 2 13020 13026
0 13028 7 1 2 12764 13027
0 13029 7 1 2 12674 13028
0 13030 5 1 1 13029
0 13031 7 1 2 72599 13030
0 13032 5 1 1 13031
0 13033 7 1 2 79783 88328
0 13034 7 1 2 91966 13033
0 13035 5 1 1 13034
0 13036 7 1 2 64322 94457
0 13037 5 1 1 13036
0 13038 7 1 2 12717 13037
0 13039 5 1 1 13038
0 13040 7 1 2 92109 84127
0 13041 7 1 2 13039 13040
0 13042 5 1 1 13041
0 13043 7 1 2 13035 13042
0 13044 5 1 1 13043
0 13045 7 1 2 73002 13044
0 13046 5 1 1 13045
0 13047 7 1 2 64650 93998
0 13048 7 1 2 91841 13047
0 13049 7 1 2 74160 13048
0 13050 7 1 2 93408 13049
0 13051 5 1 1 13050
0 13052 7 1 2 13046 13051
0 13053 5 1 1 13052
0 13054 7 1 2 72600 13053
0 13055 5 1 1 13054
0 13056 7 1 2 77657 87921
0 13057 7 1 2 91601 13056
0 13058 7 3 2 68809 84016
0 13059 7 2 2 69060 84455
0 13060 7 5 2 70378 70665
0 13061 5 1 1 94667
0 13062 7 3 2 94668 86087
0 13063 7 1 2 94665 94672
0 13064 7 1 2 94662 13063
0 13065 7 1 2 13057 13064
0 13066 5 1 1 13065
0 13067 7 1 2 13055 13066
0 13068 5 1 1 13067
0 13069 7 1 2 72134 84750
0 13070 5 1 1 13069
0 13071 7 1 2 89293 13070
0 13072 7 1 2 13068 13071
0 13073 5 1 1 13072
0 13074 7 1 2 65031 87150
0 13075 5 3 1 13074
0 13076 7 1 2 73003 88471
0 13077 5 1 1 13076
0 13078 7 1 2 94675 13077
0 13079 5 1 1 13078
0 13080 7 1 2 88179 13079
0 13081 5 1 1 13080
0 13082 7 2 2 71790 89670
0 13083 5 1 1 94678
0 13084 7 2 2 77826 94679
0 13085 5 1 1 94680
0 13086 7 1 2 66495 94681
0 13087 5 1 1 13086
0 13088 7 1 2 76566 89342
0 13089 5 1 1 13088
0 13090 7 1 2 13087 13089
0 13091 5 1 1 13090
0 13092 7 1 2 77552 13091
0 13093 5 1 1 13092
0 13094 7 1 2 13081 13093
0 13095 5 1 1 13094
0 13096 7 1 2 70379 13095
0 13097 5 1 1 13096
0 13098 7 1 2 76463 86106
0 13099 5 1 1 13098
0 13100 7 1 2 73004 13099
0 13101 5 1 1 13100
0 13102 7 1 2 94676 13101
0 13103 5 1 1 13102
0 13104 7 1 2 13103 90538
0 13105 5 1 1 13104
0 13106 7 1 2 13097 13105
0 13107 5 1 1 13106
0 13108 7 1 2 92508 79784
0 13109 7 1 2 92370 13108
0 13110 7 1 2 13107 13109
0 13111 5 1 1 13110
0 13112 7 1 2 13073 13111
0 13113 7 1 2 13032 13112
0 13114 7 1 2 12043 13113
0 13115 5 1 1 13114
0 13116 7 1 2 64051 13115
0 13117 5 1 1 13116
0 13118 7 6 2 72601 77319
0 13119 7 6 2 72026 93696
0 13120 7 3 2 81705 86340
0 13121 5 2 1 94694
0 13122 7 4 2 94646 89347
0 13123 5 1 1 94699
0 13124 7 1 2 94695 94700
0 13125 5 1 1 13124
0 13126 7 1 2 88549 94302
0 13127 5 1 1 13126
0 13128 7 1 2 65348 88791
0 13129 5 1 1 13128
0 13130 7 2 2 80533 13129
0 13131 5 1 1 94703
0 13132 7 1 2 78689 94704
0 13133 5 1 1 13132
0 13134 7 1 2 88180 13133
0 13135 5 1 1 13134
0 13136 7 1 2 13127 13135
0 13137 5 1 1 13136
0 13138 7 1 2 65032 13137
0 13139 5 1 1 13138
0 13140 7 1 2 80399 88181
0 13141 5 2 1 13140
0 13142 7 1 2 93992 94705
0 13143 5 1 1 13142
0 13144 7 1 2 73412 13143
0 13145 5 1 1 13144
0 13146 7 1 2 89294 13083
0 13147 7 1 2 93926 13146
0 13148 5 1 1 13147
0 13149 7 1 2 13145 13148
0 13150 5 1 1 13149
0 13151 7 1 2 66496 13150
0 13152 5 1 1 13151
0 13153 7 1 2 13152 6811
0 13154 7 1 2 13139 13153
0 13155 5 1 1 13154
0 13156 7 1 2 73005 13155
0 13157 5 1 1 13156
0 13158 7 1 2 13125 13157
0 13159 5 1 1 13158
0 13160 7 1 2 94688 13159
0 13161 5 1 1 13160
0 13162 7 1 2 80865 87178
0 13163 5 1 1 13162
0 13164 7 1 2 66681 13163
0 13165 5 1 1 13164
0 13166 7 1 2 86934 13165
0 13167 5 1 1 13166
0 13168 7 1 2 65349 13167
0 13169 5 1 1 13168
0 13170 7 1 2 86929 13169
0 13171 5 1 1 13170
0 13172 7 1 2 73006 13171
0 13173 5 1 1 13172
0 13174 7 1 2 83368 94481
0 13175 5 1 1 13174
0 13176 7 1 2 78933 10847
0 13177 7 1 2 13175 13176
0 13178 5 1 1 13177
0 13179 7 1 2 85675 13178
0 13180 5 1 1 13179
0 13181 7 1 2 81841 79229
0 13182 5 2 1 13181
0 13183 7 1 2 74752 94707
0 13184 5 1 1 13183
0 13185 7 1 2 88364 80926
0 13186 7 1 2 13184 13185
0 13187 5 1 1 13186
0 13188 7 1 2 13180 13187
0 13189 7 1 2 13173 13188
0 13190 5 1 1 13189
0 13191 7 1 2 88182 13190
0 13192 5 1 1 13191
0 13193 7 2 2 81590 87451
0 13194 5 1 1 94709
0 13195 7 2 2 80091 94710
0 13196 5 2 1 94711
0 13197 7 1 2 94713 9991
0 13198 5 1 1 13197
0 13199 7 1 2 73701 13198
0 13200 5 1 1 13199
0 13201 7 1 2 69109 94287
0 13202 5 1 1 13201
0 13203 7 1 2 13200 13202
0 13204 5 1 1 13203
0 13205 7 1 2 73007 13204
0 13206 5 1 1 13205
0 13207 7 5 2 69110 66682
0 13208 7 3 2 75100 94715
0 13209 5 1 1 94720
0 13210 7 6 2 67980 81842
0 13211 5 4 1 94723
0 13212 7 1 2 93794 94724
0 13213 5 1 1 13212
0 13214 7 1 2 13209 13213
0 13215 5 1 1 13214
0 13216 7 1 2 78635 13215
0 13217 5 1 1 13216
0 13218 7 1 2 13206 13217
0 13219 5 1 1 13218
0 13220 7 1 2 88550 13219
0 13221 5 1 1 13220
0 13222 7 5 2 65350 67079
0 13223 7 1 2 93842 94733
0 13224 5 2 1 13223
0 13225 7 1 2 77827 94495
0 13226 5 2 1 13225
0 13227 7 1 2 94738 94740
0 13228 5 2 1 13227
0 13229 7 1 2 75101 94739
0 13230 5 1 1 13229
0 13231 7 1 2 84540 13230
0 13232 7 1 2 94742 13231
0 13233 5 1 1 13232
0 13234 7 1 2 13221 13233
0 13235 7 1 2 13192 13234
0 13236 5 1 1 13235
0 13237 7 1 2 85251 13236
0 13238 5 1 1 13237
0 13239 7 1 2 13161 13238
0 13240 5 1 1 13239
0 13241 7 1 2 88977 13240
0 13242 5 1 1 13241
0 13243 7 3 2 73413 87508
0 13244 7 2 2 75102 94744
0 13245 5 1 1 94747
0 13246 7 6 2 80521 93928
0 13247 5 7 1 94749
0 13248 7 2 2 71603 94044
0 13249 5 1 1 94762
0 13250 7 4 2 94755 13249
0 13251 5 1 1 94764
0 13252 7 1 2 65033 94765
0 13253 5 1 1 13252
0 13254 7 1 2 13245 13253
0 13255 5 3 1 13254
0 13256 7 1 2 94768 88183
0 13257 5 1 1 13256
0 13258 7 2 2 78636 88551
0 13259 7 1 2 94696 94771
0 13260 5 1 1 13259
0 13261 7 1 2 13257 13260
0 13262 5 1 1 13261
0 13263 7 12 2 69111 70621
0 13264 7 3 2 63762 94773
0 13265 7 2 2 94785 94079
0 13266 7 1 2 94634 94788
0 13267 7 1 2 13262 13266
0 13268 5 1 1 13267
0 13269 7 1 2 13242 13268
0 13270 5 1 1 13269
0 13271 7 1 2 76199 13270
0 13272 5 1 1 13271
0 13273 7 2 2 93725 84593
0 13274 5 1 1 94790
0 13275 7 2 2 79326 84643
0 13276 5 1 1 94792
0 13277 7 1 2 13274 13276
0 13278 5 1 1 13277
0 13279 7 1 2 85252 13278
0 13280 5 1 1 13279
0 13281 7 3 2 68810 93101
0 13282 7 1 2 94794 94515
0 13283 5 1 1 13282
0 13284 7 1 2 13280 13283
0 13285 5 1 1 13284
0 13286 7 1 2 65351 13285
0 13287 5 1 1 13286
0 13288 7 9 2 66683 67080
0 13289 7 4 2 82769 94797
0 13290 7 1 2 79803 94806
0 13291 5 1 1 13290
0 13292 7 1 2 13287 13291
0 13293 5 1 1 13292
0 13294 7 3 2 66855 73702
0 13295 7 7 2 63971 73008
0 13296 7 1 2 94810 94813
0 13297 7 1 2 93341 13296
0 13298 7 1 2 92229 13297
0 13299 7 1 2 13293 13298
0 13300 5 1 1 13299
0 13301 7 1 2 13272 13300
0 13302 5 1 1 13301
0 13303 7 1 2 94682 13302
0 13304 5 1 1 13303
0 13305 7 1 2 13117 13304
0 13306 5 1 1 13305
0 13307 7 1 2 65746 13306
0 13308 5 1 1 13307
0 13309 7 3 2 76200 74165
0 13310 7 2 2 77024 86424
0 13311 7 2 2 87730 76883
0 13312 7 2 2 94823 94825
0 13313 7 1 2 94820 94827
0 13314 5 1 1 13313
0 13315 7 1 2 85 94714
0 13316 5 1 1 13315
0 13317 7 1 2 13316 75209
0 13318 5 1 1 13317
0 13319 7 5 2 70771 67081
0 13320 7 1 2 74297 94829
0 13321 7 1 2 87489 13320
0 13322 5 1 1 13321
0 13323 7 1 2 13318 13322
0 13324 5 1 1 13323
0 13325 7 1 2 73703 13324
0 13326 5 1 1 13325
0 13327 7 8 2 70772 66497
0 13328 7 2 2 77828 76839
0 13329 5 1 1 94842
0 13330 7 1 2 74274 13329
0 13331 5 2 1 13330
0 13332 7 2 2 73414 94844
0 13333 7 1 2 94834 94846
0 13334 5 1 1 13333
0 13335 7 3 2 74236 90635
0 13336 5 1 1 94848
0 13337 7 1 2 83527 94250
0 13338 7 1 2 94849 13337
0 13339 5 1 1 13338
0 13340 7 1 2 13334 13339
0 13341 7 1 2 13326 13340
0 13342 5 1 1 13341
0 13343 7 1 2 73009 13342
0 13344 5 1 1 13343
0 13345 7 3 2 72027 73704
0 13346 7 1 2 94851 94798
0 13347 7 2 2 76001 13346
0 13348 5 1 1 94854
0 13349 7 1 2 74166 94855
0 13350 5 1 1 13349
0 13351 7 1 2 86867 83119
0 13352 5 2 1 13351
0 13353 7 9 2 70773 66684
0 13354 7 3 2 73705 94858
0 13355 7 1 2 65352 94867
0 13356 5 1 1 13355
0 13357 7 1 2 94856 13356
0 13358 5 1 1 13357
0 13359 7 1 2 75210 13358
0 13360 5 1 1 13359
0 13361 7 1 2 13350 13360
0 13362 5 1 1 13361
0 13363 7 1 2 78637 13362
0 13364 5 1 1 13363
0 13365 7 1 2 13344 13364
0 13366 5 1 1 13365
0 13367 7 1 2 76201 13366
0 13368 5 1 1 13367
0 13369 7 2 2 89348 74298
0 13370 5 1 1 94870
0 13371 7 1 2 74275 13370
0 13372 5 2 1 13371
0 13373 7 1 2 78820 89618
0 13374 7 1 2 84346 13373
0 13375 7 1 2 94872 13374
0 13376 5 1 1 13375
0 13377 7 1 2 13368 13376
0 13378 5 1 1 13377
0 13379 7 1 2 78854 13378
0 13380 5 1 1 13379
0 13381 7 1 2 13314 13380
0 13382 5 1 1 13381
0 13383 7 1 2 94683 13382
0 13384 5 1 1 13383
0 13385 7 2 2 90026 87494
0 13386 5 1 1 94874
0 13387 7 1 2 79454 94875
0 13388 5 1 1 13387
0 13389 7 1 2 83528 76763
0 13390 5 1 1 13389
0 13391 7 1 2 75123 75211
0 13392 5 1 1 13391
0 13393 7 1 2 13390 13392
0 13394 5 1 1 13393
0 13395 7 1 2 71791 13394
0 13396 5 1 1 13395
0 13397 7 2 2 65034 79804
0 13398 5 1 1 94876
0 13399 7 1 2 81706 86958
0 13400 5 3 1 13399
0 13401 7 1 2 13398 94878
0 13402 5 1 1 13401
0 13403 7 1 2 76764 13402
0 13404 5 1 1 13403
0 13405 7 1 2 13396 13404
0 13406 5 1 1 13405
0 13407 7 1 2 73010 13406
0 13408 5 1 1 13407
0 13409 7 1 2 79312 91081
0 13410 5 1 1 13409
0 13411 7 1 2 806 13410
0 13412 5 1 1 13411
0 13413 7 1 2 81707 13412
0 13414 5 1 1 13413
0 13415 7 1 2 86415 75877
0 13416 7 1 2 89167 13415
0 13417 5 1 1 13416
0 13418 7 1 2 13414 13417
0 13419 5 1 1 13418
0 13420 7 1 2 65035 13419
0 13421 5 1 1 13420
0 13422 7 1 2 13408 13421
0 13423 5 1 1 13422
0 13424 7 1 2 66214 13423
0 13425 5 1 1 13424
0 13426 7 1 2 66215 86041
0 13427 5 1 1 13426
0 13428 7 1 2 83419 85764
0 13429 5 2 1 13428
0 13430 7 1 2 13427 94881
0 13431 5 1 1 13430
0 13432 7 1 2 75212 13431
0 13433 5 1 1 13432
0 13434 7 1 2 84973 89150
0 13435 7 1 2 84146 13434
0 13436 5 1 1 13435
0 13437 7 1 2 13433 13436
0 13438 5 1 1 13437
0 13439 7 1 2 74631 13438
0 13440 5 1 1 13439
0 13441 7 2 2 73011 94184
0 13442 5 2 1 94883
0 13443 7 1 2 78934 94885
0 13444 5 1 1 13443
0 13445 7 1 2 76840 90027
0 13446 7 1 2 13444 13445
0 13447 5 1 1 13446
0 13448 7 1 2 79564 78935
0 13449 5 1 1 13448
0 13450 7 3 2 75192 84594
0 13451 5 1 1 94887
0 13452 7 1 2 65353 94888
0 13453 7 1 2 13449 13452
0 13454 5 1 1 13453
0 13455 7 1 2 13447 13454
0 13456 7 1 2 13440 13455
0 13457 5 1 1 13456
0 13458 7 1 2 73415 13457
0 13459 5 1 1 13458
0 13460 7 2 2 72135 86416
0 13461 7 1 2 92057 94890
0 13462 7 1 2 89219 13461
0 13463 5 1 1 13462
0 13464 7 1 2 13459 13463
0 13465 7 1 2 13425 13464
0 13466 5 1 1 13465
0 13467 7 1 2 64651 13466
0 13468 5 1 1 13467
0 13469 7 1 2 66216 89220
0 13470 5 2 1 13469
0 13471 7 1 2 71327 77007
0 13472 5 4 1 13471
0 13473 7 3 2 75967 94894
0 13474 7 1 2 85734 94898
0 13475 5 1 1 13474
0 13476 7 1 2 94892 13475
0 13477 5 1 1 13476
0 13478 7 1 2 66498 13477
0 13479 5 1 1 13478
0 13480 7 6 2 71792 79065
0 13481 7 1 2 90189 94901
0 13482 5 1 1 13481
0 13483 7 1 2 13479 13482
0 13484 5 1 1 13483
0 13485 7 1 2 65036 13484
0 13486 5 1 1 13485
0 13487 7 2 2 70380 77043
0 13488 7 1 2 83420 77658
0 13489 7 1 2 94907 13488
0 13490 5 1 1 13489
0 13491 7 1 2 13486 13490
0 13492 5 1 1 13491
0 13493 7 1 2 75213 13492
0 13494 5 1 1 13493
0 13495 7 1 2 13468 13494
0 13496 5 1 1 13495
0 13497 7 1 2 79132 13496
0 13498 5 1 1 13497
0 13499 7 1 2 13388 13498
0 13500 5 1 1 13499
0 13501 7 1 2 69452 13500
0 13502 5 1 1 13501
0 13503 7 2 2 73706 79836
0 13504 7 4 2 78984 92492
0 13505 7 1 2 94909 94911
0 13506 5 1 1 13505
0 13507 7 1 2 75472 78855
0 13508 5 1 1 13507
0 13509 7 1 2 13506 13508
0 13510 5 1 1 13509
0 13511 7 1 2 13510 79333
0 13512 5 1 1 13511
0 13513 7 2 2 74632 82104
0 13514 7 2 2 94915 75214
0 13515 5 1 1 94917
0 13516 7 1 2 94912 94918
0 13517 5 1 1 13516
0 13518 7 1 2 13512 13517
0 13519 5 1 1 13518
0 13520 7 1 2 66217 13519
0 13521 5 1 1 13520
0 13522 7 1 2 76678 78560
0 13523 5 1 1 13522
0 13524 7 1 2 13515 13523
0 13525 5 1 1 13524
0 13526 7 3 2 71920 89080
0 13527 7 1 2 94134 94919
0 13528 7 1 2 13525 13527
0 13529 5 1 1 13528
0 13530 7 1 2 13521 13529
0 13531 5 1 1 13530
0 13532 7 1 2 73012 13531
0 13533 5 1 1 13532
0 13534 7 1 2 83901 79653
0 13535 5 1 1 13534
0 13536 7 2 2 76679 78346
0 13537 7 1 2 89081 86501
0 13538 7 1 2 94922 13537
0 13539 5 1 1 13538
0 13540 7 1 2 13535 13539
0 13541 5 1 1 13540
0 13542 7 1 2 76841 92519
0 13543 7 1 2 13541 13542
0 13544 5 1 1 13543
0 13545 7 1 2 13533 13544
0 13546 5 1 1 13545
0 13547 7 1 2 84822 13546
0 13548 5 1 1 13547
0 13549 7 2 2 68340 88334
0 13550 5 5 1 94924
0 13551 7 1 2 80799 94926
0 13552 5 5 1 13551
0 13553 7 2 2 70381 94931
0 13554 5 1 1 94936
0 13555 7 3 2 77084 74900
0 13556 5 1 1 94938
0 13557 7 1 2 13554 13556
0 13558 5 1 1 13557
0 13559 7 1 2 71793 13558
0 13560 5 1 1 13559
0 13561 7 1 2 65354 75027
0 13562 5 1 1 13561
0 13563 7 1 2 13560 13562
0 13564 5 1 1 13563
0 13565 7 1 2 75908 79399
0 13566 7 1 2 13564 13565
0 13567 5 1 1 13566
0 13568 7 1 2 13548 13567
0 13569 7 1 2 13502 13568
0 13570 5 1 1 13569
0 13571 7 1 2 65953 13570
0 13572 5 1 1 13571
0 13573 7 1 2 77418 87179
0 13574 5 1 1 13573
0 13575 7 1 2 94257 13574
0 13576 5 1 1 13575
0 13577 7 1 2 73013 13576
0 13578 5 1 1 13577
0 13579 7 1 2 12325 94857
0 13580 5 1 1 13579
0 13581 7 1 2 78638 13580
0 13582 5 1 1 13581
0 13583 7 1 2 13578 13582
0 13584 5 1 1 13583
0 13585 7 1 2 78856 13584
0 13586 5 1 1 13585
0 13587 7 1 2 79166 90190
0 13588 5 1 1 13587
0 13589 7 1 2 82794 13588
0 13590 5 1 1 13589
0 13591 7 1 2 81708 13590
0 13592 5 1 1 13591
0 13593 7 1 2 64323 73956
0 13594 7 1 2 89168 13593
0 13595 5 1 1 13594
0 13596 7 1 2 13592 13595
0 13597 5 1 1 13596
0 13598 7 1 2 65037 13597
0 13599 5 1 1 13598
0 13600 7 1 2 82678 93905
0 13601 5 1 1 13600
0 13602 7 1 2 13599 13601
0 13603 5 1 1 13602
0 13604 7 1 2 78985 91634
0 13605 7 1 2 13603 13604
0 13606 5 1 1 13605
0 13607 7 1 2 13586 13606
0 13608 5 1 1 13607
0 13609 7 1 2 64652 13608
0 13610 5 1 1 13609
0 13611 7 1 2 75270 86042
0 13612 5 1 1 13611
0 13613 7 2 2 70382 84755
0 13614 5 3 1 94941
0 13615 7 2 2 85596 94943
0 13616 5 2 1 94946
0 13617 7 3 2 73416 94948
0 13618 7 2 2 74633 94950
0 13619 5 1 1 94953
0 13620 7 1 2 13612 13619
0 13621 5 1 1 13620
0 13622 7 1 2 71024 79013
0 13623 7 1 2 13621 13622
0 13624 5 1 1 13623
0 13625 7 1 2 75271 78857
0 13626 7 1 2 94329 13625
0 13627 5 1 1 13626
0 13628 7 1 2 13624 13627
0 13629 5 1 1 13628
0 13630 7 1 2 73014 13629
0 13631 5 1 1 13630
0 13632 7 2 2 79100 76884
0 13633 7 1 2 89596 94955
0 13634 7 1 2 87004 13633
0 13635 5 1 1 13634
0 13636 7 1 2 13631 13635
0 13637 7 1 2 13610 13636
0 13638 5 1 1 13637
0 13639 7 1 2 75215 13638
0 13640 5 1 1 13639
0 13641 7 1 2 86244 79455
0 13642 5 1 1 13641
0 13643 7 1 2 86979 79014
0 13644 5 1 1 13643
0 13645 7 1 2 82632 79654
0 13646 5 2 1 13645
0 13647 7 2 2 75602 78858
0 13648 5 1 1 94959
0 13649 7 1 2 94957 13648
0 13650 7 1 2 13644 13649
0 13651 5 1 1 13650
0 13652 7 1 2 66499 82738
0 13653 7 1 2 13651 13652
0 13654 5 1 1 13653
0 13655 7 1 2 13642 13654
0 13656 5 1 1 13655
0 13657 7 1 2 65038 13656
0 13658 5 1 1 13657
0 13659 7 1 2 87470 94960
0 13660 5 1 1 13659
0 13661 7 1 2 13658 13660
0 13662 5 1 1 13661
0 13663 7 1 2 73707 13662
0 13664 5 1 1 13663
0 13665 7 3 2 69453 86263
0 13666 5 3 1 94961
0 13667 7 2 2 73015 94964
0 13668 7 1 2 94967 79456
0 13669 5 1 1 13668
0 13670 7 1 2 13664 13669
0 13671 5 1 1 13670
0 13672 7 1 2 71025 13671
0 13673 5 1 1 13672
0 13674 7 5 2 93642 77896
0 13675 7 1 2 64324 89751
0 13676 7 1 2 94969 13675
0 13677 5 1 1 13676
0 13678 7 1 2 13673 13677
0 13679 5 1 1 13678
0 13680 7 1 2 76765 13679
0 13681 5 1 1 13680
0 13682 7 1 2 13640 13681
0 13683 5 1 1 13682
0 13684 7 1 2 66218 13683
0 13685 5 1 1 13684
0 13686 7 4 2 87404 87955
0 13687 7 2 2 71921 79327
0 13688 7 1 2 91864 94978
0 13689 7 1 2 94974 13688
0 13690 5 1 1 13689
0 13691 7 1 2 66685 79655
0 13692 7 1 2 94873 13691
0 13693 5 1 1 13692
0 13694 7 1 2 13690 13693
0 13695 5 1 1 13694
0 13696 7 1 2 65355 13695
0 13697 5 1 1 13696
0 13698 7 4 2 64325 87405
0 13699 7 2 2 70383 83392
0 13700 5 2 1 94984
0 13701 7 2 2 76798 76842
0 13702 7 1 2 94985 94988
0 13703 7 1 2 94980 13702
0 13704 5 1 1 13703
0 13705 7 1 2 13697 13704
0 13706 5 1 1 13705
0 13707 7 1 2 73708 13706
0 13708 5 1 1 13707
0 13709 7 4 2 87731 87956
0 13710 7 1 2 94519 94990
0 13711 5 1 1 13710
0 13712 7 1 2 13708 13711
0 13713 5 1 1 13712
0 13714 7 1 2 75272 13713
0 13715 5 1 1 13714
0 13716 7 1 2 89896 94991
0 13717 7 1 2 94954 13716
0 13718 5 1 1 13717
0 13719 7 1 2 13715 13718
0 13720 5 1 1 13719
0 13721 7 1 2 73016 13720
0 13722 5 1 1 13721
0 13723 7 2 2 66500 86397
0 13724 7 1 2 94994 94104
0 13725 7 6 2 65039 76885
0 13726 7 2 2 68811 91149
0 13727 7 1 2 94996 95002
0 13728 7 1 2 13724 13727
0 13729 5 1 1 13728
0 13730 7 1 2 13722 13729
0 13731 5 1 1 13730
0 13732 7 1 2 71026 13731
0 13733 5 1 1 13732
0 13734 7 1 2 84569 93667
0 13735 7 1 2 86575 13734
0 13736 7 2 2 73017 90146
0 13737 7 2 2 65356 89863
0 13738 7 1 2 95004 95006
0 13739 7 1 2 13735 13738
0 13740 5 1 1 13739
0 13741 7 1 2 13733 13740
0 13742 5 1 1 13741
0 13743 7 1 2 64653 13742
0 13744 5 1 1 13743
0 13745 7 1 2 78799 78375
0 13746 7 1 2 94828 13745
0 13747 5 1 1 13746
0 13748 7 1 2 13744 13747
0 13749 7 1 2 13685 13748
0 13750 7 1 2 13572 13749
0 13751 5 1 1 13750
0 13752 7 1 2 72602 13751
0 13753 5 1 1 13752
0 13754 7 1 2 86833 89958
0 13755 5 1 1 13754
0 13756 7 2 2 78639 87010
0 13757 5 3 1 95008
0 13758 7 1 2 73709 87536
0 13759 5 1 1 13758
0 13760 7 2 2 95010 13759
0 13761 5 1 1 95013
0 13762 7 1 2 93331 94763
0 13763 5 1 1 13762
0 13764 7 2 2 81843 85588
0 13765 5 1 1 95015
0 13766 7 1 2 13763 13765
0 13767 5 1 1 13766
0 13768 7 1 2 70133 13767
0 13769 5 1 1 13768
0 13770 7 1 2 71604 95016
0 13771 5 1 1 13770
0 13772 7 1 2 76567 13771
0 13773 7 1 2 13769 13772
0 13774 5 1 1 13773
0 13775 7 1 2 76299 13774
0 13776 7 1 2 95014 13775
0 13777 5 1 1 13776
0 13778 7 1 2 67589 13777
0 13779 5 1 1 13778
0 13780 7 1 2 13755 13779
0 13781 5 1 1 13780
0 13782 7 1 2 78859 13781
0 13783 5 1 1 13782
0 13784 7 1 2 81962 92645
0 13785 5 2 1 13784
0 13786 7 2 2 73018 78147
0 13787 5 2 1 95019
0 13788 7 1 2 79862 95020
0 13789 5 1 1 13788
0 13790 7 1 2 95017 13789
0 13791 5 1 1 13790
0 13792 7 1 2 86990 13791
0 13793 5 1 1 13792
0 13794 7 4 2 65357 84736
0 13795 5 1 1 95023
0 13796 7 2 2 71605 95024
0 13797 5 1 1 95027
0 13798 7 1 2 70134 95028
0 13799 5 1 1 13798
0 13800 7 1 2 87065 13799
0 13801 5 1 1 13800
0 13802 7 1 2 84999 13801
0 13803 5 1 1 13802
0 13804 7 4 2 73019 82316
0 13805 5 2 1 95029
0 13806 7 1 2 95030 86284
0 13807 5 1 1 13806
0 13808 7 1 2 84788 86465
0 13809 5 1 1 13808
0 13810 7 1 2 13807 13809
0 13811 5 1 1 13810
0 13812 7 1 2 82132 13811
0 13813 5 1 1 13812
0 13814 7 1 2 13803 13813
0 13815 5 1 1 13814
0 13816 7 1 2 68341 13815
0 13817 5 1 1 13816
0 13818 7 1 2 85000 83518
0 13819 5 1 1 13818
0 13820 7 1 2 73020 94192
0 13821 5 1 1 13820
0 13822 7 4 2 67981 86264
0 13823 5 2 1 95035
0 13824 7 1 2 93930 88840
0 13825 5 1 1 13824
0 13826 7 1 2 95036 13825
0 13827 5 1 1 13826
0 13828 7 1 2 82133 13827
0 13829 7 1 2 13821 13828
0 13830 5 1 1 13829
0 13831 7 1 2 13819 13830
0 13832 7 1 2 13817 13831
0 13833 5 1 1 13832
0 13834 7 1 2 66219 13833
0 13835 5 1 1 13834
0 13836 7 1 2 13793 13835
0 13837 5 1 1 13836
0 13838 7 1 2 79133 13837
0 13839 5 1 1 13838
0 13840 7 1 2 13783 13839
0 13841 5 1 1 13840
0 13842 7 1 2 76766 13841
0 13843 5 1 1 13842
0 13844 7 2 2 73710 89042
0 13845 5 1 1 95041
0 13846 7 1 2 80176 13845
0 13847 5 1 1 13846
0 13848 7 1 2 67590 13847
0 13849 5 1 1 13848
0 13850 7 1 2 89438 89950
0 13851 5 1 1 13850
0 13852 7 7 2 74826 87243
0 13853 7 3 2 73711 85676
0 13854 5 2 1 95050
0 13855 7 1 2 95043 95053
0 13856 5 1 1 13855
0 13857 7 1 2 67591 13856
0 13858 5 1 1 13857
0 13859 7 1 2 13858 86690
0 13860 5 1 1 13859
0 13861 7 1 2 80158 13860
0 13862 5 1 1 13861
0 13863 7 1 2 13851 13862
0 13864 7 1 2 13849 13863
0 13865 5 1 1 13864
0 13866 7 1 2 78860 13865
0 13867 5 1 1 13866
0 13868 7 1 2 76070 94217
0 13869 5 1 1 13868
0 13870 7 1 2 94893 13869
0 13871 5 1 1 13870
0 13872 7 1 2 65040 13871
0 13873 5 1 1 13872
0 13874 7 2 2 79504 94482
0 13875 5 1 1 95055
0 13876 7 2 2 81280 84252
0 13877 5 3 1 95057
0 13878 7 1 2 95059 86043
0 13879 5 1 1 13878
0 13880 7 1 2 13875 13879
0 13881 5 1 1 13880
0 13882 7 1 2 64654 13881
0 13883 5 1 1 13882
0 13884 7 1 2 87074 93984
0 13885 5 1 1 13884
0 13886 7 1 2 75909 13885
0 13887 5 1 1 13886
0 13888 7 1 2 67592 13887
0 13889 7 1 2 13883 13888
0 13890 7 1 2 13873 13889
0 13891 5 1 1 13890
0 13892 7 2 2 74634 74944
0 13893 7 1 2 86044 95062
0 13894 5 1 1 13893
0 13895 7 8 2 66686 79022
0 13896 5 1 1 95064
0 13897 7 1 2 95065 93301
0 13898 5 1 1 13897
0 13899 7 1 2 72603 13898
0 13900 7 1 2 13894 13899
0 13901 5 1 1 13900
0 13902 7 1 2 73417 13901
0 13903 7 1 2 13891 13902
0 13904 5 1 1 13903
0 13905 7 1 2 76643 87019
0 13906 5 1 1 13905
0 13907 7 1 2 88865 13906
0 13908 5 1 1 13907
0 13909 7 2 2 75124 83470
0 13910 5 1 1 95072
0 13911 7 1 2 64655 95073
0 13912 5 1 1 13911
0 13913 7 1 2 13908 13912
0 13914 5 1 1 13913
0 13915 7 1 2 67593 13914
0 13916 5 1 1 13915
0 13917 7 1 2 75137 93161
0 13918 5 1 1 13917
0 13919 7 1 2 13916 13918
0 13920 5 1 1 13919
0 13921 7 1 2 66220 13920
0 13922 5 1 1 13921
0 13923 7 1 2 80970 92753
0 13924 5 1 1 13923
0 13925 7 1 2 87681 13924
0 13926 5 1 1 13925
0 13927 7 1 2 86045 13926
0 13928 5 1 1 13927
0 13929 7 1 2 91460 86712
0 13930 5 1 1 13929
0 13931 7 1 2 88866 13930
0 13932 5 1 1 13931
0 13933 7 1 2 13928 13932
0 13934 7 1 2 13922 13933
0 13935 7 1 2 13904 13934
0 13936 5 1 1 13935
0 13937 7 1 2 79134 13936
0 13938 5 1 1 13937
0 13939 7 1 2 13867 13938
0 13940 5 1 1 13939
0 13941 7 1 2 75216 13940
0 13942 5 1 1 13941
0 13943 7 1 2 13843 13942
0 13944 5 1 1 13943
0 13945 7 1 2 64326 13944
0 13946 5 1 1 13945
0 13947 7 1 2 77014 94135
0 13948 7 1 2 94465 13947
0 13949 7 2 2 83844 87791
0 13950 5 1 1 95074
0 13951 7 1 2 86425 95075
0 13952 7 1 2 13948 13951
0 13953 5 1 1 13952
0 13954 7 1 2 13946 13953
0 13955 5 1 1 13954
0 13956 7 1 2 65954 13955
0 13957 5 1 1 13956
0 13958 7 2 2 70622 71027
0 13959 7 1 2 74919 87612
0 13960 7 1 2 95076 13959
0 13961 7 2 2 87732 84456
0 13962 7 1 2 92254 94132
0 13963 7 1 2 95078 13962
0 13964 7 1 2 13960 13963
0 13965 5 1 1 13964
0 13966 7 1 2 13957 13965
0 13967 7 1 2 13753 13966
0 13968 5 1 1 13967
0 13969 7 1 2 65747 13968
0 13970 5 1 1 13969
0 13971 7 1 2 13384 13970
0 13972 5 1 1 13971
0 13973 7 1 2 64052 13972
0 13974 5 1 1 13973
0 13975 7 1 2 67982 78833
0 13976 5 1 1 13975
0 13977 7 1 2 82060 13976
0 13978 5 1 1 13977
0 13979 7 1 2 85677 13978
0 13980 5 1 1 13979
0 13981 7 1 2 86667 80967
0 13982 5 1 1 13981
0 13983 7 2 2 73418 13982
0 13984 5 1 1 95080
0 13985 7 6 2 64656 80583
0 13986 5 3 1 95082
0 13987 7 1 2 75359 95083
0 13988 5 2 1 13987
0 13989 7 1 2 81709 76644
0 13990 5 1 1 13989
0 13991 7 1 2 95091 13990
0 13992 5 1 1 13991
0 13993 7 1 2 68617 13992
0 13994 5 1 1 13993
0 13995 7 1 2 82306 92401
0 13996 5 1 1 13995
0 13997 7 1 2 13994 13996
0 13998 5 1 1 13997
0 13999 7 1 2 66221 13998
0 14000 5 1 1 13999
0 14001 7 3 2 81844 76300
0 14002 5 3 1 95093
0 14003 7 1 2 64327 95094
0 14004 5 1 1 14003
0 14005 7 1 2 68342 14004
0 14006 7 1 2 14000 14005
0 14007 5 1 1 14006
0 14008 7 1 2 13984 14007
0 14009 5 1 1 14008
0 14010 7 1 2 69454 89651
0 14011 5 1 1 14010
0 14012 7 1 2 73021 14011
0 14013 7 1 2 14009 14012
0 14014 5 1 1 14013
0 14015 7 4 2 70135 77962
0 14016 5 2 1 95099
0 14017 7 1 2 82795 95103
0 14018 5 1 1 14017
0 14019 7 1 2 64657 14018
0 14020 5 1 1 14019
0 14021 7 1 2 68343 81621
0 14022 5 1 1 14021
0 14023 7 1 2 14020 14022
0 14024 5 1 1 14023
0 14025 7 1 2 81845 14024
0 14026 5 1 1 14025
0 14027 7 3 2 81710 76202
0 14028 7 1 2 71606 95105
0 14029 5 1 1 14028
0 14030 7 1 2 94179 14029
0 14031 5 1 1 14030
0 14032 7 1 2 68344 14031
0 14033 5 1 1 14032
0 14034 7 2 2 82370 86550
0 14035 5 1 1 95108
0 14036 7 5 2 84803 95109
0 14037 7 3 2 68618 76203
0 14038 5 1 1 95115
0 14039 7 1 2 95110 95116
0 14040 5 1 1 14039
0 14041 7 1 2 67983 14040
0 14042 7 1 2 14033 14041
0 14043 7 1 2 14026 14042
0 14044 5 1 1 14043
0 14045 7 1 2 14014 14044
0 14046 5 1 1 14045
0 14047 7 1 2 13980 14046
0 14048 5 1 1 14047
0 14049 7 1 2 76726 14048
0 14050 5 1 1 14049
0 14051 7 1 2 76204 80796
0 14052 5 1 1 14051
0 14053 7 1 2 79252 14052
0 14054 5 1 1 14053
0 14055 7 1 2 81317 14054
0 14056 5 1 1 14055
0 14057 7 1 2 82964 14056
0 14058 5 1 1 14057
0 14059 7 1 2 77925 92100
0 14060 5 1 1 14059
0 14061 7 2 2 76301 83632
0 14062 5 1 1 95118
0 14063 7 1 2 82902 14062
0 14064 7 1 2 14060 14063
0 14065 5 1 1 14064
0 14066 7 1 2 14058 14065
0 14067 5 1 1 14066
0 14068 7 4 2 66222 82292
0 14069 5 5 1 95120
0 14070 7 1 2 95121 93032
0 14071 5 1 1 14070
0 14072 7 1 2 65358 14071
0 14073 7 1 2 14067 14072
0 14074 5 1 1 14073
0 14075 7 1 2 84717 86935
0 14076 5 1 1 14075
0 14077 7 1 2 74635 14076
0 14078 5 1 1 14077
0 14079 7 1 2 82347 79505
0 14080 5 1 1 14079
0 14081 7 1 2 14078 14080
0 14082 5 1 1 14081
0 14083 7 1 2 64328 14082
0 14084 5 1 1 14083
0 14085 7 1 2 79248 91755
0 14086 5 1 1 14085
0 14087 7 2 2 70136 94390
0 14088 5 1 1 95129
0 14089 7 1 2 76205 95130
0 14090 5 1 1 14089
0 14091 7 1 2 14086 14090
0 14092 5 1 1 14091
0 14093 7 1 2 73419 14092
0 14094 5 1 1 14093
0 14095 7 1 2 70384 14094
0 14096 7 1 2 14084 14095
0 14097 5 1 1 14096
0 14098 7 1 2 14074 14097
0 14099 5 1 1 14098
0 14100 7 8 2 64658 79554
0 14101 7 1 2 95131 94381
0 14102 5 1 1 14101
0 14103 7 1 2 14099 14102
0 14104 5 1 1 14103
0 14105 7 1 2 67984 14104
0 14106 5 1 1 14105
0 14107 7 1 2 88859 94154
0 14108 5 2 1 14107
0 14109 7 1 2 76568 95139
0 14110 5 1 1 14109
0 14111 7 1 2 83060 91587
0 14112 5 1 1 14111
0 14113 7 2 2 14110 14112
0 14114 7 1 2 84092 95141
0 14115 5 1 1 14114
0 14116 7 1 2 69455 14115
0 14117 5 1 1 14116
0 14118 7 1 2 77932 83633
0 14119 5 1 1 14118
0 14120 7 1 2 82061 14119
0 14121 5 1 1 14120
0 14122 7 1 2 75125 14121
0 14123 5 1 1 14122
0 14124 7 1 2 93433 94157
0 14125 5 1 1 14124
0 14126 7 1 2 14123 14125
0 14127 7 1 2 14117 14126
0 14128 5 1 1 14127
0 14129 7 1 2 73022 14128
0 14130 5 1 1 14129
0 14131 7 3 2 78592 87140
0 14132 5 3 1 95143
0 14133 7 1 2 70385 95146
0 14134 5 1 1 14133
0 14135 7 1 2 73957 83005
0 14136 5 1 1 14135
0 14137 7 1 2 14134 14136
0 14138 5 1 1 14137
0 14139 7 1 2 82055 14138
0 14140 5 1 1 14139
0 14141 7 1 2 14130 14140
0 14142 7 1 2 14106 14141
0 14143 5 1 1 14142
0 14144 7 1 2 14143 74111
0 14145 5 1 1 14144
0 14146 7 1 2 14050 14145
0 14147 5 1 1 14146
0 14148 7 1 2 65955 14147
0 14149 5 1 1 14148
0 14150 7 5 2 68345 94725
0 14151 5 1 1 95149
0 14152 7 1 2 95150 76727
0 14153 5 1 1 14152
0 14154 7 1 2 75739 85404
0 14155 7 1 2 90136 14154
0 14156 5 1 1 14155
0 14157 7 1 2 14153 14156
0 14158 5 1 1 14157
0 14159 7 1 2 66501 14158
0 14160 5 1 1 14159
0 14161 7 3 2 68966 94095
0 14162 7 1 2 71028 86871
0 14163 5 1 1 14162
0 14164 7 2 2 84789 83902
0 14165 7 1 2 71607 95157
0 14166 5 1 1 14165
0 14167 7 1 2 14163 14166
0 14168 5 1 1 14167
0 14169 7 1 2 95154 14168
0 14170 5 1 1 14169
0 14171 7 1 2 14160 14170
0 14172 5 1 1 14171
0 14173 7 1 2 66223 14172
0 14174 5 1 1 14173
0 14175 7 4 2 66687 92364
0 14176 7 8 2 73712 74734
0 14177 7 1 2 95159 95163
0 14178 7 1 2 77643 14177
0 14179 5 1 1 14178
0 14180 7 1 2 14174 14179
0 14181 5 1 1 14180
0 14182 7 1 2 64659 14181
0 14183 5 1 1 14182
0 14184 7 2 2 86476 95164
0 14185 5 2 1 95171
0 14186 7 1 2 71029 90028
0 14187 7 1 2 77839 14186
0 14188 7 1 2 95172 14187
0 14189 5 1 1 14188
0 14190 7 1 2 14183 14189
0 14191 5 1 1 14190
0 14192 7 1 2 64329 14191
0 14193 5 1 1 14192
0 14194 7 1 2 70137 89169
0 14195 5 1 1 14194
0 14196 7 1 2 77792 76901
0 14197 7 1 2 14195 14196
0 14198 5 1 1 14197
0 14199 7 3 2 70386 80440
0 14200 5 2 1 95175
0 14201 7 1 2 90469 11320
0 14202 7 2 2 82903 83289
0 14203 5 1 1 95180
0 14204 7 1 2 74112 14203
0 14205 7 1 2 14201 14204
0 14206 7 1 2 95178 14205
0 14207 5 1 1 14206
0 14208 7 1 2 14198 14207
0 14209 5 1 1 14208
0 14210 7 1 2 66502 14209
0 14211 5 1 1 14210
0 14212 7 1 2 65041 87608
0 14213 7 1 2 94500 14212
0 14214 5 1 1 14213
0 14215 7 1 2 14211 14214
0 14216 5 1 1 14215
0 14217 7 1 2 66224 14216
0 14218 5 1 1 14217
0 14219 7 2 2 80341 83149
0 14220 5 2 1 95182
0 14221 7 1 2 86776 95184
0 14222 7 1 2 74113 14221
0 14223 5 1 1 14222
0 14224 7 1 2 76740 14223
0 14225 5 1 1 14224
0 14226 7 1 2 78376 14225
0 14227 5 1 1 14226
0 14228 7 1 2 14218 14227
0 14229 5 1 1 14228
0 14230 7 1 2 73420 14229
0 14231 5 1 1 14230
0 14232 7 1 2 89059 82283
0 14233 5 1 1 14232
0 14234 7 1 2 77044 14233
0 14235 5 1 1 14234
0 14236 7 4 2 71328 81846
0 14237 5 1 1 95186
0 14238 7 1 2 64330 14237
0 14239 5 1 1 14238
0 14240 7 5 2 65042 84974
0 14241 7 2 2 82904 95190
0 14242 5 1 1 95195
0 14243 7 1 2 14239 14242
0 14244 7 1 2 14235 14243
0 14245 5 1 1 14244
0 14246 7 1 2 76728 14245
0 14247 5 1 1 14246
0 14248 7 1 2 70387 80400
0 14249 5 3 1 14248
0 14250 7 2 2 83011 95197
0 14251 5 4 1 95200
0 14252 7 1 2 68967 82679
0 14253 7 1 2 75768 14252
0 14254 7 1 2 95202 14253
0 14255 5 1 1 14254
0 14256 7 1 2 14247 14255
0 14257 5 1 1 14256
0 14258 7 1 2 71030 14257
0 14259 5 1 1 14258
0 14260 7 1 2 14231 14259
0 14261 5 1 1 14260
0 14262 7 1 2 64660 14261
0 14263 5 1 1 14262
0 14264 7 1 2 95140 74114
0 14265 5 1 1 14264
0 14266 7 1 2 85678 76729
0 14267 5 1 1 14266
0 14268 7 1 2 14265 14267
0 14269 5 1 1 14268
0 14270 7 1 2 66225 14269
0 14271 5 1 1 14270
0 14272 7 3 2 71329 82905
0 14273 7 1 2 95206 78640
0 14274 7 1 2 77644 14273
0 14275 5 1 1 14274
0 14276 7 1 2 14271 14275
0 14277 5 1 1 14276
0 14278 7 1 2 78377 14277
0 14279 5 1 1 14278
0 14280 7 1 2 14263 14279
0 14281 5 1 1 14280
0 14282 7 1 2 73023 14281
0 14283 5 1 1 14282
0 14284 7 1 2 14193 14283
0 14285 7 1 2 14149 14284
0 14286 5 1 1 14285
0 14287 7 1 2 72604 14286
0 14288 5 1 1 14287
0 14289 7 9 2 67594 77320
0 14290 5 1 1 95209
0 14291 7 1 2 92802 87585
0 14292 5 1 1 14291
0 14293 7 1 2 86565 77635
0 14294 5 1 1 14293
0 14295 7 1 2 76741 14294
0 14296 5 1 1 14295
0 14297 7 2 2 71330 12201
0 14298 5 3 1 95218
0 14299 7 1 2 69773 95219
0 14300 5 1 1 14299
0 14301 7 1 2 14296 14300
0 14302 5 1 1 14301
0 14303 7 1 2 14292 14302
0 14304 5 1 1 14303
0 14305 7 1 2 80094 14304
0 14306 5 1 1 14305
0 14307 7 1 2 76206 76730
0 14308 5 1 1 14307
0 14309 7 3 2 76569 86585
0 14310 7 2 2 95223 77938
0 14311 7 1 2 95226 74115
0 14312 5 1 1 14311
0 14313 7 1 2 14308 14312
0 14314 7 1 2 14306 14313
0 14315 5 1 1 14314
0 14316 7 1 2 73024 14315
0 14317 5 1 1 14316
0 14318 7 1 2 92058 76380
0 14319 7 1 2 74220 14318
0 14320 5 1 1 14319
0 14321 7 8 2 71922 91066
0 14322 7 1 2 95228 74451
0 14323 5 1 1 14322
0 14324 7 1 2 14320 14323
0 14325 5 1 1 14324
0 14326 7 1 2 76570 14325
0 14327 5 1 1 14326
0 14328 7 1 2 92059 74221
0 14329 7 1 2 87944 14328
0 14330 5 1 1 14329
0 14331 7 1 2 14327 14330
0 14332 5 1 1 14331
0 14333 7 1 2 73958 14332
0 14334 5 1 1 14333
0 14335 7 2 2 75664 90261
0 14336 5 2 1 95236
0 14337 7 1 2 95238 77846
0 14338 5 1 1 14337
0 14339 7 1 2 89975 14338
0 14340 5 1 1 14339
0 14341 7 1 2 95237 89285
0 14342 5 1 1 14341
0 14343 7 1 2 76302 83366
0 14344 5 2 1 14343
0 14345 7 1 2 95240 95155
0 14346 5 1 1 14345
0 14347 7 1 2 14342 14346
0 14348 7 1 2 14340 14347
0 14349 7 1 2 14334 14348
0 14350 5 1 1 14349
0 14351 7 1 2 80681 14350
0 14352 5 1 1 14351
0 14353 7 1 2 64661 95220
0 14354 5 1 1 14353
0 14355 7 2 2 65359 77045
0 14356 7 1 2 66688 95242
0 14357 5 1 1 14356
0 14358 7 1 2 14354 14357
0 14359 5 2 1 14358
0 14360 7 1 2 80095 76731
0 14361 5 1 1 14360
0 14362 7 1 2 86942 74116
0 14363 5 1 1 14362
0 14364 7 1 2 14361 14363
0 14365 5 1 1 14364
0 14366 7 1 2 95244 14365
0 14367 5 1 1 14366
0 14368 7 1 2 77553 83369
0 14369 5 1 1 14368
0 14370 7 1 2 79945 14369
0 14371 5 1 1 14370
0 14372 7 1 2 83933 74117
0 14373 5 1 1 14372
0 14374 7 1 2 76742 14373
0 14375 5 1 1 14374
0 14376 7 1 2 87452 14375
0 14377 7 1 2 14371 14376
0 14378 5 1 1 14377
0 14379 7 1 2 14367 14378
0 14380 7 1 2 14352 14379
0 14381 7 1 2 14317 14380
0 14382 5 1 1 14381
0 14383 7 1 2 95210 14382
0 14384 5 1 1 14383
0 14385 7 1 2 14288 14384
0 14386 5 1 1 14385
0 14387 7 1 2 65748 14386
0 14388 5 1 1 14387
0 14389 7 1 2 94297 76732
0 14390 5 1 1 14389
0 14391 7 1 2 86398 76002
0 14392 7 1 2 94040 14391
0 14393 5 1 1 14392
0 14394 7 1 2 14390 14393
0 14395 5 1 1 14394
0 14396 7 1 2 66503 14395
0 14397 5 1 1 14396
0 14398 7 1 2 93947 74118
0 14399 5 1 1 14398
0 14400 7 1 2 66689 77096
0 14401 5 3 1 14400
0 14402 7 1 2 95246 80522
0 14403 5 1 1 14402
0 14404 7 1 2 76733 14403
0 14405 5 1 1 14404
0 14406 7 1 2 14399 14405
0 14407 5 1 1 14406
0 14408 7 1 2 65360 14407
0 14409 5 1 1 14408
0 14410 7 2 2 82592 94811
0 14411 7 1 2 87621 95249
0 14412 5 1 1 14411
0 14413 7 1 2 74876 76734
0 14414 5 1 1 14413
0 14415 7 1 2 80504 74119
0 14416 5 1 1 14415
0 14417 7 1 2 14414 14416
0 14418 5 1 1 14417
0 14419 7 1 2 66504 14418
0 14420 5 1 1 14419
0 14421 7 1 2 14412 14420
0 14422 7 1 2 14409 14421
0 14423 5 1 1 14422
0 14424 7 1 2 65043 14423
0 14425 5 1 1 14424
0 14426 7 1 2 14397 14425
0 14427 5 1 1 14426
0 14428 7 2 2 65956 74330
0 14429 7 6 2 64331 73025
0 14430 5 1 1 95253
0 14431 7 1 2 93085 95254
0 14432 7 1 2 95251 14431
0 14433 7 1 2 14427 14432
0 14434 5 1 1 14433
0 14435 7 1 2 14388 14434
0 14436 5 1 1 14435
0 14437 7 1 2 64053 14436
0 14438 5 1 1 14437
0 14439 7 1 2 88291 90411
0 14440 5 2 1 14439
0 14441 7 12 2 71794 67595
0 14442 7 6 2 69774 70774
0 14443 7 7 2 69112 71031
0 14444 7 1 2 95273 95279
0 14445 7 1 2 95261 14444
0 14446 7 1 2 90002 14445
0 14447 7 1 2 95259 14446
0 14448 5 1 1 14447
0 14449 7 1 2 67082 74147
0 14450 7 1 2 83663 14449
0 14451 7 10 2 72605 73713
0 14452 5 2 1 95286
0 14453 7 3 2 66690 95287
0 14454 7 1 2 95298 84442
0 14455 7 1 2 14450 14454
0 14456 5 1 1 14455
0 14457 7 1 2 14448 14456
0 14458 5 1 1 14457
0 14459 7 1 2 69456 14458
0 14460 5 1 1 14459
0 14461 7 1 2 81328 84392
0 14462 5 1 1 14461
0 14463 7 4 2 64332 93137
0 14464 7 18 2 66691 72606
0 14465 5 1 1 95305
0 14466 7 1 2 84317 95306
0 14467 7 1 2 74284 14466
0 14468 7 1 2 95301 14467
0 14469 7 1 2 14462 14468
0 14470 5 1 1 14469
0 14471 7 1 2 14460 14470
0 14472 5 1 1 14471
0 14473 7 1 2 75740 14472
0 14474 5 1 1 14473
0 14475 7 1 2 84961 78109
0 14476 7 1 2 84268 14475
0 14477 7 2 2 87880 92407
0 14478 7 1 2 86375 95323
0 14479 7 1 2 14476 14478
0 14480 5 1 1 14479
0 14481 7 1 2 14474 14480
0 14482 5 1 1 14481
0 14483 7 1 2 78690 14482
0 14484 5 1 1 14483
0 14485 7 2 2 92336 83618
0 14486 7 1 2 95325 93495
0 14487 7 1 2 94769 14486
0 14488 5 1 1 14487
0 14489 7 1 2 89022 79946
0 14490 5 1 1 14489
0 14491 7 1 2 66505 11478
0 14492 5 1 1 14491
0 14493 7 1 2 80149 14492
0 14494 5 1 1 14493
0 14495 7 1 2 14490 14494
0 14496 5 1 1 14495
0 14497 7 1 2 70138 14496
0 14498 5 1 1 14497
0 14499 7 4 2 69775 86693
0 14500 7 1 2 95327 76752
0 14501 5 1 1 14500
0 14502 7 1 2 14498 14501
0 14503 5 1 1 14502
0 14504 7 16 2 70775 71032
0 14505 5 1 1 95331
0 14506 7 7 2 69457 95332
0 14507 5 1 1 95347
0 14508 7 3 2 63884 67596
0 14509 7 1 2 95348 95354
0 14510 7 1 2 14503 14509
0 14511 5 1 1 14510
0 14512 7 1 2 14488 14511
0 14513 5 1 1 14512
0 14514 7 1 2 67083 14513
0 14515 5 1 1 14514
0 14516 7 3 2 88377 87446
0 14517 5 2 1 95357
0 14518 7 1 2 70139 78014
0 14519 5 2 1 14518
0 14520 7 1 2 95360 95362
0 14521 5 1 1 14520
0 14522 7 9 2 69458 70776
0 14523 7 5 2 71033 95364
0 14524 7 2 2 68968 76464
0 14525 7 2 2 95373 95378
0 14526 7 7 2 67597 75556
0 14527 7 1 2 72136 95382
0 14528 7 1 2 95380 14527
0 14529 7 1 2 14521 14528
0 14530 5 1 1 14529
0 14531 7 1 2 14515 14530
0 14532 5 1 1 14531
0 14533 7 1 2 75741 14532
0 14534 5 1 1 14533
0 14535 7 2 2 74311 85427
0 14536 7 3 2 73026 91482
0 14537 7 1 2 92337 91150
0 14538 7 1 2 95391 14537
0 14539 7 1 2 95389 14538
0 14540 7 1 2 94304 14539
0 14541 5 1 1 14540
0 14542 7 1 2 14534 14541
0 14543 5 1 1 14542
0 14544 7 1 2 69113 14543
0 14545 5 1 1 14544
0 14546 7 1 2 14484 14545
0 14547 7 1 2 14438 14546
0 14548 5 1 1 14547
0 14549 7 1 2 74027 14548
0 14550 5 1 1 14549
0 14551 7 2 2 72607 79543
0 14552 5 1 1 95394
0 14553 7 2 2 78148 79863
0 14554 5 2 1 95396
0 14555 7 1 2 14552 95398
0 14556 5 1 1 14555
0 14557 7 1 2 67985 14556
0 14558 5 2 1 14557
0 14559 7 2 2 72608 83321
0 14560 5 1 1 95402
0 14561 7 1 2 92639 14560
0 14562 5 1 1 14561
0 14563 7 1 2 71331 14562
0 14564 5 1 1 14563
0 14565 7 2 2 79555 87792
0 14566 5 1 1 95404
0 14567 7 1 2 73421 14566
0 14568 7 1 2 14564 14567
0 14569 7 1 2 95400 14568
0 14570 5 1 1 14569
0 14571 7 2 2 69776 78958
0 14572 5 1 1 95406
0 14573 7 2 2 79620 14572
0 14574 7 1 2 95408 86707
0 14575 5 1 1 14574
0 14576 7 1 2 68346 91461
0 14577 7 1 2 14575 14576
0 14578 5 1 1 14577
0 14579 7 1 2 79486 14578
0 14580 7 1 2 14570 14579
0 14581 5 1 1 14580
0 14582 7 1 2 77534 86265
0 14583 5 1 1 14582
0 14584 7 3 2 79628 84583
0 14585 7 1 2 75044 95410
0 14586 7 1 2 14583 14585
0 14587 5 1 1 14586
0 14588 7 1 2 14581 14587
0 14589 5 1 1 14588
0 14590 7 1 2 75217 14589
0 14591 5 1 1 14590
0 14592 7 5 2 66856 72609
0 14593 7 6 2 79629 95413
0 14594 7 1 2 79616 95418
0 14595 5 1 1 14594
0 14596 7 2 2 71332 79826
0 14597 5 4 1 95424
0 14598 7 2 2 95425 87244
0 14599 5 2 1 95430
0 14600 7 1 2 73027 95432
0 14601 5 1 1 14600
0 14602 7 2 2 9089 88312
0 14603 5 1 1 95434
0 14604 7 1 2 74636 14603
0 14605 5 1 1 14604
0 14606 7 1 2 14601 14605
0 14607 5 1 1 14606
0 14608 7 1 2 78861 14607
0 14609 5 1 1 14608
0 14610 7 2 2 79409 79135
0 14611 7 2 2 73422 81275
0 14612 5 1 1 95438
0 14613 7 1 2 73714 95439
0 14614 7 1 2 95436 14613
0 14615 5 1 1 14614
0 14616 7 1 2 14609 14615
0 14617 5 1 1 14616
0 14618 7 1 2 67598 14617
0 14619 5 1 1 14618
0 14620 7 1 2 14595 14619
0 14621 5 1 1 14620
0 14622 7 1 2 76767 14621
0 14623 5 1 1 14622
0 14624 7 1 2 14591 14623
0 14625 5 1 1 14624
0 14626 7 1 2 64333 14625
0 14627 5 1 1 14626
0 14628 7 1 2 86502 86430
0 14629 7 2 2 91116 14628
0 14630 7 1 2 81260 87733
0 14631 7 1 2 95440 14630
0 14632 5 1 1 14631
0 14633 7 1 2 14627 14632
0 14634 5 1 1 14633
0 14635 7 1 2 65957 14634
0 14636 5 1 1 14635
0 14637 7 5 2 73028 76381
0 14638 7 1 2 95442 80187
0 14639 5 2 1 14638
0 14640 7 1 2 95165 91117
0 14641 7 2 2 87970 14640
0 14642 5 1 1 95449
0 14643 7 1 2 95447 14642
0 14644 5 2 1 14643
0 14645 7 1 2 80018 95451
0 14646 5 1 1 14645
0 14647 7 1 2 64334 82044
0 14648 5 1 1 14647
0 14649 7 1 2 79400 14648
0 14650 5 1 1 14649
0 14651 7 1 2 87376 94871
0 14652 5 1 1 14651
0 14653 7 2 2 72137 83561
0 14654 7 1 2 75193 95453
0 14655 5 1 1 14654
0 14656 7 1 2 14652 14655
0 14657 5 1 1 14656
0 14658 7 1 2 69459 79487
0 14659 7 1 2 14657 14658
0 14660 5 1 1 14659
0 14661 7 1 2 14650 14660
0 14662 5 1 1 14661
0 14663 7 1 2 64662 14662
0 14664 5 1 1 14663
0 14665 7 1 2 87852 87936
0 14666 5 1 1 14665
0 14667 7 1 2 69460 95450
0 14668 5 1 1 14667
0 14669 7 1 2 14666 14668
0 14670 7 1 2 14664 14669
0 14671 5 1 1 14670
0 14672 7 1 2 66226 14671
0 14673 5 1 1 14672
0 14674 7 1 2 14646 14673
0 14675 5 1 1 14674
0 14676 7 1 2 65958 14675
0 14677 5 1 1 14676
0 14678 7 5 2 66227 78378
0 14679 7 1 2 95455 95452
0 14680 5 1 1 14679
0 14681 7 1 2 77598 79656
0 14682 5 1 1 14681
0 14683 7 1 2 86341 82788
0 14684 7 1 2 79789 14683
0 14685 5 1 1 14684
0 14686 7 1 2 14682 14685
0 14687 5 1 1 14686
0 14688 7 1 2 66228 14687
0 14689 5 1 1 14688
0 14690 7 2 2 83370 79755
0 14691 5 1 1 95460
0 14692 7 1 2 95461 79015
0 14693 5 1 1 14692
0 14694 7 1 2 14689 14693
0 14695 5 1 1 14694
0 14696 7 1 2 75218 14695
0 14697 5 1 1 14696
0 14698 7 1 2 87942 14697
0 14699 5 1 1 14698
0 14700 7 1 2 71034 14699
0 14701 5 1 1 14700
0 14702 7 3 2 73029 77625
0 14703 5 2 1 95462
0 14704 7 2 2 72138 92509
0 14705 7 3 2 79630 89864
0 14706 7 1 2 95467 95469
0 14707 7 1 2 95463 14706
0 14708 5 1 1 14707
0 14709 7 1 2 14701 14708
0 14710 5 1 1 14709
0 14711 7 1 2 64663 14710
0 14712 5 1 1 14711
0 14713 7 1 2 14680 14712
0 14714 7 1 2 14677 14713
0 14715 5 1 1 14714
0 14716 7 1 2 72610 14715
0 14717 5 1 1 14716
0 14718 7 1 2 76869 95079
0 14719 7 1 2 95441 14718
0 14720 5 1 1 14719
0 14721 7 1 2 14717 14720
0 14722 7 1 2 14636 14721
0 14723 5 1 1 14722
0 14724 7 1 2 65749 14723
0 14725 5 1 1 14724
0 14726 7 1 2 73959 94845
0 14727 5 1 1 14726
0 14728 7 1 2 14727 1047
0 14729 5 1 1 14728
0 14730 7 6 2 66229 82239
0 14731 7 1 2 95472 74312
0 14732 7 2 2 14729 14731
0 14733 7 1 2 63763 77985
0 14734 7 1 2 94071 14733
0 14735 7 1 2 95478 14734
0 14736 5 1 1 14735
0 14737 7 1 2 14725 14736
0 14738 5 1 1 14737
0 14739 7 1 2 64054 14738
0 14740 5 1 1 14739
0 14741 7 5 2 65585 65750
0 14742 7 1 2 95480 84467
0 14743 7 1 2 95479 14742
0 14744 5 1 1 14743
0 14745 7 1 2 14740 14744
0 14746 5 1 1 14745
0 14747 7 1 2 80682 14746
0 14748 5 1 1 14747
0 14749 7 1 2 73030 88830
0 14750 5 6 1 14749
0 14751 7 1 2 75487 95485
0 14752 5 1 1 14751
0 14753 7 1 2 84253 83162
0 14754 5 1 1 14753
0 14755 7 1 2 87837 14754
0 14756 7 1 2 14752 14755
0 14757 5 1 1 14756
0 14758 7 1 2 84017 95381
0 14759 7 1 2 14757 14758
0 14760 5 1 1 14759
0 14761 7 1 2 86342 95221
0 14762 5 1 1 14761
0 14763 7 1 2 82230 14762
0 14764 5 1 1 14763
0 14765 7 1 2 73031 14764
0 14766 5 1 1 14765
0 14767 7 5 2 65361 88703
0 14768 5 1 1 95491
0 14769 7 1 2 95492 86804
0 14770 5 1 1 14769
0 14771 7 1 2 14766 14770
0 14772 5 1 1 14771
0 14773 7 1 2 64664 14772
0 14774 5 1 1 14773
0 14775 7 1 2 77867 95196
0 14776 5 1 1 14775
0 14777 7 1 2 14774 14776
0 14778 5 1 1 14777
0 14779 7 2 2 93247 78361
0 14780 7 1 2 91151 95496
0 14781 7 1 2 14778 14780
0 14782 5 1 1 14781
0 14783 7 1 2 14760 14782
0 14784 5 1 1 14783
0 14785 7 1 2 78862 14784
0 14786 5 1 1 14785
0 14787 7 2 2 68969 76954
0 14788 7 1 2 95498 92954
0 14789 7 2 2 71608 91865
0 14790 7 9 2 70777 71333
0 14791 5 1 1 95502
0 14792 7 5 2 70140 71035
0 14793 5 1 1 95511
0 14794 7 4 2 95503 95512
0 14795 7 1 2 95500 95516
0 14796 7 1 2 14788 14795
0 14797 5 1 1 14796
0 14798 7 8 2 64335 65751
0 14799 7 3 2 82527 95520
0 14800 7 2 2 95528 92800
0 14801 7 2 2 76994 92575
0 14802 7 1 2 88704 86417
0 14803 7 1 2 95533 14802
0 14804 7 1 2 95531 14803
0 14805 5 1 1 14804
0 14806 7 1 2 14797 14805
0 14807 5 1 1 14806
0 14808 7 1 2 79136 14807
0 14809 5 1 1 14808
0 14810 7 1 2 14786 14809
0 14811 5 1 1 14810
0 14812 7 1 2 72139 14811
0 14813 5 1 1 14812
0 14814 7 1 2 66230 13761
0 14815 5 1 1 14814
0 14816 7 2 2 86343 77659
0 14817 7 1 2 94218 95535
0 14818 5 1 1 14817
0 14819 7 1 2 14815 14818
0 14820 5 1 1 14819
0 14821 7 1 2 64665 14820
0 14822 5 1 1 14821
0 14823 7 2 2 83664 94009
0 14824 7 1 2 79537 95537
0 14825 5 1 1 14824
0 14826 7 1 2 14822 14825
0 14827 5 1 1 14826
0 14828 7 4 2 72611 78159
0 14829 7 2 2 68970 77321
0 14830 7 1 2 95543 95481
0 14831 7 1 2 95539 14830
0 14832 7 1 2 14827 14831
0 14833 5 1 1 14832
0 14834 7 1 2 78863 95486
0 14835 5 1 1 14834
0 14836 7 5 2 68812 80584
0 14837 7 1 2 95545 76799
0 14838 7 1 2 76753 14837
0 14839 5 1 1 14838
0 14840 7 1 2 14835 14839
0 14841 5 1 1 14840
0 14842 7 1 2 75360 14841
0 14843 5 1 1 14842
0 14844 7 1 2 84254 94970
0 14845 5 1 1 14844
0 14846 7 3 2 74528 76800
0 14847 7 1 2 68813 75557
0 14848 7 1 2 95550 14847
0 14849 5 1 1 14848
0 14850 7 1 2 14845 14849
0 14851 5 1 1 14850
0 14852 7 1 2 75126 14851
0 14853 5 1 1 14852
0 14854 7 1 2 14843 14853
0 14855 5 1 1 14854
0 14856 7 2 2 95274 89865
0 14857 7 1 2 93076 95553
0 14858 7 1 2 14855 14857
0 14859 5 1 1 14858
0 14860 7 1 2 14833 14859
0 14861 5 1 1 14860
0 14862 7 1 2 76843 14861
0 14863 5 1 1 14862
0 14864 7 1 2 14813 14863
0 14865 5 1 1 14864
0 14866 7 1 2 69114 14865
0 14867 5 1 1 14866
0 14868 7 1 2 87358 76768
0 14869 5 1 1 14868
0 14870 7 1 2 71795 74263
0 14871 5 1 1 14870
0 14872 7 1 2 14869 14871
0 14873 5 1 1 14872
0 14874 7 1 2 71609 14873
0 14875 5 1 1 14874
0 14876 7 1 2 85650 74264
0 14877 5 1 1 14876
0 14878 7 1 2 14875 14877
0 14879 5 1 1 14878
0 14880 7 1 2 68619 14879
0 14881 5 1 1 14880
0 14882 7 4 2 80585 75219
0 14883 5 1 1 95555
0 14884 7 1 2 78691 95556
0 14885 5 1 1 14884
0 14886 7 1 2 14881 14885
0 14887 5 1 1 14886
0 14888 7 1 2 73032 14887
0 14889 5 1 1 14888
0 14890 7 1 2 94105 90051
0 14891 5 1 1 14890
0 14892 7 1 2 14889 14891
0 14893 5 1 1 14892
0 14894 7 2 2 93040 93248
0 14895 7 1 2 87957 93568
0 14896 7 1 2 95559 14895
0 14897 7 1 2 14893 14896
0 14898 5 1 1 14897
0 14899 7 1 2 90968 89766
0 14900 5 1 1 14899
0 14901 7 1 2 75127 14900
0 14902 5 1 1 14901
0 14903 7 1 2 78015 91812
0 14904 5 1 1 14903
0 14905 7 1 2 14902 14904
0 14906 5 1 1 14905
0 14907 7 1 2 68347 14906
0 14908 5 1 1 14907
0 14909 7 1 2 86107 89761
0 14910 5 1 1 14909
0 14911 7 1 2 14908 14910
0 14912 5 1 1 14911
0 14913 7 5 2 69461 65586
0 14914 7 2 2 95333 95561
0 14915 7 2 2 69115 67986
0 14916 7 3 2 78160 84018
0 14917 7 1 2 95568 95570
0 14918 7 1 2 95566 14917
0 14919 7 1 2 14912 14918
0 14920 5 1 1 14919
0 14921 7 1 2 14898 14920
0 14922 5 1 1 14921
0 14923 7 1 2 70141 14922
0 14924 5 1 1 14923
0 14925 7 5 2 63764 93726
0 14926 7 2 2 95573 75831
0 14927 7 4 2 71610 82348
0 14928 7 1 2 90988 95580
0 14929 7 1 2 95567 14928
0 14930 7 1 2 95578 14929
0 14931 5 1 1 14930
0 14932 7 6 2 64336 65587
0 14933 7 1 2 74313 89690
0 14934 7 1 2 95584 14933
0 14935 7 4 2 65752 93763
0 14936 7 2 2 74210 91238
0 14937 7 1 2 95590 95594
0 14938 7 1 2 14934 14937
0 14939 5 1 1 14938
0 14940 7 1 2 14931 14939
0 14941 5 1 1 14940
0 14942 7 1 2 70388 14941
0 14943 5 1 1 14942
0 14944 7 2 2 69116 79631
0 14945 7 2 2 95365 95596
0 14946 7 1 2 71036 93173
0 14947 7 1 2 76427 14946
0 14948 7 1 2 95598 14947
0 14949 5 1 1 14948
0 14950 7 3 2 65753 78986
0 14951 7 2 2 84523 95600
0 14952 7 3 2 65959 75742
0 14953 7 1 2 95605 95392
0 14954 7 1 2 95603 14953
0 14955 5 1 1 14954
0 14956 7 1 2 14949 14955
0 14957 5 1 1 14956
0 14958 7 1 2 70389 88786
0 14959 5 1 1 14958
0 14960 7 1 2 80816 14959
0 14961 5 1 1 14960
0 14962 7 1 2 63885 14961
0 14963 7 1 2 14957 14962
0 14964 5 1 1 14963
0 14965 7 1 2 14943 14964
0 14966 7 1 2 14924 14965
0 14967 5 1 1 14966
0 14968 7 1 2 76303 14967
0 14969 5 1 1 14968
0 14970 7 2 2 66231 86418
0 14971 7 2 2 74735 91483
0 14972 7 1 2 95608 95610
0 14973 7 1 2 95532 14972
0 14974 5 1 1 14973
0 14975 7 1 2 68348 89792
0 14976 5 1 1 14975
0 14977 7 1 2 7203 14976
0 14978 5 1 1 14977
0 14979 7 4 2 69117 76955
0 14980 7 9 2 70778 72028
0 14981 7 1 2 85076 95616
0 14982 7 1 2 95612 14981
0 14983 7 1 2 78052 14982
0 14984 7 1 2 14978 14983
0 14985 5 1 1 14984
0 14986 7 1 2 14974 14985
0 14987 5 1 1 14986
0 14988 7 1 2 78864 14987
0 14989 5 1 1 14988
0 14990 7 2 2 95383 84221
0 14991 7 3 2 84062 93592
0 14992 7 3 2 70390 75818
0 14993 7 14 2 69118 69462
0 14994 7 1 2 95633 91876
0 14995 7 1 2 95630 14994
0 14996 7 1 2 95627 14995
0 14997 7 1 2 95625 14996
0 14998 5 1 1 14997
0 14999 7 1 2 14989 14998
0 15000 5 1 1 14999
0 15001 7 1 2 82965 15000
0 15002 5 1 1 15001
0 15003 7 1 2 81432 80449
0 15004 5 1 1 15003
0 15005 7 1 2 73033 94255
0 15006 5 1 1 15005
0 15007 7 1 2 15004 15006
0 15008 5 1 1 15007
0 15009 7 6 2 65754 72140
0 15010 7 2 2 77897 95647
0 15011 7 1 2 82760 78362
0 15012 7 1 2 92522 15011
0 15013 7 1 2 95653 15012
0 15014 7 1 2 15008 15013
0 15015 5 1 1 15014
0 15016 7 1 2 15002 15015
0 15017 7 1 2 14969 15016
0 15018 7 1 2 14867 15017
0 15019 7 1 2 14748 15018
0 15020 7 1 2 14550 15019
0 15021 7 1 2 13974 15020
0 15022 5 1 1 15021
0 15023 7 1 2 73837 15022
0 15024 5 1 1 15023
0 15025 7 4 2 69061 76801
0 15026 7 1 2 86694 91167
0 15027 7 1 2 95655 15026
0 15028 5 1 1 15027
0 15029 7 1 2 89012 15028
0 15030 5 1 1 15029
0 15031 7 1 2 79334 15030
0 15032 5 1 1 15031
0 15033 7 1 2 79690 91933
0 15034 7 1 2 88041 15033
0 15035 5 1 1 15034
0 15036 7 1 2 89013 15035
0 15037 5 1 1 15036
0 15038 7 1 2 75220 15037
0 15039 5 1 1 15038
0 15040 7 1 2 15032 15039
0 15041 5 1 1 15040
0 15042 7 1 2 69777 15041
0 15043 5 1 1 15042
0 15044 7 4 2 66857 92029
0 15045 7 1 2 74276 1056
0 15046 5 2 1 15045
0 15047 7 1 2 95659 95663
0 15048 5 1 1 15047
0 15049 7 1 2 15043 15048
0 15050 5 1 1 15049
0 15051 7 1 2 63765 15050
0 15052 5 1 1 15051
0 15053 7 3 2 84485 90949
0 15054 7 1 2 74100 95665
0 15055 5 1 1 15054
0 15056 7 1 2 77933 89138
0 15057 7 1 2 75832 15056
0 15058 5 1 1 15057
0 15059 7 1 2 15055 15058
0 15060 5 1 1 15059
0 15061 7 1 2 90330 15060
0 15062 5 1 1 15061
0 15063 7 1 2 15052 15062
0 15064 5 1 1 15063
0 15065 7 1 2 68620 15064
0 15066 5 1 1 15065
0 15067 7 6 2 78161 75878
0 15068 5 1 1 95668
0 15069 7 4 2 71334 87406
0 15070 7 1 2 69778 92118
0 15071 7 1 2 95674 15070
0 15072 5 1 1 15071
0 15073 7 1 2 15068 15072
0 15074 5 1 1 15073
0 15075 7 1 2 76304 91532
0 15076 7 1 2 86618 15075
0 15077 7 1 2 15074 15076
0 15078 5 1 1 15077
0 15079 7 1 2 15066 15078
0 15080 5 1 1 15079
0 15081 7 1 2 67987 15080
0 15082 5 1 1 15081
0 15083 7 1 2 63766 95664
0 15084 5 1 1 15083
0 15085 7 4 2 72029 87734
0 15086 7 1 2 70391 77724
0 15087 7 1 2 95678 15086
0 15088 5 1 1 15087
0 15089 7 1 2 15084 15088
0 15090 5 1 1 15089
0 15091 7 1 2 94545 95660
0 15092 7 1 2 15090 15091
0 15093 5 1 1 15092
0 15094 7 1 2 15082 15093
0 15095 5 1 1 15094
0 15096 7 1 2 71796 15095
0 15097 5 1 1 15096
0 15098 7 1 2 67084 79369
0 15099 5 2 1 15098
0 15100 7 1 2 83055 87760
0 15101 5 1 1 15100
0 15102 7 1 2 95682 15101
0 15103 5 1 1 15102
0 15104 7 4 2 69779 92030
0 15105 7 1 2 76428 95684
0 15106 7 1 2 15103 15105
0 15107 5 1 1 15106
0 15108 7 1 2 15097 15107
0 15109 5 1 1 15108
0 15110 7 1 2 75361 15109
0 15111 5 1 1 15110
0 15112 7 5 2 80342 75558
0 15113 5 2 1 95688
0 15114 7 1 2 81281 95487
0 15115 5 1 1 15114
0 15116 7 1 2 95693 15115
0 15117 5 1 1 15116
0 15118 7 1 2 90209 15117
0 15119 5 1 1 15118
0 15120 7 3 2 92278 92514
0 15121 7 1 2 86606 95695
0 15122 5 1 1 15121
0 15123 7 5 2 67988 85887
0 15124 7 7 2 68621 82349
0 15125 5 1 1 95703
0 15126 7 1 2 71923 95704
0 15127 7 1 2 90533 15126
0 15128 5 1 1 15127
0 15129 7 1 2 89014 15128
0 15130 5 1 1 15129
0 15131 7 1 2 95698 15130
0 15132 5 1 1 15131
0 15133 7 1 2 15122 15132
0 15134 5 1 1 15133
0 15135 7 1 2 81608 15134
0 15136 5 1 1 15135
0 15137 7 1 2 15119 15136
0 15138 5 1 1 15137
0 15139 7 1 2 69780 15138
0 15140 5 1 1 15139
0 15141 7 2 2 88821 74945
0 15142 5 1 1 95710
0 15143 7 1 2 71335 95488
0 15144 5 1 1 15143
0 15145 7 1 2 95694 15144
0 15146 5 1 1 15145
0 15147 7 1 2 74529 15146
0 15148 5 1 1 15147
0 15149 7 1 2 15142 15148
0 15150 5 3 1 15149
0 15151 7 1 2 90210 95712
0 15152 5 1 1 15151
0 15153 7 1 2 15140 15152
0 15154 5 1 1 15153
0 15155 7 1 2 75879 15154
0 15156 5 1 1 15155
0 15157 7 1 2 79370 89754
0 15158 5 1 1 15157
0 15159 7 1 2 68349 87761
0 15160 5 1 1 15159
0 15161 7 1 2 15158 15160
0 15162 5 2 1 15161
0 15163 7 1 2 94630 95715
0 15164 5 1 1 15163
0 15165 7 9 2 68971 88020
0 15166 7 3 2 95717 91898
0 15167 7 1 2 67085 75559
0 15168 7 1 2 91680 15167
0 15169 7 1 2 95726 15168
0 15170 5 1 1 15169
0 15171 7 1 2 15164 15170
0 15172 5 1 1 15171
0 15173 7 1 2 72030 15172
0 15174 5 1 1 15173
0 15175 7 4 2 63767 91556
0 15176 7 4 2 67989 74237
0 15177 7 1 2 95729 95733
0 15178 7 1 2 91978 15177
0 15179 5 1 1 15178
0 15180 7 1 2 15174 15179
0 15181 5 1 1 15180
0 15182 7 1 2 91429 15181
0 15183 5 1 1 15182
0 15184 7 9 2 72031 67990
0 15185 7 2 2 95737 95661
0 15186 7 1 2 76645 95716
0 15187 7 1 2 95746 15186
0 15188 5 1 1 15187
0 15189 7 1 2 15183 15188
0 15190 5 1 1 15189
0 15191 7 1 2 75128 15190
0 15192 5 1 1 15191
0 15193 7 1 2 69781 95713
0 15194 5 1 1 15193
0 15195 7 3 2 75560 81609
0 15196 5 1 1 95748
0 15197 7 1 2 80343 95749
0 15198 5 1 1 15197
0 15199 7 1 2 15194 15198
0 15200 5 1 1 15199
0 15201 7 1 2 75769 90435
0 15202 7 1 2 15200 15201
0 15203 5 1 1 15202
0 15204 7 1 2 15192 15203
0 15205 7 1 2 15156 15204
0 15206 7 1 2 15111 15205
0 15207 5 1 1 15206
0 15208 7 1 2 67599 15207
0 15209 5 1 1 15208
0 15210 7 3 2 69782 86607
0 15211 7 1 2 90646 90285
0 15212 7 2 2 95751 15211
0 15213 7 2 2 77710 87102
0 15214 7 3 2 76821 95756
0 15215 7 3 2 74238 89541
0 15216 7 1 2 95758 95761
0 15217 7 1 2 95754 15216
0 15218 5 1 1 15217
0 15219 7 1 2 15209 15218
0 15220 5 1 1 15219
0 15221 7 1 2 71037 15220
0 15222 5 1 1 15221
0 15223 7 1 2 84053 84617
0 15224 7 1 2 90286 15223
0 15225 7 2 2 71797 89542
0 15226 7 1 2 76822 95764
0 15227 7 2 2 15224 15226
0 15228 7 1 2 70142 86197
0 15229 7 1 2 90256 15228
0 15230 7 1 2 95766 15229
0 15231 5 1 1 15230
0 15232 7 1 2 15222 15231
0 15233 5 1 1 15232
0 15234 7 1 2 69463 15233
0 15235 5 1 1 15234
0 15236 7 2 2 66858 74530
0 15237 7 1 2 76932 82820
0 15238 7 1 2 95768 15237
0 15239 7 1 2 95767 15238
0 15240 5 1 1 15239
0 15241 7 1 2 15235 15240
0 15242 5 1 1 15241
0 15243 7 1 2 69119 15242
0 15244 5 1 1 15243
0 15245 7 1 2 87256 91984
0 15246 5 1 1 15245
0 15247 7 1 2 89015 15246
0 15248 5 1 1 15247
0 15249 7 1 2 85253 15248
0 15250 5 1 1 15249
0 15251 7 5 2 71611 85622
0 15252 5 1 1 95770
0 15253 7 1 2 81847 95771
0 15254 5 1 1 15253
0 15255 7 1 2 90911 15254
0 15256 5 1 1 15255
0 15257 7 1 2 15250 15256
0 15258 5 1 1 15257
0 15259 7 1 2 73715 15258
0 15260 5 1 1 15259
0 15261 7 1 2 87471 90912
0 15262 5 1 1 15261
0 15263 7 1 2 15260 15262
0 15264 5 1 1 15263
0 15265 7 1 2 65044 15264
0 15266 5 1 1 15265
0 15267 7 1 2 85888 94298
0 15268 5 1 1 15267
0 15269 7 8 2 70392 82350
0 15270 5 5 1 95775
0 15271 7 1 2 85254 95783
0 15272 5 1 1 15271
0 15273 7 1 2 15268 15272
0 15274 5 1 1 15273
0 15275 7 1 2 66506 15274
0 15276 5 1 1 15275
0 15277 7 1 2 85255 85610
0 15278 5 1 1 15277
0 15279 7 1 2 15276 15278
0 15280 5 1 1 15279
0 15281 7 1 2 88978 15280
0 15282 5 1 1 15281
0 15283 7 1 2 15266 15282
0 15284 5 1 1 15283
0 15285 7 1 2 88552 15284
0 15286 5 1 1 15285
0 15287 7 3 2 75362 90111
0 15288 5 3 1 95788
0 15289 7 2 2 72032 95791
0 15290 7 1 2 68814 95794
0 15291 5 1 1 15290
0 15292 7 1 2 94022 15291
0 15293 5 1 1 15292
0 15294 7 1 2 88979 15293
0 15295 5 1 1 15294
0 15296 7 6 2 74637 78571
0 15297 5 3 1 95796
0 15298 7 1 2 95797 94581
0 15299 7 1 2 90384 15298
0 15300 5 1 1 15299
0 15301 7 1 2 15295 15300
0 15302 5 1 1 15301
0 15303 7 1 2 65362 15302
0 15304 5 1 1 15303
0 15305 7 2 2 86419 91404
0 15306 7 1 2 93483 95805
0 15307 5 1 1 15306
0 15308 7 1 2 11683 15307
0 15309 5 1 1 15308
0 15310 7 1 2 94756 15309
0 15311 5 1 1 15310
0 15312 7 1 2 3561 94019
0 15313 5 1 1 15312
0 15314 7 1 2 15125 88980
0 15315 7 1 2 15313 15314
0 15316 5 1 1 15315
0 15317 7 1 2 15311 15316
0 15318 7 1 2 15304 15317
0 15319 5 1 1 15318
0 15320 7 1 2 88184 15319
0 15321 5 1 1 15320
0 15322 7 1 2 15286 15321
0 15323 5 1 1 15322
0 15324 7 1 2 73034 15323
0 15325 5 1 1 15324
0 15326 7 2 2 65045 89188
0 15327 5 1 1 95807
0 15328 7 1 2 89324 15327
0 15329 5 1 1 15328
0 15330 7 1 2 65588 81586
0 15331 7 1 2 90313 15330
0 15332 7 1 2 95250 15331
0 15333 7 1 2 15329 15332
0 15334 5 1 1 15333
0 15335 7 1 2 15325 15334
0 15336 5 1 1 15335
0 15337 7 1 2 76207 15336
0 15338 5 1 1 15337
0 15339 7 2 2 72033 89349
0 15340 7 1 2 87735 95809
0 15341 5 1 1 15340
0 15342 7 1 2 89325 15341
0 15343 5 2 1 15342
0 15344 7 2 2 86209 93342
0 15345 5 1 1 95813
0 15346 7 5 2 65363 90582
0 15347 7 1 2 88915 94812
0 15348 7 1 2 95815 15347
0 15349 7 1 2 95814 15348
0 15350 7 1 2 95811 15349
0 15351 5 1 1 15350
0 15352 7 1 2 15338 15351
0 15353 5 1 1 15352
0 15354 7 1 2 83722 84524
0 15355 7 1 2 15353 15354
0 15356 5 1 1 15355
0 15357 7 1 2 15244 15356
0 15358 5 1 1 15357
0 15359 7 1 2 70779 15358
0 15360 5 1 1 15359
0 15361 7 2 2 90191 86477
0 15362 7 6 2 67086 92060
0 15363 7 1 2 78207 95822
0 15364 7 1 2 95820 15363
0 15365 5 2 1 15364
0 15366 7 1 2 90118 88185
0 15367 5 1 1 15366
0 15368 7 1 2 66692 90126
0 15369 5 1 1 15368
0 15370 7 1 2 15367 15369
0 15371 5 1 1 15370
0 15372 7 1 2 65364 15371
0 15373 5 1 1 15372
0 15374 7 1 2 89368 6781
0 15375 5 2 1 15374
0 15376 7 1 2 73035 95830
0 15377 5 1 1 15376
0 15378 7 1 2 15373 15377
0 15379 5 1 1 15378
0 15380 7 1 2 75273 15379
0 15381 5 1 1 15380
0 15382 7 3 2 76995 89350
0 15383 7 1 2 90052 95832
0 15384 5 1 1 15383
0 15385 7 1 2 15381 15384
0 15386 5 1 1 15385
0 15387 7 1 2 78208 15386
0 15388 5 1 1 15387
0 15389 7 1 2 65046 95821
0 15390 7 1 2 89907 15389
0 15391 5 1 1 15390
0 15392 7 1 2 15388 15391
0 15393 5 1 1 15392
0 15394 7 1 2 64666 15393
0 15395 5 1 1 15394
0 15396 7 1 2 95828 15395
0 15397 5 1 1 15396
0 15398 7 1 2 77986 15397
0 15399 5 1 1 15398
0 15400 7 1 2 66507 78016
0 15401 5 1 1 15400
0 15402 7 1 2 86641 15401
0 15403 5 1 1 15402
0 15404 7 1 2 65047 15403
0 15405 5 1 1 15404
0 15406 7 1 2 82045 93877
0 15407 5 1 1 15406
0 15408 7 1 2 15405 15407
0 15409 5 1 1 15408
0 15410 7 1 2 85118 15409
0 15411 5 1 1 15410
0 15412 7 1 2 94729 78209
0 15413 5 1 1 15412
0 15414 7 2 2 71924 86566
0 15415 7 1 2 68815 86528
0 15416 7 1 2 95835 15415
0 15417 5 1 1 15416
0 15418 7 1 2 91027 15417
0 15419 5 1 1 15418
0 15420 7 1 2 73423 15419
0 15421 5 1 1 15420
0 15422 7 1 2 15413 15421
0 15423 7 1 2 15411 15422
0 15424 5 1 1 15423
0 15425 7 1 2 69464 15424
0 15426 5 1 1 15425
0 15427 7 1 2 75645 86961
0 15428 5 1 1 15427
0 15429 7 2 2 80586 83347
0 15430 5 1 1 95837
0 15431 7 1 2 74847 95838
0 15432 5 1 1 15431
0 15433 7 1 2 94185 81372
0 15434 5 1 1 15433
0 15435 7 1 2 15432 15434
0 15436 7 1 2 15428 15435
0 15437 5 1 1 15436
0 15438 7 1 2 78210 15437
0 15439 5 1 1 15438
0 15440 7 1 2 15426 15439
0 15441 5 1 1 15440
0 15442 7 1 2 64667 15441
0 15443 5 1 1 15442
0 15444 7 3 2 81208 85119
0 15445 5 1 1 95839
0 15446 7 1 2 89373 95840
0 15447 5 1 1 15446
0 15448 7 4 2 73036 76646
0 15449 5 2 1 95842
0 15450 7 3 2 81711 90997
0 15451 5 1 1 95848
0 15452 7 1 2 95843 95849
0 15453 5 1 1 15452
0 15454 7 1 2 15447 15453
0 15455 5 1 1 15454
0 15456 7 1 2 68622 15455
0 15457 5 1 1 15456
0 15458 7 2 2 81848 78162
0 15459 7 2 2 72034 95851
0 15460 5 2 1 95853
0 15461 7 1 2 83025 90065
0 15462 5 1 1 15461
0 15463 7 1 2 95855 15462
0 15464 5 1 1 15463
0 15465 7 1 2 81209 15464
0 15466 5 1 1 15465
0 15467 7 1 2 15457 15466
0 15468 5 1 1 15467
0 15469 7 1 2 68350 15468
0 15470 5 1 1 15469
0 15471 7 1 2 83520 89854
0 15472 5 1 1 15471
0 15473 7 1 2 89774 15472
0 15474 5 1 1 15473
0 15475 7 1 2 87387 14430
0 15476 7 3 2 78064 15475
0 15477 7 1 2 93878 95857
0 15478 5 1 1 15477
0 15479 7 1 2 65365 86730
0 15480 5 1 1 15479
0 15481 7 2 2 66508 87996
0 15482 7 1 2 95860 86735
0 15483 7 1 2 15480 15482
0 15484 5 1 1 15483
0 15485 7 1 2 15478 15484
0 15486 5 1 1 15485
0 15487 7 1 2 85120 15486
0 15488 5 1 1 15487
0 15489 7 1 2 15474 15488
0 15490 7 1 2 15470 15489
0 15491 7 1 2 15443 15490
0 15492 5 1 1 15491
0 15493 7 1 2 88553 15492
0 15494 5 1 1 15493
0 15495 7 1 2 79422 83797
0 15496 5 1 1 15495
0 15497 7 1 2 79051 78163
0 15498 7 1 2 15496 15497
0 15499 5 1 1 15498
0 15500 7 3 2 69465 73960
0 15501 5 1 1 95862
0 15502 7 1 2 82739 95863
0 15503 5 1 1 15502
0 15504 7 2 2 64668 83542
0 15505 5 1 1 95865
0 15506 7 1 2 87147 95866
0 15507 5 1 1 15506
0 15508 7 1 2 15503 15507
0 15509 5 1 1 15508
0 15510 7 1 2 85121 15509
0 15511 5 1 1 15510
0 15512 7 1 2 65366 15511
0 15513 7 1 2 15499 15512
0 15514 5 1 1 15513
0 15515 7 2 2 93383 78164
0 15516 5 3 1 95867
0 15517 7 1 2 77110 85122
0 15518 5 1 1 15517
0 15519 7 1 2 95869 15518
0 15520 5 1 1 15519
0 15521 7 1 2 75603 15520
0 15522 5 1 1 15521
0 15523 7 1 2 15445 15522
0 15524 5 1 1 15523
0 15525 7 1 2 68351 15524
0 15526 5 1 1 15525
0 15527 7 1 2 73424 74493
0 15528 5 1 1 15527
0 15529 7 1 2 81220 15528
0 15530 5 1 1 15529
0 15531 7 1 2 78211 15530
0 15532 5 1 1 15531
0 15533 7 1 2 70393 15532
0 15534 7 1 2 15526 15533
0 15535 5 1 1 15534
0 15536 7 1 2 15514 15535
0 15537 5 1 1 15536
0 15538 7 2 2 68816 80019
0 15539 7 1 2 95229 95872
0 15540 5 1 1 15539
0 15541 7 1 2 15537 15540
0 15542 5 1 1 15541
0 15543 7 1 2 71798 15542
0 15544 5 1 1 15543
0 15545 7 1 2 64337 87845
0 15546 5 4 1 15545
0 15547 7 1 2 83698 95874
0 15548 5 1 1 15547
0 15549 7 1 2 67991 80848
0 15550 5 1 1 15549
0 15551 7 1 2 64338 15550
0 15552 5 1 1 15551
0 15553 7 1 2 84128 15552
0 15554 5 1 1 15553
0 15555 7 1 2 15548 15554
0 15556 5 1 1 15555
0 15557 7 1 2 73425 15556
0 15558 5 1 1 15557
0 15559 7 1 2 75129 94259
0 15560 5 1 1 15559
0 15561 7 1 2 86910 15560
0 15562 5 1 1 15561
0 15563 7 1 2 69466 15562
0 15564 5 1 1 15563
0 15565 7 1 2 15558 15564
0 15566 5 1 1 15565
0 15567 7 1 2 64669 15566
0 15568 5 1 1 15567
0 15569 7 2 2 69467 74736
0 15570 5 1 1 95878
0 15571 7 3 2 75103 87509
0 15572 5 2 1 95880
0 15573 7 1 2 95879 95881
0 15574 5 1 1 15573
0 15575 7 1 2 15568 15574
0 15576 5 1 1 15575
0 15577 7 1 2 85123 15576
0 15578 5 1 1 15577
0 15579 7 1 2 66693 90090
0 15580 5 1 1 15579
0 15581 7 1 2 82128 15580
0 15582 5 1 1 15581
0 15583 7 1 2 65367 15582
0 15584 5 1 1 15583
0 15585 7 1 2 66509 86193
0 15586 5 1 1 15585
0 15587 7 1 2 64670 75130
0 15588 5 1 1 15587
0 15589 7 1 2 15586 15588
0 15590 7 1 2 15584 15589
0 15591 5 1 1 15590
0 15592 7 1 2 91103 15591
0 15593 5 1 1 15592
0 15594 7 1 2 80683 79344
0 15595 7 1 2 80227 15594
0 15596 7 1 2 93937 15595
0 15597 5 1 1 15596
0 15598 7 1 2 80039 15597
0 15599 5 1 1 15598
0 15600 7 1 2 78212 15599
0 15601 5 1 1 15600
0 15602 7 1 2 15593 15601
0 15603 5 1 1 15602
0 15604 7 1 2 73037 15603
0 15605 5 1 1 15604
0 15606 7 1 2 78213 87854
0 15607 5 1 1 15606
0 15608 7 1 2 94395 75743
0 15609 7 1 2 81354 15608
0 15610 5 1 1 15609
0 15611 7 1 2 15607 15610
0 15612 5 1 1 15611
0 15613 7 1 2 80684 15612
0 15614 5 1 1 15613
0 15615 7 1 2 89612 95158
0 15616 5 1 1 15615
0 15617 7 1 2 15614 15616
0 15618 7 1 2 15605 15617
0 15619 7 1 2 15578 15618
0 15620 7 1 2 15544 15619
0 15621 5 1 1 15620
0 15622 7 1 2 88186 15621
0 15623 5 1 1 15622
0 15624 7 1 2 15494 15623
0 15625 5 1 1 15624
0 15626 7 1 2 65755 15625
0 15627 5 1 1 15626
0 15628 7 1 2 15399 15627
0 15629 5 1 1 15628
0 15630 7 1 2 66232 15629
0 15631 5 1 1 15630
0 15632 7 1 2 81433 83577
0 15633 5 1 1 15632
0 15634 7 7 2 67992 80685
0 15635 5 1 1 95885
0 15636 7 1 2 83483 15635
0 15637 5 1 1 15636
0 15638 7 1 2 76305 15637
0 15639 5 1 1 15638
0 15640 7 1 2 15633 15639
0 15641 5 1 1 15640
0 15642 7 1 2 88187 15641
0 15643 5 1 1 15642
0 15644 7 1 2 87096 87219
0 15645 7 1 2 84924 15644
0 15646 5 1 1 15645
0 15647 7 1 2 73038 95096
0 15648 5 1 1 15647
0 15649 7 1 2 68352 15648
0 15650 7 1 2 15646 15649
0 15651 5 1 1 15650
0 15652 7 1 2 89965 15651
0 15653 5 1 1 15652
0 15654 7 1 2 88554 15653
0 15655 5 1 1 15654
0 15656 7 1 2 15643 15655
0 15657 5 1 1 15656
0 15658 7 1 2 78214 15657
0 15659 5 1 1 15658
0 15660 7 3 2 71336 79899
0 15661 5 2 1 95892
0 15662 7 1 2 86766 95893
0 15663 5 2 1 15662
0 15664 7 1 2 95897 86629
0 15665 5 1 1 15664
0 15666 7 1 2 76306 15665
0 15667 5 1 1 15666
0 15668 7 1 2 83529 86307
0 15669 5 3 1 15668
0 15670 7 1 2 87331 76348
0 15671 5 1 1 15670
0 15672 7 1 2 82966 75073
0 15673 5 1 1 15672
0 15674 7 1 2 15671 15673
0 15675 5 1 1 15674
0 15676 7 1 2 65368 15675
0 15677 5 1 1 15676
0 15678 7 1 2 95899 15677
0 15679 5 1 1 15678
0 15680 7 1 2 67993 15679
0 15681 5 1 1 15680
0 15682 7 1 2 15667 15681
0 15683 5 1 1 15682
0 15684 7 1 2 88188 15683
0 15685 5 1 1 15684
0 15686 7 1 2 75561 78800
0 15687 5 3 1 15686
0 15688 7 1 2 79206 93302
0 15689 5 1 1 15688
0 15690 7 1 2 95902 15689
0 15691 5 1 1 15690
0 15692 7 1 2 82906 15691
0 15693 5 1 1 15692
0 15694 7 3 2 71612 83471
0 15695 7 1 2 75131 95905
0 15696 5 1 1 15695
0 15697 7 1 2 86731 15696
0 15698 5 1 1 15697
0 15699 7 1 2 86583 15698
0 15700 5 1 1 15699
0 15701 7 4 2 75363 74775
0 15702 5 3 1 95908
0 15703 7 1 2 76307 95909
0 15704 5 1 1 15703
0 15705 7 1 2 92945 15704
0 15706 5 1 1 15705
0 15707 7 1 2 86046 15706
0 15708 5 1 1 15707
0 15709 7 1 2 15700 15708
0 15710 7 1 2 15693 15709
0 15711 5 1 1 15710
0 15712 7 1 2 88555 15711
0 15713 5 1 1 15712
0 15714 7 1 2 15685 15713
0 15715 5 1 1 15714
0 15716 7 1 2 90066 15715
0 15717 5 1 1 15716
0 15718 7 1 2 15659 15717
0 15719 5 1 1 15718
0 15720 7 1 2 65756 15719
0 15721 5 1 1 15720
0 15722 7 3 2 82410 83599
0 15723 5 1 1 95915
0 15724 7 2 2 66510 74167
0 15725 7 1 2 95538 95918
0 15726 5 1 1 15725
0 15727 7 1 2 15723 15726
0 15728 5 1 1 15727
0 15729 7 2 2 82761 92234
0 15730 7 1 2 77028 95920
0 15731 7 1 2 15728 15730
0 15732 5 1 1 15731
0 15733 7 1 2 15721 15732
0 15734 5 1 1 15733
0 15735 7 1 2 64339 15734
0 15736 5 1 1 15735
0 15737 7 2 2 64671 82967
0 15738 5 1 1 95922
0 15739 7 1 2 86738 15738
0 15740 5 1 1 15739
0 15741 7 1 2 88189 15740
0 15742 5 1 1 15741
0 15743 7 1 2 78801 94048
0 15744 5 1 1 15743
0 15745 7 1 2 15742 15744
0 15746 5 1 1 15745
0 15747 7 1 2 65369 15746
0 15748 5 1 1 15747
0 15749 7 1 2 89139 89351
0 15750 5 2 1 15749
0 15751 7 1 2 77829 93898
0 15752 5 1 1 15751
0 15753 7 1 2 95924 15752
0 15754 5 2 1 15753
0 15755 7 1 2 64672 95926
0 15756 5 1 1 15755
0 15757 7 1 2 15748 15756
0 15758 5 1 1 15757
0 15759 7 1 2 66511 15758
0 15760 5 1 1 15759
0 15761 7 1 2 89629 94734
0 15762 7 1 2 83174 15761
0 15763 5 1 1 15762
0 15764 7 1 2 15760 15763
0 15765 5 1 1 15764
0 15766 7 1 2 85124 15765
0 15767 5 1 1 15766
0 15768 7 1 2 79447 94454
0 15769 5 1 1 15768
0 15770 7 1 2 15767 15769
0 15771 5 1 1 15770
0 15772 7 1 2 73039 15771
0 15773 5 1 1 15772
0 15774 7 2 2 86490 86426
0 15775 7 1 2 89995 90178
0 15776 5 1 1 15775
0 15777 7 2 2 95166 15776
0 15778 7 1 2 95928 95930
0 15779 5 1 1 15778
0 15780 7 1 2 15773 15779
0 15781 5 1 1 15780
0 15782 7 1 2 93053 15781
0 15783 5 1 1 15782
0 15784 7 1 2 15736 15783
0 15785 7 1 2 15631 15784
0 15786 5 1 1 15785
0 15787 7 1 2 65960 15786
0 15788 5 1 1 15787
0 15789 7 5 2 76382 94641
0 15790 5 1 1 95932
0 15791 7 2 2 81849 92699
0 15792 5 1 1 95937
0 15793 7 1 2 95933 95938
0 15794 5 1 1 15793
0 15795 7 5 2 66694 75744
0 15796 7 4 2 87736 95939
0 15797 7 2 2 70394 82105
0 15798 7 1 2 83956 95948
0 15799 7 1 2 95944 15798
0 15800 5 1 1 15799
0 15801 7 1 2 15794 15800
0 15802 5 1 1 15801
0 15803 7 1 2 81210 15802
0 15804 5 1 1 15803
0 15805 7 2 2 81587 95833
0 15806 7 1 2 83182 95950
0 15807 7 1 2 95945 15806
0 15808 5 1 1 15807
0 15809 7 1 2 15804 15808
0 15810 5 1 1 15809
0 15811 7 1 2 64673 15810
0 15812 5 1 1 15811
0 15813 7 2 2 71799 77660
0 15814 5 1 1 95952
0 15815 7 1 2 80893 95953
0 15816 7 4 2 63768 91152
0 15817 7 1 2 79351 95954
0 15818 7 1 2 15815 15817
0 15819 5 1 1 15818
0 15820 7 1 2 15812 15819
0 15821 5 1 1 15820
0 15822 7 1 2 66233 15821
0 15823 5 1 1 15822
0 15824 7 2 2 76571 82968
0 15825 7 1 2 73961 95958
0 15826 5 1 1 15825
0 15827 7 3 2 73716 88705
0 15828 7 1 2 78692 95960
0 15829 5 1 1 15828
0 15830 7 1 2 15826 15829
0 15831 5 1 1 15830
0 15832 7 1 2 93189 15831
0 15833 5 1 1 15832
0 15834 7 3 2 65048 82969
0 15835 5 1 1 95963
0 15836 7 1 2 95964 89649
0 15837 5 1 1 15836
0 15838 7 1 2 82907 79896
0 15839 7 1 2 93228 15838
0 15840 7 1 2 90182 15839
0 15841 5 1 1 15840
0 15842 7 1 2 15837 15841
0 15843 5 1 1 15842
0 15844 7 1 2 78641 15843
0 15845 5 1 1 15844
0 15846 7 1 2 15833 15845
0 15847 5 1 1 15846
0 15848 7 1 2 85125 15847
0 15849 5 1 1 15848
0 15850 7 1 2 86344 94745
0 15851 5 1 1 15850
0 15852 7 1 2 69468 15851
0 15853 5 1 1 15852
0 15854 7 1 2 88190 15853
0 15855 5 1 1 15854
0 15856 7 3 2 83619 84595
0 15857 5 1 1 95966
0 15858 7 1 2 15855 15857
0 15859 5 1 1 15858
0 15860 7 1 2 76572 15859
0 15861 5 1 1 15860
0 15862 7 1 2 95792 88191
0 15863 5 1 1 15862
0 15864 7 1 2 84596 92047
0 15865 5 1 1 15864
0 15866 7 1 2 15863 15865
0 15867 5 1 1 15866
0 15868 7 1 2 76208 15867
0 15869 5 1 1 15868
0 15870 7 1 2 15861 15869
0 15871 5 1 1 15870
0 15872 7 1 2 78215 15871
0 15873 5 1 1 15872
0 15874 7 1 2 15849 15873
0 15875 5 1 1 15874
0 15876 7 1 2 65370 15875
0 15877 5 1 1 15876
0 15878 7 1 2 91050 95927
0 15879 5 1 1 15878
0 15880 7 7 2 63886 94799
0 15881 5 2 1 95969
0 15882 7 1 2 89830 95976
0 15883 5 1 1 15882
0 15884 7 1 2 78216 15883
0 15885 5 1 1 15884
0 15886 7 1 2 15879 15885
0 15887 5 1 1 15886
0 15888 7 1 2 76573 15887
0 15889 5 1 1 15888
0 15890 7 2 2 78217 89295
0 15891 5 1 1 95978
0 15892 7 1 2 76209 95979
0 15893 5 1 1 15892
0 15894 7 1 2 15889 15893
0 15895 5 1 1 15894
0 15896 7 1 2 64340 15895
0 15897 5 1 1 15896
0 15898 7 2 2 76210 84570
0 15899 7 1 2 95980 90662
0 15900 7 1 2 95831 15899
0 15901 5 1 1 15900
0 15902 7 1 2 15897 15901
0 15903 7 1 2 15877 15902
0 15904 5 1 1 15903
0 15905 7 1 2 73040 15904
0 15906 5 1 1 15905
0 15907 7 1 2 79075 88809
0 15908 5 1 1 15907
0 15909 7 1 2 88192 15908
0 15910 5 1 1 15909
0 15911 7 1 2 88457 90172
0 15912 5 1 1 15911
0 15913 7 1 2 15910 15912
0 15914 5 1 1 15913
0 15915 7 1 2 66695 15914
0 15916 5 1 1 15915
0 15917 7 1 2 82970 94463
0 15918 5 1 1 15917
0 15919 7 1 2 13085 95925
0 15920 7 1 2 15918 15919
0 15921 5 1 1 15920
0 15922 7 1 2 66234 15921
0 15923 5 1 1 15922
0 15924 7 1 2 15916 15923
0 15925 5 1 1 15924
0 15926 7 1 2 66512 15925
0 15927 5 1 1 15926
0 15928 7 1 2 88193 86875
0 15929 5 1 1 15928
0 15930 7 1 2 86637 90173
0 15931 5 1 1 15930
0 15932 7 1 2 15929 15931
0 15933 5 1 1 15932
0 15934 7 1 2 66235 15933
0 15935 5 1 1 15934
0 15936 7 1 2 15927 15935
0 15937 5 1 1 15936
0 15938 7 1 2 64674 15937
0 15939 5 1 1 15938
0 15940 7 1 2 89938 95931
0 15941 5 1 1 15940
0 15942 7 1 2 15939 15941
0 15943 5 1 1 15942
0 15944 7 1 2 79119 15943
0 15945 5 1 1 15944
0 15946 7 1 2 89638 95191
0 15947 7 1 2 89625 15946
0 15948 5 1 1 15947
0 15949 7 1 2 15945 15948
0 15950 7 1 2 15906 15949
0 15951 5 1 1 15950
0 15952 7 1 2 71038 15951
0 15953 5 1 1 15952
0 15954 7 1 2 15823 15953
0 15955 5 1 1 15954
0 15956 7 1 2 65757 15955
0 15957 5 1 1 15956
0 15958 7 1 2 15788 15957
0 15959 5 1 1 15958
0 15960 7 1 2 72612 15959
0 15961 5 1 1 15960
0 15962 7 1 2 85126 79308
0 15963 5 1 1 15962
0 15964 7 1 2 15790 15963
0 15965 5 1 1 15964
0 15966 7 1 2 65049 15965
0 15967 5 1 1 15966
0 15968 7 3 2 76574 78218
0 15969 5 1 1 95982
0 15970 7 1 2 95100 85127
0 15971 5 1 1 15970
0 15972 7 1 2 15969 15971
0 15973 7 1 2 15967 15972
0 15974 5 1 1 15973
0 15975 7 1 2 82543 92614
0 15976 7 1 2 15974 15975
0 15977 5 1 1 15976
0 15978 7 1 2 95426 82544
0 15979 5 1 1 15978
0 15980 7 1 2 93117 94821
0 15981 5 1 1 15980
0 15982 7 1 2 15979 15981
0 15983 5 2 1 15982
0 15984 7 3 2 83215 85100
0 15985 5 1 1 95987
0 15986 7 1 2 91028 15985
0 15987 5 1 1 15986
0 15988 7 1 2 88194 15987
0 15989 7 1 2 95985 15988
0 15990 5 1 1 15989
0 15991 7 1 2 15977 15990
0 15992 5 1 1 15991
0 15993 7 1 2 73041 15992
0 15994 5 1 1 15993
0 15995 7 1 2 95401 83923
0 15996 5 1 1 15995
0 15997 7 1 2 92615 15996
0 15998 5 1 1 15997
0 15999 7 2 2 86695 85001
0 16000 5 1 1 95990
0 16001 7 1 2 95399 16000
0 16002 5 1 1 16001
0 16003 7 1 2 88195 16002
0 16004 5 1 1 16003
0 16005 7 1 2 15998 16004
0 16006 5 1 1 16005
0 16007 7 1 2 73426 16006
0 16008 5 1 1 16007
0 16009 7 1 2 84027 93171
0 16010 5 1 1 16009
0 16011 7 1 2 16008 16010
0 16012 5 1 1 16011
0 16013 7 1 2 85128 16012
0 16014 5 1 1 16013
0 16015 7 2 2 76902 95397
0 16016 7 1 2 65371 79371
0 16017 7 1 2 95992 16016
0 16018 5 1 1 16017
0 16019 7 1 2 16014 16018
0 16020 5 1 1 16019
0 16021 7 1 2 65758 16020
0 16022 5 1 1 16021
0 16023 7 1 2 15994 16022
0 16024 5 1 1 16023
0 16025 7 1 2 64341 16024
0 16026 5 1 1 16025
0 16027 7 1 2 77599 89793
0 16028 5 1 1 16027
0 16029 7 1 2 83643 90550
0 16030 5 1 1 16029
0 16031 7 1 2 16028 16030
0 16032 5 1 1 16031
0 16033 7 1 2 76575 16032
0 16034 5 2 1 16033
0 16035 7 12 2 64675 65372
0 16036 5 1 1 95996
0 16037 7 2 2 95997 90029
0 16038 7 1 2 95454 96008
0 16039 5 1 1 16038
0 16040 7 1 2 95994 16039
0 16041 5 1 1 16040
0 16042 7 1 2 72613 16041
0 16043 5 1 1 16042
0 16044 7 2 2 84975 91998
0 16045 7 1 2 92255 88556
0 16046 7 1 2 96010 16045
0 16047 5 2 1 16046
0 16048 7 1 2 16043 96012
0 16049 5 1 1 16048
0 16050 7 1 2 93054 85129
0 16051 7 1 2 16049 16050
0 16052 5 1 1 16051
0 16053 7 1 2 16026 16052
0 16054 5 1 1 16053
0 16055 7 1 2 65961 16054
0 16056 5 1 1 16055
0 16057 7 3 2 68972 78309
0 16058 7 1 2 75057 78110
0 16059 7 1 2 96014 16058
0 16060 5 1 1 16059
0 16061 7 1 2 95995 16060
0 16062 5 1 1 16061
0 16063 7 1 2 72614 16062
0 16064 5 1 1 16063
0 16065 7 1 2 96013 16064
0 16066 5 1 1 16065
0 16067 7 1 2 64342 16066
0 16068 5 1 1 16067
0 16069 7 1 2 66236 91999
0 16070 7 7 2 72615 77661
0 16071 7 1 2 96017 89794
0 16072 7 1 2 16069 16071
0 16073 5 1 1 16072
0 16074 7 1 2 16068 16073
0 16075 5 1 1 16074
0 16076 7 1 2 85130 16075
0 16077 5 1 1 16076
0 16078 7 6 2 64676 75274
0 16079 5 1 1 96024
0 16080 7 1 2 95473 96025
0 16081 7 1 2 91038 16080
0 16082 5 1 1 16081
0 16083 7 1 2 16077 16082
0 16084 5 1 1 16083
0 16085 7 1 2 74058 16084
0 16086 5 1 1 16085
0 16087 7 1 2 16056 16086
0 16088 5 1 1 16087
0 16089 7 1 2 80401 16088
0 16090 5 1 1 16089
0 16091 7 7 2 66696 67600
0 16092 7 1 2 92110 89987
0 16093 5 1 1 16092
0 16094 7 1 2 64677 92708
0 16095 5 1 1 16094
0 16096 7 1 2 16093 16095
0 16097 5 1 1 16096
0 16098 7 1 2 96030 16097
0 16099 5 1 1 16098
0 16100 7 4 2 70395 85002
0 16101 5 1 1 96037
0 16102 7 1 2 94793 96038
0 16103 5 1 1 16102
0 16104 7 1 2 16099 16103
0 16105 5 1 1 16104
0 16106 7 1 2 73717 16105
0 16107 5 1 1 16106
0 16108 7 1 2 88196 95991
0 16109 5 1 1 16108
0 16110 7 1 2 83947 86718
0 16111 5 3 1 16110
0 16112 7 2 2 89691 89671
0 16113 7 1 2 96041 96044
0 16114 5 1 1 16113
0 16115 7 1 2 16109 16114
0 16116 5 1 1 16115
0 16117 7 1 2 73427 16116
0 16118 5 1 1 16117
0 16119 7 5 2 67994 91239
0 16120 7 1 2 65373 90266
0 16121 7 1 2 96046 16120
0 16122 5 1 1 16121
0 16123 7 1 2 75709 77015
0 16124 7 1 2 96042 16123
0 16125 5 1 1 16124
0 16126 7 1 2 16122 16125
0 16127 5 1 1 16126
0 16128 7 1 2 82971 16127
0 16129 5 1 1 16128
0 16130 7 2 2 74946 95307
0 16131 5 1 1 96051
0 16132 7 1 2 70396 96052
0 16133 5 1 1 16132
0 16134 7 1 2 92723 16133
0 16135 5 1 1 16134
0 16136 7 1 2 88197 16135
0 16137 5 1 1 16136
0 16138 7 1 2 16129 16137
0 16139 7 1 2 16118 16138
0 16140 7 1 2 16107 16139
0 16141 5 1 1 16140
0 16142 7 1 2 65962 16141
0 16143 5 1 1 16142
0 16144 7 2 2 92073 93906
0 16145 7 1 2 87881 85405
0 16146 7 1 2 96053 16145
0 16147 5 1 1 16146
0 16148 7 1 2 16143 16147
0 16149 5 1 1 16148
0 16150 7 1 2 64343 16149
0 16151 5 1 1 16150
0 16152 7 1 2 87909 93513
0 16153 7 1 2 96054 16152
0 16154 5 1 1 16153
0 16155 7 1 2 16151 16154
0 16156 5 1 1 16155
0 16157 7 1 2 85131 16156
0 16158 5 1 1 16157
0 16159 7 4 2 63769 64344
0 16160 7 2 2 86857 96055
0 16161 7 1 2 11761 11809
0 16162 5 1 1 16161
0 16163 7 1 2 76576 16162
0 16164 5 1 1 16163
0 16165 7 1 2 16164 5233
0 16166 5 1 1 16165
0 16167 7 1 2 67601 16166
0 16168 5 1 1 16167
0 16169 7 1 2 15792 5982
0 16170 5 1 1 16169
0 16171 7 1 2 85003 16170
0 16172 5 1 1 16171
0 16173 7 1 2 16168 16172
0 16174 5 1 1 16173
0 16175 7 1 2 96059 16174
0 16176 5 1 1 16175
0 16177 7 1 2 93907 89908
0 16178 5 1 1 16177
0 16179 7 1 2 15891 16178
0 16180 5 1 1 16179
0 16181 7 1 2 78434 16180
0 16182 5 1 1 16181
0 16183 7 1 2 72616 89897
0 16184 7 2 2 94951 16183
0 16185 7 1 2 89338 96061
0 16186 5 1 1 16185
0 16187 7 1 2 16182 16186
0 16188 5 1 1 16187
0 16189 7 1 2 64345 16188
0 16190 5 1 1 16189
0 16191 7 1 2 96062 90667
0 16192 5 1 1 16191
0 16193 7 1 2 16190 16192
0 16194 5 1 1 16193
0 16195 7 1 2 76577 16194
0 16196 5 1 1 16195
0 16197 7 3 2 85826 78165
0 16198 5 2 1 96063
0 16199 7 1 2 82167 85132
0 16200 5 1 1 16199
0 16201 7 1 2 96066 16200
0 16202 5 1 1 16201
0 16203 7 1 2 88557 16202
0 16204 5 1 1 16203
0 16205 7 1 2 90067 93960
0 16206 5 1 1 16205
0 16207 7 1 2 16204 16206
0 16208 5 1 1 16207
0 16209 7 4 2 64346 73718
0 16210 5 1 1 96068
0 16211 7 6 2 67602 84962
0 16212 5 1 1 96072
0 16213 7 1 2 96069 96073
0 16214 7 1 2 16208 16213
0 16215 5 1 1 16214
0 16216 7 1 2 16196 16215
0 16217 5 1 1 16216
0 16218 7 1 2 73042 16217
0 16219 5 1 1 16218
0 16220 7 1 2 16176 16219
0 16221 7 1 2 16158 16220
0 16222 5 1 1 16221
0 16223 7 1 2 65759 16222
0 16224 5 1 1 16223
0 16225 7 1 2 74059 95474
0 16226 5 1 1 16225
0 16227 7 9 2 70780 72617
0 16228 5 4 1 96078
0 16229 7 1 2 96087 82556
0 16230 5 2 1 16229
0 16231 7 1 2 77322 6005
0 16232 7 1 2 96091 16231
0 16233 5 1 1 16232
0 16234 7 1 2 16226 16233
0 16235 5 1 1 16234
0 16236 7 1 2 64678 16235
0 16237 5 1 1 16236
0 16238 7 3 2 77323 82545
0 16239 7 1 2 75007 96093
0 16240 5 1 1 16239
0 16241 7 1 2 16237 16240
0 16242 5 1 1 16241
0 16243 7 1 2 93869 16242
0 16244 5 1 1 16243
0 16245 7 2 2 67603 92803
0 16246 7 14 2 65963 95521
0 16247 7 1 2 96098 77500
0 16248 7 1 2 96096 16247
0 16249 5 1 1 16248
0 16250 7 1 2 16244 16249
0 16251 5 1 1 16250
0 16252 7 1 2 78219 16251
0 16253 5 1 1 16252
0 16254 7 1 2 76578 88198
0 16255 5 2 1 16254
0 16256 7 1 2 79195 89770
0 16257 5 1 1 16256
0 16258 7 1 2 96112 16257
0 16259 5 1 1 16258
0 16260 7 1 2 73043 16259
0 16261 5 1 1 16260
0 16262 7 1 2 77725 96009
0 16263 5 1 1 16262
0 16264 7 1 2 16261 16263
0 16265 5 1 1 16264
0 16266 7 1 2 96094 85133
0 16267 7 1 2 16265 16266
0 16268 5 1 1 16267
0 16269 7 1 2 16253 16268
0 16270 5 1 1 16269
0 16271 7 1 2 80402 16270
0 16272 5 1 1 16271
0 16273 7 3 2 87737 84436
0 16274 7 3 2 77324 82773
0 16275 7 1 2 96114 96117
0 16276 5 1 1 16275
0 16277 7 2 2 64347 77060
0 16278 5 4 1 96120
0 16279 7 2 2 69 96122
0 16280 5 2 1 96126
0 16281 7 1 2 96128 95961
0 16282 7 1 2 91492 16281
0 16283 5 1 1 16282
0 16284 7 1 2 16276 16283
0 16285 5 1 1 16284
0 16286 7 1 2 64679 16285
0 16287 5 1 1 16286
0 16288 7 1 2 87922 96099
0 16289 7 1 2 96115 16288
0 16290 5 1 1 16289
0 16291 7 1 2 16287 16290
0 16292 5 1 1 16291
0 16293 7 1 2 79821 16292
0 16294 5 1 1 16293
0 16295 7 1 2 89255 84976
0 16296 7 1 2 96079 16295
0 16297 7 5 2 67087 86399
0 16298 7 2 2 66961 81103
0 16299 7 1 2 96135 95003
0 16300 7 1 2 96130 16299
0 16301 7 1 2 16296 16300
0 16302 5 1 1 16301
0 16303 7 1 2 16294 16302
0 16304 5 1 1 16303
0 16305 7 1 2 73044 16304
0 16306 5 1 1 16305
0 16307 7 1 2 16272 16306
0 16308 7 1 2 16224 16307
0 16309 5 1 1 16308
0 16310 7 1 2 74638 16309
0 16311 5 1 1 16310
0 16312 7 1 2 67995 93873
0 16313 5 1 1 16312
0 16314 7 1 2 88199 16313
0 16315 5 2 1 16314
0 16316 7 1 2 94050 96137
0 16317 5 1 1 16316
0 16318 7 1 2 66237 16317
0 16319 5 1 1 16318
0 16320 7 2 2 64680 78017
0 16321 5 1 1 96139
0 16322 7 1 2 86739 16321
0 16323 5 1 1 16322
0 16324 7 1 2 90127 16323
0 16325 5 1 1 16324
0 16326 7 1 2 16319 16325
0 16327 5 1 1 16326
0 16328 7 1 2 66513 16327
0 16329 5 1 1 16328
0 16330 7 1 2 92053 86241
0 16331 5 1 1 16330
0 16332 7 1 2 16329 16331
0 16333 5 1 1 16332
0 16334 7 1 2 65050 16333
0 16335 5 1 1 16334
0 16336 7 1 2 86529 90030
0 16337 7 1 2 77025 16336
0 16338 5 1 1 16337
0 16339 7 1 2 16335 16338
0 16340 5 1 1 16339
0 16341 7 1 2 85134 16340
0 16342 5 1 1 16341
0 16343 7 2 2 86491 75745
0 16344 7 1 2 86732 13910
0 16345 5 1 1 16344
0 16346 7 1 2 88558 16345
0 16347 5 1 1 16346
0 16348 7 1 2 96138 16347
0 16349 5 1 1 16348
0 16350 7 1 2 96141 16349
0 16351 5 1 1 16350
0 16352 7 1 2 65374 90119
0 16353 5 3 1 16352
0 16354 7 1 2 69783 77687
0 16355 7 1 2 96143 16354
0 16356 5 1 1 16355
0 16357 7 1 2 91039 16356
0 16358 5 1 1 16357
0 16359 7 1 2 16351 16358
0 16360 5 1 1 16359
0 16361 7 1 2 79506 16360
0 16362 5 1 1 16361
0 16363 7 1 2 90998 90139
0 16364 5 1 1 16363
0 16365 7 2 2 87923 74239
0 16366 7 1 2 89934 96146
0 16367 7 1 2 89170 16366
0 16368 5 1 1 16367
0 16369 7 1 2 16364 16368
0 16370 5 1 1 16369
0 16371 7 1 2 82740 16370
0 16372 5 1 1 16371
0 16373 7 2 2 92061 84022
0 16374 5 2 1 96148
0 16375 7 1 2 64681 90128
0 16376 5 1 1 16375
0 16377 7 1 2 96150 16376
0 16378 5 1 1 16377
0 16379 7 1 2 66238 16378
0 16380 5 1 1 16379
0 16381 7 1 2 75604 93901
0 16382 5 1 1 16381
0 16383 7 1 2 16380 16382
0 16384 5 1 1 16383
0 16385 7 1 2 78220 16384
0 16386 5 1 1 16385
0 16387 7 1 2 16372 16386
0 16388 7 1 2 16362 16387
0 16389 7 1 2 16342 16388
0 16390 5 1 1 16389
0 16391 7 1 2 65964 16390
0 16392 5 1 1 16391
0 16393 7 1 2 90192 89898
0 16394 7 1 2 95160 16393
0 16395 7 1 2 90165 16394
0 16396 5 1 1 16395
0 16397 7 1 2 16392 16396
0 16398 5 1 1 16397
0 16399 7 1 2 64348 16398
0 16400 5 1 1 16399
0 16401 7 1 2 94143 90682
0 16402 7 1 2 94824 16401
0 16403 5 1 1 16402
0 16404 7 1 2 16400 16403
0 16405 5 1 1 16404
0 16406 7 1 2 82546 16405
0 16407 5 1 1 16406
0 16408 7 1 2 85135 95986
0 16409 5 1 1 16408
0 16410 7 4 2 74639 90999
0 16411 5 2 1 96152
0 16412 7 1 2 5851 96092
0 16413 7 1 2 96153 16412
0 16414 5 1 1 16413
0 16415 7 1 2 16409 16414
0 16416 5 1 1 16415
0 16417 7 1 2 77325 16416
0 16418 5 1 1 16417
0 16419 7 2 2 72618 96154
0 16420 7 3 2 64682 92408
0 16421 7 1 2 71039 96160
0 16422 7 1 2 96158 16421
0 16423 5 1 1 16422
0 16424 7 1 2 16418 16423
0 16425 5 1 1 16424
0 16426 7 1 2 89988 16425
0 16427 5 1 1 16426
0 16428 7 2 2 79372 74314
0 16429 7 3 2 67604 75819
0 16430 7 1 2 95522 96165
0 16431 7 1 2 96163 16430
0 16432 7 1 2 95427 16431
0 16433 5 1 1 16432
0 16434 7 1 2 16427 16433
0 16435 5 1 1 16434
0 16436 7 1 2 73045 16435
0 16437 5 1 1 16436
0 16438 7 1 2 79373 96100
0 16439 7 1 2 95993 16438
0 16440 5 1 1 16439
0 16441 7 1 2 16437 16440
0 16442 5 1 1 16441
0 16443 7 1 2 87637 16442
0 16444 5 1 1 16443
0 16445 7 1 2 64055 16444
0 16446 7 1 2 16407 16445
0 16447 7 1 2 16311 16446
0 16448 7 1 2 16090 16447
0 16449 7 1 2 15961 16448
0 16450 5 1 1 16449
0 16451 7 2 2 83723 95523
0 16452 7 4 2 68817 66697
0 16453 7 4 2 75746 96170
0 16454 7 1 2 95798 96174
0 16455 5 1 1 16454
0 16456 7 1 2 78166 95795
0 16457 5 1 1 16456
0 16458 7 1 2 16455 16457
0 16459 5 1 1 16458
0 16460 7 1 2 65375 16459
0 16461 5 1 1 16460
0 16462 7 1 2 96156 7797
0 16463 5 1 1 16462
0 16464 7 1 2 94757 16463
0 16465 5 1 1 16464
0 16466 7 2 2 66514 84571
0 16467 7 1 2 88831 76383
0 16468 7 1 2 96178 16467
0 16469 5 1 1 16468
0 16470 7 1 2 16465 16469
0 16471 7 1 2 16461 16470
0 16472 5 1 1 16471
0 16473 7 1 2 88200 16472
0 16474 5 1 1 16473
0 16475 7 1 2 74888 78221
0 16476 5 1 1 16475
0 16477 7 1 2 86805 85136
0 16478 5 1 1 16477
0 16479 7 1 2 16476 16478
0 16480 5 1 1 16479
0 16481 7 1 2 66698 16480
0 16482 5 1 1 16481
0 16483 7 1 2 78572 78222
0 16484 5 1 1 16483
0 16485 7 1 2 16482 16484
0 16486 5 1 1 16485
0 16487 7 1 2 75505 16486
0 16488 5 1 1 16487
0 16489 7 1 2 65051 86948
0 16490 7 1 2 83833 16489
0 16491 5 1 1 16490
0 16492 7 1 2 94300 16491
0 16493 5 1 1 16492
0 16494 7 1 2 91000 16493
0 16495 5 1 1 16494
0 16496 7 1 2 16488 16495
0 16497 5 1 1 16496
0 16498 7 1 2 88559 16497
0 16499 5 1 1 16498
0 16500 7 1 2 16474 16499
0 16501 5 1 1 16500
0 16502 7 1 2 73046 16501
0 16503 5 1 1 16502
0 16504 7 3 2 90104 81594
0 16505 5 1 1 96180
0 16506 7 1 2 96181 91040
0 16507 5 1 1 16506
0 16508 7 1 2 16503 16507
0 16509 5 1 1 16508
0 16510 7 1 2 66239 16509
0 16511 5 1 1 16510
0 16512 7 1 2 16511 95829
0 16513 5 1 1 16512
0 16514 7 1 2 64683 16513
0 16515 5 1 1 16514
0 16516 7 3 2 94030 76384
0 16517 7 1 2 66240 92062
0 16518 7 1 2 96183 16517
0 16519 7 1 2 95951 16518
0 16520 5 1 1 16519
0 16521 7 1 2 16515 16520
0 16522 5 1 1 16521
0 16523 7 1 2 96168 16522
0 16524 5 1 1 16523
0 16525 7 1 2 75770 89692
0 16526 5 1 1 16525
0 16527 7 1 2 76743 16526
0 16528 5 1 1 16527
0 16529 7 3 2 63770 16528
0 16530 5 2 1 96186
0 16531 7 1 2 94623 89921
0 16532 5 1 1 16531
0 16533 7 1 2 96189 16532
0 16534 5 1 1 16533
0 16535 7 1 2 75132 16534
0 16536 5 1 1 16535
0 16537 7 1 2 82623 78223
0 16538 5 1 1 16537
0 16539 7 1 2 75886 90068
0 16540 5 1 1 16539
0 16541 7 1 2 16538 16540
0 16542 5 1 1 16541
0 16543 7 1 2 75880 16542
0 16544 5 1 1 16543
0 16545 7 3 2 79691 74452
0 16546 7 1 2 94618 96191
0 16547 5 1 1 16546
0 16548 7 1 2 16544 16547
0 16549 7 1 2 16536 16548
0 16550 5 1 1 16549
0 16551 7 1 2 67996 16550
0 16552 5 1 1 16551
0 16553 7 2 2 72141 74848
0 16554 7 6 2 63887 80587
0 16555 7 1 2 78224 96196
0 16556 7 1 2 96194 16555
0 16557 5 1 1 16556
0 16558 7 1 2 16552 16557
0 16559 5 1 1 16558
0 16560 7 1 2 71337 16559
0 16561 5 1 1 16560
0 16562 7 1 2 78167 84644
0 16563 7 1 2 76823 16562
0 16564 7 1 2 95631 16563
0 16565 5 1 1 16564
0 16566 7 1 2 16561 16565
0 16567 5 1 1 16566
0 16568 7 1 2 69784 16567
0 16569 5 1 1 16568
0 16570 7 1 2 94562 96197
0 16571 7 1 2 76909 16570
0 16572 5 1 1 16571
0 16573 7 1 2 16569 16572
0 16574 5 1 1 16573
0 16575 7 1 2 75364 16574
0 16576 5 1 1 16575
0 16577 7 1 2 95699 77636
0 16578 5 1 1 16577
0 16579 7 1 2 96190 16578
0 16580 5 1 1 16579
0 16581 7 1 2 68353 16580
0 16582 5 1 1 16581
0 16583 7 3 2 75747 89394
0 16584 7 1 2 94624 96202
0 16585 5 1 1 16584
0 16586 7 1 2 16582 16585
0 16587 5 1 1 16586
0 16588 7 1 2 81610 16587
0 16589 5 1 1 16588
0 16590 7 1 2 75562 81282
0 16591 7 1 2 96187 16590
0 16592 5 1 1 16591
0 16593 7 1 2 16589 16592
0 16594 5 1 1 16593
0 16595 7 1 2 69785 16594
0 16596 5 1 1 16595
0 16597 7 1 2 95750 96188
0 16598 5 1 1 16597
0 16599 7 1 2 16596 16598
0 16600 5 1 1 16599
0 16601 7 1 2 75133 16600
0 16602 5 1 1 16601
0 16603 7 1 2 75008 75890
0 16604 5 1 1 16603
0 16605 7 1 2 91046 16604
0 16606 5 1 1 16605
0 16607 7 3 2 68623 81434
0 16608 7 1 2 75690 96205
0 16609 5 1 1 16608
0 16610 7 1 2 16606 16609
0 16611 5 1 1 16610
0 16612 7 1 2 69786 16611
0 16613 5 1 1 16612
0 16614 7 1 2 83209 76754
0 16615 5 1 1 16614
0 16616 7 1 2 16613 16615
0 16617 5 1 1 16616
0 16618 7 1 2 74120 16617
0 16619 5 1 1 16618
0 16620 7 1 2 77788 90799
0 16621 5 1 1 16620
0 16622 7 1 2 16619 16621
0 16623 5 1 1 16622
0 16624 7 1 2 63771 16623
0 16625 5 1 1 16624
0 16626 7 1 2 16602 16625
0 16627 7 1 2 16576 16626
0 16628 5 1 1 16627
0 16629 7 1 2 95366 78476
0 16630 7 1 2 16628 16629
0 16631 5 1 1 16630
0 16632 7 1 2 69120 16631
0 16633 7 1 2 16524 16632
0 16634 5 1 1 16633
0 16635 7 1 2 16634 89572
0 16636 7 1 2 16450 16635
0 16637 5 1 1 16636
0 16638 7 3 2 67605 82423
0 16639 5 1 1 96208
0 16640 7 2 2 95679 88981
0 16641 7 1 2 89395 96211
0 16642 5 1 1 16641
0 16643 7 1 2 76844 91362
0 16644 5 1 1 16643
0 16645 7 2 2 88053 91515
0 16646 7 1 2 95734 96213
0 16647 5 1 1 16646
0 16648 7 1 2 16644 16647
0 16649 5 1 1 16648
0 16650 7 1 2 63772 79805
0 16651 7 1 2 16649 16650
0 16652 5 1 1 16651
0 16653 7 1 2 16642 16652
0 16654 5 1 1 16653
0 16655 7 1 2 71338 16654
0 16656 5 1 1 16655
0 16657 7 2 2 90314 76009
0 16658 7 3 2 70397 79374
0 16659 7 1 2 96217 76401
0 16660 7 1 2 96215 16659
0 16661 5 1 1 16660
0 16662 7 1 2 16656 16661
0 16663 5 1 1 16662
0 16664 7 1 2 69787 16663
0 16665 5 1 1 16664
0 16666 7 1 2 94417 96218
0 16667 7 1 2 95662 16666
0 16668 5 1 1 16667
0 16669 7 1 2 16665 16668
0 16670 5 1 1 16669
0 16671 7 1 2 75365 16670
0 16672 5 1 1 16671
0 16673 7 1 2 86116 95669
0 16674 5 1 1 16673
0 16675 7 1 2 76647 95670
0 16676 5 1 1 16675
0 16677 7 2 2 94342 90974
0 16678 7 1 2 87407 96220
0 16679 5 1 1 16678
0 16680 7 1 2 16676 16679
0 16681 5 1 1 16680
0 16682 7 1 2 75968 16681
0 16683 5 1 1 16682
0 16684 7 1 2 75009 86848
0 16685 5 1 1 16684
0 16686 7 1 2 95671 16685
0 16687 5 1 1 16686
0 16688 7 6 2 71925 77746
0 16689 7 1 2 76648 95675
0 16690 7 1 2 96222 16689
0 16691 5 1 1 16690
0 16692 7 1 2 16687 16691
0 16693 7 1 2 16683 16692
0 16694 5 1 1 16693
0 16695 7 1 2 79806 16694
0 16696 5 1 1 16695
0 16697 7 1 2 16674 16696
0 16698 5 1 1 16697
0 16699 7 1 2 16698 90751
0 16700 5 1 1 16699
0 16701 7 1 2 72035 94673
0 16702 7 1 2 87762 91663
0 16703 7 1 2 92019 16702
0 16704 7 1 2 16701 16703
0 16705 5 1 1 16704
0 16706 7 1 2 16700 16705
0 16707 7 1 2 16672 16706
0 16708 5 1 1 16707
0 16709 7 1 2 71040 16708
0 16710 5 1 1 16709
0 16711 7 2 2 65629 95755
0 16712 7 2 2 91828 74240
0 16713 7 1 2 75563 92026
0 16714 7 1 2 96230 16713
0 16715 7 1 2 96228 16714
0 16716 5 1 1 16715
0 16717 7 1 2 16710 16716
0 16718 5 1 1 16717
0 16719 7 1 2 69469 16718
0 16720 5 1 1 16719
0 16721 7 2 2 89273 76933
0 16722 5 1 1 96232
0 16723 7 1 2 77769 90606
0 16724 7 1 2 96233 16723
0 16725 7 1 2 96229 16724
0 16726 5 1 1 16725
0 16727 7 1 2 16720 16726
0 16728 5 1 1 16727
0 16729 7 1 2 96209 16728
0 16730 5 1 1 16729
0 16731 7 1 2 74920 91281
0 16732 7 1 2 93637 16731
0 16733 7 4 2 87984 85415
0 16734 7 1 2 92434 96234
0 16735 7 1 2 82156 94099
0 16736 7 1 2 16734 16735
0 16737 7 1 2 16732 16736
0 16738 5 1 1 16737
0 16739 7 1 2 16730 16738
0 16740 5 1 1 16739
0 16741 7 1 2 82972 16740
0 16742 5 1 1 16741
0 16743 7 1 2 88560 94253
0 16744 5 1 1 16743
0 16745 7 1 2 88201 94165
0 16746 5 1 1 16745
0 16747 7 1 2 16744 16746
0 16748 5 1 1 16747
0 16749 7 1 2 73047 16748
0 16750 5 1 1 16749
0 16751 7 1 2 92038 87591
0 16752 5 1 1 16751
0 16753 7 1 2 16750 16752
0 16754 5 1 1 16753
0 16755 7 1 2 68354 16754
0 16756 5 1 1 16755
0 16757 7 1 2 86598 88561
0 16758 5 1 1 16757
0 16759 7 1 2 74640 89989
0 16760 5 1 1 16759
0 16761 7 1 2 16758 16760
0 16762 5 1 1 16761
0 16763 7 1 2 80403 16762
0 16764 5 1 1 16763
0 16765 7 1 2 93863 88202
0 16766 5 1 1 16765
0 16767 7 1 2 16764 16766
0 16768 5 1 1 16767
0 16769 7 1 2 73428 16768
0 16770 5 1 1 16769
0 16771 7 1 2 81595 95970
0 16772 5 1 1 16771
0 16773 7 1 2 16770 16772
0 16774 5 1 1 16773
0 16775 7 1 2 67997 16774
0 16776 5 1 1 16775
0 16777 7 1 2 16756 16776
0 16778 5 1 1 16777
0 16779 7 1 2 76211 16778
0 16780 5 1 1 16779
0 16781 7 2 2 88728 96149
0 16782 5 1 1 96238
0 16783 7 5 2 68355 76579
0 16784 7 2 2 73719 96240
0 16785 7 1 2 96239 96245
0 16786 5 1 1 16785
0 16787 7 1 2 16780 16786
0 16788 5 1 1 16787
0 16789 7 2 2 65965 90419
0 16790 7 1 2 72619 92510
0 16791 7 8 2 63972 64349
0 16792 7 1 2 93764 96249
0 16793 7 1 2 16790 16792
0 16794 7 1 2 96247 16793
0 16795 7 1 2 16788 16794
0 16796 5 1 1 16795
0 16797 7 1 2 16742 16796
0 16798 7 1 2 16637 16797
0 16799 7 1 2 15360 16798
0 16800 7 1 2 15024 16799
0 16801 7 1 2 13308 16800
0 16802 5 1 1 16801
0 16803 7 1 2 67252 16802
0 16804 5 1 1 16803
0 16805 7 1 2 81329 1618
0 16806 5 4 1 16805
0 16807 7 7 2 64056 72298
0 16808 5 1 1 96261
0 16809 7 15 2 65630 67088
0 16810 5 6 1 96268
0 16811 7 2 2 79657 96269
0 16812 7 4 2 73720 84666
0 16813 7 1 2 96289 96291
0 16814 5 1 1 16813
0 16815 7 10 2 70781 72142
0 16816 7 2 2 96295 93569
0 16817 7 1 2 88021 79101
0 16818 7 1 2 96305 16817
0 16819 5 1 1 16818
0 16820 7 1 2 16814 16819
0 16821 5 1 1 16820
0 16822 7 1 2 88916 16821
0 16823 5 1 1 16822
0 16824 7 2 2 92312 93472
0 16825 7 9 2 70623 65631
0 16826 5 1 1 96309
0 16827 7 1 2 91484 96310
0 16828 7 1 2 79008 16827
0 16829 7 1 2 96307 16828
0 16830 5 1 1 16829
0 16831 7 1 2 16823 16830
0 16832 5 1 1 16831
0 16833 7 1 2 80686 16832
0 16834 5 1 1 16833
0 16835 7 2 2 93668 92279
0 16836 7 1 2 91842 96318
0 16837 7 1 2 84695 16836
0 16838 5 1 1 16837
0 16839 7 1 2 16834 16838
0 16840 5 1 1 16839
0 16841 7 1 2 63888 16840
0 16842 5 1 1 16841
0 16843 7 1 2 80687 83620
0 16844 7 1 2 96306 16843
0 16845 7 1 2 90395 16844
0 16846 5 1 1 16845
0 16847 7 1 2 16842 16846
0 16848 5 1 1 16847
0 16849 7 1 2 66962 16848
0 16850 5 1 1 16849
0 16851 7 2 2 68973 73838
0 16852 5 1 1 96320
0 16853 7 1 2 8232 16852
0 16854 5 13 1 16853
0 16855 7 6 2 67089 96322
0 16856 7 4 2 72620 92304
0 16857 7 2 2 93593 87958
0 16858 7 1 2 88365 96345
0 16859 7 1 2 96341 16858
0 16860 7 1 2 96335 16859
0 16861 5 1 1 16860
0 16862 7 1 2 16850 16861
0 16863 5 1 1 16862
0 16864 7 1 2 73429 16863
0 16865 5 1 1 16864
0 16866 7 1 2 92305 95308
0 16867 7 1 2 78293 16866
0 16868 7 1 2 94956 16867
0 16869 7 1 2 96336 16868
0 16870 5 1 1 16869
0 16871 7 1 2 16865 16870
0 16872 5 1 1 16871
0 16873 7 1 2 67998 16872
0 16874 5 1 1 16873
0 16875 7 5 2 91270 89506
0 16876 5 1 1 96347
0 16877 7 1 2 65589 16876
0 16878 5 1 1 16877
0 16879 7 3 2 63889 73839
0 16880 5 1 1 96352
0 16881 7 3 2 90424 89543
0 16882 5 1 1 96355
0 16883 7 2 2 16880 16882
0 16884 5 22 1 96358
0 16885 7 1 2 70624 96359
0 16886 5 1 1 16885
0 16887 7 6 2 16878 16886
0 16888 7 1 2 68818 96382
0 16889 5 1 1 16888
0 16890 7 1 2 7917 16889
0 16891 5 3 1 16890
0 16892 7 2 2 72621 74241
0 16893 7 11 2 70782 71926
0 16894 7 1 2 80588 96393
0 16895 7 1 2 96391 16894
0 16896 7 1 2 96388 16895
0 16897 5 1 1 16896
0 16898 7 1 2 67606 92471
0 16899 5 2 1 16898
0 16900 7 9 2 71927 88022
0 16901 7 1 2 96406 84369
0 16902 7 2 2 96308 16901
0 16903 5 1 1 96415
0 16904 7 1 2 96404 16903
0 16905 5 1 1 16904
0 16906 7 1 2 63890 16905
0 16907 5 1 1 16906
0 16908 7 2 2 72622 73840
0 16909 7 1 2 92306 95628
0 16910 7 1 2 96417 16909
0 16911 5 1 1 16910
0 16912 7 1 2 16907 16911
0 16913 5 1 1 16912
0 16914 7 1 2 67090 85651
0 16915 7 1 2 16913 16914
0 16916 5 1 1 16915
0 16917 7 1 2 16897 16916
0 16918 5 1 1 16917
0 16919 7 1 2 95255 16918
0 16920 5 1 1 16919
0 16921 7 1 2 16874 16920
0 16922 5 1 1 16921
0 16923 7 1 2 74641 16922
0 16924 5 1 1 16923
0 16925 7 23 2 70666 72143
0 16926 5 1 1 96419
0 16927 7 7 2 70143 80688
0 16928 5 5 1 96442
0 16929 7 5 2 71613 80689
0 16930 5 1 1 96454
0 16931 7 5 2 96449 16930
0 16932 5 2 1 96459
0 16933 7 1 2 94947 96460
0 16934 5 2 1 16933
0 16935 7 1 2 96420 96466
0 16936 5 1 1 16935
0 16937 7 1 2 86777 96270
0 16938 5 1 1 16937
0 16939 7 1 2 16936 16938
0 16940 5 1 1 16939
0 16941 7 1 2 73048 16940
0 16942 5 1 1 16941
0 16943 7 2 2 68356 96271
0 16944 5 2 1 96468
0 16945 7 2 2 70667 77016
0 16946 5 2 1 96472
0 16947 7 1 2 96283 96474
0 16948 5 2 1 16947
0 16949 7 1 2 67999 96476
0 16950 5 1 1 16949
0 16951 7 1 2 96470 16950
0 16952 5 1 1 16951
0 16953 7 1 2 83061 16952
0 16954 5 1 1 16953
0 16955 7 1 2 16942 16954
0 16956 5 1 1 16955
0 16957 7 1 2 89507 16956
0 16958 5 1 1 16957
0 16959 7 1 2 77662 83062
0 16960 5 1 1 16959
0 16961 7 1 2 67091 86788
0 16962 7 3 2 16960 16961
0 16963 7 1 2 73817 96478
0 16964 5 1 1 16963
0 16965 7 1 2 16958 16964
0 16966 5 1 1 16965
0 16967 7 1 2 68974 16966
0 16968 5 1 1 16967
0 16969 7 1 2 91567 96479
0 16970 5 1 1 16969
0 16971 7 1 2 16968 16970
0 16972 5 1 1 16971
0 16973 7 1 2 66963 16972
0 16974 5 1 1 16973
0 16975 7 1 2 79003 16974
0 16976 5 1 1 16975
0 16977 7 5 2 72144 96360
0 16978 7 1 2 73049 96467
0 16979 5 1 1 16978
0 16980 7 1 2 85760 16979
0 16981 5 1 1 16980
0 16982 7 1 2 96481 16981
0 16983 5 1 1 16982
0 16984 7 4 2 89544 90287
0 16985 7 1 2 96486 96480
0 16986 5 1 1 16985
0 16987 7 1 2 66964 16986
0 16988 7 1 2 16983 16987
0 16989 5 1 1 16988
0 16990 7 1 2 87453 83120
0 16991 5 2 1 16990
0 16992 7 1 2 88424 96490
0 16993 5 1 1 16992
0 16994 7 1 2 73430 16993
0 16995 5 1 1 16994
0 16996 7 2 2 83808 96455
0 16997 5 2 1 96492
0 16998 7 1 2 86302 96494
0 16999 5 1 1 16998
0 17000 7 1 2 83348 16999
0 17001 5 1 1 17000
0 17002 7 1 2 16995 17001
0 17003 5 1 1 17002
0 17004 7 1 2 96337 17003
0 17005 5 1 1 17004
0 17006 7 1 2 73050 89723
0 17007 7 1 2 79313 17006
0 17008 7 1 2 91185 95949
0 17009 7 1 2 17007 17008
0 17010 5 1 1 17009
0 17011 7 1 2 72036 17010
0 17012 7 1 2 17005 17011
0 17013 5 1 1 17012
0 17014 7 1 2 68819 17013
0 17015 7 1 2 16989 17014
0 17016 5 1 1 17015
0 17017 7 1 2 74011 17016
0 17018 5 1 1 17017
0 17019 7 1 2 96080 79009
0 17020 7 1 2 17018 17019
0 17021 7 1 2 16976 17020
0 17022 5 1 1 17021
0 17023 7 1 2 64350 96416
0 17024 5 2 1 17023
0 17025 7 1 2 84667 92299
0 17026 5 1 1 17025
0 17027 7 1 2 96496 17026
0 17028 5 1 1 17027
0 17029 7 1 2 84823 17028
0 17030 5 1 1 17029
0 17031 7 1 2 83699 96081
0 17032 7 1 2 92484 17031
0 17033 5 1 1 17032
0 17034 7 1 2 17030 17033
0 17035 5 1 1 17034
0 17036 7 1 2 65052 17035
0 17037 5 1 1 17036
0 17038 7 4 2 70668 72037
0 17039 7 4 2 76802 96498
0 17040 7 1 2 70719 94859
0 17041 7 2 2 96502 17040
0 17042 7 9 2 69062 64351
0 17043 7 1 2 95288 96508
0 17044 7 1 2 92218 17043
0 17045 7 1 2 96506 17044
0 17046 5 1 1 17045
0 17047 7 1 2 17037 17046
0 17048 5 1 1 17047
0 17049 7 1 2 88562 17048
0 17050 5 1 1 17049
0 17051 7 1 2 84824 84785
0 17052 7 1 2 96292 17051
0 17053 5 1 1 17052
0 17054 7 5 2 64352 72038
0 17055 7 1 2 70783 95309
0 17056 7 1 2 96517 17055
0 17057 7 1 2 84504 77637
0 17058 7 1 2 17056 17057
0 17059 5 1 1 17058
0 17060 7 1 2 17053 17059
0 17061 5 1 1 17060
0 17062 7 1 2 73841 17061
0 17063 5 1 1 17062
0 17064 7 10 2 65376 72623
0 17065 5 1 1 96522
0 17066 7 2 2 64353 67092
0 17067 7 1 2 96523 96532
0 17068 7 1 2 94412 17067
0 17069 7 1 2 96507 17068
0 17070 5 1 1 17069
0 17071 7 1 2 17063 17070
0 17072 7 1 2 17050 17071
0 17073 5 1 1 17072
0 17074 7 1 2 84541 17073
0 17075 5 1 1 17074
0 17076 7 1 2 84370 96296
0 17077 7 1 2 96383 17076
0 17078 5 1 1 17077
0 17079 7 2 2 86420 91293
0 17080 7 1 2 90288 84311
0 17081 7 1 2 96534 17080
0 17082 5 1 1 17081
0 17083 7 1 2 17078 17082
0 17084 5 1 1 17083
0 17085 7 1 2 64354 17084
0 17086 5 1 1 17085
0 17087 7 2 2 67093 85004
0 17088 7 1 2 63973 89866
0 17089 7 1 2 96536 17088
0 17090 7 1 2 96535 17089
0 17091 5 1 1 17090
0 17092 7 1 2 17086 17091
0 17093 5 1 1 17092
0 17094 7 1 2 63773 17093
0 17095 5 1 1 17094
0 17096 7 4 2 68820 84371
0 17097 7 1 2 96297 95585
0 17098 7 1 2 96538 17097
0 17099 7 1 2 96361 17098
0 17100 5 1 1 17099
0 17101 7 1 2 17095 17100
0 17102 5 1 1 17101
0 17103 7 1 2 85679 17102
0 17104 5 1 1 17103
0 17105 7 2 2 64355 95617
0 17106 7 1 2 96323 96542
0 17107 5 1 1 17106
0 17108 7 2 2 77605 87151
0 17109 7 1 2 92063 90597
0 17110 7 1 2 92321 17109
0 17111 7 1 2 96544 17110
0 17112 5 1 1 17111
0 17113 7 1 2 17107 17112
0 17114 5 1 1 17113
0 17115 7 1 2 65590 17114
0 17116 5 1 1 17115
0 17117 7 6 2 70625 70784
0 17118 7 1 2 96546 96518
0 17119 7 1 2 96487 17118
0 17120 5 1 1 17119
0 17121 7 1 2 17116 17120
0 17122 5 1 1 17121
0 17123 7 1 2 63774 17122
0 17124 5 1 1 17123
0 17125 7 1 2 91209 96543
0 17126 5 1 1 17125
0 17127 7 1 2 17124 17126
0 17128 5 1 1 17127
0 17129 7 1 2 80690 17128
0 17130 5 1 1 17129
0 17131 7 4 2 71614 81712
0 17132 5 3 1 96552
0 17133 7 8 2 71800 79764
0 17134 5 1 1 96559
0 17135 7 1 2 96556 17134
0 17136 5 10 1 17135
0 17137 7 2 2 73721 96567
0 17138 7 2 2 63891 90890
0 17139 7 1 2 74776 96579
0 17140 7 1 2 90752 17139
0 17141 7 1 2 96577 17140
0 17142 5 1 1 17141
0 17143 7 1 2 17130 17142
0 17144 5 1 1 17143
0 17145 7 1 2 91240 17144
0 17146 5 1 1 17145
0 17147 7 1 2 17104 17146
0 17148 5 1 1 17147
0 17149 7 1 2 66859 17148
0 17150 5 1 1 17149
0 17151 7 1 2 17075 17150
0 17152 7 1 2 17022 17151
0 17153 7 1 2 16924 17152
0 17154 5 1 1 17153
0 17155 7 1 2 96262 17154
0 17156 5 1 1 17155
0 17157 7 1 2 83497 82689
0 17158 5 1 1 17157
0 17159 7 1 2 69470 80437
0 17160 7 1 2 84542 17159
0 17161 5 1 1 17160
0 17162 7 1 2 17158 17161
0 17163 5 1 1 17162
0 17164 7 1 2 96421 17163
0 17165 5 1 1 17164
0 17166 7 5 2 69471 65632
0 17167 7 1 2 78722 96581
0 17168 7 1 2 86919 17167
0 17169 5 1 1 17168
0 17170 7 1 2 17165 17169
0 17171 5 1 1 17170
0 17172 7 1 2 70398 17171
0 17173 5 1 1 17172
0 17174 7 2 2 87562 87377
0 17175 5 3 1 96586
0 17176 7 1 2 79923 96272
0 17177 7 1 2 96587 17176
0 17178 5 1 1 17177
0 17179 7 1 2 17173 17178
0 17180 5 1 1 17179
0 17181 7 1 2 89508 17180
0 17182 5 1 1 17181
0 17183 7 3 2 80589 79719
0 17184 5 3 1 96591
0 17185 7 1 2 96594 96588
0 17186 5 1 1 17185
0 17187 7 1 2 73431 17186
0 17188 5 1 1 17187
0 17189 7 1 2 84790 85821
0 17190 5 1 1 17189
0 17191 7 1 2 17188 17190
0 17192 5 2 1 17191
0 17193 7 2 2 67094 96597
0 17194 7 2 2 73808 96599
0 17195 7 1 2 90598 96601
0 17196 5 1 1 17195
0 17197 7 1 2 17182 17196
0 17198 5 1 1 17197
0 17199 7 1 2 68975 17198
0 17200 5 1 1 17199
0 17201 7 1 2 91336 91649
0 17202 7 1 2 96598 17201
0 17203 5 1 1 17202
0 17204 7 1 2 17200 17203
0 17205 5 1 1 17204
0 17206 7 1 2 74466 17205
0 17207 5 1 1 17206
0 17208 7 3 2 69472 86210
0 17209 5 1 1 96603
0 17210 7 1 2 83688 17209
0 17211 5 2 1 17210
0 17212 7 1 2 74242 96606
0 17213 7 1 2 96384 17212
0 17214 5 1 1 17213
0 17215 7 2 2 80590 74467
0 17216 7 1 2 90224 96608
0 17217 7 1 2 96338 17216
0 17218 5 1 1 17217
0 17219 7 1 2 17214 17218
0 17220 5 1 1 17219
0 17221 7 1 2 75366 17220
0 17222 5 1 1 17221
0 17223 7 12 2 73051 80691
0 17224 5 2 1 96610
0 17225 7 1 2 68000 82624
0 17226 5 3 1 17225
0 17227 7 1 2 74642 96624
0 17228 7 1 2 96622 17227
0 17229 5 1 1 17228
0 17230 7 1 2 73052 94942
0 17231 5 1 1 17230
0 17232 7 1 2 17229 17231
0 17233 5 2 1 17232
0 17234 7 2 2 72145 96627
0 17235 5 1 1 96629
0 17236 7 1 2 75155 96630
0 17237 5 1 1 17236
0 17238 7 1 2 92034 78070
0 17239 5 1 1 17238
0 17240 7 1 2 17237 17239
0 17241 5 1 1 17240
0 17242 7 1 2 69473 17241
0 17243 5 1 1 17242
0 17244 7 2 2 71801 75532
0 17245 7 2 2 84543 96631
0 17246 7 2 2 87597 86608
0 17247 7 1 2 96633 96635
0 17248 5 1 1 17247
0 17249 7 1 2 17243 17248
0 17250 5 1 1 17249
0 17251 7 1 2 73842 17250
0 17252 5 1 1 17251
0 17253 7 1 2 70144 89140
0 17254 7 1 2 96634 17253
0 17255 5 1 1 17254
0 17256 7 4 2 63892 79720
0 17257 5 1 1 96637
0 17258 7 1 2 17235 17257
0 17259 5 1 1 17258
0 17260 7 1 2 69474 308
0 17261 7 1 2 17259 17260
0 17262 5 1 1 17261
0 17263 7 1 2 17255 17262
0 17264 5 1 1 17263
0 17265 7 1 2 89573 17264
0 17266 5 1 1 17265
0 17267 7 1 2 17252 17266
0 17268 5 1 1 17267
0 17269 7 1 2 66965 17268
0 17270 5 1 1 17269
0 17271 7 1 2 17222 17270
0 17272 7 1 2 17207 17271
0 17273 5 1 1 17272
0 17274 7 1 2 68821 17273
0 17275 5 1 1 17274
0 17276 7 1 2 75367 96607
0 17277 5 1 1 17276
0 17278 7 1 2 69475 96628
0 17279 5 1 1 17278
0 17280 7 1 2 17277 17279
0 17281 5 1 1 17280
0 17282 7 1 2 96422 17281
0 17283 5 1 1 17282
0 17284 7 2 2 68624 96273
0 17285 5 1 1 96641
0 17286 7 10 2 71802 80291
0 17287 5 2 1 96643
0 17288 7 4 2 84544 96644
0 17289 5 3 1 96655
0 17290 7 1 2 96659 81249
0 17291 5 2 1 17290
0 17292 7 1 2 96642 96662
0 17293 5 1 1 17292
0 17294 7 1 2 17283 17293
0 17295 5 1 1 17294
0 17296 7 1 2 89509 17295
0 17297 5 1 1 17296
0 17298 7 2 2 75533 96663
0 17299 7 1 2 73818 96664
0 17300 5 1 1 17299
0 17301 7 1 2 17297 17300
0 17302 5 1 1 17301
0 17303 7 1 2 68976 17302
0 17304 5 1 1 17303
0 17305 7 1 2 91568 96665
0 17306 5 1 1 17305
0 17307 7 1 2 17304 17306
0 17308 5 1 1 17307
0 17309 7 1 2 83105 17308
0 17310 5 1 1 17309
0 17311 7 1 2 17275 17310
0 17312 5 1 1 17311
0 17313 7 1 2 71928 17312
0 17314 5 1 1 17313
0 17315 7 3 2 70720 91557
0 17316 5 1 1 96666
0 17317 7 1 2 91358 17316
0 17318 5 5 1 17317
0 17319 7 3 2 80591 74777
0 17320 5 3 1 96674
0 17321 7 1 2 96311 89672
0 17322 7 1 2 96675 17321
0 17323 5 1 1 17322
0 17324 7 1 2 73053 83683
0 17325 5 3 1 17324
0 17326 7 2 2 83607 96680
0 17327 7 2 2 70669 67095
0 17328 7 1 2 65591 96685
0 17329 7 1 2 96683 17328
0 17330 5 1 1 17329
0 17331 7 1 2 17323 17330
0 17332 5 1 1 17331
0 17333 7 1 2 75368 17332
0 17334 5 1 1 17333
0 17335 7 1 2 77017 96312
0 17336 5 1 1 17335
0 17337 7 1 2 94800 89495
0 17338 5 2 1 17337
0 17339 7 1 2 17336 96687
0 17340 5 2 1 17339
0 17341 7 1 2 66699 96688
0 17342 5 1 1 17341
0 17343 7 1 2 96206 17342
0 17344 5 1 1 17343
0 17345 7 1 2 64356 17344
0 17346 5 1 1 17345
0 17347 7 1 2 96689 17346
0 17348 5 1 1 17347
0 17349 7 1 2 17334 17348
0 17350 5 1 1 17349
0 17351 7 1 2 63775 17350
0 17352 5 1 1 17351
0 17353 7 1 2 74753 95912
0 17354 5 1 1 17353
0 17355 7 1 2 86668 17354
0 17356 5 1 1 17355
0 17357 7 1 2 79929 17356
0 17358 5 1 1 17357
0 17359 7 3 2 65633 72146
0 17360 5 1 1 96691
0 17361 7 2 2 73999 96692
0 17362 7 1 2 17358 96694
0 17363 5 1 1 17362
0 17364 7 1 2 17352 17363
0 17365 5 1 1 17364
0 17366 7 1 2 96669 17365
0 17367 5 1 1 17366
0 17368 7 6 2 68977 69063
0 17369 7 3 2 65592 70721
0 17370 7 1 2 96696 96702
0 17371 5 1 1 17370
0 17372 7 1 2 7051 17371
0 17373 5 3 1 17372
0 17374 7 1 2 63776 96705
0 17375 5 1 1 17374
0 17376 7 2 2 65684 91721
0 17377 7 1 2 87738 96708
0 17378 5 1 1 17377
0 17379 7 1 2 17375 17378
0 17380 5 2 1 17379
0 17381 7 2 2 65634 94801
0 17382 5 1 1 96712
0 17383 7 1 2 96475 17382
0 17384 5 2 1 17383
0 17385 7 1 2 66700 96284
0 17386 5 1 1 17385
0 17387 7 1 2 96207 17386
0 17388 5 1 1 17387
0 17389 7 1 2 64357 17388
0 17390 5 1 1 17389
0 17391 7 1 2 96714 17390
0 17392 5 1 1 17391
0 17393 7 3 2 70670 89673
0 17394 5 1 1 96716
0 17395 7 1 2 96676 96717
0 17396 5 1 1 17395
0 17397 7 1 2 96274 96684
0 17398 5 1 1 17397
0 17399 7 1 2 17396 17398
0 17400 5 1 1 17399
0 17401 7 1 2 75369 17400
0 17402 5 1 1 17401
0 17403 7 1 2 17392 17402
0 17404 5 1 1 17403
0 17405 7 1 2 96710 17404
0 17406 5 1 1 17405
0 17407 7 1 2 17367 17406
0 17408 5 1 1 17407
0 17409 7 1 2 76385 17408
0 17410 5 1 1 17409
0 17411 7 1 2 17314 17410
0 17412 5 1 1 17411
0 17413 7 1 2 67607 17412
0 17414 5 1 1 17413
0 17415 7 1 2 96499 75534
0 17416 5 1 1 17415
0 17417 7 1 2 65635 74243
0 17418 5 1 1 17417
0 17419 7 1 2 17416 17418
0 17420 5 1 1 17419
0 17421 7 1 2 96670 17420
0 17422 5 1 1 17421
0 17423 7 1 2 73830 83925
0 17424 5 1 1 17423
0 17425 7 1 2 17422 17424
0 17426 5 1 1 17425
0 17427 7 1 2 70626 17426
0 17428 5 1 1 17427
0 17429 7 1 2 66966 96423
0 17430 7 1 2 96706 17429
0 17431 5 1 1 17430
0 17432 7 1 2 17428 17431
0 17433 5 1 1 17432
0 17434 7 1 2 68822 17433
0 17435 5 1 1 17434
0 17436 7 1 2 89310 90534
0 17437 5 1 1 17436
0 17438 7 1 2 17435 17437
0 17439 5 1 1 17438
0 17440 7 1 2 75370 17439
0 17441 5 1 1 17440
0 17442 7 2 2 85889 89683
0 17443 7 1 2 91189 96719
0 17444 5 1 1 17443
0 17445 7 1 2 17441 17444
0 17446 5 1 1 17445
0 17447 7 2 2 71929 85005
0 17448 7 9 2 69476 70399
0 17449 7 1 2 82351 96723
0 17450 7 1 2 96721 17449
0 17451 7 1 2 17446 17450
0 17452 5 1 1 17451
0 17453 7 1 2 17414 17452
0 17454 5 1 1 17453
0 17455 7 1 2 72299 17454
0 17456 5 1 1 17455
0 17457 7 53 2 67253 72624
0 17458 5 2 1 96732
0 17459 7 5 2 64358 96733
0 17460 5 3 1 96787
0 17461 7 1 2 96711 96715
0 17462 5 1 1 17461
0 17463 7 1 2 63777 96690
0 17464 5 1 1 17463
0 17465 7 1 2 73432 96695
0 17466 5 1 1 17465
0 17467 7 1 2 17464 17466
0 17468 5 1 1 17467
0 17469 7 1 2 96671 17468
0 17470 5 1 1 17469
0 17471 7 1 2 17462 17470
0 17472 5 1 1 17471
0 17473 7 1 2 76386 17472
0 17474 5 1 1 17473
0 17475 7 3 2 2235 2243
0 17476 5 8 1 96795
0 17477 7 1 2 93881 96798
0 17478 5 3 1 17477
0 17479 7 1 2 66515 82352
0 17480 5 3 1 17479
0 17481 7 2 2 71615 86365
0 17482 5 2 1 96812
0 17483 7 1 2 96813 80505
0 17484 5 2 1 17483
0 17485 7 1 2 96809 96816
0 17486 5 1 1 17485
0 17487 7 1 2 70400 17486
0 17488 5 1 1 17487
0 17489 7 1 2 96806 17488
0 17490 5 1 1 17489
0 17491 7 1 2 96424 17490
0 17492 5 1 1 17491
0 17493 7 1 2 86923 96275
0 17494 5 1 1 17493
0 17495 7 1 2 17492 17494
0 17496 5 1 1 17495
0 17497 7 1 2 73054 17496
0 17498 5 1 1 17497
0 17499 7 1 2 80490 96425
0 17500 5 1 1 17499
0 17501 7 1 2 65636 93987
0 17502 5 1 1 17501
0 17503 7 1 2 17500 17502
0 17504 5 1 1 17503
0 17505 7 1 2 65053 17504
0 17506 5 1 1 17505
0 17507 7 2 2 65637 74285
0 17508 7 1 2 87510 96818
0 17509 5 1 1 17508
0 17510 7 1 2 17506 17509
0 17511 5 1 1 17510
0 17512 7 1 2 74737 17511
0 17513 5 1 1 17512
0 17514 7 1 2 17498 17513
0 17515 5 1 1 17514
0 17516 7 1 2 89510 17515
0 17517 5 1 1 17516
0 17518 7 1 2 63974 96602
0 17519 5 1 1 17518
0 17520 7 1 2 17517 17519
0 17521 5 1 1 17520
0 17522 7 1 2 68978 17521
0 17523 5 1 1 17522
0 17524 7 1 2 91569 96600
0 17525 5 1 1 17524
0 17526 7 1 2 72039 17525
0 17527 7 1 2 17523 17526
0 17528 5 1 1 17527
0 17529 7 3 2 73055 85623
0 17530 5 3 1 96820
0 17531 7 1 2 73433 93976
0 17532 5 1 1 17531
0 17533 7 1 2 96823 17532
0 17534 5 1 1 17533
0 17535 7 1 2 96482 17534
0 17536 5 1 1 17535
0 17537 7 3 2 96276 88917
0 17538 7 1 2 96638 96826
0 17539 5 1 1 17538
0 17540 7 1 2 66967 17539
0 17541 7 1 2 17536 17540
0 17542 5 1 1 17541
0 17543 7 1 2 68823 17542
0 17544 7 1 2 17528 17543
0 17545 5 1 1 17544
0 17546 7 1 2 74012 17545
0 17547 5 1 1 17546
0 17548 7 3 2 96426 89511
0 17549 7 1 2 85624 96829
0 17550 5 1 1 17549
0 17551 7 2 2 73843 75535
0 17552 5 1 1 96832
0 17553 7 1 2 17550 17552
0 17554 5 1 1 17553
0 17555 7 1 2 73056 17554
0 17556 5 1 1 17555
0 17557 7 1 2 82908 77018
0 17558 7 1 2 91186 17557
0 17559 5 1 1 17558
0 17560 7 1 2 17556 17559
0 17561 5 1 1 17560
0 17562 7 1 2 68979 17561
0 17563 5 1 1 17562
0 17564 7 1 2 92035 91570
0 17565 5 1 1 17564
0 17566 7 1 2 17563 17565
0 17567 5 1 1 17566
0 17568 7 1 2 66968 17567
0 17569 5 1 1 17568
0 17570 7 1 2 79004 17569
0 17571 5 1 1 17570
0 17572 7 1 2 71930 17571
0 17573 7 1 2 17547 17572
0 17574 5 1 1 17573
0 17575 7 1 2 17474 17574
0 17576 5 1 1 17575
0 17577 7 1 2 96788 17576
0 17578 5 1 1 17577
0 17579 7 1 2 17456 17578
0 17580 5 1 1 17579
0 17581 7 1 2 64057 17580
0 17582 5 1 1 17581
0 17583 7 4 2 72625 74183
0 17584 5 2 1 96834
0 17585 7 3 2 67608 78121
0 17586 5 1 1 96840
0 17587 7 1 2 96838 17586
0 17588 5 1 1 17587
0 17589 7 1 2 74761 92916
0 17590 5 1 1 17589
0 17591 7 1 2 17590 96830
0 17592 5 1 1 17591
0 17593 7 1 2 89512 96477
0 17594 5 1 1 17593
0 17595 7 3 2 63975 67096
0 17596 7 1 2 73809 96843
0 17597 5 1 1 17596
0 17598 7 1 2 17594 17597
0 17599 5 1 1 17598
0 17600 7 1 2 88467 17599
0 17601 5 1 1 17600
0 17602 7 1 2 17592 17601
0 17603 5 1 1 17602
0 17604 7 1 2 68980 17603
0 17605 5 1 1 17604
0 17606 7 3 2 86895 74286
0 17607 7 1 2 91571 96846
0 17608 5 2 1 17607
0 17609 7 1 2 17605 96849
0 17610 5 1 1 17609
0 17611 7 1 2 83106 17610
0 17612 5 1 1 17611
0 17613 7 1 2 93956 75221
0 17614 5 1 1 17613
0 17615 7 1 2 82803 76769
0 17616 5 1 1 17615
0 17617 7 1 2 17614 17616
0 17618 5 1 1 17617
0 17619 7 1 2 74738 17618
0 17620 5 1 1 17619
0 17621 7 1 2 83393 76770
0 17622 5 1 1 17621
0 17623 7 1 2 75240 17622
0 17624 5 1 1 17623
0 17625 7 1 2 80498 75222
0 17626 5 1 1 17625
0 17627 7 1 2 65054 17626
0 17628 5 1 1 17627
0 17629 7 1 2 73057 17628
0 17630 7 1 2 17624 17629
0 17631 5 1 1 17630
0 17632 7 1 2 17620 17631
0 17633 5 1 1 17632
0 17634 7 1 2 70627 17633
0 17635 5 1 1 17634
0 17636 7 1 2 84147 86561
0 17637 5 1 1 17636
0 17638 7 1 2 17635 17637
0 17639 5 1 1 17638
0 17640 7 1 2 73844 17639
0 17641 5 1 1 17640
0 17642 7 2 2 75145 74287
0 17643 7 1 2 93843 96851
0 17644 5 1 1 17643
0 17645 7 2 2 73434 93957
0 17646 7 1 2 68001 96853
0 17647 5 1 1 17646
0 17648 7 1 2 92917 17647
0 17649 5 1 1 17648
0 17650 7 1 2 66969 88563
0 17651 7 1 2 17649 17650
0 17652 5 1 1 17651
0 17653 7 1 2 17644 17652
0 17654 5 1 1 17653
0 17655 7 1 2 89574 17654
0 17656 5 1 1 17655
0 17657 7 1 2 80506 87378
0 17658 5 2 1 17657
0 17659 7 1 2 66701 74813
0 17660 5 1 1 17659
0 17661 7 1 2 96855 17660
0 17662 5 1 1 17661
0 17663 7 1 2 88203 17662
0 17664 5 1 1 17663
0 17665 7 1 2 93978 15835
0 17666 5 3 1 17665
0 17667 7 2 2 84545 88564
0 17668 5 1 1 96860
0 17669 7 1 2 96857 96861
0 17670 5 1 1 17669
0 17671 7 1 2 17664 17670
0 17672 5 1 1 17671
0 17673 7 1 2 74468 94080
0 17674 7 1 2 17672 17673
0 17675 5 1 1 17674
0 17676 7 1 2 17656 17675
0 17677 7 1 2 17641 17676
0 17678 5 1 1 17677
0 17679 7 1 2 68824 17678
0 17680 5 1 1 17679
0 17681 7 1 2 17612 17680
0 17682 5 1 1 17681
0 17683 7 1 2 17588 17682
0 17684 5 1 1 17683
0 17685 7 8 2 64058 70145
0 17686 7 2 2 71616 96862
0 17687 7 1 2 84285 96870
0 17688 5 1 1 17687
0 17689 7 1 2 96839 17688
0 17690 5 1 1 17689
0 17691 7 2 2 68357 17690
0 17692 7 1 2 83201 96872
0 17693 5 1 1 17692
0 17694 7 2 2 87379 84372
0 17695 7 2 2 93697 87959
0 17696 7 1 2 96874 96876
0 17697 5 1 1 17696
0 17698 7 1 2 17693 17697
0 17699 5 1 1 17698
0 17700 7 1 2 73722 17699
0 17701 5 1 1 17700
0 17702 7 2 2 73058 77097
0 17703 5 1 1 96878
0 17704 7 1 2 82046 96841
0 17705 7 1 2 17703 17704
0 17706 5 1 1 17705
0 17707 7 1 2 83380 74184
0 17708 7 1 2 87899 17707
0 17709 5 1 1 17708
0 17710 7 1 2 17706 17709
0 17711 5 1 1 17710
0 17712 7 1 2 83880 17711
0 17713 5 1 1 17712
0 17714 7 1 2 17701 17713
0 17715 5 1 1 17714
0 17716 7 1 2 66702 17715
0 17717 5 1 1 17716
0 17718 7 1 2 74185 90931
0 17719 5 2 1 17718
0 17720 7 2 2 71803 92347
0 17721 7 1 2 78122 96882
0 17722 5 1 1 17721
0 17723 7 1 2 96880 17722
0 17724 5 1 1 17723
0 17725 7 1 2 83881 76996
0 17726 7 1 2 17724 17725
0 17727 5 1 1 17726
0 17728 7 1 2 17717 17727
0 17729 5 1 1 17728
0 17730 7 1 2 96324 17729
0 17731 5 1 1 17730
0 17732 7 2 2 87739 89559
0 17733 5 1 1 96884
0 17734 7 2 2 66970 96885
0 17735 5 1 1 96886
0 17736 7 1 2 82909 96887
0 17737 7 1 2 96873 17736
0 17738 5 1 1 17737
0 17739 7 1 2 17731 17738
0 17740 5 1 1 17739
0 17741 7 1 2 67097 17740
0 17742 5 1 1 17741
0 17743 7 1 2 17684 17742
0 17744 5 1 1 17743
0 17745 7 1 2 72300 17744
0 17746 5 1 1 17745
0 17747 7 2 2 73059 86936
0 17748 5 2 1 96888
0 17749 7 1 2 77098 80096
0 17750 5 3 1 17749
0 17751 7 1 2 66703 96892
0 17752 5 1 1 17751
0 17753 7 1 2 96889 17752
0 17754 5 1 1 17753
0 17755 7 4 2 65055 87511
0 17756 5 3 1 96895
0 17757 7 2 2 68002 96899
0 17758 5 1 1 96902
0 17759 7 1 2 74643 80507
0 17760 5 1 1 17759
0 17761 7 1 2 96903 17760
0 17762 5 1 1 17761
0 17763 7 1 2 67098 17762
0 17764 7 2 2 17754 17763
0 17765 7 1 2 73819 96904
0 17766 5 1 1 17765
0 17767 7 1 2 77085 96427
0 17768 5 1 1 17767
0 17769 7 1 2 96471 17768
0 17770 5 1 1 17769
0 17771 7 1 2 70146 17770
0 17772 5 1 1 17771
0 17773 7 2 2 70671 77726
0 17774 5 1 1 96906
0 17775 7 1 2 17774 17285
0 17776 5 1 1 17775
0 17777 7 1 2 71617 17776
0 17778 5 1 1 17777
0 17779 7 1 2 17772 17778
0 17780 5 1 1 17779
0 17781 7 1 2 73060 17780
0 17782 5 1 1 17781
0 17783 7 1 2 70672 92
0 17784 5 1 1 17783
0 17785 7 1 2 17360 17784
0 17786 7 1 2 88443 17785
0 17787 5 1 1 17786
0 17788 7 1 2 17782 17787
0 17789 5 1 1 17788
0 17790 7 1 2 66704 17789
0 17791 5 1 1 17790
0 17792 7 1 2 74644 96819
0 17793 5 1 1 17792
0 17794 7 2 2 70673 90147
0 17795 7 1 2 65056 96908
0 17796 5 1 1 17795
0 17797 7 1 2 17793 17796
0 17798 5 1 1 17797
0 17799 7 1 2 68003 17798
0 17800 5 1 1 17799
0 17801 7 1 2 80463 79721
0 17802 7 1 2 96428 17801
0 17803 5 1 1 17802
0 17804 7 1 2 17800 17803
0 17805 5 1 1 17804
0 17806 7 1 2 73435 17805
0 17807 5 1 1 17806
0 17808 7 2 2 65638 89755
0 17809 5 1 1 96910
0 17810 7 1 2 85822 96911
0 17811 5 1 1 17810
0 17812 7 1 2 17807 17811
0 17813 7 1 2 17791 17812
0 17814 5 1 1 17813
0 17815 7 1 2 89513 17814
0 17816 5 1 1 17815
0 17817 7 1 2 17766 17816
0 17818 5 1 1 17817
0 17819 7 1 2 68981 17818
0 17820 5 1 1 17819
0 17821 7 1 2 91572 96905
0 17822 5 1 1 17821
0 17823 7 1 2 72040 17822
0 17824 7 1 2 17820 17823
0 17825 5 1 1 17824
0 17826 7 1 2 77019 88428
0 17827 7 1 2 96362 17826
0 17828 5 1 1 17827
0 17829 7 1 2 96488 96847
0 17830 5 1 1 17829
0 17831 7 1 2 66971 17830
0 17832 7 1 2 17828 17831
0 17833 5 1 1 17832
0 17834 7 1 2 68825 17833
0 17835 7 1 2 17825 17834
0 17836 5 1 1 17835
0 17837 7 1 2 74013 17836
0 17838 5 1 1 17837
0 17839 7 1 2 76155 96713
0 17840 5 1 1 17839
0 17841 7 1 2 88429 96473
0 17842 5 1 1 17841
0 17843 7 1 2 17840 17842
0 17844 5 1 1 17843
0 17845 7 1 2 89514 17844
0 17846 5 1 1 17845
0 17847 7 1 2 73820 96848
0 17848 5 1 1 17847
0 17849 7 1 2 17846 17848
0 17850 5 1 1 17849
0 17851 7 1 2 68982 17850
0 17852 5 1 1 17851
0 17853 7 1 2 96850 17852
0 17854 5 1 1 17853
0 17855 7 1 2 66972 17854
0 17856 5 1 1 17855
0 17857 7 1 2 79005 17856
0 17858 5 1 1 17857
0 17859 7 1 2 64359 17858
0 17860 7 1 2 17838 17859
0 17861 5 1 1 17860
0 17862 7 1 2 74028 96325
0 17863 5 1 1 17862
0 17864 7 1 2 17733 17863
0 17865 5 2 1 17864
0 17866 7 1 2 82839 86556
0 17867 7 1 2 95834 17866
0 17868 7 1 2 96912 17867
0 17869 5 1 1 17868
0 17870 7 1 2 17861 17869
0 17871 5 1 1 17870
0 17872 7 1 2 64059 96734
0 17873 7 1 2 17871 17872
0 17874 5 1 1 17873
0 17875 7 1 2 17746 17874
0 17876 5 1 1 17875
0 17877 7 1 2 71931 17876
0 17878 5 1 1 17877
0 17879 7 37 2 69121 72301
0 17880 5 2 1 96914
0 17881 7 38 2 64060 67254
0 17882 5 2 1 96953
0 17883 7 2 2 96951 96991
0 17884 5 9 1 96993
0 17885 7 1 2 84935 96995
0 17886 5 3 1 17885
0 17887 7 3 2 67609 96263
0 17888 7 2 2 68004 92906
0 17889 5 1 1 97010
0 17890 7 1 2 64360 17889
0 17891 5 1 1 17890
0 17892 7 1 2 97007 17891
0 17893 5 1 1 17892
0 17894 7 1 2 97004 17893
0 17895 5 1 1 17894
0 17896 7 1 2 80188 17895
0 17897 5 1 1 17896
0 17898 7 1 2 68005 96893
0 17899 5 1 1 17898
0 17900 7 1 2 64361 17899
0 17901 5 1 1 17900
0 17902 7 1 2 97008 17901
0 17903 5 1 1 17902
0 17904 7 1 2 97005 17903
0 17905 5 1 1 17904
0 17906 7 1 2 66705 81339
0 17907 7 1 2 17905 17906
0 17908 5 1 1 17907
0 17909 7 1 2 17897 17908
0 17910 5 1 1 17909
0 17911 7 1 2 73845 17910
0 17912 5 1 1 17911
0 17913 7 7 2 68983 84597
0 17914 5 1 1 97012
0 17915 7 1 2 88292 17914
0 17916 5 2 1 17915
0 17917 7 49 2 72302 67610
0 17918 5 1 1 97021
0 17919 7 8 2 69477 97022
0 17920 5 2 1 97070
0 17921 7 1 2 97071 96994
0 17922 5 1 1 17921
0 17923 7 1 2 97006 17922
0 17924 5 1 1 17923
0 17925 7 1 2 97019 17924
0 17926 5 1 1 17925
0 17927 7 1 2 92907 88204
0 17928 5 1 1 17927
0 17929 7 1 2 96894 97013
0 17930 5 1 1 17929
0 17931 7 1 2 17928 17930
0 17932 5 1 1 17931
0 17933 7 11 2 68006 97023
0 17934 7 1 2 64061 97080
0 17935 7 1 2 17932 17934
0 17936 5 1 1 17935
0 17937 7 1 2 17926 17936
0 17938 5 1 1 17937
0 17939 7 1 2 90334 17938
0 17940 5 1 1 17939
0 17941 7 1 2 17912 17940
0 17942 5 1 1 17941
0 17943 7 1 2 72041 17942
0 17944 5 1 1 17943
0 17945 7 1 2 68007 94202
0 17946 5 1 1 17945
0 17947 7 1 2 73902 90470
0 17948 5 1 1 17947
0 17949 7 1 2 73061 83514
0 17950 7 1 2 17948 17949
0 17951 5 1 1 17950
0 17952 7 1 2 81464 17951
0 17953 7 1 2 17946 17952
0 17954 5 1 1 17953
0 17955 7 1 2 74817 78936
0 17956 5 1 1 17955
0 17957 7 1 2 66706 17956
0 17958 5 1 1 17957
0 17959 7 1 2 74763 17958
0 17960 5 1 1 17959
0 17961 7 1 2 80404 81526
0 17962 7 1 2 17960 17961
0 17963 5 1 1 17962
0 17964 7 1 2 17954 17963
0 17965 5 1 1 17964
0 17966 7 1 2 96277 17965
0 17967 5 1 1 17966
0 17968 7 4 2 65057 70674
0 17969 5 1 1 97091
0 17970 7 1 2 72147 84756
0 17971 7 1 2 84668 17970
0 17972 7 3 2 84546 17971
0 17973 7 1 2 97092 97095
0 17974 5 1 1 17973
0 17975 7 1 2 17967 17974
0 17976 5 1 1 17975
0 17977 7 1 2 88918 17976
0 17978 5 1 1 17977
0 17979 7 1 2 91266 73825
0 17980 7 1 2 97096 17979
0 17981 5 1 1 17980
0 17982 7 1 2 17978 17981
0 17983 5 1 1 17982
0 17984 7 1 2 63893 17983
0 17985 5 1 1 17984
0 17986 7 1 2 91547 97097
0 17987 5 1 1 17986
0 17988 7 1 2 17985 17987
0 17989 5 1 1 17988
0 17990 7 12 2 66973 72303
0 17991 7 1 2 97098 79632
0 17992 7 1 2 17989 17991
0 17993 5 1 1 17992
0 17994 7 1 2 17944 17993
0 17995 5 1 1 17994
0 17996 7 1 2 66860 17995
0 17997 5 1 1 17996
0 17998 7 3 2 64062 72042
0 17999 7 2 2 88023 91127
0 18000 7 1 2 89724 89515
0 18001 7 1 2 97113 18000
0 18002 7 23 2 67255 73062
0 18003 7 2 2 92576 97115
0 18004 7 2 2 68826 74087
0 18005 7 1 2 97138 97140
0 18006 7 1 2 18001 18005
0 18007 5 1 1 18006
0 18008 7 1 2 89121 91619
0 18009 5 1 1 18008
0 18010 7 1 2 76915 91421
0 18011 5 1 1 18010
0 18012 7 1 2 18009 18011
0 18013 5 1 1 18012
0 18014 7 1 2 68827 18013
0 18015 5 1 1 18014
0 18016 7 2 2 63894 74005
0 18017 7 1 2 77783 97142
0 18018 5 1 1 18017
0 18019 7 1 2 18015 18018
0 18020 5 1 1 18019
0 18021 7 1 2 97024 18020
0 18022 5 1 1 18021
0 18023 7 4 2 67256 82240
0 18024 5 1 1 97144
0 18025 7 6 2 74088 84194
0 18026 7 2 2 79102 97148
0 18027 7 1 2 97145 97154
0 18028 5 1 1 18027
0 18029 7 1 2 18022 18028
0 18030 5 1 1 18029
0 18031 7 1 2 73846 18030
0 18032 5 1 1 18031
0 18033 7 2 2 91849 88565
0 18034 7 1 2 90335 97156
0 18035 5 1 1 18034
0 18036 7 3 2 69064 87740
0 18037 7 1 2 94232 97158
0 18038 7 1 2 91338 18037
0 18039 5 1 1 18038
0 18040 7 1 2 18035 18039
0 18041 5 1 1 18040
0 18042 7 1 2 97025 18041
0 18043 5 1 1 18042
0 18044 7 8 2 73063 96735
0 18045 5 1 1 97161
0 18046 7 1 2 97162 91511
0 18047 7 1 2 92148 97159
0 18048 7 1 2 18046 18047
0 18049 5 1 1 18048
0 18050 7 1 2 18043 18049
0 18051 7 1 2 18032 18050
0 18052 5 1 1 18051
0 18053 7 1 2 66707 83381
0 18054 7 1 2 18052 18053
0 18055 5 1 1 18054
0 18056 7 1 2 18007 18055
0 18057 5 1 1 18056
0 18058 7 1 2 97110 18057
0 18059 5 1 1 18058
0 18060 7 4 2 64362 65685
0 18061 7 3 2 94636 97169
0 18062 7 3 2 74778 97026
0 18063 7 1 2 86557 92235
0 18064 7 1 2 97176 18063
0 18065 7 1 2 97173 18064
0 18066 5 1 1 18065
0 18067 7 1 2 18059 18066
0 18068 5 1 1 18067
0 18069 7 1 2 77293 18068
0 18070 5 1 1 18069
0 18071 7 1 2 17997 18070
0 18072 7 1 2 17878 18071
0 18073 5 1 1 18072
0 18074 7 1 2 65377 18073
0 18075 5 1 1 18074
0 18076 7 3 2 93698 90371
0 18077 7 4 2 91168 96342
0 18078 7 1 2 97179 97182
0 18079 5 1 1 18078
0 18080 7 1 2 96405 18079
0 18081 5 2 1 18080
0 18082 7 1 2 63895 97186
0 18083 5 1 1 18082
0 18084 7 2 2 84063 93699
0 18085 7 1 2 92307 97188
0 18086 7 2 2 73847 18085
0 18087 7 1 2 72626 97190
0 18088 5 1 1 18087
0 18089 7 1 2 18083 18088
0 18090 5 1 1 18089
0 18091 7 1 2 83020 18090
0 18092 5 1 1 18091
0 18093 7 2 2 75748 96913
0 18094 7 1 2 93348 97192
0 18095 5 1 1 18094
0 18096 7 1 2 18092 18095
0 18097 5 1 1 18096
0 18098 7 1 2 72304 18097
0 18099 5 1 1 18098
0 18100 7 1 2 83882 83562
0 18101 5 1 1 18100
0 18102 7 1 2 2373 18101
0 18103 5 1 1 18102
0 18104 7 1 2 96326 18103
0 18105 5 1 1 18104
0 18106 7 1 2 17735 18105
0 18107 5 2 1 18106
0 18108 7 1 2 96954 93570
0 18109 7 1 2 97194 18108
0 18110 5 1 1 18109
0 18111 7 1 2 18099 18110
0 18112 5 1 1 18111
0 18113 7 1 2 64363 18112
0 18114 5 1 1 18113
0 18115 7 5 2 71932 72305
0 18116 7 1 2 97196 96842
0 18117 7 1 2 97195 18116
0 18118 5 1 1 18117
0 18119 7 1 2 18114 18118
0 18120 5 1 1 18119
0 18121 7 1 2 67099 18120
0 18122 5 1 1 18121
0 18123 7 12 2 67257 68625
0 18124 7 1 2 84936 97201
0 18125 7 1 2 85573 18124
0 18126 5 1 1 18125
0 18127 7 4 2 71618 92348
0 18128 7 4 2 72306 77898
0 18129 7 1 2 91819 97217
0 18130 7 1 2 97213 18129
0 18131 5 1 1 18130
0 18132 7 1 2 18126 18131
0 18133 5 2 1 18132
0 18134 7 1 2 68828 97221
0 18135 5 1 1 18134
0 18136 7 4 2 72307 92349
0 18137 7 1 2 86523 90653
0 18138 7 1 2 97223 18137
0 18139 5 1 1 18138
0 18140 7 1 2 18135 18139
0 18141 5 1 1 18140
0 18142 7 1 2 96363 18141
0 18143 5 1 1 18142
0 18144 7 1 2 63778 97222
0 18145 5 1 1 18144
0 18146 7 1 2 82835 3873
0 18147 5 1 1 18146
0 18148 7 4 2 67258 83986
0 18149 7 1 2 71933 79103
0 18150 7 1 2 97227 18149
0 18151 7 1 2 18147 18150
0 18152 5 1 1 18151
0 18153 7 1 2 18145 18152
0 18154 5 1 1 18153
0 18155 7 1 2 96348 18154
0 18156 5 1 1 18155
0 18157 7 1 2 18143 18156
0 18158 5 1 1 18157
0 18159 7 1 2 92858 18158
0 18160 5 1 1 18159
0 18161 7 1 2 18122 18160
0 18162 5 1 1 18161
0 18163 7 1 2 73064 18162
0 18164 5 1 1 18163
0 18165 7 5 2 72308 83135
0 18166 7 4 2 68984 87960
0 18167 7 2 2 73903 97236
0 18168 7 1 2 97240 92119
0 18169 5 1 1 18168
0 18170 7 1 2 77020 77032
0 18171 5 1 1 18170
0 18172 7 1 2 18169 18171
0 18173 5 1 1 18172
0 18174 7 1 2 68829 18173
0 18175 5 1 1 18174
0 18176 7 2 2 73436 75175
0 18177 5 1 1 97242
0 18178 7 1 2 78168 97243
0 18179 5 1 1 18178
0 18180 7 1 2 18175 18179
0 18181 5 1 1 18180
0 18182 7 1 2 73848 18181
0 18183 5 1 1 18182
0 18184 7 1 2 92690 90344
0 18185 5 1 1 18184
0 18186 7 1 2 71619 87741
0 18187 7 1 2 91169 18186
0 18188 7 1 2 94979 91408
0 18189 7 1 2 18187 18188
0 18190 5 1 1 18189
0 18191 7 1 2 18185 18190
0 18192 7 1 2 18183 18191
0 18193 5 1 1 18192
0 18194 7 1 2 67611 18193
0 18195 5 1 1 18194
0 18196 7 2 2 67100 81412
0 18197 7 4 2 69478 88024
0 18198 7 1 2 97244 97246
0 18199 7 1 2 94415 18198
0 18200 5 1 1 18199
0 18201 7 3 2 67101 91877
0 18202 7 2 2 81413 97250
0 18203 7 5 2 89082 84064
0 18204 7 1 2 73849 97255
0 18205 7 1 2 97253 18204
0 18206 5 1 1 18205
0 18207 7 1 2 18200 18206
0 18208 7 1 2 18195 18207
0 18209 5 1 1 18208
0 18210 7 1 2 97111 18209
0 18211 5 1 1 18210
0 18212 7 2 2 78363 92236
0 18213 7 1 2 89251 97260
0 18214 7 1 2 97174 18213
0 18215 5 1 1 18214
0 18216 7 1 2 18211 18215
0 18217 5 1 1 18216
0 18218 7 1 2 97231 18217
0 18219 5 1 1 18218
0 18220 7 1 2 18164 18219
0 18221 5 1 1 18220
0 18222 7 1 2 81850 18221
0 18223 5 1 1 18222
0 18224 7 1 2 81451 92250
0 18225 5 8 1 18224
0 18226 7 2 2 68626 97262
0 18227 7 2 2 77899 90647
0 18228 7 1 2 97270 97272
0 18229 5 1 1 18228
0 18230 7 2 2 79790 93349
0 18231 7 1 2 96879 97274
0 18232 5 1 1 18231
0 18233 7 1 2 18229 18232
0 18234 5 1 1 18233
0 18235 7 1 2 64364 18234
0 18236 5 1 1 18235
0 18237 7 10 2 70147 72627
0 18238 5 1 1 97276
0 18239 7 4 2 66516 82106
0 18240 5 1 1 97286
0 18241 7 2 2 97277 97287
0 18242 7 2 2 90891 77900
0 18243 7 1 2 73065 97292
0 18244 7 1 2 97290 18243
0 18245 5 1 1 18244
0 18246 7 1 2 18236 18245
0 18247 5 1 1 18246
0 18248 7 1 2 71804 18247
0 18249 5 1 1 18248
0 18250 7 5 2 72628 79722
0 18251 7 1 2 86400 97294
0 18252 7 1 2 96877 18251
0 18253 5 1 1 18252
0 18254 7 1 2 18249 18253
0 18255 5 1 1 18254
0 18256 7 1 2 96364 18255
0 18257 5 1 1 18256
0 18258 7 1 2 71934 82973
0 18259 7 1 2 96835 18258
0 18260 7 1 2 90249 18259
0 18261 7 3 2 73066 83587
0 18262 5 1 1 97299
0 18263 7 1 2 97300 83659
0 18264 7 1 2 18260 18263
0 18265 5 1 1 18264
0 18266 7 1 2 18257 18265
0 18267 5 1 1 18266
0 18268 7 1 2 66974 18267
0 18269 5 1 1 18268
0 18270 7 2 2 66975 91496
0 18271 7 1 2 97302 90420
0 18272 7 1 2 96319 18271
0 18273 5 1 1 18272
0 18274 7 1 2 80405 94774
0 18275 7 1 2 92313 18274
0 18276 7 1 2 97183 18275
0 18277 5 1 1 18276
0 18278 7 1 2 18273 18277
0 18279 5 1 1 18278
0 18280 7 1 2 68985 18279
0 18281 5 1 1 18280
0 18282 7 2 2 79633 93844
0 18283 7 1 2 86567 84584
0 18284 7 1 2 97304 18283
0 18285 7 1 2 73850 18284
0 18286 5 1 1 18285
0 18287 7 1 2 18281 18286
0 18288 5 1 1 18287
0 18289 7 1 2 64365 18288
0 18290 5 1 1 18289
0 18291 7 3 2 69479 66976
0 18292 7 1 2 82910 97306
0 18293 7 1 2 95419 18292
0 18294 7 1 2 96365 18293
0 18295 5 1 1 18294
0 18296 7 1 2 18290 18295
0 18297 5 1 1 18296
0 18298 7 1 2 84547 18297
0 18299 5 1 1 18298
0 18300 7 2 2 73067 78364
0 18301 7 1 2 86095 74186
0 18302 7 1 2 97309 18301
0 18303 7 1 2 96389 18302
0 18304 5 1 1 18303
0 18305 7 1 2 18299 18304
0 18306 5 1 1 18305
0 18307 7 1 2 65058 18306
0 18308 5 1 1 18307
0 18309 7 5 2 73068 82107
0 18310 7 1 2 97311 96343
0 18311 7 2 2 70722 86134
0 18312 7 3 2 93727 92314
0 18313 7 1 2 97114 97318
0 18314 7 1 2 97316 18313
0 18315 7 1 2 18310 18314
0 18316 5 1 1 18315
0 18317 7 1 2 18308 18316
0 18318 7 1 2 18269 18317
0 18319 5 1 1 18318
0 18320 7 1 2 70401 18319
0 18321 5 1 1 18320
0 18322 7 1 2 70628 87380
0 18323 7 1 2 95940 18322
0 18324 5 1 1 18323
0 18325 7 1 2 85792 18324
0 18326 5 1 1 18325
0 18327 7 1 2 68830 18326
0 18328 5 1 1 18327
0 18329 7 1 2 3603 18328
0 18330 5 1 1 18329
0 18331 7 1 2 73437 18330
0 18332 5 1 1 18331
0 18333 7 1 2 78987 87548
0 18334 7 1 2 94582 18333
0 18335 5 1 1 18334
0 18336 7 1 2 18332 18335
0 18337 5 1 1 18336
0 18338 7 1 2 96366 18337
0 18339 5 1 1 18338
0 18340 7 1 2 85827 79658
0 18341 5 1 1 18340
0 18342 7 1 2 86401 83202
0 18343 7 1 2 87683 18342
0 18344 5 1 1 18343
0 18345 7 1 2 18341 18344
0 18346 5 1 1 18345
0 18347 7 1 2 96349 18346
0 18348 5 1 1 18347
0 18349 7 1 2 18339 18348
0 18350 5 1 1 18349
0 18351 7 1 2 96836 18350
0 18352 5 1 1 18351
0 18353 7 1 2 72148 18352
0 18354 7 1 2 18321 18353
0 18355 5 1 1 18354
0 18356 7 1 2 89151 94775
0 18357 5 1 1 18356
0 18358 7 4 2 71805 66977
0 18359 7 2 2 79807 97321
0 18360 7 1 2 83136 76976
0 18361 7 1 2 97325 18360
0 18362 5 1 1 18361
0 18363 7 1 2 18357 18362
0 18364 5 1 1 18363
0 18365 7 1 2 90315 18364
0 18366 5 1 1 18365
0 18367 7 6 2 69122 65593
0 18368 7 1 2 89152 97327
0 18369 7 1 2 94081 18368
0 18370 5 1 1 18369
0 18371 7 1 2 18366 18370
0 18372 5 1 1 18371
0 18373 7 1 2 66861 18372
0 18374 5 1 1 18373
0 18375 7 2 2 66978 79723
0 18376 7 1 2 94776 94240
0 18377 7 1 2 97333 18376
0 18378 5 1 1 18377
0 18379 7 1 2 18374 18378
0 18380 5 1 1 18379
0 18381 7 1 2 64366 18380
0 18382 5 1 1 18381
0 18383 7 1 2 84751 86143
0 18384 5 6 1 18383
0 18385 7 5 2 73069 80292
0 18386 7 1 2 97335 97341
0 18387 5 1 1 18386
0 18388 7 1 2 96589 18387
0 18389 5 1 1 18388
0 18390 7 1 2 73438 18389
0 18391 5 1 1 18390
0 18392 7 1 2 79808 87089
0 18393 5 2 1 18392
0 18394 7 1 2 66708 96545
0 18395 5 1 1 18394
0 18396 7 1 2 97346 18395
0 18397 5 1 1 18396
0 18398 7 1 2 65059 18397
0 18399 5 1 1 18398
0 18400 7 1 2 18391 18399
0 18401 5 1 1 18400
0 18402 7 1 2 88982 97307
0 18403 7 1 2 18401 18402
0 18404 5 1 1 18403
0 18405 7 1 2 18382 18404
0 18406 5 1 1 18405
0 18407 7 1 2 63779 18406
0 18408 5 1 1 18407
0 18409 7 1 2 73070 83026
0 18410 5 1 1 18409
0 18411 7 1 2 96590 18410
0 18412 5 1 1 18411
0 18413 7 1 2 73439 18412
0 18414 5 1 1 18413
0 18415 7 1 2 88439 18414
0 18416 5 2 1 18415
0 18417 7 1 2 74469 97348
0 18418 5 1 1 18417
0 18419 7 1 2 79724 82821
0 18420 5 1 1 18419
0 18421 7 1 2 18418 18420
0 18422 5 2 1 18421
0 18423 7 1 2 94241 97350
0 18424 5 1 1 18423
0 18425 7 1 2 76803 97334
0 18426 5 1 1 18425
0 18427 7 1 2 66709 85790
0 18428 5 1 1 18427
0 18429 7 1 2 18426 18428
0 18430 5 2 1 18429
0 18431 7 1 2 90316 97352
0 18432 5 1 1 18431
0 18433 7 1 2 18424 18432
0 18434 5 1 1 18433
0 18435 7 1 2 64367 93700
0 18436 7 1 2 18434 18435
0 18437 5 1 1 18436
0 18438 7 1 2 18408 18437
0 18439 5 1 1 18438
0 18440 7 1 2 63896 18439
0 18441 5 1 1 18440
0 18442 7 1 2 63780 97353
0 18443 5 1 1 18442
0 18444 7 1 2 85101 97351
0 18445 5 1 1 18444
0 18446 7 1 2 18443 18445
0 18447 5 1 1 18446
0 18448 7 1 2 74187 96321
0 18449 7 1 2 18447 18448
0 18450 5 1 1 18449
0 18451 7 1 2 18441 18450
0 18452 5 1 1 18451
0 18453 7 1 2 72629 18452
0 18454 5 1 1 18453
0 18455 7 2 2 63897 81527
0 18456 7 1 2 92472 97354
0 18457 7 1 2 97349 18456
0 18458 5 1 1 18457
0 18459 7 1 2 67102 18458
0 18460 7 1 2 18454 18459
0 18461 5 1 1 18460
0 18462 7 1 2 72309 18461
0 18463 7 1 2 18355 18462
0 18464 5 1 1 18463
0 18465 7 1 2 18223 18464
0 18466 7 1 2 18075 18465
0 18467 7 1 2 17582 18466
0 18468 5 1 1 18467
0 18469 7 1 2 65760 18468
0 18470 5 1 1 18469
0 18471 7 1 2 17156 18470
0 18472 5 1 1 18471
0 18473 7 1 2 96257 18472
0 18474 5 1 1 18473
0 18475 7 10 2 64684 71339
0 18476 5 6 1 97356
0 18477 7 2 2 92930 97366
0 18478 5 58 1 97372
0 18479 7 1 2 91850 87982
0 18480 5 1 1 18479
0 18481 7 2 2 78723 93318
0 18482 7 1 2 97256 97432
0 18483 5 1 1 18482
0 18484 7 1 2 18480 18483
0 18485 5 1 1 18484
0 18486 7 1 2 97027 18485
0 18487 5 1 1 18486
0 18488 7 2 2 73723 82241
0 18489 7 11 2 67103 67259
0 18490 7 2 2 76804 97436
0 18491 7 2 2 94981 97447
0 18492 7 1 2 97434 97449
0 18493 5 1 1 18492
0 18494 7 1 2 18487 18493
0 18495 5 1 1 18494
0 18496 7 1 2 71041 18495
0 18497 5 1 1 18496
0 18498 7 2 2 73071 96293
0 18499 7 2 2 65966 87408
0 18500 7 1 2 97448 97453
0 18501 7 1 2 97451 18500
0 18502 5 1 1 18501
0 18503 7 1 2 18497 18502
0 18504 5 1 1 18503
0 18505 7 1 2 65761 18504
0 18506 5 1 1 18505
0 18507 7 2 2 76997 93524
0 18508 7 2 2 72310 92120
0 18509 7 2 2 97455 97457
0 18510 7 1 2 95629 97459
0 18511 5 1 1 18510
0 18512 7 1 2 18506 18511
0 18513 5 1 1 18512
0 18514 7 1 2 64063 18513
0 18515 5 1 1 18514
0 18516 7 1 2 85431 87426
0 18517 7 1 2 97460 18516
0 18518 5 1 1 18517
0 18519 7 1 2 18515 18518
0 18520 5 1 1 18519
0 18521 7 1 2 66710 18520
0 18522 5 1 1 18521
0 18523 7 1 2 76133 92237
0 18524 7 1 2 85406 18523
0 18525 7 7 2 72311 84286
0 18526 7 1 2 97461 95591
0 18527 7 1 2 18524 18526
0 18528 5 1 1 18527
0 18529 7 1 2 18522 18528
0 18530 5 1 1 18529
0 18531 7 1 2 73440 18530
0 18532 5 1 1 18531
0 18533 7 2 2 70402 93643
0 18534 7 1 2 78477 93237
0 18535 7 1 2 97468 18534
0 18536 7 17 2 67104 72312
0 18537 7 5 2 66862 97470
0 18538 7 5 2 65594 84318
0 18539 7 1 2 97487 97492
0 18540 7 1 2 18535 18539
0 18541 5 1 1 18540
0 18542 7 1 2 18532 18541
0 18543 5 1 1 18542
0 18544 7 1 2 74645 18543
0 18545 5 1 1 18544
0 18546 7 2 2 82848 94879
0 18547 5 4 1 97497
0 18548 7 1 2 87049 97499
0 18549 5 1 1 18548
0 18550 7 1 2 68627 89073
0 18551 5 3 1 18550
0 18552 7 1 2 85680 93447
0 18553 5 1 1 18552
0 18554 7 1 2 97503 18553
0 18555 5 1 1 18554
0 18556 7 1 2 73072 18555
0 18557 5 1 1 18556
0 18558 7 1 2 18549 18557
0 18559 5 1 1 18558
0 18560 7 1 2 69480 18559
0 18561 5 1 1 18560
0 18562 7 1 2 81713 95044
0 18563 5 1 1 18562
0 18564 7 2 2 82849 18563
0 18565 5 3 1 97506
0 18566 7 2 2 66711 78593
0 18567 7 3 2 65378 75371
0 18568 5 1 1 97513
0 18569 7 1 2 97511 97514
0 18570 5 1 1 18569
0 18571 7 1 2 97507 18570
0 18572 5 1 1 18571
0 18573 7 1 2 68008 18572
0 18574 5 1 1 18573
0 18575 7 4 2 88675 74779
0 18576 5 1 1 97516
0 18577 7 1 2 75372 97517
0 18578 5 1 1 18577
0 18579 7 1 2 18574 18578
0 18580 5 1 1 18579
0 18581 7 1 2 78379 18580
0 18582 5 1 1 18581
0 18583 7 1 2 18561 18582
0 18584 5 1 1 18583
0 18585 7 2 2 68831 97149
0 18586 7 1 2 18584 97520
0 18587 5 1 1 18586
0 18588 7 1 2 73073 97500
0 18589 5 2 1 18588
0 18590 7 1 2 85681 78929
0 18591 5 1 1 18590
0 18592 7 1 2 97522 18591
0 18593 5 1 1 18592
0 18594 7 1 2 71042 18593
0 18595 5 1 1 18594
0 18596 7 1 2 81234 97508
0 18597 5 2 1 18596
0 18598 7 2 2 73074 78594
0 18599 7 1 2 94656 97526
0 18600 5 1 1 18599
0 18601 7 1 2 87171 18600
0 18602 5 1 1 18601
0 18603 7 1 2 75373 18602
0 18604 5 1 1 18603
0 18605 7 1 2 97524 18604
0 18606 7 1 2 18595 18605
0 18607 5 1 1 18606
0 18608 7 1 2 81340 18607
0 18609 5 1 1 18608
0 18610 7 1 2 77419 96611
0 18611 5 1 1 18610
0 18612 7 1 2 75564 87164
0 18613 5 1 1 18612
0 18614 7 1 2 18611 18613
0 18615 5 1 1 18614
0 18616 7 1 2 75374 18615
0 18617 5 1 1 18616
0 18618 7 7 2 65379 94468
0 18619 5 2 1 97528
0 18620 7 1 2 88458 97529
0 18621 5 2 1 18620
0 18622 7 7 2 68358 80692
0 18623 5 4 1 97539
0 18624 7 1 2 69481 97540
0 18625 5 2 1 18624
0 18626 7 7 2 71043 71806
0 18627 5 1 1 97552
0 18628 7 6 2 70403 97553
0 18629 7 1 2 73724 97559
0 18630 5 1 1 18629
0 18631 7 1 2 97550 18630
0 18632 5 1 1 18631
0 18633 7 1 2 73075 18632
0 18634 5 1 1 18633
0 18635 7 1 2 97537 18634
0 18636 7 1 2 18617 18635
0 18637 5 1 1 18636
0 18638 7 1 2 80189 18637
0 18639 5 1 1 18638
0 18640 7 1 2 18609 18639
0 18641 5 1 1 18640
0 18642 7 1 2 66863 18641
0 18643 5 1 1 18642
0 18644 7 1 2 18587 18643
0 18645 5 1 1 18644
0 18646 7 1 2 67612 18645
0 18647 5 1 1 18646
0 18648 7 5 2 72313 74380
0 18649 5 1 1 97565
0 18650 7 2 2 68628 75176
0 18651 5 1 1 97570
0 18652 7 1 2 78104 18651
0 18653 5 2 1 18652
0 18654 7 1 2 63781 97572
0 18655 5 1 1 18654
0 18656 7 1 2 87768 89674
0 18657 5 1 1 18656
0 18658 7 1 2 18655 18657
0 18659 5 1 1 18658
0 18660 7 2 2 87103 18659
0 18661 7 1 2 79809 97574
0 18662 5 1 1 18661
0 18663 7 1 2 80050 97530
0 18664 7 1 2 97521 18663
0 18665 5 1 1 18664
0 18666 7 1 2 18662 18665
0 18667 5 1 1 18666
0 18668 7 1 2 82577 18667
0 18669 5 1 1 18668
0 18670 7 3 2 77143 87427
0 18671 7 1 2 92121 97518
0 18672 7 1 2 97576 18671
0 18673 5 1 1 18672
0 18674 7 1 2 18669 18673
0 18675 5 1 1 18674
0 18676 7 1 2 75375 18675
0 18677 5 1 1 18676
0 18678 7 1 2 87351 82850
0 18679 5 2 1 18678
0 18680 7 1 2 71044 96223
0 18681 7 1 2 97257 18680
0 18682 7 1 2 97579 18681
0 18683 5 1 1 18682
0 18684 7 1 2 18677 18683
0 18685 5 1 1 18684
0 18686 7 1 2 72630 18685
0 18687 5 1 1 18686
0 18688 7 1 2 97566 18687
0 18689 7 1 2 18647 18688
0 18690 5 1 1 18689
0 18691 7 2 2 79516 94975
0 18692 7 2 2 96047 97581
0 18693 7 1 2 97501 97583
0 18694 5 1 1 18693
0 18695 7 8 2 70629 72149
0 18696 7 3 2 97585 93845
0 18697 7 1 2 78595 97593
0 18698 5 1 1 18697
0 18699 7 1 2 78105 18698
0 18700 5 1 1 18699
0 18701 7 1 2 65380 18700
0 18702 5 1 1 18701
0 18703 7 3 2 94802 78071
0 18704 5 1 1 97596
0 18705 7 1 2 18702 18704
0 18706 5 1 1 18705
0 18707 7 1 2 75376 18706
0 18708 5 1 1 18707
0 18709 7 1 2 75177 97580
0 18710 5 1 1 18709
0 18711 7 1 2 18708 18710
0 18712 5 1 1 18711
0 18713 7 1 2 95540 18712
0 18714 5 1 1 18713
0 18715 7 5 2 81714 75377
0 18716 5 2 1 97599
0 18717 7 1 2 97600 95802
0 18718 5 1 1 18717
0 18719 7 2 2 82851 18718
0 18720 5 3 1 97606
0 18721 7 2 2 91485 77033
0 18722 7 1 2 68832 97611
0 18723 7 1 2 97608 18722
0 18724 5 1 1 18723
0 18725 7 1 2 18714 18724
0 18726 5 1 1 18725
0 18727 7 1 2 65967 18726
0 18728 5 1 1 18727
0 18729 7 1 2 86669 84937
0 18730 7 2 2 80228 18729
0 18731 5 1 1 97613
0 18732 7 1 2 65968 97614
0 18733 5 1 1 18732
0 18734 7 4 2 66517 85682
0 18735 5 2 1 97615
0 18736 7 1 2 65060 97616
0 18737 7 1 2 93525 18736
0 18738 5 1 1 18737
0 18739 7 1 2 18733 18738
0 18740 5 1 1 18739
0 18741 7 2 2 97150 18740
0 18742 5 1 1 97621
0 18743 7 1 2 68833 97622
0 18744 5 1 1 18743
0 18745 7 1 2 18728 18744
0 18746 5 1 1 18745
0 18747 7 1 2 73076 18746
0 18748 5 1 1 18747
0 18749 7 1 2 18694 18748
0 18750 5 1 1 18749
0 18751 7 1 2 74381 18750
0 18752 5 1 1 18751
0 18753 7 1 2 68359 82680
0 18754 5 1 1 18753
0 18755 7 1 2 81117 18754
0 18756 5 6 1 18755
0 18757 7 1 2 80592 97623
0 18758 5 2 1 18757
0 18759 7 2 2 66712 93441
0 18760 7 1 2 83787 97631
0 18761 5 1 1 18760
0 18762 7 1 2 97629 18761
0 18763 5 1 1 18762
0 18764 7 1 2 97612 18763
0 18765 5 1 1 18764
0 18766 7 1 2 18742 18765
0 18767 5 1 1 18766
0 18768 7 1 2 68834 18767
0 18769 5 1 1 18768
0 18770 7 1 2 76680 97594
0 18771 5 1 1 18770
0 18772 7 1 2 94435 78072
0 18773 5 1 1 18772
0 18774 7 1 2 18771 18773
0 18775 5 1 1 18774
0 18776 7 1 2 75378 18775
0 18777 5 1 1 18776
0 18778 7 1 2 83455 88436
0 18779 5 1 1 18778
0 18780 7 1 2 75803 97586
0 18781 7 1 2 18779 18780
0 18782 5 1 1 18781
0 18783 7 1 2 18777 18782
0 18784 5 1 1 18783
0 18785 7 1 2 65969 18784
0 18786 5 1 1 18785
0 18787 7 1 2 77727 96198
0 18788 7 1 2 87968 18787
0 18789 5 1 1 18788
0 18790 7 1 2 18786 18789
0 18791 5 1 1 18790
0 18792 7 1 2 95541 18791
0 18793 5 1 1 18792
0 18794 7 1 2 18769 18793
0 18795 5 1 1 18794
0 18796 7 1 2 73077 18795
0 18797 5 1 1 18796
0 18798 7 1 2 97609 97584
0 18799 5 1 1 18798
0 18800 7 1 2 74420 18799
0 18801 7 1 2 18797 18800
0 18802 5 1 1 18801
0 18803 7 1 2 72314 18802
0 18804 5 1 1 18803
0 18805 7 1 2 18752 18804
0 18806 5 1 1 18805
0 18807 7 1 2 82486 18806
0 18808 7 1 2 18690 18807
0 18809 5 1 1 18808
0 18810 7 2 2 84065 91128
0 18811 7 2 2 68360 82381
0 18812 7 2 2 97635 92122
0 18813 7 1 2 97633 97637
0 18814 5 1 1 18813
0 18815 7 1 2 89675 77034
0 18816 7 1 2 97624 18815
0 18817 5 1 1 18816
0 18818 7 1 2 18814 18817
0 18819 5 1 1 18818
0 18820 7 1 2 73078 18819
0 18821 5 1 1 18820
0 18822 7 1 2 83555 2886
0 18823 5 1 1 18822
0 18824 7 2 2 65970 87961
0 18825 7 1 2 97639 77760
0 18826 7 1 2 18823 18825
0 18827 5 1 1 18826
0 18828 7 1 2 18821 18827
0 18829 5 1 1 18828
0 18830 7 1 2 85481 18829
0 18831 5 1 1 18830
0 18832 7 2 2 77420 77770
0 18833 7 1 2 76981 97641
0 18834 5 1 1 18833
0 18835 7 2 2 77144 84066
0 18836 7 1 2 80866 92123
0 18837 7 1 2 97643 18836
0 18838 5 1 1 18837
0 18839 7 1 2 18834 18838
0 18840 5 1 1 18839
0 18841 7 1 2 68361 18840
0 18842 5 1 1 18841
0 18843 7 2 2 83183 84067
0 18844 7 1 2 89352 91635
0 18845 7 1 2 97645 18844
0 18846 5 1 1 18845
0 18847 7 1 2 18842 18846
0 18848 5 1 1 18847
0 18849 7 1 2 68009 18848
0 18850 5 1 1 18849
0 18851 7 3 2 80881 95513
0 18852 7 1 2 97647 75864
0 18853 7 1 2 96192 18852
0 18854 5 1 1 18853
0 18855 7 1 2 18850 18854
0 18856 5 1 1 18855
0 18857 7 1 2 74382 18856
0 18858 5 1 1 18857
0 18859 7 1 2 18831 18858
0 18860 5 1 1 18859
0 18861 7 1 2 72631 18860
0 18862 5 1 1 18861
0 18863 7 1 2 87050 81307
0 18864 5 2 1 18863
0 18865 7 2 2 65061 76619
0 18866 5 2 1 97652
0 18867 7 2 2 73441 77421
0 18868 7 1 2 65062 80888
0 18869 5 2 1 18868
0 18870 7 1 2 97656 97658
0 18871 5 1 1 18870
0 18872 7 1 2 97654 18871
0 18873 5 5 1 18872
0 18874 7 1 2 73079 97660
0 18875 5 1 1 18874
0 18876 7 1 2 97650 18875
0 18877 5 1 1 18876
0 18878 7 1 2 75678 18877
0 18879 5 1 1 18878
0 18880 7 1 2 2324 81381
0 18881 5 2 1 18880
0 18882 7 1 2 81023 97151
0 18883 7 1 2 97665 18882
0 18884 5 1 1 18883
0 18885 7 1 2 18879 18884
0 18886 5 1 1 18885
0 18887 7 1 2 78536 18886
0 18888 5 1 1 18887
0 18889 7 1 2 18862 18888
0 18890 5 1 1 18889
0 18891 7 1 2 68835 18890
0 18892 5 1 1 18891
0 18893 7 5 2 68629 85482
0 18894 7 2 2 72632 97625
0 18895 7 1 2 97667 97672
0 18896 5 1 1 18895
0 18897 7 2 2 67613 97661
0 18898 7 1 2 74383 97674
0 18899 5 1 1 18898
0 18900 7 1 2 18896 18899
0 18901 5 1 1 18900
0 18902 7 1 2 73080 18901
0 18903 5 1 1 18902
0 18904 7 2 2 96863 92418
0 18905 7 1 2 10221 78445
0 18906 5 6 1 18905
0 18907 7 4 2 68362 97678
0 18908 7 2 2 68010 97684
0 18909 7 1 2 97676 97688
0 18910 5 1 1 18909
0 18911 7 1 2 18903 18910
0 18912 5 1 1 18911
0 18913 7 3 2 63782 75665
0 18914 7 1 2 97690 97587
0 18915 7 1 2 18912 18914
0 18916 5 1 1 18915
0 18917 7 1 2 18892 18916
0 18918 5 1 1 18917
0 18919 7 1 2 72315 18918
0 18920 5 1 1 18919
0 18921 7 8 2 67260 74384
0 18922 7 2 2 72633 97693
0 18923 7 4 2 66864 81341
0 18924 7 1 2 97626 97703
0 18925 5 1 1 18924
0 18926 7 2 2 97237 79680
0 18927 7 1 2 97638 97707
0 18928 5 1 1 18927
0 18929 7 1 2 18925 18928
0 18930 5 1 1 18929
0 18931 7 1 2 73081 18930
0 18932 5 1 1 18931
0 18933 7 1 2 83563 77747
0 18934 7 1 2 97582 18933
0 18935 5 1 1 18934
0 18936 7 1 2 18932 18935
0 18937 5 1 1 18936
0 18938 7 1 2 97701 18937
0 18939 5 1 1 18938
0 18940 7 1 2 18920 18939
0 18941 5 1 1 18940
0 18942 7 1 2 81851 18941
0 18943 5 1 1 18942
0 18944 7 1 2 92598 97155
0 18945 5 1 1 18944
0 18946 7 2 2 65595 87578
0 18947 5 1 1 97709
0 18948 7 1 2 76681 75178
0 18949 5 1 1 18948
0 18950 7 1 2 18947 18949
0 18951 5 1 1 18950
0 18952 7 1 2 63783 18951
0 18953 5 1 1 18952
0 18954 7 1 2 68363 87772
0 18955 5 1 1 18954
0 18956 7 1 2 18953 18955
0 18957 5 1 1 18956
0 18958 7 1 2 85842 18957
0 18959 5 1 1 18958
0 18960 7 1 2 18945 18959
0 18961 5 1 1 18960
0 18962 7 1 2 71045 18961
0 18963 5 1 1 18962
0 18964 7 2 2 67105 89122
0 18965 7 1 2 79725 79659
0 18966 5 2 1 18965
0 18967 7 13 2 71935 68011
0 18968 7 2 2 76682 97715
0 18969 7 1 2 68836 79676
0 18970 7 1 2 97728 18969
0 18971 5 1 1 18970
0 18972 7 1 2 97713 18971
0 18973 5 1 1 18972
0 18974 7 1 2 97711 18973
0 18975 5 1 1 18974
0 18976 7 1 2 18963 18975
0 18977 5 1 1 18976
0 18978 7 1 2 97028 18977
0 18979 5 1 1 18978
0 18980 7 1 2 92477 97729
0 18981 5 1 1 18980
0 18982 7 1 2 97714 18981
0 18983 5 1 1 18982
0 18984 7 19 2 65971 67261
0 18985 5 1 1 97730
0 18986 7 9 2 72634 97731
0 18987 5 1 1 97749
0 18988 7 1 2 97750 74453
0 18989 7 1 2 18983 18988
0 18990 5 1 1 18989
0 18991 7 1 2 18979 18990
0 18992 5 1 1 18991
0 18993 7 1 2 65762 18992
0 18994 5 1 1 18993
0 18995 7 2 2 97295 97488
0 18996 7 1 2 77061 79388
0 18997 7 1 2 97758 18996
0 18998 5 1 1 18997
0 18999 7 1 2 18994 18998
0 19000 5 1 1 18999
0 19001 7 1 2 64064 19000
0 19002 5 1 1 19001
0 19003 7 1 2 65596 93249
0 19004 7 1 2 95574 19003
0 19005 7 1 2 97759 19004
0 19006 5 1 1 19005
0 19007 7 1 2 19002 19006
0 19008 5 1 1 19007
0 19009 7 1 2 84825 19008
0 19010 5 1 1 19009
0 19011 7 1 2 72043 19010
0 19012 7 1 2 18943 19011
0 19013 7 1 2 18809 19012
0 19014 7 1 2 18545 19013
0 19015 5 1 1 19014
0 19016 7 2 2 75506 84548
0 19017 5 2 1 97760
0 19018 7 1 2 84142 97312
0 19019 5 1 1 19018
0 19020 7 1 2 97762 19019
0 19021 5 1 1 19020
0 19022 7 1 2 67614 19021
0 19023 5 1 1 19022
0 19024 7 1 2 77111 79810
0 19025 5 1 1 19024
0 19026 7 1 2 64368 19025
0 19027 5 1 1 19026
0 19028 7 1 2 85006 19027
0 19029 5 1 1 19028
0 19030 7 1 2 19023 19029
0 19031 5 1 1 19030
0 19032 7 1 2 71807 19031
0 19033 5 1 1 19032
0 19034 7 2 2 68012 75134
0 19035 7 1 2 81465 97764
0 19036 5 1 1 19035
0 19037 7 7 2 65381 67615
0 19038 5 1 1 97766
0 19039 7 1 2 76998 88877
0 19040 5 1 1 19039
0 19041 7 1 2 86366 90471
0 19042 7 1 2 84549 19041
0 19043 5 1 1 19042
0 19044 7 1 2 19040 19043
0 19045 5 1 1 19044
0 19046 7 1 2 97767 19045
0 19047 5 1 1 19046
0 19048 7 1 2 19036 19047
0 19049 7 1 2 19033 19048
0 19050 5 1 1 19049
0 19051 7 1 2 71046 19050
0 19052 5 1 1 19051
0 19053 7 5 2 70404 80464
0 19054 5 4 1 97773
0 19055 7 2 2 74849 85007
0 19056 7 1 2 97774 97782
0 19057 5 2 1 19056
0 19058 7 2 2 80593 78642
0 19059 5 1 1 97786
0 19060 7 1 2 79726 97787
0 19061 5 1 1 19060
0 19062 7 4 2 73725 84550
0 19063 7 1 2 81715 97788
0 19064 5 1 1 19063
0 19065 7 1 2 19061 19064
0 19066 5 2 1 19065
0 19067 7 1 2 67616 97792
0 19068 5 1 1 19067
0 19069 7 1 2 97784 19068
0 19070 5 1 1 19069
0 19071 7 1 2 83184 19070
0 19072 5 1 1 19071
0 19073 7 1 2 19052 19072
0 19074 5 1 1 19073
0 19075 7 1 2 74385 19074
0 19076 5 1 1 19075
0 19077 7 2 2 83498 79727
0 19078 7 1 2 78643 97794
0 19079 5 1 1 19078
0 19080 7 1 2 81221 19079
0 19081 5 1 1 19080
0 19082 7 1 2 70405 19081
0 19083 5 2 1 19082
0 19084 7 1 2 64369 93966
0 19085 5 1 1 19084
0 19086 7 1 2 97796 19085
0 19087 5 1 1 19086
0 19088 7 1 2 72635 19087
0 19089 5 1 1 19088
0 19090 7 2 2 64370 87793
0 19091 5 1 1 97798
0 19092 7 1 2 83092 85008
0 19093 5 1 1 19092
0 19094 7 1 2 19091 19093
0 19095 5 1 1 19094
0 19096 7 1 2 83063 19095
0 19097 5 1 1 19096
0 19098 7 1 2 19089 19097
0 19099 5 1 1 19098
0 19100 7 1 2 85483 19099
0 19101 5 1 1 19100
0 19102 7 5 2 80344 81435
0 19103 5 1 1 97800
0 19104 7 2 2 68364 97801
0 19105 5 2 1 97805
0 19106 7 1 2 67617 97677
0 19107 7 1 2 97806 19106
0 19108 5 1 1 19107
0 19109 7 1 2 19101 19108
0 19110 5 1 1 19109
0 19111 7 1 2 65972 19110
0 19112 5 1 1 19111
0 19113 7 1 2 19076 19112
0 19114 5 1 1 19113
0 19115 7 1 2 72316 19114
0 19116 5 1 1 19115
0 19117 7 2 2 83724 97694
0 19118 7 1 2 70148 97793
0 19119 5 1 1 19118
0 19120 7 1 2 64371 86785
0 19121 5 1 1 19120
0 19122 7 1 2 19119 19121
0 19123 5 1 1 19122
0 19124 7 1 2 97809 19123
0 19125 5 1 1 19124
0 19126 7 1 2 19116 19125
0 19127 5 1 1 19126
0 19128 7 1 2 87267 19127
0 19129 5 1 1 19128
0 19130 7 1 2 80594 77121
0 19131 5 2 1 19130
0 19132 7 2 2 88769 97811
0 19133 5 2 1 97813
0 19134 7 1 2 68013 97815
0 19135 5 1 1 19134
0 19136 7 3 2 80693 82025
0 19137 5 1 1 97817
0 19138 7 1 2 87556 19137
0 19139 7 1 2 19135 19138
0 19140 5 3 1 19139
0 19141 7 1 2 78537 97820
0 19142 5 1 1 19141
0 19143 7 3 2 93808 94263
0 19144 5 4 1 97823
0 19145 7 1 2 83077 97824
0 19146 5 2 1 19145
0 19147 7 4 2 73442 97830
0 19148 7 2 2 85484 82242
0 19149 7 1 2 97832 97836
0 19150 5 1 1 19149
0 19151 7 1 2 19142 19150
0 19152 5 2 1 19151
0 19153 7 1 2 75179 97838
0 19154 5 1 1 19153
0 19155 7 2 2 73443 85485
0 19156 7 2 2 86211 96524
0 19157 7 1 2 97840 97842
0 19158 5 1 1 19157
0 19159 7 1 2 86786 78538
0 19160 5 1 1 19159
0 19161 7 1 2 19158 19160
0 19162 5 2 1 19161
0 19163 7 1 2 78088 97844
0 19164 5 1 1 19163
0 19165 7 1 2 19154 19164
0 19166 5 1 1 19165
0 19167 7 1 2 68837 19166
0 19168 5 1 1 19167
0 19169 7 2 2 79375 84195
0 19170 5 1 1 97846
0 19171 7 1 2 97845 97847
0 19172 5 1 1 19171
0 19173 7 1 2 19168 19172
0 19174 5 1 1 19173
0 19175 7 1 2 72317 19174
0 19176 5 1 1 19175
0 19177 7 3 2 86212 95289
0 19178 7 2 2 97695 97848
0 19179 7 1 2 78106 18177
0 19180 5 1 1 19179
0 19181 7 1 2 68838 19180
0 19182 5 1 1 19181
0 19183 7 1 2 19170 19182
0 19184 5 1 1 19183
0 19185 7 1 2 65382 19184
0 19186 5 1 1 19185
0 19187 7 1 2 74646 87275
0 19188 5 1 1 19187
0 19189 7 1 2 19186 19188
0 19190 5 1 1 19189
0 19191 7 1 2 97851 19190
0 19192 5 1 1 19191
0 19193 7 1 2 19176 19192
0 19194 5 1 1 19193
0 19195 7 1 2 81024 19194
0 19196 5 1 1 19195
0 19197 7 4 2 70785 77422
0 19198 5 5 1 97853
0 19199 7 3 2 65763 77208
0 19200 5 6 1 97862
0 19201 7 18 2 97857 97865
0 19202 7 3 2 72318 97871
0 19203 7 1 2 97889 97821
0 19204 5 1 1 19203
0 19205 7 25 2 65764 67262
0 19206 5 9 1 97892
0 19207 7 3 2 97893 77326
0 19208 7 8 2 86022 80508
0 19209 5 4 1 97929
0 19210 7 4 2 68014 97937
0 19211 5 2 1 97941
0 19212 7 1 2 97926 97942
0 19213 5 1 1 19212
0 19214 7 1 2 19204 19213
0 19215 5 1 1 19214
0 19216 7 1 2 72636 19215
0 19217 5 1 1 19216
0 19218 7 2 2 66713 75139
0 19219 5 1 1 97947
0 19220 7 1 2 93938 19219
0 19221 5 1 1 19220
0 19222 7 1 2 97890 19221
0 19223 5 1 1 19222
0 19224 7 10 2 67263 73726
0 19225 5 1 1 97949
0 19226 7 1 2 66714 97950
0 19227 7 1 2 96101 19226
0 19228 5 1 1 19227
0 19229 7 1 2 19223 19228
0 19230 5 1 1 19229
0 19231 7 1 2 92256 19230
0 19232 5 1 1 19231
0 19233 7 1 2 19217 19232
0 19234 5 1 1 19233
0 19235 7 1 2 64065 19234
0 19236 5 1 1 19235
0 19237 7 10 2 65765 72319
0 19238 5 1 1 97959
0 19239 7 3 2 97960 78288
0 19240 5 1 1 97969
0 19241 7 1 2 72637 97822
0 19242 5 1 1 19241
0 19243 7 1 2 97831 92257
0 19244 5 1 1 19243
0 19245 7 1 2 19242 19244
0 19246 5 2 1 19245
0 19247 7 1 2 97970 97972
0 19248 5 1 1 19247
0 19249 7 1 2 19236 19248
0 19250 5 1 1 19249
0 19251 7 1 2 87276 19250
0 19252 5 1 1 19251
0 19253 7 1 2 19196 19252
0 19254 7 1 2 19129 19253
0 19255 5 1 1 19254
0 19256 7 1 2 71936 19255
0 19257 5 1 1 19256
0 19258 7 1 2 97263 81025
0 19259 5 1 1 19258
0 19260 7 2 2 72638 92365
0 19261 7 1 2 90216 97974
0 19262 5 1 1 19261
0 19263 7 2 2 19259 19262
0 19264 7 1 2 81528 87161
0 19265 5 1 1 19264
0 19266 7 1 2 97976 19265
0 19267 5 1 1 19266
0 19268 7 1 2 65766 19267
0 19269 5 1 1 19268
0 19270 7 4 2 66518 92577
0 19271 7 2 2 77062 95256
0 19272 5 1 1 97982
0 19273 7 1 2 97978 97983
0 19274 5 1 1 19273
0 19275 7 1 2 19269 19274
0 19276 5 1 1 19275
0 19277 7 1 2 84774 19276
0 19278 5 1 1 19277
0 19279 7 2 2 64066 84900
0 19280 5 1 1 97984
0 19281 7 1 2 75565 82215
0 19282 7 1 2 97858 19281
0 19283 5 1 1 19282
0 19284 7 1 2 97977 19283
0 19285 5 1 1 19284
0 19286 7 1 2 97985 19285
0 19287 5 1 1 19286
0 19288 7 2 2 65383 80314
0 19289 7 1 2 74188 95310
0 19290 7 1 2 97986 19289
0 19291 7 1 2 97313 19290
0 19292 5 1 1 19291
0 19293 7 1 2 19287 19292
0 19294 7 1 2 19278 19293
0 19295 5 1 1 19294
0 19296 7 1 2 65063 19295
0 19297 5 1 1 19296
0 19298 7 4 2 64372 84174
0 19299 7 1 2 80808 97988
0 19300 5 1 1 19299
0 19301 7 1 2 82701 19300
0 19302 5 1 1 19301
0 19303 7 1 2 73082 19302
0 19304 5 1 1 19303
0 19305 7 1 2 91129 80315
0 19306 7 1 2 83613 19305
0 19307 5 1 1 19306
0 19308 7 1 2 19304 19307
0 19309 5 1 1 19308
0 19310 7 1 2 70406 19309
0 19311 5 1 1 19310
0 19312 7 1 2 82593 75652
0 19313 5 1 1 19312
0 19314 7 1 2 82693 96625
0 19315 7 1 2 19313 19314
0 19316 5 1 1 19315
0 19317 7 1 2 19311 19316
0 19318 5 1 1 19317
0 19319 7 1 2 67618 19318
0 19320 5 1 1 19319
0 19321 7 2 2 83987 81026
0 19322 5 1 1 97992
0 19323 7 1 2 96656 97993
0 19324 5 1 1 19323
0 19325 7 1 2 19320 19324
0 19326 5 1 1 19325
0 19327 7 1 2 65767 19326
0 19328 5 1 1 19327
0 19329 7 1 2 19297 19328
0 19330 5 1 1 19329
0 19331 7 1 2 72320 19330
0 19332 5 1 1 19331
0 19333 7 2 2 96736 83360
0 19334 5 1 1 97994
0 19335 7 2 2 64067 97859
0 19336 5 1 1 97996
0 19337 7 5 2 64373 93250
0 19338 5 1 1 97998
0 19339 7 1 2 19336 19338
0 19340 5 5 1 19339
0 19341 7 1 2 89787 98003
0 19342 5 1 1 19341
0 19343 7 2 2 82911 79785
0 19344 7 1 2 95302 98008
0 19345 5 1 1 19344
0 19346 7 1 2 19342 19345
0 19347 5 1 1 19346
0 19348 7 1 2 97995 19347
0 19349 5 1 1 19348
0 19350 7 1 2 19332 19349
0 19351 5 1 1 19350
0 19352 7 7 2 65597 77771
0 19353 7 1 2 82762 98010
0 19354 7 1 2 19351 19353
0 19355 5 1 1 19354
0 19356 7 1 2 66979 19355
0 19357 7 1 2 19257 19356
0 19358 5 1 1 19357
0 19359 7 1 2 73851 19358
0 19360 7 1 2 19015 19359
0 19361 5 1 1 19360
0 19362 7 25 2 72321 68015
0 19363 7 2 2 73444 86421
0 19364 7 1 2 63898 89575
0 19365 5 1 1 19364
0 19366 7 1 2 73852 78073
0 19367 5 1 1 19366
0 19368 7 1 2 19365 19367
0 19369 5 4 1 19368
0 19370 7 3 2 67106 98044
0 19371 7 2 2 67619 98048
0 19372 7 1 2 98042 98051
0 19373 5 1 1 19372
0 19374 7 3 2 81414 75820
0 19375 7 1 2 91659 96697
0 19376 7 1 2 97247 19375
0 19377 7 1 2 98053 19376
0 19378 5 1 1 19377
0 19379 7 1 2 19373 19378
0 19380 5 1 1 19379
0 19381 7 1 2 74060 19380
0 19382 5 1 1 19381
0 19383 7 3 2 70786 82382
0 19384 7 1 2 98056 96509
0 19385 7 1 2 91276 98054
0 19386 7 1 2 19384 19385
0 19387 5 1 1 19386
0 19388 7 1 2 19382 19387
0 19389 5 1 1 19388
0 19390 7 1 2 64068 19389
0 19391 5 1 1 19390
0 19392 7 1 2 93728 92419
0 19393 7 1 2 94148 19392
0 19394 7 1 2 91409 98055
0 19395 7 1 2 19393 19394
0 19396 5 1 1 19395
0 19397 7 1 2 19391 19396
0 19398 5 1 1 19397
0 19399 7 1 2 84448 19398
0 19400 5 1 1 19399
0 19401 7 2 2 93138 92556
0 19402 7 1 2 76903 92904
0 19403 7 1 2 98059 19402
0 19404 7 1 2 96367 19403
0 19405 5 1 1 19404
0 19406 7 1 2 19400 19405
0 19407 5 1 1 19406
0 19408 7 1 2 68839 19407
0 19409 5 1 1 19408
0 19410 7 2 2 75749 89420
0 19411 7 2 2 70675 66519
0 19412 7 1 2 98061 98063
0 19413 5 1 1 19412
0 19414 7 2 2 88890 78111
0 19415 7 1 2 72044 98065
0 19416 5 1 1 19415
0 19417 7 1 2 19413 19416
0 19418 5 1 1 19417
0 19419 7 1 2 96672 19418
0 19420 5 1 1 19419
0 19421 7 2 2 75821 91255
0 19422 7 3 2 63976 70676
0 19423 7 1 2 77501 98069
0 19424 7 1 2 98067 19423
0 19425 5 1 1 19424
0 19426 7 3 2 69065 70407
0 19427 7 1 2 73826 79314
0 19428 7 1 2 98072 19427
0 19429 7 1 2 75771 19428
0 19430 5 1 1 19429
0 19431 7 1 2 19425 19430
0 19432 7 1 2 19420 19431
0 19433 5 1 1 19432
0 19434 7 1 2 70630 19433
0 19435 5 1 1 19434
0 19436 7 1 2 76904 85187
0 19437 7 1 2 90250 19436
0 19438 5 1 1 19437
0 19439 7 1 2 19435 19438
0 19440 5 1 1 19439
0 19441 7 2 2 74061 81395
0 19442 7 1 2 93765 98075
0 19443 7 1 2 19440 19442
0 19444 5 1 1 19443
0 19445 7 1 2 19409 19444
0 19446 5 1 1 19445
0 19447 7 1 2 65064 19446
0 19448 5 1 1 19447
0 19449 7 1 2 74029 96368
0 19450 5 2 1 19449
0 19451 7 1 2 79634 96350
0 19452 5 1 1 19451
0 19453 7 1 2 98077 19452
0 19454 5 6 1 19453
0 19455 7 1 2 65384 92859
0 19456 7 1 2 90663 19455
0 19457 7 1 2 98076 19456
0 19458 7 1 2 98079 19457
0 19459 5 1 1 19458
0 19460 7 1 2 19448 19459
0 19461 5 1 1 19460
0 19462 7 1 2 98017 19461
0 19463 5 1 1 19462
0 19464 7 1 2 87830 90211
0 19465 5 1 1 19464
0 19466 7 4 2 74647 77663
0 19467 7 1 2 68840 93574
0 19468 7 1 2 98085 19467
0 19469 7 1 2 92459 19468
0 19470 5 1 1 19469
0 19471 7 1 2 19465 19470
0 19472 5 1 1 19471
0 19473 7 1 2 63899 19472
0 19474 5 1 1 19473
0 19475 7 1 2 97191 98086
0 19476 5 1 1 19475
0 19477 7 1 2 19474 19476
0 19478 5 1 1 19477
0 19479 7 1 2 72322 19478
0 19480 5 1 1 19479
0 19481 7 2 2 96327 98087
0 19482 7 4 2 72045 67264
0 19483 7 5 2 85102 93306
0 19484 7 1 2 98091 98095
0 19485 7 1 2 98089 19484
0 19486 5 1 1 19485
0 19487 7 1 2 19480 19486
0 19488 5 1 1 19487
0 19489 7 1 2 67107 19488
0 19490 5 1 1 19489
0 19491 7 5 2 67265 74648
0 19492 7 1 2 95230 92860
0 19493 7 1 2 98100 19492
0 19494 7 1 2 96390 19493
0 19495 5 1 1 19494
0 19496 7 1 2 19490 19495
0 19497 5 1 1 19496
0 19498 7 1 2 65768 19497
0 19499 5 1 1 19498
0 19500 7 2 2 93594 93307
0 19501 7 1 2 92308 97471
0 19502 7 1 2 98105 19501
0 19503 7 1 2 98090 19502
0 19504 5 1 1 19503
0 19505 7 1 2 19499 19504
0 19506 5 1 1 19505
0 19507 7 1 2 72639 19506
0 19508 5 1 1 19507
0 19509 7 1 2 66980 82487
0 19510 7 1 2 97489 19509
0 19511 7 1 2 84265 19510
0 19512 7 1 2 93544 19511
0 19513 5 1 1 19512
0 19514 7 1 2 19508 19513
0 19515 5 1 1 19514
0 19516 7 1 2 65385 19515
0 19517 5 1 1 19516
0 19518 7 1 2 78644 97163
0 19519 5 1 1 19518
0 19520 7 1 2 89274 97029
0 19521 5 1 1 19520
0 19522 7 1 2 19519 19521
0 19523 5 3 1 19522
0 19524 7 1 2 64069 98107
0 19525 5 1 1 19524
0 19526 7 1 2 85475 19525
0 19527 5 1 1 19526
0 19528 7 8 2 72323 73083
0 19529 7 4 2 98110 97979
0 19530 5 1 1 98118
0 19531 7 1 2 74421 19530
0 19532 5 1 1 19531
0 19533 7 4 2 68986 96429
0 19534 7 5 2 98122 89516
0 19535 7 2 2 74470 85103
0 19536 7 1 2 79765 98131
0 19537 7 1 2 98126 19536
0 19538 7 1 2 19532 19537
0 19539 7 1 2 19527 19538
0 19540 5 1 1 19539
0 19541 7 1 2 19517 19540
0 19542 5 1 1 19541
0 19543 7 1 2 81027 19542
0 19544 5 1 1 19543
0 19545 7 2 2 85486 80935
0 19546 7 6 2 72046 72324
0 19547 7 2 2 98135 91282
0 19548 7 2 2 98133 98141
0 19549 7 1 2 76886 73853
0 19550 7 1 2 98143 19549
0 19551 5 1 1 19550
0 19552 7 6 2 64070 65386
0 19553 7 4 2 65769 98145
0 19554 5 1 1 98151
0 19555 7 1 2 77973 93389
0 19556 5 1 1 19555
0 19557 7 1 2 19554 19556
0 19558 5 1 1 19557
0 19559 7 1 2 98101 19558
0 19560 5 1 1 19559
0 19561 7 7 2 66520 72325
0 19562 7 2 2 82488 77145
0 19563 5 1 1 98162
0 19564 7 1 2 96123 19563
0 19565 5 3 1 19564
0 19566 7 2 2 65065 98164
0 19567 7 1 2 98155 98167
0 19568 5 1 1 19567
0 19569 7 1 2 19560 19568
0 19570 5 1 1 19569
0 19571 7 2 2 73445 74101
0 19572 7 1 2 98169 90788
0 19573 7 1 2 19570 19572
0 19574 5 1 1 19573
0 19575 7 1 2 19551 19574
0 19576 5 1 1 19575
0 19577 7 1 2 63900 19576
0 19578 5 1 1 19577
0 19579 7 1 2 76003 89576
0 19580 7 1 2 98144 19579
0 19581 5 1 1 19580
0 19582 7 1 2 19578 19581
0 19583 5 1 1 19582
0 19584 7 1 2 63784 19583
0 19585 5 1 1 19584
0 19586 7 1 2 72326 75822
0 19587 7 1 2 79611 19586
0 19588 7 1 2 98134 19587
0 19589 7 1 2 96369 19588
0 19590 5 1 1 19589
0 19591 7 1 2 19585 19590
0 19592 5 1 1 19591
0 19593 7 1 2 95414 19592
0 19594 5 1 1 19593
0 19595 7 1 2 68841 96707
0 19596 5 1 1 19595
0 19597 7 1 2 90513 91921
0 19598 5 1 1 19597
0 19599 7 1 2 19596 19598
0 19600 5 1 1 19599
0 19601 7 12 2 67266 73446
0 19602 7 2 2 98171 91283
0 19603 7 1 2 64374 91773
0 19604 7 1 2 98183 19603
0 19605 5 1 1 19604
0 19606 7 1 2 72327 82870
0 19607 7 1 2 77519 19606
0 19608 7 1 2 96469 19607
0 19609 5 1 1 19608
0 19610 7 1 2 19605 19609
0 19611 5 1 1 19610
0 19612 7 1 2 19600 19611
0 19613 5 1 1 19612
0 19614 7 10 2 72328 68365
0 19615 7 5 2 71620 98185
0 19616 7 8 2 71047 67108
0 19617 7 2 2 98195 98200
0 19618 7 1 2 79766 89496
0 19619 7 1 2 98208 19618
0 19620 5 1 1 19619
0 19621 7 1 2 83290 96313
0 19622 7 1 2 98184 19621
0 19623 5 1 1 19622
0 19624 7 1 2 19620 19623
0 19625 5 1 1 19624
0 19626 7 1 2 68842 19625
0 19627 5 1 1 19626
0 19628 7 8 2 63785 70408
0 19629 7 1 2 98210 91386
0 19630 7 1 2 98209 19629
0 19631 5 1 1 19630
0 19632 7 1 2 19627 19631
0 19633 5 1 1 19632
0 19634 7 1 2 96673 19633
0 19635 5 1 1 19634
0 19636 7 1 2 19613 19635
0 19637 5 1 1 19636
0 19638 7 1 2 66981 19637
0 19639 5 1 1 19638
0 19640 7 8 2 64375 97732
0 19641 5 6 1 98218
0 19642 7 14 2 71048 72329
0 19643 7 5 2 69482 98232
0 19644 5 3 1 98246
0 19645 7 1 2 98226 98251
0 19646 5 10 1 19645
0 19647 7 2 2 66521 98254
0 19648 5 1 1 98264
0 19649 7 17 2 67267 77327
0 19650 5 2 1 98266
0 19651 7 9 2 72330 77146
0 19652 7 1 2 65387 96285
0 19653 5 1 1 19652
0 19654 7 1 2 98285 19653
0 19655 5 1 1 19654
0 19656 7 1 2 98283 19655
0 19657 5 1 1 19656
0 19658 7 2 2 65066 19657
0 19659 5 1 1 98294
0 19660 7 1 2 19648 19659
0 19661 5 1 1 19660
0 19662 7 1 2 65639 94735
0 19663 7 1 2 19661 19662
0 19664 5 1 1 19663
0 19665 7 1 2 96909 98295
0 19666 5 1 1 19665
0 19667 7 1 2 19664 19666
0 19668 5 1 1 19667
0 19669 7 1 2 89517 19668
0 19670 5 1 1 19669
0 19671 7 2 2 98255 90673
0 19672 7 1 2 65388 73821
0 19673 7 1 2 98296 19672
0 19674 5 1 1 19673
0 19675 7 1 2 19670 19674
0 19676 5 1 1 19675
0 19677 7 1 2 68987 19676
0 19678 5 1 1 19677
0 19679 7 1 2 91774 96667
0 19680 7 1 2 98297 19679
0 19681 5 1 1 19680
0 19682 7 1 2 19678 19681
0 19683 5 1 1 19682
0 19684 7 1 2 85828 78988
0 19685 7 1 2 19683 19684
0 19686 5 1 1 19685
0 19687 7 1 2 19639 19686
0 19688 5 1 1 19687
0 19689 7 1 2 74386 19688
0 19690 5 1 1 19689
0 19691 7 1 2 93931 96339
0 19692 5 1 1 19691
0 19693 7 1 2 86599 98127
0 19694 5 1 1 19693
0 19695 7 1 2 19692 19694
0 19696 5 1 1 19695
0 19697 7 1 2 81104 98136
0 19698 7 1 2 85487 19697
0 19699 7 1 2 92478 19698
0 19700 7 1 2 19696 19699
0 19701 5 1 1 19700
0 19702 7 1 2 19690 19701
0 19703 5 1 1 19702
0 19704 7 1 2 91702 19703
0 19705 5 1 1 19704
0 19706 7 1 2 19594 19705
0 19707 5 1 1 19706
0 19708 7 1 2 73084 19707
0 19709 5 1 1 19708
0 19710 7 1 2 19544 19709
0 19711 7 1 2 19463 19710
0 19712 5 1 1 19711
0 19713 7 1 2 80406 19712
0 19714 5 1 1 19713
0 19715 7 1 2 72640 94306
0 19716 5 2 1 19715
0 19717 7 1 2 97617 92627
0 19718 5 1 1 19717
0 19719 7 1 2 98298 19718
0 19720 5 1 1 19719
0 19721 7 1 2 71049 19720
0 19722 5 1 1 19721
0 19723 7 1 2 94307 92731
0 19724 5 1 1 19723
0 19725 7 1 2 19722 19724
0 19726 5 1 1 19725
0 19727 7 1 2 85890 19726
0 19728 5 1 1 19727
0 19729 7 5 2 68366 82871
0 19730 7 2 2 84901 98300
0 19731 5 1 1 98305
0 19732 7 1 2 82594 94321
0 19733 5 1 1 19732
0 19734 7 1 2 19731 19733
0 19735 5 1 1 19734
0 19736 7 1 2 92181 19735
0 19737 5 1 1 19736
0 19738 7 1 2 19728 19737
0 19739 5 1 1 19738
0 19740 7 1 2 64071 19739
0 19741 5 1 1 19740
0 19742 7 3 2 83078 83809
0 19743 7 2 2 93802 98307
0 19744 5 1 1 98310
0 19745 7 1 2 73904 98311
0 19746 5 1 1 19745
0 19747 7 1 2 82860 19746
0 19748 5 1 1 19747
0 19749 7 1 2 85256 93526
0 19750 7 1 2 19748 19749
0 19751 5 1 1 19750
0 19752 7 1 2 19741 19751
0 19753 5 1 1 19752
0 19754 7 1 2 88566 19753
0 19755 5 1 1 19754
0 19756 7 1 2 86463 96557
0 19757 5 2 1 19756
0 19758 7 1 2 98312 77328
0 19759 5 1 1 19758
0 19760 7 1 2 19280 19759
0 19761 5 1 1 19760
0 19762 7 1 2 68367 19761
0 19763 5 1 1 19762
0 19764 7 1 2 68630 87068
0 19765 5 1 1 19764
0 19766 7 1 2 94189 19765
0 19767 5 1 1 19766
0 19768 7 1 2 77329 19767
0 19769 5 1 1 19768
0 19770 7 1 2 19763 19769
0 19771 5 1 1 19770
0 19772 7 1 2 85257 19771
0 19773 5 1 1 19772
0 19774 7 2 2 92866 83064
0 19775 5 1 1 98314
0 19776 7 1 2 19775 89076
0 19777 5 1 1 19776
0 19778 7 1 2 93454 19777
0 19779 5 1 1 19778
0 19780 7 1 2 67620 19779
0 19781 7 1 2 19773 19780
0 19782 5 1 1 19781
0 19783 7 1 2 87332 76683
0 19784 5 3 1 19783
0 19785 7 1 2 88378 83569
0 19786 5 3 1 19785
0 19787 7 1 2 98316 98319
0 19788 5 1 1 19787
0 19789 7 1 2 85258 81028
0 19790 7 1 2 19788 19789
0 19791 5 1 1 19790
0 19792 7 3 2 75379 83680
0 19793 5 1 1 98322
0 19794 7 1 2 85891 82694
0 19795 7 1 2 98323 19794
0 19796 5 1 1 19795
0 19797 7 1 2 72641 19796
0 19798 7 1 2 19791 19797
0 19799 5 1 1 19798
0 19800 7 1 2 88205 19799
0 19801 7 1 2 19782 19800
0 19802 5 1 1 19801
0 19803 7 1 2 19755 19802
0 19804 5 1 1 19803
0 19805 7 1 2 65770 19804
0 19806 5 1 1 19805
0 19807 7 5 2 71621 66982
0 19808 7 3 2 63786 98325
0 19809 5 1 1 98330
0 19810 7 4 2 64072 65067
0 19811 7 1 2 98331 98333
0 19812 7 1 2 89458 19811
0 19813 7 1 2 86980 19812
0 19814 7 1 2 93527 19813
0 19815 5 1 1 19814
0 19816 7 1 2 19806 19815
0 19817 5 1 1 19816
0 19818 7 1 2 98018 19817
0 19819 5 1 1 19818
0 19820 7 13 2 69123 65973
0 19821 5 1 1 98337
0 19822 7 1 2 98338 95290
0 19823 5 1 1 19822
0 19824 7 1 2 82695 97768
0 19825 5 1 1 19824
0 19826 7 1 2 19823 19825
0 19827 5 1 1 19826
0 19828 7 2 2 73085 89333
0 19829 7 1 2 19827 98350
0 19830 5 1 1 19829
0 19831 7 1 2 95291 80992
0 19832 5 1 1 19831
0 19833 7 2 2 664 95296
0 19834 5 1 1 98352
0 19835 7 1 2 64376 83737
0 19836 7 1 2 19834 19835
0 19837 5 1 1 19836
0 19838 7 1 2 19832 19837
0 19839 5 1 1 19838
0 19840 7 1 2 93373 19839
0 19841 5 1 1 19840
0 19842 7 1 2 19830 19841
0 19843 5 1 1 19842
0 19844 7 1 2 70149 19843
0 19845 5 1 1 19844
0 19846 7 1 2 93455 81235
0 19847 5 1 1 19846
0 19848 7 1 2 75646 88302
0 19849 7 1 2 89433 19848
0 19850 5 1 1 19849
0 19851 7 1 2 19847 19850
0 19852 5 1 1 19851
0 19853 7 1 2 88206 19852
0 19854 5 1 1 19853
0 19855 7 1 2 80059 98146
0 19856 7 1 2 98351 19855
0 19857 5 1 1 19856
0 19858 7 1 2 19854 19857
0 19859 5 1 1 19858
0 19860 7 1 2 67621 19859
0 19861 5 1 1 19860
0 19862 7 1 2 19845 19861
0 19863 5 1 1 19862
0 19864 7 1 2 72331 19863
0 19865 5 1 1 19864
0 19866 7 1 2 96737 89114
0 19867 7 1 2 74915 92853
0 19868 7 1 2 19866 19867
0 19869 5 1 1 19868
0 19870 7 1 2 19865 19869
0 19871 5 1 1 19870
0 19872 7 1 2 66715 19871
0 19873 5 1 1 19872
0 19874 7 2 2 72332 87794
0 19875 7 1 2 78123 98354
0 19876 7 1 2 92210 19875
0 19877 5 1 1 19876
0 19878 7 1 2 19873 19877
0 19879 5 1 1 19878
0 19880 7 1 2 65771 19879
0 19881 5 1 1 19880
0 19882 7 1 2 96864 87526
0 19883 7 1 2 93595 19882
0 19884 7 5 2 72333 82243
0 19885 7 1 2 98356 93990
0 19886 7 1 2 19883 19885
0 19887 5 1 1 19886
0 19888 7 1 2 19881 19887
0 19889 5 1 1 19888
0 19890 7 1 2 78693 19889
0 19891 5 1 1 19890
0 19892 7 4 2 72642 85488
0 19893 7 1 2 71622 98009
0 19894 5 1 1 19893
0 19895 7 1 2 97630 19894
0 19896 5 1 1 19895
0 19897 7 1 2 98361 19896
0 19898 5 1 1 19897
0 19899 7 1 2 84902 76620
0 19900 5 3 1 19899
0 19901 7 1 2 80959 94230
0 19902 5 2 1 19901
0 19903 7 1 2 82852 98368
0 19904 5 1 1 19903
0 19905 7 1 2 77423 19904
0 19906 5 1 1 19905
0 19907 7 1 2 98365 19906
0 19908 5 1 1 19907
0 19909 7 1 2 78539 19908
0 19910 5 1 1 19909
0 19911 7 1 2 19898 19910
0 19912 5 1 1 19911
0 19913 7 1 2 72334 19912
0 19914 5 1 1 19913
0 19915 7 11 2 72335 68631
0 19916 7 1 2 70787 98370
0 19917 5 1 1 19916
0 19918 7 1 2 97917 19917
0 19919 5 8 1 19918
0 19920 7 1 2 64073 98381
0 19921 5 1 1 19920
0 19922 7 1 2 85432 98371
0 19923 5 1 1 19922
0 19924 7 1 2 19921 19923
0 19925 5 1 1 19924
0 19926 7 1 2 97673 19925
0 19927 5 1 1 19926
0 19928 7 1 2 97567 97675
0 19929 5 1 1 19928
0 19930 7 1 2 19927 19929
0 19931 5 1 1 19930
0 19932 7 1 2 81852 19931
0 19933 5 1 1 19932
0 19934 7 1 2 66716 80960
0 19935 7 1 2 86748 19934
0 19936 5 1 1 19935
0 19937 7 1 2 82853 19936
0 19938 5 1 1 19937
0 19939 7 1 2 19938 97810
0 19940 5 1 1 19939
0 19941 7 1 2 19933 19940
0 19942 7 1 2 19914 19941
0 19943 5 1 1 19942
0 19944 7 1 2 88567 19943
0 19945 5 1 1 19944
0 19946 7 3 2 65974 96738
0 19947 5 4 1 98389
0 19948 7 5 2 71050 97030
0 19949 5 2 1 98396
0 19950 7 1 2 98392 98401
0 19951 5 15 1 19950
0 19952 7 1 2 65772 98403
0 19953 5 1 1 19952
0 19954 7 28 2 70788 72336
0 19955 5 2 1 98418
0 19956 7 7 2 72643 98419
0 19957 5 1 1 98448
0 19958 7 1 2 65975 98449
0 19959 5 1 1 19958
0 19960 7 1 2 19953 19959
0 19961 5 1 1 19960
0 19962 7 1 2 64074 19961
0 19963 5 1 1 19962
0 19964 7 12 2 65976 72337
0 19965 7 2 2 85433 98455
0 19966 7 1 2 72644 98467
0 19967 5 2 1 19966
0 19968 7 1 2 19963 98469
0 19969 5 1 1 19968
0 19970 7 1 2 75380 19969
0 19971 5 1 1 19970
0 19972 7 7 2 72338 83185
0 19973 7 1 2 98471 78540
0 19974 5 1 1 19973
0 19975 7 1 2 19971 19974
0 19976 5 1 1 19975
0 19977 7 1 2 80694 19976
0 19978 5 1 1 19977
0 19979 7 5 2 67622 97961
0 19980 7 1 2 77424 98478
0 19981 5 1 1 19980
0 19982 7 1 2 98446 97918
0 19983 5 33 1 19982
0 19984 7 1 2 98483 83725
0 19985 5 1 1 19984
0 19986 7 1 2 19981 19985
0 19987 5 1 1 19986
0 19988 7 1 2 64075 19987
0 19989 5 1 1 19988
0 19990 7 1 2 98470 19989
0 19991 5 1 1 19990
0 19992 7 1 2 88758 19991
0 19993 5 1 1 19992
0 19994 7 2 2 71808 97031
0 19995 7 1 2 79338 84500
0 19996 7 1 2 98516 19995
0 19997 5 1 1 19996
0 19998 7 1 2 19993 19997
0 19999 7 1 2 19978 19998
0 20000 5 1 1 19999
0 20001 7 1 2 88207 20000
0 20002 5 1 1 20001
0 20003 7 1 2 19945 20002
0 20004 5 1 1 20003
0 20005 7 1 2 85892 20004
0 20006 5 1 1 20005
0 20007 7 1 2 89693 78602
0 20008 5 1 1 20007
0 20009 7 1 2 11535 20008
0 20010 5 1 1 20009
0 20011 7 1 2 65389 20010
0 20012 5 1 1 20011
0 20013 7 1 2 84765 92691
0 20014 5 1 1 20013
0 20015 7 1 2 20012 20014
0 20016 5 1 1 20015
0 20017 7 1 2 20016 98165
0 20018 5 1 1 20017
0 20019 7 10 2 71051 93055
0 20020 5 1 1 98518
0 20021 7 1 2 74422 77330
0 20022 5 1 1 20021
0 20023 7 1 2 20020 20022
0 20024 5 3 1 20023
0 20025 7 1 2 82108 94526
0 20026 7 1 2 98528 20025
0 20027 5 1 1 20026
0 20028 7 1 2 20018 20027
0 20029 5 1 1 20028
0 20030 7 1 2 72645 20029
0 20031 5 1 1 20030
0 20032 7 1 2 85683 88208
0 20033 5 3 1 20032
0 20034 7 1 2 84903 89827
0 20035 5 1 1 20034
0 20036 7 1 2 98531 20035
0 20037 5 1 1 20036
0 20038 7 1 2 82489 20037
0 20039 5 1 1 20038
0 20040 7 2 2 82109 97014
0 20041 7 1 2 93139 98534
0 20042 5 1 1 20041
0 20043 7 1 2 20039 20042
0 20044 5 1 1 20043
0 20045 7 1 2 92893 20044
0 20046 5 1 1 20045
0 20047 7 1 2 20031 20046
0 20048 5 1 1 20047
0 20049 7 1 2 75275 20048
0 20050 5 1 1 20049
0 20051 7 1 2 82399 88303
0 20052 5 1 1 20051
0 20053 7 1 2 82646 82696
0 20054 5 2 1 20053
0 20055 7 1 2 20052 98536
0 20056 5 1 1 20055
0 20057 7 1 2 88568 20056
0 20058 5 1 1 20057
0 20059 7 1 2 65977 93190
0 20060 7 1 2 94308 20059
0 20061 5 1 1 20060
0 20062 7 1 2 20058 20061
0 20063 5 1 1 20062
0 20064 7 1 2 67623 20063
0 20065 5 1 1 20064
0 20066 7 1 2 86670 88569
0 20067 5 1 1 20066
0 20068 7 1 2 88383 88209
0 20069 5 1 1 20068
0 20070 7 1 2 20067 20069
0 20071 5 2 1 20070
0 20072 7 7 2 72646 81029
0 20073 7 1 2 81308 98540
0 20074 7 1 2 98538 20073
0 20075 5 1 1 20074
0 20076 7 1 2 20065 20075
0 20077 5 1 1 20076
0 20078 7 1 2 65773 20077
0 20079 5 1 1 20078
0 20080 7 1 2 20050 20079
0 20081 5 1 1 20080
0 20082 7 1 2 72339 20081
0 20083 5 1 1 20082
0 20084 7 1 2 89788 88570
0 20085 5 1 1 20084
0 20086 7 1 2 98532 20085
0 20087 5 1 1 20086
0 20088 7 1 2 20087 98004
0 20089 5 1 1 20088
0 20090 7 2 2 83394 89459
0 20091 5 1 1 98547
0 20092 7 1 2 77331 93140
0 20093 7 1 2 98548 20092
0 20094 5 1 1 20093
0 20095 7 1 2 20089 20094
0 20096 5 1 1 20095
0 20097 7 7 2 66522 67268
0 20098 7 5 2 65068 72647
0 20099 7 1 2 98549 98556
0 20100 7 1 2 20096 20099
0 20101 5 1 1 20100
0 20102 7 1 2 20083 20101
0 20103 5 1 1 20102
0 20104 7 1 2 85259 20103
0 20105 5 1 1 20104
0 20106 7 1 2 20006 20105
0 20107 5 1 1 20106
0 20108 7 1 2 73086 20107
0 20109 5 1 1 20108
0 20110 7 1 2 19891 20109
0 20111 7 1 2 19819 20110
0 20112 5 1 1 20111
0 20113 7 1 2 88983 20112
0 20114 5 1 1 20113
0 20115 7 1 2 87512 95808
0 20116 5 2 1 20115
0 20117 7 1 2 94225 96858
0 20118 5 1 1 20117
0 20119 7 1 2 11770 20118
0 20120 5 1 1 20119
0 20121 7 1 2 92692 20120
0 20122 5 1 1 20121
0 20123 7 1 2 98561 20122
0 20124 5 1 1 20123
0 20125 7 1 2 84669 20124
0 20126 5 1 1 20125
0 20127 7 2 2 69483 92578
0 20128 5 2 1 98563
0 20129 7 1 2 98565 6043
0 20130 5 1 1 20129
0 20131 7 1 2 94807 20130
0 20132 5 1 1 20131
0 20133 7 1 2 20126 20132
0 20134 5 1 1 20133
0 20135 7 1 2 73087 20134
0 20136 5 1 1 20135
0 20137 7 1 2 88571 96859
0 20138 5 1 1 20137
0 20139 7 1 2 95977 20138
0 20140 5 1 1 20139
0 20141 7 1 2 68368 20140
0 20142 5 1 1 20141
0 20143 7 1 2 86367 93854
0 20144 5 1 1 20143
0 20145 7 1 2 20142 20144
0 20146 5 1 1 20145
0 20147 7 1 2 71623 20146
0 20148 5 1 1 20147
0 20149 7 1 2 86939 95971
0 20150 5 1 1 20149
0 20151 7 1 2 20148 20150
0 20152 5 1 1 20151
0 20153 7 1 2 85893 20152
0 20154 5 1 1 20153
0 20155 7 1 2 92908 89311
0 20156 5 1 1 20155
0 20157 7 1 2 20154 20156
0 20158 5 1 1 20157
0 20159 7 1 2 64377 20158
0 20160 5 1 1 20159
0 20161 7 1 2 94808 87326
0 20162 5 1 1 20161
0 20163 7 1 2 20160 20162
0 20164 5 1 1 20163
0 20165 7 1 2 85009 20164
0 20166 5 1 1 20165
0 20167 7 1 2 20136 20166
0 20168 5 1 1 20167
0 20169 7 1 2 65978 20168
0 20170 5 1 1 20169
0 20171 7 1 2 85260 89470
0 20172 5 1 1 20171
0 20173 7 1 2 91824 89656
0 20174 5 1 1 20173
0 20175 7 1 2 20172 20174
0 20176 5 1 1 20175
0 20177 7 1 2 66717 20176
0 20178 5 1 1 20177
0 20179 7 1 2 66523 85894
0 20180 7 1 2 77830 20179
0 20181 7 1 2 90545 20180
0 20182 5 1 1 20181
0 20183 7 1 2 20178 20182
0 20184 5 1 1 20183
0 20185 7 1 2 73447 20184
0 20186 5 1 1 20185
0 20187 7 1 2 20186 98562
0 20188 5 1 1 20187
0 20189 7 1 2 82565 84938
0 20190 7 1 2 20188 20189
0 20191 5 1 1 20190
0 20192 7 1 2 74423 20191
0 20193 7 1 2 20170 20192
0 20194 5 1 1 20193
0 20195 7 1 2 90546 90258
0 20196 5 1 1 20195
0 20197 7 1 2 7001 20196
0 20198 5 1 1 20197
0 20199 7 2 2 75566 97032
0 20200 7 1 2 20198 98567
0 20201 5 1 1 20200
0 20202 7 1 2 95045 88210
0 20203 5 1 1 20202
0 20204 7 1 2 92700 75639
0 20205 5 1 1 20204
0 20206 7 1 2 20203 20205
0 20207 5 1 1 20206
0 20208 7 1 2 97081 20207
0 20209 5 1 1 20208
0 20210 7 2 2 96739 84378
0 20211 7 1 2 92048 98569
0 20212 5 1 1 20211
0 20213 7 1 2 97082 89883
0 20214 5 1 1 20213
0 20215 7 1 2 20212 20214
0 20216 5 1 1 20215
0 20217 7 1 2 78596 20216
0 20218 5 1 1 20217
0 20219 7 1 2 67269 98557
0 20220 7 1 2 90193 20219
0 20221 7 1 2 90963 20220
0 20222 5 1 1 20221
0 20223 7 1 2 20218 20222
0 20224 7 1 2 20209 20223
0 20225 5 1 1 20224
0 20226 7 1 2 66718 20225
0 20227 5 1 1 20226
0 20228 7 1 2 20201 20227
0 20229 5 1 1 20228
0 20230 7 1 2 85895 20229
0 20231 5 1 1 20230
0 20232 7 2 2 79376 97033
0 20233 7 1 2 98571 95735
0 20234 7 1 2 92909 20233
0 20235 5 1 1 20234
0 20236 7 1 2 20231 20235
0 20237 5 1 1 20236
0 20238 7 1 2 69484 20237
0 20239 5 1 1 20238
0 20240 7 1 2 87638 91457
0 20241 5 1 1 20240
0 20242 7 1 2 92251 20241
0 20243 5 1 1 20242
0 20244 7 1 2 65069 20243
0 20245 5 1 1 20244
0 20246 7 1 2 83515 98317
0 20247 5 2 1 20246
0 20248 7 1 2 98573 85010
0 20249 5 1 1 20248
0 20250 7 1 2 20245 20249
0 20251 5 1 1 20250
0 20252 7 1 2 88572 20251
0 20253 5 1 1 20252
0 20254 7 1 2 92636 95972
0 20255 5 1 1 20254
0 20256 7 1 2 20253 20255
0 20257 5 1 1 20256
0 20258 7 1 2 79104 98092
0 20259 7 1 2 20257 20258
0 20260 5 1 1 20259
0 20261 7 1 2 65979 20260
0 20262 7 1 2 20239 20261
0 20263 5 1 1 20262
0 20264 7 8 2 65070 71809
0 20265 5 2 1 98575
0 20266 7 1 2 93979 98583
0 20267 5 2 1 20266
0 20268 7 14 2 64378 67270
0 20269 5 1 1 98587
0 20270 7 1 2 77698 98588
0 20271 5 1 1 20270
0 20272 7 5 2 72340 75567
0 20273 7 1 2 80882 98601
0 20274 5 1 1 20273
0 20275 7 1 2 20271 20274
0 20276 5 1 1 20275
0 20277 7 1 2 98585 20276
0 20278 5 1 1 20277
0 20279 7 16 2 69485 72341
0 20280 7 2 2 77086 75568
0 20281 7 1 2 98606 98622
0 20282 5 1 1 20281
0 20283 7 2 2 86213 98589
0 20284 7 1 2 86809 86949
0 20285 7 1 2 98624 20284
0 20286 5 1 1 20285
0 20287 7 1 2 20282 20286
0 20288 5 1 1 20287
0 20289 7 1 2 65071 20288
0 20290 5 1 1 20289
0 20291 7 1 2 20278 20290
0 20292 5 1 1 20291
0 20293 7 1 2 88573 20292
0 20294 5 1 1 20293
0 20295 7 1 2 97116 88750
0 20296 5 1 1 20295
0 20297 7 1 2 82026 98607
0 20298 7 1 2 95803 20297
0 20299 5 1 1 20298
0 20300 7 1 2 20296 20299
0 20301 5 1 1 20300
0 20302 7 1 2 93855 20301
0 20303 5 1 1 20302
0 20304 7 1 2 20294 20303
0 20305 5 1 1 20304
0 20306 7 1 2 85896 20305
0 20307 5 1 1 20306
0 20308 7 6 2 72150 72342
0 20309 7 1 2 89123 98626
0 20310 7 1 2 97011 20309
0 20311 5 1 1 20310
0 20312 7 1 2 73727 98625
0 20313 7 1 2 89832 20312
0 20314 5 1 1 20313
0 20315 7 1 2 20311 20314
0 20316 5 1 1 20315
0 20317 7 1 2 85261 20316
0 20318 5 1 1 20317
0 20319 7 1 2 20307 20318
0 20320 5 1 1 20319
0 20321 7 1 2 72648 20320
0 20322 5 1 1 20321
0 20323 7 2 2 89381 77728
0 20324 7 1 2 83634 98632
0 20325 5 1 1 20324
0 20326 7 1 2 85262 94701
0 20327 5 1 1 20326
0 20328 7 1 2 20325 20327
0 20329 5 1 1 20328
0 20330 7 1 2 95965 20329
0 20331 5 1 1 20330
0 20332 7 1 2 92910 90490
0 20333 7 1 2 85356 8548
0 20334 5 2 1 20333
0 20335 7 1 2 85357 98318
0 20336 5 1 1 20335
0 20337 7 1 2 98634 20336
0 20338 7 1 2 20332 20337
0 20339 5 1 1 20338
0 20340 7 1 2 20331 20339
0 20341 5 1 1 20340
0 20342 7 1 2 68016 20341
0 20343 5 1 1 20342
0 20344 7 1 2 98332 90000
0 20345 5 1 1 20344
0 20346 7 1 2 81100 96720
0 20347 5 1 1 20346
0 20348 7 1 2 20345 20347
0 20349 5 1 1 20348
0 20350 7 1 2 87011 20349
0 20351 5 1 1 20350
0 20352 7 1 2 20343 20351
0 20353 5 1 1 20352
0 20354 7 1 2 97034 20353
0 20355 5 1 1 20354
0 20356 7 1 2 71052 20355
0 20357 7 1 2 20322 20356
0 20358 5 1 1 20357
0 20359 7 1 2 20263 20358
0 20360 5 1 1 20359
0 20361 7 4 2 64379 75045
0 20362 5 3 1 98636
0 20363 7 1 2 98640 88211
0 20364 5 1 1 20363
0 20365 7 1 2 89135 20364
0 20366 5 1 1 20365
0 20367 7 1 2 73088 20366
0 20368 5 1 1 20367
0 20369 7 1 2 66524 75804
0 20370 7 1 2 91609 20369
0 20371 5 1 1 20370
0 20372 7 1 2 20368 20371
0 20373 5 1 1 20372
0 20374 7 1 2 94036 20373
0 20375 5 1 1 20374
0 20376 7 1 2 92693 98586
0 20377 5 1 1 20376
0 20378 7 1 2 66719 95823
0 20379 5 1 1 20378
0 20380 7 1 2 20377 20379
0 20381 5 1 1 20380
0 20382 7 1 2 66525 81236
0 20383 7 1 2 20381 20382
0 20384 5 1 1 20383
0 20385 7 1 2 81211 88212
0 20386 7 1 2 86963 20385
0 20387 5 1 1 20386
0 20388 7 1 2 20384 20387
0 20389 5 1 1 20388
0 20390 7 1 2 85897 20389
0 20391 5 1 1 20390
0 20392 7 1 2 20375 20391
0 20393 5 1 1 20392
0 20394 7 1 2 98404 20393
0 20395 5 1 1 20394
0 20396 7 1 2 83186 97035
0 20397 7 1 2 94809 20396
0 20398 7 1 2 97789 20397
0 20399 5 1 1 20398
0 20400 7 1 2 74387 20399
0 20401 7 1 2 20395 20400
0 20402 7 1 2 20360 20401
0 20403 5 1 1 20402
0 20404 7 3 2 67271 74424
0 20405 5 1 1 98643
0 20406 7 2 2 82490 20405
0 20407 7 1 2 65390 98646
0 20408 7 1 2 20403 20407
0 20409 7 1 2 20194 20408
0 20410 5 1 1 20409
0 20411 7 5 2 72343 85434
0 20412 5 1 1 98648
0 20413 7 1 2 81396 78724
0 20414 7 1 2 92039 20413
0 20415 5 1 1 20414
0 20416 7 2 2 74780 88213
0 20417 5 1 1 98653
0 20418 7 1 2 17668 20417
0 20419 5 1 1 20418
0 20420 7 1 2 70150 20419
0 20421 5 1 1 20420
0 20422 7 1 2 81373 88214
0 20423 5 1 1 20422
0 20424 7 1 2 20421 20423
0 20425 5 1 1 20424
0 20426 7 6 2 70409 72649
0 20427 5 2 1 98655
0 20428 7 1 2 80345 98656
0 20429 7 1 2 20425 20428
0 20430 5 1 1 20429
0 20431 7 1 2 20415 20430
0 20432 5 1 1 20431
0 20433 7 1 2 65980 20432
0 20434 5 1 1 20433
0 20435 7 2 2 93118 88215
0 20436 7 1 2 92867 87012
0 20437 7 1 2 98663 20436
0 20438 5 1 1 20437
0 20439 7 1 2 20434 20438
0 20440 5 1 1 20439
0 20441 7 1 2 85898 20440
0 20442 5 1 1 20441
0 20443 7 2 2 82047 19793
0 20444 5 1 1 98665
0 20445 7 1 2 83608 20444
0 20446 5 1 1 20445
0 20447 7 1 2 84757 81436
0 20448 5 1 1 20447
0 20449 7 1 2 20446 20448
0 20450 5 1 1 20449
0 20451 7 1 2 88574 20450
0 20452 5 1 1 20451
0 20453 7 1 2 7496 20452
0 20454 5 1 1 20453
0 20455 7 1 2 89428 78365
0 20456 7 1 2 20454 20455
0 20457 5 1 1 20456
0 20458 7 1 2 20442 20457
0 20459 5 1 1 20458
0 20460 7 1 2 64380 20459
0 20461 5 1 1 20460
0 20462 7 3 2 66983 68632
0 20463 7 3 2 63787 98667
0 20464 5 1 1 98670
0 20465 7 1 2 98671 96645
0 20466 5 1 1 20465
0 20467 7 4 2 72047 89925
0 20468 7 1 2 69486 98673
0 20469 5 1 1 20468
0 20470 7 1 2 20466 20469
0 20471 5 1 1 20470
0 20472 7 3 2 67109 94647
0 20473 7 1 2 81105 82244
0 20474 7 1 2 98677 20473
0 20475 7 1 2 20471 20474
0 20476 5 1 1 20475
0 20477 7 1 2 20461 20476
0 20478 5 1 1 20477
0 20479 7 1 2 98649 20478
0 20480 5 1 1 20479
0 20481 7 6 2 63788 75146
0 20482 5 1 1 98680
0 20483 7 1 2 92220 82077
0 20484 5 1 1 20483
0 20485 7 1 2 20482 20484
0 20486 5 1 1 20485
0 20487 7 16 2 72344 72650
0 20488 7 2 2 98686 96102
0 20489 5 1 1 98702
0 20490 7 1 2 69124 20489
0 20491 5 1 1 20490
0 20492 7 12 2 70789 77332
0 20493 7 3 2 98704 98687
0 20494 5 1 1 98716
0 20495 7 1 2 64381 98405
0 20496 5 2 1 20495
0 20497 7 2 2 98608 78456
0 20498 5 1 1 98721
0 20499 7 1 2 98719 20498
0 20500 5 2 1 20499
0 20501 7 1 2 65774 98723
0 20502 5 1 1 20501
0 20503 7 2 2 20494 20502
0 20504 5 1 1 98725
0 20505 7 1 2 64076 98726
0 20506 5 1 1 20505
0 20507 7 2 2 20491 20506
0 20508 7 1 2 88216 98727
0 20509 5 1 1 20508
0 20510 7 1 2 96103 92854
0 20511 7 1 2 97228 20510
0 20512 5 1 1 20511
0 20513 7 1 2 20509 20512
0 20514 5 1 1 20513
0 20515 7 1 2 20486 20514
0 20516 5 1 1 20515
0 20517 7 1 2 83564 98728
0 20518 5 1 1 20517
0 20519 7 6 2 93251 74189
0 20520 5 2 1 98729
0 20521 7 2 2 97866 97997
0 20522 5 1 1 98737
0 20523 7 1 2 98735 20522
0 20524 5 11 1 20523
0 20525 7 1 2 76684 98688
0 20526 7 1 2 98739 20525
0 20527 5 1 1 20526
0 20528 7 1 2 20518 20527
0 20529 5 1 1 20528
0 20530 7 1 2 95680 77748
0 20531 7 1 2 20529 20530
0 20532 5 1 1 20531
0 20533 7 1 2 20516 20532
0 20534 5 1 1 20533
0 20535 7 1 2 81853 20534
0 20536 5 1 1 20535
0 20537 7 1 2 98397 90734
0 20538 5 1 1 20537
0 20539 7 2 2 68843 96740
0 20540 7 1 2 72048 87667
0 20541 7 1 2 98750 20540
0 20542 5 1 1 20541
0 20543 7 1 2 20538 20542
0 20544 5 1 1 20543
0 20545 7 1 2 83681 20544
0 20546 5 1 1 20545
0 20547 7 28 2 67272 67624
0 20548 7 2 2 83216 98752
0 20549 7 1 2 82912 89429
0 20550 7 1 2 98780 20549
0 20551 5 1 1 20550
0 20552 7 1 2 20546 20551
0 20553 5 1 1 20552
0 20554 7 1 2 64382 20553
0 20555 5 1 1 20554
0 20556 7 1 2 95776 98722
0 20557 7 1 2 90735 20556
0 20558 5 1 1 20557
0 20559 7 1 2 20555 20558
0 20560 5 1 1 20559
0 20561 7 1 2 65775 20560
0 20562 5 1 1 20561
0 20563 7 1 2 95777 98717
0 20564 7 1 2 90736 20563
0 20565 5 1 1 20564
0 20566 7 1 2 20562 20565
0 20567 5 1 1 20566
0 20568 7 1 2 88575 20567
0 20569 5 1 1 20568
0 20570 7 1 2 5263 18731
0 20571 5 1 1 20570
0 20572 7 1 2 85899 20571
0 20573 5 1 1 20572
0 20574 7 2 2 98211 97322
0 20575 5 2 1 98782
0 20576 7 1 2 98783 97291
0 20577 5 1 1 20576
0 20578 7 1 2 20573 20577
0 20579 5 1 1 20578
0 20580 7 1 2 65981 20579
0 20581 5 1 1 20580
0 20582 7 1 2 92868 98558
0 20583 7 1 2 92083 20582
0 20584 5 1 1 20583
0 20585 7 1 2 20581 20584
0 20586 5 1 1 20585
0 20587 7 1 2 98484 20586
0 20588 5 1 1 20587
0 20589 7 1 2 77425 92158
0 20590 7 1 2 89246 20589
0 20591 5 1 1 20590
0 20592 7 1 2 92552 92902
0 20593 5 1 1 20592
0 20594 7 1 2 85900 80229
0 20595 7 1 2 20593 20594
0 20596 5 1 1 20595
0 20597 7 1 2 20591 20596
0 20598 5 1 1 20597
0 20599 7 1 2 86671 20598
0 20600 5 1 1 20599
0 20601 7 2 2 85901 92628
0 20602 7 1 2 79924 92366
0 20603 7 1 2 98786 20602
0 20604 5 1 1 20603
0 20605 7 1 2 20600 20604
0 20606 5 1 1 20605
0 20607 7 1 2 97962 20606
0 20608 5 1 1 20607
0 20609 7 1 2 20588 20608
0 20610 5 1 1 20609
0 20611 7 1 2 88217 20610
0 20612 5 1 1 20611
0 20613 7 1 2 73089 20612
0 20614 7 1 2 20569 20613
0 20615 5 1 1 20614
0 20616 7 1 2 80595 89110
0 20617 5 1 1 20616
0 20618 7 1 2 85358 20617
0 20619 5 2 1 20618
0 20620 7 1 2 98788 20504
0 20621 5 1 1 20620
0 20622 7 4 2 83499 82411
0 20623 5 1 1 98790
0 20624 7 4 2 63789 71624
0 20625 7 1 2 97099 98794
0 20626 7 1 2 98791 20625
0 20627 7 1 2 97685 20626
0 20628 5 1 1 20627
0 20629 7 1 2 20621 20628
0 20630 5 1 1 20629
0 20631 7 1 2 68633 20630
0 20632 5 1 1 20631
0 20633 7 1 2 65982 97072
0 20634 5 1 1 20633
0 20635 7 1 2 98720 20634
0 20636 5 1 1 20635
0 20637 7 1 2 82913 82412
0 20638 7 1 2 92221 20637
0 20639 7 1 2 20636 20638
0 20640 5 1 1 20639
0 20641 7 1 2 20632 20640
0 20642 5 1 1 20641
0 20643 7 1 2 88218 20642
0 20644 5 1 1 20643
0 20645 7 1 2 85902 82858
0 20646 5 1 1 20645
0 20647 7 2 2 70410 83421
0 20648 5 4 1 98798
0 20649 7 1 2 87344 98800
0 20650 5 7 1 20649
0 20651 7 1 2 85263 98804
0 20652 5 1 1 20651
0 20653 7 1 2 93797 94054
0 20654 5 1 1 20653
0 20655 7 1 2 20652 20654
0 20656 7 1 2 20646 20655
0 20657 5 1 1 20656
0 20658 7 2 2 65776 78465
0 20659 5 1 1 98811
0 20660 7 1 2 65777 78478
0 20661 5 5 1 20660
0 20662 7 1 2 98813 11152
0 20663 5 6 1 20662
0 20664 7 1 2 64383 98818
0 20665 5 1 1 20664
0 20666 7 1 2 20659 20665
0 20667 5 1 1 20666
0 20668 7 1 2 72345 20667
0 20669 7 1 2 20657 20668
0 20670 5 1 1 20669
0 20671 7 1 2 85264 85625
0 20672 5 2 1 20671
0 20673 7 6 2 68844 70411
0 20674 7 2 2 91820 98826
0 20675 5 1 1 98832
0 20676 7 3 2 73448 97336
0 20677 5 1 1 98834
0 20678 7 1 2 98833 98835
0 20679 5 1 1 20678
0 20680 7 1 2 98824 20679
0 20681 5 1 1 20680
0 20682 7 1 2 97894 94684
0 20683 7 1 2 20681 20682
0 20684 5 1 1 20683
0 20685 7 6 2 65072 65778
0 20686 5 1 1 98837
0 20687 7 1 2 64384 98838
0 20688 7 3 2 68845 68369
0 20689 7 1 2 83726 98093
0 20690 7 1 2 98843 20689
0 20691 7 1 2 20687 20690
0 20692 7 1 2 98805 20691
0 20693 5 1 1 20692
0 20694 7 1 2 20684 20693
0 20695 7 1 2 20670 20694
0 20696 5 1 1 20695
0 20697 7 1 2 88576 20696
0 20698 5 1 1 20697
0 20699 7 1 2 68017 20698
0 20700 7 1 2 20644 20699
0 20701 5 1 1 20700
0 20702 7 1 2 64077 20701
0 20703 7 1 2 20615 20702
0 20704 5 1 1 20703
0 20705 7 1 2 20536 20704
0 20706 7 1 2 20480 20705
0 20707 7 1 2 20410 20706
0 20708 5 1 1 20707
0 20709 7 1 2 88074 20708
0 20710 5 1 1 20709
0 20711 7 2 2 14290 19322
0 20712 5 1 1 98846
0 20713 7 1 2 82557 98847
0 20714 5 1 1 20713
0 20715 7 1 2 81854 20714
0 20716 5 1 1 20715
0 20717 7 1 2 80596 98541
0 20718 5 1 1 20717
0 20719 7 1 2 20716 20718
0 20720 5 1 1 20719
0 20721 7 1 2 75569 20720
0 20722 5 1 1 20721
0 20723 7 1 2 17065 81006
0 20724 5 1 1 20723
0 20725 7 4 2 72651 77209
0 20726 5 2 1 98848
0 20727 7 1 2 86915 98852
0 20728 7 1 2 20724 20727
0 20729 5 1 1 20728
0 20730 7 1 2 20722 20729
0 20731 5 1 1 20730
0 20732 7 1 2 91313 20731
0 20733 5 1 1 20732
0 20734 7 3 2 91318 91392
0 20735 7 5 2 73449 96612
0 20736 5 1 1 98857
0 20737 7 1 2 69487 98858
0 20738 5 1 1 20737
0 20739 7 1 2 5106 20738
0 20740 5 1 1 20739
0 20741 7 1 2 98819 20740
0 20742 5 1 1 20741
0 20743 7 1 2 77987 98859
0 20744 5 1 1 20743
0 20745 7 1 2 69488 95916
0 20746 5 1 1 20745
0 20747 7 1 2 20744 20746
0 20748 5 1 1 20747
0 20749 7 1 2 83747 20748
0 20750 5 1 1 20749
0 20751 7 1 2 20742 20750
0 20752 5 1 1 20751
0 20753 7 1 2 98854 20752
0 20754 5 1 1 20753
0 20755 7 1 2 20733 20754
0 20756 5 1 1 20755
0 20757 7 1 2 64078 20756
0 20758 5 1 1 20757
0 20759 7 1 2 98661 98812
0 20760 5 1 1 20759
0 20761 7 1 2 3015 78495
0 20762 5 1 1 20761
0 20763 7 2 2 70790 83738
0 20764 5 2 1 98862
0 20765 7 1 2 64385 98864
0 20766 7 1 2 20762 20765
0 20767 5 1 1 20766
0 20768 7 1 2 20760 20767
0 20769 5 1 1 20768
0 20770 7 1 2 82914 91314
0 20771 7 1 2 20769 20770
0 20772 5 1 1 20771
0 20773 7 4 2 69125 96698
0 20774 7 1 2 94496 98866
0 20775 7 1 2 93365 20774
0 20776 7 1 2 93528 20775
0 20777 5 1 1 20776
0 20778 7 1 2 20772 20777
0 20779 5 1 1 20778
0 20780 7 1 2 77664 20779
0 20781 5 1 1 20780
0 20782 7 1 2 94206 91284
0 20783 7 1 2 93361 96722
0 20784 7 1 2 98867 20783
0 20785 7 1 2 20782 20784
0 20786 5 1 1 20785
0 20787 7 1 2 20781 20786
0 20788 7 1 2 20758 20787
0 20789 5 1 1 20788
0 20790 7 1 2 85265 20789
0 20791 5 1 1 20790
0 20792 7 1 2 95886 88984
0 20793 5 1 1 20792
0 20794 7 1 2 70723 92493
0 20795 7 1 2 87302 20794
0 20796 7 1 2 88042 20795
0 20797 5 1 1 20796
0 20798 7 1 2 20793 20797
0 20799 5 1 1 20798
0 20800 7 1 2 82547 20799
0 20801 5 1 1 20800
0 20802 7 1 2 96394 97849
0 20803 7 1 2 94338 20802
0 20804 5 1 1 20803
0 20805 7 1 2 20801 20804
0 20806 5 1 1 20805
0 20807 7 1 2 71053 20806
0 20808 5 1 1 20807
0 20809 7 2 2 66720 91937
0 20810 7 3 2 70724 98870
0 20811 7 1 2 77063 98872
0 20812 7 1 2 97452 20811
0 20813 5 1 1 20812
0 20814 7 1 2 20808 20813
0 20815 5 1 1 20814
0 20816 7 1 2 64079 20815
0 20817 5 1 1 20816
0 20818 7 6 2 65779 66721
0 20819 7 3 2 71937 98875
0 20820 7 2 2 94777 94082
0 20821 7 1 2 98881 98884
0 20822 7 1 2 97456 20821
0 20823 5 1 1 20822
0 20824 7 1 2 20817 20823
0 20825 5 1 1 20824
0 20826 7 1 2 73450 20825
0 20827 5 1 1 20826
0 20828 7 1 2 67625 94814
0 20829 7 1 2 84501 20828
0 20830 7 2 2 66865 80597
0 20831 7 1 2 92230 98886
0 20832 7 1 2 20829 20831
0 20833 5 1 1 20832
0 20834 7 1 2 20827 20833
0 20835 5 1 1 20834
0 20836 7 1 2 88219 20835
0 20837 5 1 1 20836
0 20838 7 3 2 90583 92439
0 20839 7 7 2 93648 98888
0 20840 7 2 2 76156 81397
0 20841 7 4 2 71054 66866
0 20842 7 1 2 98900 97015
0 20843 7 1 2 98898 20842
0 20844 7 1 2 98891 20843
0 20845 5 1 1 20844
0 20846 7 1 2 20837 20845
0 20847 5 1 1 20846
0 20848 7 1 2 85903 20847
0 20849 5 1 1 20848
0 20850 7 1 2 20791 20849
0 20851 5 1 1 20850
0 20852 7 1 2 72346 20851
0 20853 5 1 1 20852
0 20854 7 2 2 97951 86214
0 20855 7 1 2 83217 91305
0 20856 7 1 2 94637 20855
0 20857 5 1 1 20856
0 20858 7 1 2 81030 88075
0 20859 7 1 2 95812 20858
0 20860 5 1 1 20859
0 20861 7 1 2 20857 20860
0 20862 5 1 1 20861
0 20863 7 1 2 65780 20862
0 20864 5 1 1 20863
0 20865 7 3 2 66984 90584
0 20866 7 1 2 98906 89353
0 20867 7 2 2 65686 74315
0 20868 7 1 2 92605 98909
0 20869 7 1 2 20866 20868
0 20870 5 1 1 20869
0 20871 7 1 2 20864 20870
0 20872 5 1 1 20871
0 20873 7 1 2 72652 20872
0 20874 5 1 1 20873
0 20875 7 1 2 93252 93551
0 20876 7 1 2 92625 20875
0 20877 7 1 2 92482 20876
0 20878 5 1 1 20877
0 20879 7 1 2 20874 20878
0 20880 5 1 1 20879
0 20881 7 1 2 64080 20880
0 20882 5 1 1 20881
0 20883 7 1 2 65781 81106
0 20884 7 1 2 97261 20883
0 20885 7 1 2 97175 20884
0 20886 5 1 1 20885
0 20887 7 1 2 20882 20886
0 20888 5 1 1 20887
0 20889 7 1 2 98904 20888
0 20890 5 1 1 20889
0 20891 7 1 2 20853 20890
0 20892 5 1 1 20891
0 20893 7 1 2 74649 20892
0 20894 5 1 1 20893
0 20895 7 1 2 92350 87137
0 20896 5 1 1 20895
0 20897 7 15 2 67626 80695
0 20898 7 2 2 73090 98911
0 20899 5 1 1 98926
0 20900 7 1 2 80598 92754
0 20901 5 2 1 20900
0 20902 7 1 2 20899 98928
0 20903 5 2 1 20902
0 20904 7 1 2 77426 98930
0 20905 5 1 1 20904
0 20906 7 1 2 20896 20905
0 20907 5 1 1 20906
0 20908 7 1 2 75381 20907
0 20909 5 1 1 20908
0 20910 7 1 2 71055 97816
0 20911 5 1 1 20910
0 20912 7 1 2 88770 97546
0 20913 5 2 1 20912
0 20914 7 1 2 69489 98932
0 20915 5 1 1 20914
0 20916 7 1 2 20911 20915
0 20917 5 1 1 20916
0 20918 7 1 2 73091 20917
0 20919 5 1 1 20918
0 20920 7 3 2 74650 85611
0 20921 7 9 2 71056 68018
0 20922 7 1 2 98934 98937
0 20923 5 1 1 20922
0 20924 7 1 2 97538 20923
0 20925 7 1 2 20919 20924
0 20926 5 1 1 20925
0 20927 7 1 2 67627 20926
0 20928 5 1 1 20927
0 20929 7 1 2 20909 20928
0 20930 5 1 1 20929
0 20931 7 1 2 72347 20930
0 20932 5 1 1 20931
0 20933 7 2 2 83727 97117
0 20934 7 1 2 88771 96461
0 20935 5 1 1 20934
0 20936 7 1 2 98946 20935
0 20937 5 1 1 20936
0 20938 7 1 2 20932 20937
0 20939 5 1 1 20938
0 20940 7 1 2 88220 20939
0 20941 5 1 1 20940
0 20942 7 1 2 76824 86834
0 20943 5 2 1 20942
0 20944 7 2 2 66722 87795
0 20945 5 1 1 98950
0 20946 7 1 2 86749 98951
0 20947 5 1 1 20946
0 20948 7 1 2 98948 20947
0 20949 5 1 1 20948
0 20950 7 1 2 77427 20949
0 20951 5 1 1 20950
0 20952 7 3 2 67628 74850
0 20953 7 1 2 87138 98952
0 20954 5 1 1 20953
0 20955 7 1 2 20951 20954
0 20956 5 1 1 20955
0 20957 7 1 2 75382 20956
0 20958 5 1 1 20957
0 20959 7 1 2 77428 97509
0 20960 5 1 1 20959
0 20961 7 1 2 98366 20960
0 20962 5 1 1 20961
0 20963 7 1 2 73092 20962
0 20964 5 1 1 20963
0 20965 7 1 2 86266 1820
0 20966 7 1 2 95804 20965
0 20967 5 1 1 20966
0 20968 7 2 2 71810 86267
0 20969 5 1 1 98955
0 20970 7 1 2 98938 20969
0 20971 7 1 2 20967 20970
0 20972 5 1 1 20971
0 20973 7 1 2 20964 20972
0 20974 5 1 1 20973
0 20975 7 1 2 67629 20974
0 20976 5 1 1 20975
0 20977 7 1 2 20958 20976
0 20978 5 1 1 20977
0 20979 7 1 2 72348 20978
0 20980 5 1 1 20979
0 20981 7 1 2 97610 98947
0 20982 5 1 1 20981
0 20983 7 1 2 77429 92262
0 20984 5 1 1 20983
0 20985 7 1 2 67630 87162
0 20986 5 1 1 20985
0 20987 7 1 2 20984 20986
0 20988 5 1 1 20987
0 20989 7 1 2 72349 20988
0 20990 5 1 1 20989
0 20991 7 1 2 77665 97751
0 20992 5 1 1 20991
0 20993 7 1 2 20990 20992
0 20994 5 1 1 20993
0 20995 7 1 2 70151 20994
0 20996 5 1 1 20995
0 20997 7 2 2 73451 80883
0 20998 5 1 1 98957
0 20999 7 1 2 20998 97655
0 21000 5 3 1 20999
0 21001 7 1 2 97036 98959
0 21002 5 1 1 21001
0 21003 7 1 2 79230 96789
0 21004 5 1 1 21003
0 21005 7 1 2 21002 21004
0 21006 5 1 1 21005
0 21007 7 1 2 73093 21006
0 21008 5 1 1 21007
0 21009 7 1 2 20996 21008
0 21010 5 1 1 21009
0 21011 7 1 2 81855 21010
0 21012 5 1 1 21011
0 21013 7 1 2 20982 21012
0 21014 7 1 2 20980 21013
0 21015 5 1 1 21014
0 21016 7 1 2 88577 21015
0 21017 5 1 1 21016
0 21018 7 1 2 20941 21017
0 21019 5 1 1 21018
0 21020 7 1 2 74388 21019
0 21021 5 1 1 21020
0 21022 7 1 2 83438 90404
0 21023 5 1 1 21022
0 21024 7 1 2 89848 21023
0 21025 5 1 1 21024
0 21026 7 1 2 68634 21025
0 21027 5 1 1 21026
0 21028 7 1 2 88435 90405
0 21029 5 1 1 21028
0 21030 7 1 2 94446 20091
0 21031 5 1 1 21030
0 21032 7 1 2 75383 21031
0 21033 5 1 1 21032
0 21034 7 1 2 21029 21033
0 21035 7 1 2 21027 21034
0 21036 5 1 1 21035
0 21037 7 1 2 65983 21036
0 21038 5 1 1 21037
0 21039 7 1 2 86135 82789
0 21040 7 1 2 89684 21039
0 21041 5 1 1 21040
0 21042 7 1 2 21038 21041
0 21043 5 1 1 21042
0 21044 7 6 2 73094 98689
0 21045 7 1 2 74425 98962
0 21046 7 1 2 21043 21045
0 21047 5 1 1 21046
0 21048 7 1 2 21021 21047
0 21049 5 1 1 21048
0 21050 7 1 2 82491 91001
0 21051 7 1 2 21049 21050
0 21052 5 1 1 21051
0 21053 7 2 2 73095 88687
0 21054 5 3 1 98968
0 21055 7 8 2 86789 98970
0 21056 7 1 2 67631 92539
0 21057 7 1 2 98973 21056
0 21058 5 1 1 21057
0 21059 7 3 2 71811 72653
0 21060 7 3 2 70412 98981
0 21061 7 1 2 79728 77064
0 21062 7 1 2 98984 21061
0 21063 5 1 1 21062
0 21064 7 1 2 21058 21063
0 21065 5 1 1 21064
0 21066 7 1 2 83543 21065
0 21067 5 1 1 21066
0 21068 7 1 2 76157 74168
0 21069 7 1 2 96525 21068
0 21070 7 1 2 94204 21069
0 21071 5 1 1 21070
0 21072 7 1 2 21067 21071
0 21073 5 1 1 21072
0 21074 7 1 2 66526 21073
0 21075 5 1 1 21074
0 21076 7 1 2 77430 88660
0 21077 5 1 1 21076
0 21078 7 1 2 87165 90989
0 21079 5 1 1 21078
0 21080 7 1 2 21077 21079
0 21081 5 1 1 21080
0 21082 7 1 2 80092 92420
0 21083 7 1 2 21081 21082
0 21084 5 1 1 21083
0 21085 7 1 2 21075 21084
0 21086 5 1 1 21085
0 21087 7 1 2 88221 21086
0 21088 5 1 1 21087
0 21089 7 1 2 16101 88658
0 21090 5 1 1 21089
0 21091 7 1 2 88222 21090
0 21092 5 1 1 21091
0 21093 7 1 2 88578 97973
0 21094 5 1 1 21093
0 21095 7 1 2 21092 21094
0 21096 5 2 1 21095
0 21097 7 1 2 97872 98987
0 21098 5 1 1 21097
0 21099 7 1 2 21088 21098
0 21100 5 1 1 21099
0 21101 7 1 2 72350 21100
0 21102 5 1 1 21101
0 21103 7 4 2 67273 93253
0 21104 7 1 2 87069 86806
0 21105 5 2 1 21104
0 21106 7 1 2 88358 98993
0 21107 5 1 1 21106
0 21108 7 1 2 88223 21107
0 21109 5 1 1 21108
0 21110 7 1 2 80523 90491
0 21111 5 1 1 21110
0 21112 7 1 2 21109 21111
0 21113 5 1 1 21112
0 21114 7 1 2 68019 21113
0 21115 5 1 1 21114
0 21116 7 2 2 84129 84112
0 21117 5 2 1 98995
0 21118 7 1 2 96553 76685
0 21119 5 2 1 21118
0 21120 7 1 2 98997 98999
0 21121 5 3 1 21120
0 21122 7 1 2 99001 91401
0 21123 5 1 1 21122
0 21124 7 1 2 21115 21123
0 21125 5 1 1 21124
0 21126 7 1 2 72654 21125
0 21127 5 1 1 21126
0 21128 7 1 2 86431 95967
0 21129 5 1 1 21128
0 21130 7 1 2 21127 21129
0 21131 5 1 1 21130
0 21132 7 1 2 98989 21131
0 21133 5 1 1 21132
0 21134 7 1 2 21102 21133
0 21135 5 1 1 21134
0 21136 7 1 2 64081 21135
0 21137 5 1 1 21136
0 21138 7 1 2 72351 97839
0 21139 5 1 1 21138
0 21140 7 1 2 74531 83056
0 21141 5 2 1 21140
0 21142 7 1 2 97852 99004
0 21143 5 1 1 21142
0 21144 7 1 2 21139 21143
0 21145 5 1 1 21144
0 21146 7 1 2 88579 21145
0 21147 5 1 1 21146
0 21148 7 1 2 19225 9565
0 21149 5 1 1 21148
0 21150 7 2 2 21149 98647
0 21151 7 1 2 99006 97843
0 21152 5 1 1 21151
0 21153 7 1 2 97462 84427
0 21154 5 1 1 21153
0 21155 7 1 2 21152 21154
0 21156 5 1 1 21155
0 21157 7 1 2 88224 21156
0 21158 5 1 1 21157
0 21159 7 1 2 21147 21158
0 21160 5 1 1 21159
0 21161 7 1 2 81031 21160
0 21162 5 1 1 21161
0 21163 7 1 2 64386 98988
0 21164 5 1 1 21163
0 21165 7 3 2 75570 87279
0 21166 5 2 1 99008
0 21167 7 1 2 73728 99009
0 21168 5 1 1 21167
0 21169 7 1 2 96646 97314
0 21170 5 1 1 21169
0 21171 7 1 2 21168 21170
0 21172 5 1 1 21171
0 21173 7 1 2 21172 98664
0 21174 5 1 1 21173
0 21175 7 1 2 21164 21174
0 21176 5 1 1 21175
0 21177 7 1 2 98468 21176
0 21178 5 1 1 21177
0 21179 7 1 2 21162 21178
0 21180 7 1 2 21137 21179
0 21181 5 1 1 21180
0 21182 7 1 2 85137 21181
0 21183 5 1 1 21182
0 21184 7 2 2 87742 75750
0 21185 7 1 2 77333 77749
0 21186 7 1 2 99013 21185
0 21187 5 1 1 21186
0 21188 7 1 2 97627 89808
0 21189 7 1 2 89775 21188
0 21190 5 1 1 21189
0 21191 7 1 2 21187 21190
0 21192 5 1 1 21191
0 21193 7 1 2 85489 21192
0 21194 5 1 1 21193
0 21195 7 2 2 66985 77750
0 21196 7 1 2 89083 77793
0 21197 7 1 2 82782 21196
0 21198 7 1 2 99015 21197
0 21199 5 1 1 21198
0 21200 7 1 2 21194 21199
0 21201 5 1 1 21200
0 21202 7 1 2 72655 21201
0 21203 5 1 1 21202
0 21204 7 1 2 81222 97763
0 21205 5 1 1 21204
0 21206 7 1 2 71057 21205
0 21207 5 1 1 21206
0 21208 7 1 2 7754 21207
0 21209 5 1 1 21208
0 21210 7 1 2 96116 82783
0 21211 7 1 2 21209 21210
0 21212 5 1 1 21211
0 21213 7 1 2 21203 21212
0 21214 5 1 1 21213
0 21215 7 1 2 72352 21214
0 21216 5 1 1 21215
0 21217 7 1 2 88293 6373
0 21218 5 1 1 21217
0 21219 7 6 2 67274 85011
0 21220 5 1 1 99017
0 21221 7 1 2 66986 93041
0 21222 7 1 2 99018 21221
0 21223 7 1 2 96118 21222
0 21224 7 1 2 21218 21223
0 21225 5 1 1 21224
0 21226 7 1 2 21216 21225
0 21227 5 1 1 21226
0 21228 7 1 2 82974 21227
0 21229 5 1 1 21228
0 21230 7 1 2 21183 21229
0 21231 7 1 2 21052 21230
0 21232 5 1 1 21231
0 21233 7 1 2 89577 21232
0 21234 5 1 1 21233
0 21235 7 1 2 20894 21234
0 21236 7 1 2 20710 21235
0 21237 7 1 2 20114 21236
0 21238 7 1 2 19714 21237
0 21239 7 1 2 19361 21238
0 21240 5 1 1 21239
0 21241 7 1 2 97374 21240
0 21242 5 1 1 21241
0 21243 7 3 2 95374 98753
0 21244 7 1 2 74947 85138
0 21245 5 1 1 21244
0 21246 7 1 2 72049 93644
0 21247 7 1 2 94627 21246
0 21248 5 1 1 21247
0 21249 7 1 2 21245 21248
0 21250 5 1 1 21249
0 21251 7 1 2 75881 21250
0 21252 5 1 1 21251
0 21253 7 1 2 89382 77751
0 21254 7 1 2 91975 21253
0 21255 5 1 1 21254
0 21256 7 1 2 21252 21255
0 21257 5 1 1 21256
0 21258 7 1 2 69788 21257
0 21259 5 1 1 21258
0 21260 7 1 2 72151 94563
0 21261 7 1 2 84645 21260
0 21262 7 1 2 76429 21261
0 21263 5 1 1 21262
0 21264 7 1 2 21259 21263
0 21265 5 1 1 21264
0 21266 7 1 2 99023 21265
0 21267 5 1 1 21266
0 21268 7 10 2 66723 72353
0 21269 7 3 2 72656 99026
0 21270 7 1 2 84152 96203
0 21271 5 1 1 21270
0 21272 7 1 2 7793 21271
0 21273 5 1 1 21272
0 21274 7 1 2 66241 21273
0 21275 5 1 1 21274
0 21276 7 3 2 83244 87972
0 21277 7 1 2 94982 99039
0 21278 5 1 1 21277
0 21279 7 1 2 21275 21278
0 21280 5 1 1 21279
0 21281 7 2 2 99036 21280
0 21282 7 1 2 93254 99042
0 21283 5 1 1 21282
0 21284 7 1 2 21267 21283
0 21285 5 1 1 21284
0 21286 7 1 2 89578 21285
0 21287 5 1 1 21286
0 21288 7 2 2 87271 84646
0 21289 5 1 1 99044
0 21290 7 1 2 95683 21289
0 21291 5 2 1 21290
0 21292 7 1 2 94631 99046
0 21293 5 1 1 21292
0 21294 7 4 2 68020 92124
0 21295 7 1 2 71812 91934
0 21296 7 1 2 99048 21295
0 21297 7 1 2 95727 21296
0 21298 5 1 1 21297
0 21299 7 1 2 21293 21298
0 21300 5 1 1 21299
0 21301 7 1 2 72050 21300
0 21302 5 1 1 21301
0 21303 7 1 2 74948 89899
0 21304 7 1 2 90304 21303
0 21305 5 1 1 21304
0 21306 7 1 2 21302 21305
0 21307 5 1 1 21306
0 21308 7 1 2 69789 21307
0 21309 5 1 1 21308
0 21310 7 1 2 95747 99047
0 21311 5 1 1 21310
0 21312 7 1 2 21309 21311
0 21313 5 1 1 21312
0 21314 7 1 2 21313 99024
0 21315 5 1 1 21314
0 21316 7 2 2 68021 91414
0 21317 5 1 1 99052
0 21318 7 1 2 89312 99053
0 21319 5 1 1 21318
0 21320 7 1 2 91227 21319
0 21321 5 1 1 21320
0 21322 7 1 2 66242 21321
0 21323 5 1 1 21322
0 21324 7 1 2 79377 96510
0 21325 7 1 2 91694 21324
0 21326 7 1 2 99040 21325
0 21327 5 1 1 21326
0 21328 7 1 2 21323 21327
0 21329 5 2 1 21328
0 21330 7 1 2 93255 99037
0 21331 7 1 2 99054 21330
0 21332 5 1 1 21331
0 21333 7 1 2 21315 21332
0 21334 7 1 2 21287 21333
0 21335 5 1 1 21334
0 21336 7 1 2 71625 21335
0 21337 5 1 1 21336
0 21338 7 1 2 90039 95672
0 21339 5 1 1 21338
0 21340 7 2 2 68846 77752
0 21341 7 1 2 95666 99056
0 21342 5 1 1 21341
0 21343 7 1 2 21339 21342
0 21344 5 1 1 21343
0 21345 7 3 2 65687 70791
0 21346 5 2 1 99058
0 21347 7 2 2 63977 99059
0 21348 7 5 2 71058 98754
0 21349 7 1 2 99065 91425
0 21350 7 2 2 99063 21349
0 21351 7 1 2 66987 99070
0 21352 7 1 2 21344 21351
0 21353 5 1 1 21352
0 21354 7 2 2 77147 74089
0 21355 7 2 2 94572 99072
0 21356 7 6 2 67275 68022
0 21357 7 3 2 99076 93174
0 21358 7 1 2 95275 99082
0 21359 7 1 2 99074 21358
0 21360 7 1 2 89579 21359
0 21361 5 1 1 21360
0 21362 7 1 2 21353 21361
0 21363 7 1 2 21337 21362
0 21364 5 1 1 21363
0 21365 7 1 2 70152 21364
0 21366 5 1 1 21365
0 21367 7 1 2 72051 84148
0 21368 5 1 1 21367
0 21369 7 1 2 13336 21368
0 21370 5 1 1 21369
0 21371 7 1 2 63790 21370
0 21372 5 1 1 21371
0 21373 7 1 2 95738 99045
0 21374 5 1 1 21373
0 21375 7 1 2 21372 21374
0 21376 5 1 1 21375
0 21377 7 1 2 66867 21376
0 21378 5 1 1 21377
0 21379 7 1 2 92984 84149
0 21380 5 1 1 21379
0 21381 7 1 2 21378 21380
0 21382 5 1 1 21381
0 21383 7 1 2 71340 21382
0 21384 5 1 1 21383
0 21385 7 1 2 91829 75882
0 21386 7 1 2 98681 21385
0 21387 5 1 1 21386
0 21388 7 1 2 21384 21387
0 21389 5 1 1 21388
0 21390 7 1 2 69790 21389
0 21391 5 1 1 21390
0 21392 7 1 2 94564 91851
0 21393 7 1 2 94850 21392
0 21394 5 1 1 21393
0 21395 7 1 2 21391 21394
0 21396 5 1 1 21395
0 21397 7 1 2 99071 21396
0 21398 5 1 1 21397
0 21399 7 1 2 75833 84647
0 21400 5 1 1 21399
0 21401 7 1 2 517 21400
0 21402 5 1 1 21401
0 21403 7 5 2 68023 98755
0 21404 7 5 2 95504 80829
0 21405 7 1 2 90892 99090
0 21406 7 1 2 99085 21405
0 21407 7 1 2 89580 21406
0 21408 7 1 2 21402 21407
0 21409 5 1 1 21408
0 21410 7 1 2 69126 21409
0 21411 7 1 2 21398 21410
0 21412 7 1 2 21366 21411
0 21413 5 1 1 21412
0 21414 7 1 2 99055 98820
0 21415 5 1 1 21414
0 21416 7 2 2 88891 95562
0 21417 7 3 2 88919 99095
0 21418 7 2 2 89189 99097
0 21419 7 3 2 65984 90035
0 21420 5 2 1 99102
0 21421 7 1 2 72657 99105
0 21422 5 1 1 21421
0 21423 7 1 2 90768 21422
0 21424 5 1 1 21423
0 21425 7 1 2 99100 21424
0 21426 5 1 1 21425
0 21427 7 2 2 68024 91220
0 21428 5 1 1 99107
0 21429 7 1 2 91067 97588
0 21430 7 1 2 91342 21429
0 21431 7 1 2 94102 21430
0 21432 5 1 1 21431
0 21433 7 1 2 21428 21432
0 21434 5 2 1 21433
0 21435 7 1 2 76308 99109
0 21436 5 1 1 21435
0 21437 7 3 2 69490 95728
0 21438 7 1 2 70725 87924
0 21439 7 1 2 95736 21438
0 21440 7 1 2 99111 21439
0 21441 5 1 1 21440
0 21442 7 1 2 87743 79352
0 21443 7 1 2 95685 21442
0 21444 5 1 1 21443
0 21445 7 1 2 21441 21444
0 21446 7 1 2 21436 21445
0 21447 5 1 1 21446
0 21448 7 1 2 83748 21447
0 21449 5 1 1 21448
0 21450 7 1 2 21426 21449
0 21451 5 1 1 21450
0 21452 7 1 2 65782 21451
0 21453 5 1 1 21452
0 21454 7 1 2 21415 21453
0 21455 5 1 1 21454
0 21456 7 1 2 66724 21455
0 21457 5 1 1 21456
0 21458 7 1 2 93529 89313
0 21459 5 1 1 21458
0 21460 7 1 2 87604 79105
0 21461 7 1 2 91241 84648
0 21462 7 1 2 21460 21461
0 21463 5 1 1 21462
0 21464 7 1 2 21459 21463
0 21465 5 1 1 21464
0 21466 7 1 2 92500 91669
0 21467 7 1 2 93362 21466
0 21468 7 1 2 21465 21467
0 21469 5 1 1 21468
0 21470 7 1 2 21457 21469
0 21471 5 1 1 21470
0 21472 7 1 2 70153 21471
0 21473 5 1 1 21472
0 21474 7 1 2 77535 93530
0 21475 5 1 1 21474
0 21476 7 1 2 9614 21475
0 21477 5 1 1 21476
0 21478 7 2 2 75772 90305
0 21479 7 1 2 80197 99114
0 21480 7 1 2 21477 21479
0 21481 5 1 1 21480
0 21482 7 1 2 21473 21481
0 21483 5 1 1 21482
0 21484 7 1 2 71626 21483
0 21485 5 1 1 21484
0 21486 7 2 2 84670 91230
0 21487 7 1 2 73096 87973
0 21488 7 1 2 99116 21487
0 21489 5 1 1 21488
0 21490 7 1 2 76387 96048
0 21491 7 1 2 91210 21490
0 21492 5 1 1 21491
0 21493 7 1 2 21489 21492
0 21494 5 1 1 21493
0 21495 7 1 2 71341 21494
0 21496 5 1 1 21495
0 21497 7 3 2 72658 76388
0 21498 7 1 2 69491 99118
0 21499 7 2 2 88225 93999
0 21500 7 1 2 92231 99121
0 21501 7 1 2 21498 21500
0 21502 5 1 1 21501
0 21503 7 1 2 21496 21502
0 21504 5 1 1 21503
0 21505 7 1 2 69791 21504
0 21506 5 1 1 21505
0 21507 7 1 2 89439 99101
0 21508 5 1 1 21507
0 21509 7 1 2 21506 21508
0 21510 5 1 1 21509
0 21511 7 1 2 66725 21510
0 21512 5 1 1 21511
0 21513 7 1 2 87581 89878
0 21514 7 2 2 72659 91170
0 21515 7 2 2 90648 90372
0 21516 7 1 2 99123 99125
0 21517 7 1 2 21513 21516
0 21518 7 1 2 83259 21517
0 21519 5 1 1 21518
0 21520 7 1 2 21512 21519
0 21521 5 1 1 21520
0 21522 7 1 2 71059 21521
0 21523 5 1 1 21522
0 21524 7 2 2 90810 77753
0 21525 7 1 2 89159 99098
0 21526 7 1 2 99127 21525
0 21527 5 1 1 21526
0 21528 7 1 2 21523 21527
0 21529 5 1 1 21528
0 21530 7 1 2 65783 21529
0 21531 5 1 1 21530
0 21532 7 1 2 21485 21531
0 21533 5 1 1 21532
0 21534 7 1 2 72354 21533
0 21535 5 1 1 21534
0 21536 7 7 2 70154 70792
0 21537 7 3 2 99129 82383
0 21538 7 1 2 99043 99136
0 21539 5 1 1 21538
0 21540 7 1 2 74532 90778
0 21541 5 1 1 21540
0 21542 7 1 2 91328 21541
0 21543 5 1 1 21542
0 21544 7 1 2 77431 21543
0 21545 5 1 1 21544
0 21546 7 5 2 69492 78406
0 21547 5 3 1 99139
0 21548 7 1 2 82216 81148
0 21549 5 1 1 21548
0 21550 7 1 2 99144 21549
0 21551 5 1 1 21550
0 21552 7 1 2 75969 21551
0 21553 5 1 1 21552
0 21554 7 1 2 99145 85067
0 21555 5 1 1 21554
0 21556 7 1 2 74533 21555
0 21557 5 1 1 21556
0 21558 7 3 2 69792 78407
0 21559 5 1 1 99147
0 21560 7 1 2 82153 21559
0 21561 5 1 1 21560
0 21562 7 1 2 69493 21561
0 21563 5 1 1 21562
0 21564 7 1 2 21557 21563
0 21565 7 1 2 21553 21564
0 21566 7 1 2 21545 21565
0 21567 5 1 1 21566
0 21568 7 1 2 72355 21567
0 21569 5 1 1 21568
0 21570 7 10 2 66243 67276
0 21571 7 3 2 72660 99150
0 21572 7 2 2 99160 82078
0 21573 5 1 1 99163
0 21574 7 1 2 65985 99164
0 21575 5 1 1 21574
0 21576 7 1 2 21569 21575
0 21577 5 1 1 21576
0 21578 7 2 2 66726 21577
0 21579 7 1 2 91041 99165
0 21580 5 1 1 21579
0 21581 7 4 2 76212 97118
0 21582 5 1 1 99167
0 21583 7 8 2 71342 98019
0 21584 7 1 2 99171 86841
0 21585 5 1 1 21584
0 21586 7 1 2 21582 21585
0 21587 5 1 1 21586
0 21588 7 1 2 65986 21587
0 21589 5 1 1 21588
0 21590 7 1 2 72356 94469
0 21591 7 1 2 92094 21590
0 21592 5 1 1 21591
0 21593 7 1 2 21589 21592
0 21594 5 1 1 21593
0 21595 7 1 2 88580 21594
0 21596 5 1 1 21595
0 21597 7 1 2 71060 83260
0 21598 5 1 1 21597
0 21599 7 1 2 90359 21598
0 21600 5 2 1 21599
0 21601 7 10 2 71813 72357
0 21602 7 1 2 99181 90640
0 21603 7 1 2 99179 21602
0 21604 5 1 1 21603
0 21605 7 1 2 21596 21604
0 21606 5 1 1 21605
0 21607 7 1 2 84671 21606
0 21608 5 1 1 21607
0 21609 7 3 2 69494 97554
0 21610 7 3 2 72661 97472
0 21611 7 2 2 99191 99194
0 21612 7 2 2 75805 99197
0 21613 5 1 1 99199
0 21614 7 1 2 97037 88878
0 21615 5 1 1 21614
0 21616 7 1 2 96792 21615
0 21617 5 2 1 21616
0 21618 7 1 2 90406 99201
0 21619 5 2 1 21618
0 21620 7 1 2 97078 96793
0 21621 5 9 1 21620
0 21622 7 1 2 90539 99205
0 21623 5 1 1 21622
0 21624 7 1 2 99203 21623
0 21625 5 1 1 21624
0 21626 7 1 2 82384 21625
0 21627 5 1 1 21626
0 21628 7 1 2 21613 21627
0 21629 5 1 1 21628
0 21630 7 1 2 83245 21629
0 21631 5 1 1 21630
0 21632 7 2 2 71814 97073
0 21633 5 1 1 99214
0 21634 7 1 2 96794 21633
0 21635 5 1 1 21634
0 21636 7 1 2 88226 21635
0 21637 5 1 1 21636
0 21638 7 1 2 99204 21637
0 21639 5 1 1 21638
0 21640 7 1 2 74148 21639
0 21641 5 1 1 21640
0 21642 7 1 2 98690 84726
0 21643 7 1 2 90413 21642
0 21644 5 1 1 21643
0 21645 7 1 2 21641 21644
0 21646 5 1 1 21645
0 21647 7 1 2 71627 21646
0 21648 5 1 1 21647
0 21649 7 1 2 66244 99200
0 21650 5 1 1 21649
0 21651 7 1 2 21648 21650
0 21652 5 1 1 21651
0 21653 7 1 2 68025 21652
0 21654 5 1 1 21653
0 21655 7 1 2 21631 21654
0 21656 7 1 2 21608 21655
0 21657 5 1 1 21656
0 21658 7 1 2 85139 21657
0 21659 5 1 1 21658
0 21660 7 1 2 21580 21659
0 21661 5 1 1 21660
0 21662 7 1 2 65784 21661
0 21663 5 1 1 21662
0 21664 7 1 2 21539 21663
0 21665 5 1 1 21664
0 21666 7 1 2 89581 21665
0 21667 5 1 1 21666
0 21668 7 5 2 64387 85266
0 21669 5 1 1 99216
0 21670 7 1 2 99217 92654
0 21671 5 1 1 21670
0 21672 7 1 2 68847 96796
0 21673 5 1 1 21672
0 21674 7 1 2 81261 90708
0 21675 7 1 2 21673 21674
0 21676 5 1 1 21675
0 21677 7 1 2 21671 21676
0 21678 5 1 1 21677
0 21679 7 1 2 88581 21678
0 21680 5 1 1 21679
0 21681 7 1 2 97323 96056
0 21682 7 1 2 90947 21681
0 21683 5 1 1 21682
0 21684 7 1 2 21680 21683
0 21685 5 1 1 21684
0 21686 7 1 2 73097 21685
0 21687 5 1 1 21686
0 21688 7 3 2 66245 75848
0 21689 5 1 1 99221
0 21690 7 1 2 99218 99222
0 21691 7 1 2 95260 21690
0 21692 5 1 1 21691
0 21693 7 1 2 21687 21692
0 21694 5 1 1 21693
0 21695 7 1 2 72662 21694
0 21696 5 1 1 21695
0 21697 7 3 2 73098 84618
0 21698 7 1 2 93893 88886
0 21699 7 1 2 99224 21698
0 21700 5 1 1 21699
0 21701 7 1 2 21696 21700
0 21702 5 1 1 21701
0 21703 7 1 2 88076 21702
0 21704 5 1 1 21703
0 21705 7 1 2 79556 87333
0 21706 7 1 2 91205 21705
0 21707 7 1 2 91261 95595
0 21708 7 1 2 21706 21707
0 21709 5 1 1 21708
0 21710 7 1 2 21704 21709
0 21711 5 1 1 21710
0 21712 7 1 2 98990 21711
0 21713 5 1 1 21712
0 21714 7 1 2 64082 21713
0 21715 7 1 2 21667 21714
0 21716 7 1 2 21535 21715
0 21717 5 1 1 21716
0 21718 7 1 2 21413 21717
0 21719 5 1 1 21718
0 21720 7 3 2 86088 87763
0 21721 7 5 2 68026 79467
0 21722 5 1 1 99230
0 21723 7 1 2 21722 86235
0 21724 5 1 1 21723
0 21725 7 1 2 69793 21724
0 21726 5 1 1 21725
0 21727 7 1 2 76071 94470
0 21728 5 1 1 21727
0 21729 7 1 2 21726 21728
0 21730 5 1 1 21729
0 21731 7 1 2 99227 21730
0 21732 5 1 1 21731
0 21733 7 2 2 84563 89694
0 21734 7 1 2 99180 99235
0 21735 5 1 1 21734
0 21736 7 1 2 21732 21735
0 21737 5 1 1 21736
0 21738 7 1 2 71628 21737
0 21739 5 1 1 21738
0 21740 7 2 2 66727 84379
0 21741 7 1 2 76934 83716
0 21742 7 1 2 99237 21741
0 21743 5 1 1 21742
0 21744 7 1 2 21739 21743
0 21745 5 1 1 21744
0 21746 7 1 2 72358 21745
0 21747 5 1 1 21746
0 21748 7 4 2 72152 97119
0 21749 7 3 2 66246 94136
0 21750 7 1 2 65987 87744
0 21751 7 1 2 99243 21750
0 21752 7 1 2 99239 21751
0 21753 5 1 1 21752
0 21754 7 1 2 21747 21753
0 21755 5 1 1 21754
0 21756 7 1 2 84672 21755
0 21757 5 1 1 21756
0 21758 7 1 2 99202 99228
0 21759 5 1 1 21758
0 21760 7 1 2 99206 99236
0 21761 5 1 1 21760
0 21762 7 1 2 21759 21761
0 21763 5 1 1 21762
0 21764 7 1 2 82385 21763
0 21765 5 1 1 21764
0 21766 7 1 2 74030 87598
0 21767 7 2 2 99198 21766
0 21768 5 1 1 99246
0 21769 7 1 2 21765 21768
0 21770 5 1 1 21769
0 21771 7 1 2 83246 21770
0 21772 5 1 1 21771
0 21773 7 3 2 65988 99151
0 21774 5 2 1 99248
0 21775 7 4 2 71343 80830
0 21776 7 1 2 99182 99253
0 21777 5 1 1 21776
0 21778 7 1 2 99251 21777
0 21779 5 1 1 21778
0 21780 7 1 2 84939 21779
0 21781 5 1 1 21780
0 21782 7 1 2 74149 99215
0 21783 5 1 1 21782
0 21784 7 1 2 21781 21783
0 21785 5 1 1 21784
0 21786 7 1 2 87268 21785
0 21787 5 1 1 21786
0 21788 7 3 2 76465 98233
0 21789 5 1 1 99257
0 21790 7 1 2 21789 99252
0 21791 5 1 1 21790
0 21792 7 1 2 84940 21791
0 21793 5 1 1 21792
0 21794 7 11 2 66247 72359
0 21795 5 1 1 99260
0 21796 7 1 2 69495 99261
0 21797 7 1 2 96074 21796
0 21798 5 1 1 21797
0 21799 7 1 2 21793 21798
0 21800 5 1 1 21799
0 21801 7 1 2 99229 21800
0 21802 5 1 1 21801
0 21803 7 1 2 21787 21802
0 21804 5 1 1 21803
0 21805 7 1 2 71629 21804
0 21806 5 1 1 21805
0 21807 7 1 2 66248 99247
0 21808 5 1 1 21807
0 21809 7 1 2 21806 21808
0 21810 5 1 1 21809
0 21811 7 1 2 68027 21810
0 21812 5 1 1 21811
0 21813 7 1 2 21772 21812
0 21814 7 1 2 21757 21813
0 21815 5 1 1 21814
0 21816 7 1 2 66988 21815
0 21817 5 1 1 21816
0 21818 7 7 2 69794 72360
0 21819 7 2 2 78408 99271
0 21820 7 1 2 86089 77754
0 21821 7 1 2 99278 21820
0 21822 7 1 2 84170 21821
0 21823 5 1 1 21822
0 21824 7 1 2 21817 21823
0 21825 5 1 1 21824
0 21826 7 1 2 71938 21825
0 21827 5 1 1 21826
0 21828 7 1 2 79401 99166
0 21829 5 1 1 21828
0 21830 7 1 2 21827 21829
0 21831 5 1 1 21830
0 21832 7 1 2 65785 21831
0 21833 5 1 1 21832
0 21834 7 1 2 94992 96204
0 21835 5 1 1 21834
0 21836 7 1 2 95448 21835
0 21837 5 1 1 21836
0 21838 7 1 2 66249 21837
0 21839 5 1 1 21838
0 21840 7 1 2 94993 99041
0 21841 5 1 1 21840
0 21842 7 1 2 21839 21841
0 21843 5 1 1 21842
0 21844 7 2 2 99038 21843
0 21845 7 1 2 99137 99280
0 21846 5 1 1 21845
0 21847 7 1 2 64083 21846
0 21848 7 1 2 21833 21847
0 21849 5 1 1 21848
0 21850 7 1 2 93256 99281
0 21851 5 1 1 21850
0 21852 7 3 2 76389 79635
0 21853 7 1 2 78825 99282
0 21854 7 1 2 91813 21853
0 21855 5 1 1 21854
0 21856 7 1 2 74244 78074
0 21857 5 1 1 21856
0 21858 7 1 2 74471 89762
0 21859 5 1 1 21858
0 21860 7 1 2 21857 21859
0 21861 5 1 1 21860
0 21862 7 1 2 68848 21861
0 21863 5 1 1 21862
0 21864 7 1 2 93894 97589
0 21865 5 1 1 21864
0 21866 7 1 2 21863 21865
0 21867 5 1 1 21866
0 21868 7 1 2 82724 84486
0 21869 7 1 2 21867 21868
0 21870 5 1 1 21869
0 21871 7 1 2 21855 21870
0 21872 5 1 1 21871
0 21873 7 1 2 76309 99025
0 21874 7 1 2 21872 21873
0 21875 5 1 1 21874
0 21876 7 1 2 21851 21875
0 21877 5 1 1 21876
0 21878 7 1 2 71630 21877
0 21879 5 1 1 21878
0 21880 7 1 2 74031 99083
0 21881 7 2 2 76935 75751
0 21882 7 1 2 99285 95554
0 21883 7 1 2 21880 21882
0 21884 5 1 1 21883
0 21885 7 1 2 21879 21884
0 21886 5 1 1 21885
0 21887 7 1 2 70155 21886
0 21888 5 1 1 21887
0 21889 7 1 2 71631 85574
0 21890 5 1 1 21889
0 21891 7 1 2 85793 21890
0 21892 5 1 1 21891
0 21893 7 1 2 63791 21892
0 21894 5 1 1 21893
0 21895 7 1 2 85140 76977
0 21896 5 1 1 21895
0 21897 7 1 2 21894 21896
0 21898 5 1 1 21897
0 21899 7 1 2 88227 21898
0 21900 5 1 1 21899
0 21901 7 3 2 63792 78075
0 21902 7 2 2 76390 89725
0 21903 7 1 2 99287 99290
0 21904 5 1 1 21903
0 21905 7 1 2 21900 21904
0 21906 5 1 1 21905
0 21907 7 10 2 71344 67277
0 21908 7 3 2 99292 84287
0 21909 7 3 2 95367 80831
0 21910 7 1 2 99302 99305
0 21911 7 1 2 21906 21910
0 21912 5 1 1 21911
0 21913 7 1 2 69127 21912
0 21914 7 1 2 21888 21913
0 21915 5 1 1 21914
0 21916 7 1 2 73854 21915
0 21917 7 1 2 21849 21916
0 21918 5 1 1 21917
0 21919 7 1 2 21719 21918
0 21920 5 1 1 21919
0 21921 7 1 2 93882 21920
0 21922 5 1 1 21921
0 21923 7 1 2 92881 92877
0 21924 5 1 1 21923
0 21925 7 1 2 74534 21924
0 21926 5 1 1 21925
0 21927 7 1 2 779 21926
0 21928 5 1 1 21927
0 21929 7 1 2 65786 21928
0 21930 5 1 1 21929
0 21931 7 3 2 72663 76213
0 21932 7 1 2 99308 99138
0 21933 5 1 1 21932
0 21934 7 1 2 21930 21933
0 21935 5 1 1 21934
0 21936 7 1 2 72361 21935
0 21937 5 1 1 21936
0 21938 7 2 2 76310 96741
0 21939 7 1 2 96104 99311
0 21940 5 1 1 21939
0 21941 7 1 2 21937 21940
0 21942 5 1 1 21941
0 21943 7 1 2 64084 21942
0 21944 5 1 1 21943
0 21945 7 4 2 84350 93086
0 21946 5 1 1 99313
0 21947 7 4 2 71632 92837
0 21948 7 1 2 98456 99317
0 21949 7 1 2 99314 21948
0 21950 5 1 1 21949
0 21951 7 1 2 21944 21950
0 21952 5 1 1 21951
0 21953 7 3 2 74032 73855
0 21954 7 1 2 96193 99321
0 21955 5 1 1 21954
0 21956 7 1 2 79692 88228
0 21957 7 1 2 90396 21956
0 21958 5 1 1 21957
0 21959 7 1 2 21955 21958
0 21960 5 1 1 21959
0 21961 7 1 2 21952 21960
0 21962 5 1 1 21961
0 21963 7 6 2 66868 67278
0 21964 7 1 2 99324 95482
0 21965 7 1 2 97980 21964
0 21966 7 1 2 95955 21965
0 21967 7 2 2 95132 91285
0 21968 7 1 2 73856 99330
0 21969 7 1 2 21966 21968
0 21970 5 1 1 21969
0 21971 7 2 2 80316 92409
0 21972 7 2 2 89545 99332
0 21973 7 1 2 97278 81173
0 21974 7 1 2 96250 21973
0 21975 7 2 2 67279 77772
0 21976 7 1 2 79389 99336
0 21977 7 1 2 21974 21976
0 21978 7 1 2 99334 21977
0 21979 5 1 1 21978
0 21980 7 1 2 21970 21979
0 21981 7 1 2 21962 21980
0 21982 5 1 1 21981
0 21983 7 1 2 66989 21982
0 21984 5 1 1 21983
0 21985 7 1 2 64085 92333
0 21986 5 1 1 21985
0 21987 7 1 2 85435 82537
0 21988 5 1 1 21987
0 21989 7 1 2 21986 21988
0 21990 5 1 1 21989
0 21991 7 3 2 87409 96503
0 21992 7 1 2 73452 91182
0 21993 7 1 2 91321 98156
0 21994 7 1 2 21992 21993
0 21995 7 1 2 84673 21994
0 21996 7 1 2 99338 21995
0 21997 7 1 2 21990 21996
0 21998 5 1 1 21997
0 21999 7 1 2 21984 21998
0 22000 5 1 1 21999
0 22001 7 1 2 98974 22000
0 22002 5 1 1 22001
0 22003 7 1 2 21922 22002
0 22004 7 1 2 21242 22003
0 22005 7 1 2 18474 22004
0 22006 7 1 2 16804 22005
0 22007 7 1 2 11398 22006
0 22008 5 1 1 22007
0 22009 7 1 2 67153 22008
0 22010 5 1 1 22009
0 22011 7 6 2 69066 65688
0 22012 5 1 1 99341
0 22013 7 6 2 63978 70726
0 22014 5 1 1 99347
0 22015 7 5 2 22012 22014
0 22016 5 22 1 99353
0 22017 7 19 2 72362 82424
0 22018 5 1 1 99380
0 22019 7 19 2 67280 85490
0 22020 5 3 1 99399
0 22021 7 1 2 22018 99418
0 22022 5 1 1 22021
0 22023 7 1 2 90690 85684
0 22024 7 1 2 22022 22023
0 22025 5 1 1 22024
0 22026 7 5 2 65391 94860
0 22027 7 1 2 86003 96915
0 22028 7 1 2 99421 22027
0 22029 5 1 1 22028
0 22030 7 1 2 22025 22029
0 22031 5 1 1 22030
0 22032 7 1 2 66250 22031
0 22033 5 1 1 22032
0 22034 7 3 2 73453 77099
0 22035 5 3 1 99426
0 22036 7 5 2 99429 95247
0 22037 7 4 2 66990 98212
0 22038 5 1 1 99437
0 22039 7 1 2 96955 99438
0 22040 7 1 2 93411 22039
0 22041 7 1 2 99432 22040
0 22042 5 1 1 22041
0 22043 7 1 2 22033 22042
0 22044 5 1 1 22043
0 22045 7 1 2 69496 22044
0 22046 5 1 1 22045
0 22047 7 15 2 70793 67281
0 22048 5 2 1 99441
0 22049 7 9 2 64086 99442
0 22050 5 3 1 99458
0 22051 7 2 2 69128 98485
0 22052 5 2 1 99470
0 22053 7 1 2 99467 99472
0 22054 5 15 1 22053
0 22055 7 3 2 85904 99474
0 22056 7 2 2 76466 88413
0 22057 5 1 1 99492
0 22058 7 1 2 97375 94186
0 22059 5 1 1 22058
0 22060 7 1 2 95081 22059
0 22061 7 1 2 22057 22060
0 22062 5 1 1 22061
0 22063 7 1 2 87352 95092
0 22064 5 1 1 22063
0 22065 7 2 2 68635 22064
0 22066 5 1 1 99494
0 22067 7 2 2 87334 79023
0 22068 5 2 1 99496
0 22069 7 1 2 22066 99498
0 22070 5 1 1 22069
0 22071 7 1 2 66251 22070
0 22072 5 1 1 22071
0 22073 7 1 2 81856 95224
0 22074 7 1 2 78783 22073
0 22075 5 1 1 22074
0 22076 7 2 2 71345 79837
0 22077 5 2 1 99500
0 22078 7 1 2 92931 99502
0 22079 5 2 1 22078
0 22080 7 1 2 84904 99504
0 22081 5 1 1 22080
0 22082 7 3 2 71633 84703
0 22083 7 2 2 95998 99506
0 22084 5 1 1 99509
0 22085 7 1 2 68370 22084
0 22086 7 1 2 22081 22085
0 22087 7 1 2 22075 22086
0 22088 7 1 2 22072 22087
0 22089 5 1 1 22088
0 22090 7 1 2 22062 22089
0 22091 5 1 1 22090
0 22092 7 1 2 84737 92712
0 22093 5 1 1 22092
0 22094 7 1 2 83853 22093
0 22095 5 1 1 22094
0 22096 7 1 2 64685 22095
0 22097 5 1 1 22096
0 22098 7 1 2 886 92746
0 22099 5 2 1 22098
0 22100 7 1 2 85685 99511
0 22101 5 1 1 22100
0 22102 7 3 2 70156 94546
0 22103 5 1 1 99513
0 22104 7 1 2 95493 99514
0 22105 5 1 1 22104
0 22106 7 1 2 22101 22105
0 22107 7 1 2 22097 22106
0 22108 7 1 2 22091 22107
0 22109 5 1 1 22108
0 22110 7 1 2 99489 22109
0 22111 5 1 1 22110
0 22112 7 1 2 64087 83508
0 22113 5 1 1 22112
0 22114 7 1 2 20686 22113
0 22115 5 1 1 22114
0 22116 7 1 2 71634 22115
0 22117 5 1 1 22116
0 22118 7 1 2 70157 92463
0 22119 5 2 1 22118
0 22120 7 1 2 22117 99516
0 22121 5 1 1 22120
0 22122 7 1 2 67282 22121
0 22123 5 1 1 22122
0 22124 7 1 2 69129 82840
0 22125 7 2 2 99183 22124
0 22126 5 1 1 99518
0 22127 7 1 2 22123 22126
0 22128 5 1 1 22127
0 22129 7 1 2 70413 22128
0 22130 5 1 1 22129
0 22131 7 6 2 71815 67283
0 22132 7 2 2 65787 99520
0 22133 7 1 2 74901 99526
0 22134 5 1 1 22133
0 22135 7 1 2 22130 22134
0 22136 5 1 1 22135
0 22137 7 1 2 73454 22136
0 22138 5 1 1 22137
0 22139 7 3 2 65392 87335
0 22140 5 4 1 99528
0 22141 7 2 2 96916 99529
0 22142 5 1 1 99535
0 22143 7 1 2 83530 99536
0 22144 5 1 1 22143
0 22145 7 1 2 22138 22144
0 22146 5 1 1 22145
0 22147 7 1 2 68636 22146
0 22148 5 1 1 22147
0 22149 7 1 2 82492 82872
0 22150 5 1 1 22149
0 22151 7 1 2 99517 22150
0 22152 5 1 1 22151
0 22153 7 1 2 80696 22152
0 22154 5 1 1 22153
0 22155 7 5 2 80599 80867
0 22156 5 2 1 99537
0 22157 7 2 2 82493 99538
0 22158 5 1 1 99544
0 22159 7 1 2 96814 99545
0 22160 5 1 1 22159
0 22161 7 1 2 22154 22160
0 22162 5 1 1 22161
0 22163 7 1 2 68371 22162
0 22164 5 1 1 22163
0 22165 7 2 2 75635 83544
0 22166 5 1 1 99546
0 22167 7 1 2 82413 99547
0 22168 5 1 1 22167
0 22169 7 1 2 22164 22168
0 22170 5 1 1 22169
0 22171 7 1 2 67284 22170
0 22172 5 1 1 22171
0 22173 7 1 2 22148 22172
0 22174 5 1 1 22173
0 22175 7 1 2 69497 22174
0 22176 5 1 1 22175
0 22177 7 1 2 97895 94721
0 22178 5 1 1 22177
0 22179 7 1 2 22176 22178
0 22180 5 1 1 22179
0 22181 7 1 2 69795 22180
0 22182 5 1 1 22181
0 22183 7 9 2 69130 70414
0 22184 7 1 2 97896 99548
0 22185 7 1 2 95147 22184
0 22186 5 1 1 22185
0 22187 7 1 2 22182 22186
0 22188 5 1 1 22187
0 22189 7 1 2 71346 22188
0 22190 5 1 1 22189
0 22191 7 1 2 79167 82517
0 22192 5 1 1 22191
0 22193 7 4 2 69131 81716
0 22194 5 1 1 99557
0 22195 7 1 2 22192 22194
0 22196 5 1 1 22195
0 22197 7 1 2 69796 22196
0 22198 5 1 1 22197
0 22199 7 1 2 89210 11400
0 22200 5 2 1 22199
0 22201 7 1 2 69132 99561
0 22202 5 1 1 22201
0 22203 7 1 2 22198 22202
0 22204 5 1 1 22203
0 22205 7 1 2 73455 22204
0 22206 5 1 1 22205
0 22207 7 9 2 69133 65393
0 22208 7 3 2 66728 99563
0 22209 5 1 1 99572
0 22210 7 1 2 84775 81632
0 22211 5 1 1 22210
0 22212 7 1 2 22209 22211
0 22213 5 1 1 22212
0 22214 7 1 2 68372 22213
0 22215 5 1 1 22214
0 22216 7 1 2 69134 89202
0 22217 5 1 1 22216
0 22218 7 1 2 22215 22217
0 22219 5 1 1 22218
0 22220 7 1 2 65073 22219
0 22221 5 1 1 22220
0 22222 7 1 2 22206 22221
0 22223 5 1 1 22222
0 22224 7 1 2 71347 22223
0 22225 5 1 1 22224
0 22226 7 1 2 70158 80346
0 22227 5 3 1 22226
0 22228 7 1 2 73962 99575
0 22229 5 1 1 22228
0 22230 7 1 2 70415 22229
0 22231 5 1 1 22230
0 22232 7 1 2 68373 92733
0 22233 5 1 1 22232
0 22234 7 1 2 22231 22233
0 22235 5 1 1 22234
0 22236 7 1 2 66252 22235
0 22237 5 1 1 22236
0 22238 7 2 2 69498 85801
0 22239 5 1 1 99578
0 22240 7 1 2 64686 77122
0 22241 5 1 1 22240
0 22242 7 2 2 77309 22241
0 22243 7 1 2 85735 99580
0 22244 5 1 1 22243
0 22245 7 1 2 22239 22244
0 22246 7 1 2 22237 22245
0 22247 5 1 1 22246
0 22248 7 1 2 69135 22247
0 22249 5 1 1 22248
0 22250 7 1 2 22225 22249
0 22251 5 1 1 22250
0 22252 7 1 2 72363 22251
0 22253 5 1 1 22252
0 22254 7 1 2 66253 99433
0 22255 5 2 1 22254
0 22256 7 1 2 71348 95148
0 22257 5 1 1 22256
0 22258 7 1 2 99582 22257
0 22259 5 1 1 22258
0 22260 7 1 2 70416 22259
0 22261 5 1 1 22260
0 22262 7 1 2 71349 86778
0 22263 5 2 1 22262
0 22264 7 1 2 69499 99584
0 22265 5 2 1 22264
0 22266 7 1 2 79024 95207
0 22267 5 2 1 22266
0 22268 7 1 2 91785 99588
0 22269 7 1 2 99586 22268
0 22270 7 1 2 22261 22269
0 22271 5 1 1 22270
0 22272 7 1 2 96956 22271
0 22273 5 1 1 22272
0 22274 7 1 2 22253 22273
0 22275 5 1 1 22274
0 22276 7 1 2 70794 22275
0 22277 5 1 1 22276
0 22278 7 4 2 67285 85436
0 22279 7 2 2 93683 95144
0 22280 7 1 2 66254 99594
0 22281 5 2 1 22280
0 22282 7 1 2 99587 99596
0 22283 5 1 1 22282
0 22284 7 1 2 99590 22283
0 22285 5 1 1 22284
0 22286 7 1 2 90556 95705
0 22287 5 1 1 22286
0 22288 7 1 2 65788 22287
0 22289 5 1 1 22288
0 22290 7 1 2 69136 22289
0 22291 5 1 1 22290
0 22292 7 2 2 69500 99130
0 22293 7 1 2 80809 99598
0 22294 5 1 1 22293
0 22295 7 1 2 22291 22294
0 22296 5 1 1 22295
0 22297 7 1 2 70417 22296
0 22298 5 1 1 22297
0 22299 7 1 2 82425 82625
0 22300 5 1 1 22299
0 22301 7 1 2 72364 22300
0 22302 7 1 2 22298 22301
0 22303 5 1 1 22302
0 22304 7 1 2 92848 80810
0 22305 5 1 1 22304
0 22306 7 3 2 70418 85491
0 22307 5 1 1 99600
0 22308 7 1 2 67286 22307
0 22309 7 1 2 22305 22308
0 22310 5 1 1 22309
0 22311 7 1 2 97376 22310
0 22312 7 1 2 22303 22311
0 22313 5 1 1 22312
0 22314 7 1 2 22285 22313
0 22315 7 1 2 22277 22314
0 22316 7 1 2 22190 22315
0 22317 5 1 1 22316
0 22318 7 1 2 85267 22317
0 22319 5 1 1 22318
0 22320 7 1 2 22111 22319
0 22321 5 1 1 22320
0 22322 7 1 2 73099 22321
0 22323 5 1 1 22322
0 22324 7 1 2 22046 22323
0 22325 5 1 1 22324
0 22326 7 1 2 67154 22325
0 22327 5 1 1 22326
0 22328 7 2 2 70419 70795
0 22329 5 1 1 99603
0 22330 7 1 2 3218 22329
0 22331 5 1 1 22330
0 22332 7 1 2 97377 93795
0 22333 7 1 2 22331 22332
0 22334 5 1 1 22333
0 22335 7 1 2 66729 22334
0 22336 5 1 1 22335
0 22337 7 2 2 86345 76410
0 22338 5 1 1 99605
0 22339 7 1 2 68637 81564
0 22340 5 1 1 22339
0 22341 7 1 2 22338 22340
0 22342 5 1 1 22341
0 22343 7 1 2 64687 22342
0 22344 5 1 1 22343
0 22345 7 2 2 66255 75507
0 22346 7 1 2 83409 99607
0 22347 5 1 1 22346
0 22348 7 1 2 22344 22347
0 22349 5 1 1 22348
0 22350 7 1 2 70796 22349
0 22351 5 1 1 22350
0 22352 7 2 2 85492 76311
0 22353 5 1 1 99609
0 22354 7 2 2 69137 82005
0 22355 7 3 2 70420 82403
0 22356 5 1 1 99613
0 22357 7 1 2 99611 99614
0 22358 5 1 1 22357
0 22359 7 1 2 71816 22358
0 22360 7 1 2 22353 22359
0 22361 7 1 2 22351 22360
0 22362 5 1 1 22361
0 22363 7 1 2 22336 22362
0 22364 5 1 1 22363
0 22365 7 1 2 72365 22364
0 22366 5 1 1 22365
0 22367 7 3 2 82494 93818
0 22368 5 1 1 99616
0 22369 7 1 2 97378 99617
0 22370 5 1 1 22369
0 22371 7 3 2 66256 80347
0 22372 5 3 1 99619
0 22373 7 2 2 70159 92338
0 22374 7 1 2 99620 99625
0 22375 5 1 1 22374
0 22376 7 1 2 67287 22375
0 22377 7 1 2 22370 22376
0 22378 5 1 1 22377
0 22379 7 1 2 67155 22378
0 22380 7 1 2 22366 22379
0 22381 5 1 1 22380
0 22382 7 9 2 72210 72366
0 22383 5 1 1 99627
0 22384 7 5 2 72367 85493
0 22385 5 1 1 99636
0 22386 7 23 2 72211 82426
0 22387 5 1 1 99641
0 22388 7 1 2 22385 22387
0 22389 5 1 1 22388
0 22390 7 2 2 22383 22389
0 22391 7 1 2 75514 79534
0 22392 7 1 2 99664 22391
0 22393 5 1 1 22392
0 22394 7 1 2 22381 22393
0 22395 5 1 1 22394
0 22396 7 1 2 85268 22395
0 22397 5 1 1 22396
0 22398 7 1 2 71350 99665
0 22399 5 1 1 22398
0 22400 7 3 2 69138 99131
0 22401 7 9 2 72212 68638
0 22402 5 1 1 99669
0 22403 7 3 2 99521 99670
0 22404 7 1 2 99666 99678
0 22405 5 1 1 22404
0 22406 7 1 2 22399 22405
0 22407 5 1 1 22406
0 22408 7 6 2 72052 90714
0 22409 5 1 1 99681
0 22410 7 1 2 22038 22409
0 22411 5 1 1 22410
0 22412 7 1 2 22407 22411
0 22413 5 1 1 22412
0 22414 7 1 2 99637 80441
0 22415 5 1 1 22414
0 22416 7 1 2 97897 96865
0 22417 5 1 1 22416
0 22418 7 1 2 22415 22417
0 22419 5 1 1 22418
0 22420 7 1 2 89960 22419
0 22421 5 1 1 22420
0 22422 7 3 2 93604 99293
0 22423 7 1 2 65789 99687
0 22424 5 1 1 22423
0 22425 7 1 2 22421 22424
0 22426 5 1 1 22425
0 22427 7 1 2 67156 22426
0 22428 5 1 1 22427
0 22429 7 7 2 69139 70160
0 22430 7 1 2 95505 99690
0 22431 7 1 2 99679 22430
0 22432 5 1 1 22431
0 22433 7 1 2 22428 22432
0 22434 5 1 1 22433
0 22435 7 1 2 85905 22434
0 22436 5 1 1 22435
0 22437 7 1 2 22413 22436
0 22438 7 1 2 22397 22437
0 22439 5 1 1 22438
0 22440 7 1 2 71635 22439
0 22441 5 1 1 22440
0 22442 7 4 2 66991 97379
0 22443 7 2 2 67157 97952
0 22444 7 1 2 82495 80600
0 22445 7 1 2 84572 22444
0 22446 7 1 2 99701 22445
0 22447 7 1 2 99697 22446
0 22448 5 1 1 22447
0 22449 7 1 2 22441 22448
0 22450 5 1 1 22449
0 22451 7 1 2 69501 22450
0 22452 5 1 1 22451
0 22453 7 1 2 76214 98313
0 22454 5 1 1 22453
0 22455 7 1 2 84905 87201
0 22456 5 1 1 22455
0 22457 7 1 2 22454 22456
0 22458 5 1 1 22457
0 22459 7 1 2 99490 22458
0 22460 5 1 1 22459
0 22461 7 3 2 72368 85269
0 22462 7 2 2 82427 99703
0 22463 7 1 2 76312 78962
0 22464 5 1 1 22463
0 22465 7 2 2 95097 22464
0 22466 7 1 2 99706 99708
0 22467 5 1 1 22466
0 22468 7 1 2 22460 22467
0 22469 5 1 1 22468
0 22470 7 1 2 67158 22469
0 22471 5 1 1 22470
0 22472 7 5 2 66992 67288
0 22473 7 2 2 99671 99710
0 22474 7 1 2 70797 99549
0 22475 7 1 2 99715 22474
0 22476 7 3 2 71351 80465
0 22477 7 2 2 70161 84054
0 22478 7 1 2 99717 99720
0 22479 7 1 2 22475 22478
0 22480 5 1 1 22479
0 22481 7 1 2 22471 22480
0 22482 7 1 2 22452 22481
0 22483 5 1 1 22482
0 22484 7 1 2 68374 22483
0 22485 5 1 1 22484
0 22486 7 2 2 68639 79557
0 22487 5 1 1 99722
0 22488 7 1 2 64688 79587
0 22489 7 1 2 22487 22488
0 22490 5 1 1 22489
0 22491 7 1 2 69797 79541
0 22492 5 1 1 22491
0 22493 7 1 2 81717 22492
0 22494 7 1 2 22490 22493
0 22495 5 1 1 22494
0 22496 7 1 2 76313 88416
0 22497 5 1 1 22496
0 22498 7 1 2 94182 76215
0 22499 5 1 1 22498
0 22500 7 1 2 22499 92111
0 22501 7 1 2 22497 22500
0 22502 5 1 1 22501
0 22503 7 1 2 22495 22502
0 22504 5 1 1 22503
0 22505 7 1 2 99491 22504
0 22506 5 1 1 22505
0 22507 7 1 2 66730 84631
0 22508 5 1 1 22507
0 22509 7 3 2 97380 84826
0 22510 7 1 2 80849 99724
0 22511 5 1 1 22510
0 22512 7 1 2 22508 22511
0 22513 5 1 1 22512
0 22514 7 1 2 65790 22513
0 22515 5 1 1 22514
0 22516 7 3 2 64088 91443
0 22517 7 1 2 99727 90142
0 22518 5 1 1 22517
0 22519 7 1 2 22515 22518
0 22520 5 1 1 22519
0 22521 7 1 2 67289 22520
0 22522 5 1 1 22521
0 22523 7 1 2 76411 86539
0 22524 5 3 1 22523
0 22525 7 2 2 80293 84079
0 22526 5 2 1 99733
0 22527 7 1 2 99730 99735
0 22528 5 2 1 22527
0 22529 7 1 2 69798 99737
0 22530 5 1 1 22529
0 22531 7 2 2 70421 84159
0 22532 7 1 2 82006 99739
0 22533 5 1 1 22532
0 22534 7 1 2 22530 22533
0 22535 5 1 1 22534
0 22536 7 1 2 84952 22535
0 22537 5 1 1 22536
0 22538 7 5 2 69799 95506
0 22539 7 1 2 99741 87317
0 22540 5 1 1 22539
0 22541 7 1 2 72369 22540
0 22542 7 1 2 22537 22541
0 22543 5 1 1 22542
0 22544 7 3 2 65394 90472
0 22545 5 1 1 99746
0 22546 7 1 2 80442 22545
0 22547 5 1 1 22546
0 22548 7 1 2 82496 76467
0 22549 7 1 2 22547 22548
0 22550 5 1 1 22549
0 22551 7 1 2 97381 98792
0 22552 5 1 1 22551
0 22553 7 1 2 67290 22552
0 22554 7 1 2 22550 22553
0 22555 5 1 1 22554
0 22556 7 1 2 66527 22555
0 22557 7 1 2 22543 22556
0 22558 5 1 1 22557
0 22559 7 1 2 22522 22558
0 22560 5 1 1 22559
0 22561 7 1 2 69502 22560
0 22562 5 1 1 22561
0 22563 7 11 2 69140 98420
0 22564 5 2 1 99749
0 22565 7 2 2 81857 76580
0 22566 5 1 1 99762
0 22567 7 1 2 74651 99763
0 22568 5 1 1 22567
0 22569 7 2 2 78953 89256
0 22570 5 1 1 99764
0 22571 7 1 2 81718 22570
0 22572 7 1 2 95428 22571
0 22573 5 1 1 22572
0 22574 7 1 2 22568 22573
0 22575 5 1 1 22574
0 22576 7 1 2 99750 22575
0 22577 5 1 1 22576
0 22578 7 3 2 85494 76581
0 22579 7 1 2 67291 97778
0 22580 7 1 2 99766 22579
0 22581 5 1 1 22580
0 22582 7 1 2 22577 22581
0 22583 7 1 2 22562 22582
0 22584 5 1 1 22583
0 22585 7 1 2 73456 22584
0 22586 5 1 1 22585
0 22587 7 4 2 72370 81858
0 22588 7 1 2 82428 99769
0 22589 5 1 1 22588
0 22590 7 1 2 99419 22589
0 22591 5 1 1 22590
0 22592 7 1 2 76216 22591
0 22593 5 1 1 22592
0 22594 7 1 2 80697 99767
0 22595 5 1 1 22594
0 22596 7 8 2 73729 82497
0 22597 7 1 2 99773 77515
0 22598 7 1 2 94657 22597
0 22599 5 1 1 22598
0 22600 7 1 2 22595 22599
0 22601 5 1 1 22600
0 22602 7 1 2 67292 22601
0 22603 5 1 1 22602
0 22604 7 1 2 99381 76582
0 22605 7 1 2 86458 22604
0 22606 5 1 1 22605
0 22607 7 1 2 22603 22606
0 22608 5 1 1 22607
0 22609 7 1 2 66528 22608
0 22610 5 1 1 22609
0 22611 7 1 2 22593 22610
0 22612 7 1 2 22586 22611
0 22613 5 1 1 22612
0 22614 7 1 2 85270 22613
0 22615 5 1 1 22614
0 22616 7 1 2 22506 22615
0 22617 5 1 1 22616
0 22618 7 1 2 67159 22617
0 22619 5 1 1 22618
0 22620 7 1 2 22485 22619
0 22621 5 1 1 22620
0 22622 7 1 2 68028 22621
0 22623 5 1 1 22622
0 22624 7 1 2 63793 95276
0 22625 7 1 2 95634 22624
0 22626 7 3 2 80601 77803
0 22627 7 1 2 99716 99781
0 22628 7 1 2 22625 22627
0 22629 5 1 1 22628
0 22630 7 1 2 22623 22629
0 22631 7 1 2 22327 22630
0 22632 5 1 1 22631
0 22633 7 1 2 71061 22632
0 22634 5 1 1 22633
0 22635 7 1 2 64388 77577
0 22636 5 1 1 22635
0 22637 7 2 2 76217 89911
0 22638 5 1 1 99784
0 22639 7 1 2 22636 22638
0 22640 5 2 1 22639
0 22641 7 1 2 86023 94200
0 22642 5 1 1 22641
0 22643 7 1 2 86268 22642
0 22644 5 3 1 22643
0 22645 7 1 2 99786 99788
0 22646 5 1 1 22645
0 22647 7 1 2 90880 89028
0 22648 5 1 1 22647
0 22649 7 2 2 76583 77334
0 22650 7 1 2 79621 99791
0 22651 7 1 2 22648 22650
0 22652 5 1 1 22651
0 22653 7 1 2 22646 22652
0 22654 5 1 1 22653
0 22655 7 1 2 82429 22654
0 22656 5 1 1 22655
0 22657 7 7 2 73730 77210
0 22658 5 1 1 99793
0 22659 7 3 2 84827 99794
0 22660 5 3 1 99800
0 22661 7 8 2 65395 84963
0 22662 7 1 2 71636 99806
0 22663 5 1 1 22662
0 22664 7 1 2 99803 22663
0 22665 5 1 1 22664
0 22666 7 1 2 71352 22665
0 22667 5 1 1 22666
0 22668 7 4 2 80602 80076
0 22669 5 2 1 99814
0 22670 7 3 2 66257 80603
0 22671 5 3 1 99820
0 22672 7 1 2 99531 99823
0 22673 5 1 1 22672
0 22674 7 1 2 70162 22673
0 22675 5 1 1 22674
0 22676 7 1 2 99818 22675
0 22677 5 1 1 22676
0 22678 7 1 2 91675 22677
0 22679 5 1 1 22678
0 22680 7 1 2 22667 22679
0 22681 5 1 1 22680
0 22682 7 1 2 69800 22681
0 22683 5 1 1 22682
0 22684 7 1 2 99495 79468
0 22685 5 1 1 22684
0 22686 7 1 2 99530 81262
0 22687 5 1 1 22686
0 22688 7 1 2 68029 22687
0 22689 7 1 2 22685 22688
0 22690 7 1 2 22683 22689
0 22691 5 1 1 22690
0 22692 7 2 2 87347 83845
0 22693 5 1 1 99826
0 22694 7 1 2 81267 81330
0 22695 5 4 1 22694
0 22696 7 1 2 83027 99828
0 22697 5 1 1 22696
0 22698 7 1 2 22693 22697
0 22699 5 1 1 22698
0 22700 7 1 2 68640 22699
0 22701 5 1 1 22700
0 22702 7 3 2 81719 97382
0 22703 5 1 1 99832
0 22704 7 1 2 80884 99833
0 22705 5 1 1 22704
0 22706 7 1 2 73100 22705
0 22707 7 1 2 22701 22706
0 22708 5 1 1 22707
0 22709 7 1 2 68375 22708
0 22710 7 1 2 22691 22709
0 22711 5 1 1 22710
0 22712 7 2 2 71353 77688
0 22713 5 1 1 99835
0 22714 7 1 2 69503 75587
0 22715 7 2 2 22713 22714
0 22716 5 1 1 99837
0 22717 7 1 2 95465 99838
0 22718 5 1 1 22717
0 22719 7 1 2 79469 89275
0 22720 5 1 1 22719
0 22721 7 1 2 22718 22720
0 22722 5 1 1 22721
0 22723 7 1 2 70163 22722
0 22724 5 1 1 22723
0 22725 7 1 2 76072 98958
0 22726 5 1 1 22725
0 22727 7 1 2 22724 22726
0 22728 5 1 1 22727
0 22729 7 1 2 64689 22728
0 22730 5 1 1 22729
0 22731 7 3 2 65074 77211
0 22732 5 2 1 99839
0 22733 7 1 2 1939 99842
0 22734 5 1 1 22733
0 22735 7 1 2 68376 22734
0 22736 5 1 1 22735
0 22737 7 1 2 81118 22736
0 22738 5 1 1 22737
0 22739 7 1 2 68030 22738
0 22740 5 1 1 22739
0 22741 7 1 2 82386 74814
0 22742 5 2 1 22741
0 22743 7 1 2 71354 99844
0 22744 7 1 2 22740 22743
0 22745 5 1 1 22744
0 22746 7 1 2 75384 90217
0 22747 5 1 1 22746
0 22748 7 1 2 66258 97651
0 22749 7 1 2 22747 22748
0 22750 5 1 1 22749
0 22751 7 1 2 69801 22750
0 22752 7 1 2 22745 22751
0 22753 5 1 1 22752
0 22754 7 1 2 22730 22753
0 22755 5 1 1 22754
0 22756 7 1 2 81859 22755
0 22757 5 1 1 22756
0 22758 7 6 2 69802 75910
0 22759 5 3 1 99846
0 22760 7 2 2 90921 99852
0 22761 5 11 1 99855
0 22762 7 1 2 99857 95111
0 22763 5 1 1 22762
0 22764 7 3 2 70164 77666
0 22765 5 1 1 99868
0 22766 7 1 2 99869 99815
0 22767 5 1 1 22766
0 22768 7 1 2 22763 22767
0 22769 5 1 1 22768
0 22770 7 1 2 69504 22769
0 22771 5 1 1 22770
0 22772 7 1 2 77804 75849
0 22773 5 2 1 22772
0 22774 7 4 2 75970 95058
0 22775 7 1 2 69803 99873
0 22776 5 1 1 22775
0 22777 7 3 2 99871 22776
0 22778 5 2 1 99877
0 22779 7 2 2 82669 80481
0 22780 5 1 1 99882
0 22781 7 1 2 99880 99883
0 22782 5 1 1 22781
0 22783 7 1 2 22771 22782
0 22784 5 1 1 22783
0 22785 7 1 2 68641 22784
0 22786 5 1 1 22785
0 22787 7 1 2 22757 22786
0 22788 7 1 2 22711 22787
0 22789 5 1 1 22788
0 22790 7 1 2 85495 22789
0 22791 5 1 1 22790
0 22792 7 1 2 22656 22791
0 22793 5 1 1 22792
0 22794 7 1 2 85906 22793
0 22795 5 1 1 22794
0 22796 7 1 2 64089 99434
0 22797 5 1 1 22796
0 22798 7 1 2 65075 77087
0 22799 5 1 1 22798
0 22800 7 1 2 14088 22799
0 22801 5 2 1 22800
0 22802 7 1 2 73457 99884
0 22803 5 1 1 22802
0 22804 7 1 2 71817 94555
0 22805 5 3 1 22804
0 22806 7 1 2 22803 99886
0 22807 5 1 1 22806
0 22808 7 1 2 89912 22807
0 22809 5 1 1 22808
0 22810 7 1 2 22797 22809
0 22811 5 1 1 22810
0 22812 7 1 2 70422 22811
0 22813 5 1 1 22812
0 22814 7 1 2 81368 88447
0 22815 5 1 1 22814
0 22816 7 1 2 82915 22815
0 22817 5 1 1 22816
0 22818 7 1 2 80348 99870
0 22819 5 1 1 22818
0 22820 7 1 2 22817 22819
0 22821 5 1 1 22820
0 22822 7 1 2 65396 22821
0 22823 5 1 1 22822
0 22824 7 1 2 22823 14691
0 22825 5 1 1 22824
0 22826 7 1 2 65989 22825
0 22827 5 1 1 22826
0 22828 7 1 2 22813 22827
0 22829 5 1 1 22828
0 22830 7 1 2 71355 22829
0 22831 5 1 1 22830
0 22832 7 2 2 75571 93487
0 22833 5 1 1 99889
0 22834 7 2 2 65397 98574
0 22835 5 1 1 99891
0 22836 7 2 2 83545 97337
0 22837 5 1 1 99893
0 22838 7 1 2 65076 86931
0 22839 5 1 1 22838
0 22840 7 1 2 22837 22839
0 22841 5 2 1 22840
0 22842 7 1 2 70423 99895
0 22843 5 1 1 22842
0 22844 7 1 2 22835 22843
0 22845 5 2 1 22844
0 22846 7 1 2 68031 99897
0 22847 5 1 1 22846
0 22848 7 1 2 88822 74494
0 22849 5 1 1 22848
0 22850 7 1 2 22847 22849
0 22851 5 1 1 22850
0 22852 7 1 2 74150 22851
0 22853 5 1 1 22852
0 22854 7 1 2 22833 22853
0 22855 7 1 2 22831 22854
0 22856 5 1 1 22855
0 22857 7 1 2 69804 22856
0 22858 5 1 1 22857
0 22859 7 2 2 68642 83150
0 22860 5 1 1 99899
0 22861 7 1 2 77667 22860
0 22862 5 1 1 22861
0 22863 7 1 2 93288 22862
0 22864 5 1 1 22863
0 22865 7 1 2 69141 22864
0 22866 5 1 1 22865
0 22867 7 1 2 99898 74949
0 22868 5 1 1 22867
0 22869 7 1 2 71356 87026
0 22870 5 2 1 22869
0 22871 7 1 2 69142 99901
0 22872 5 1 1 22871
0 22873 7 3 2 74535 88823
0 22874 5 2 1 99903
0 22875 7 1 2 76073 99904
0 22876 5 1 1 22875
0 22877 7 1 2 22872 22876
0 22878 7 1 2 22868 22877
0 22879 5 1 1 22878
0 22880 7 1 2 64690 22879
0 22881 5 1 1 22880
0 22882 7 1 2 22866 22881
0 22883 5 1 1 22882
0 22884 7 1 2 65990 22883
0 22885 5 1 1 22884
0 22886 7 1 2 71357 99890
0 22887 5 1 1 22886
0 22888 7 1 2 65398 88318
0 22889 5 1 1 22888
0 22890 7 2 2 64691 77100
0 22891 5 1 1 99908
0 22892 7 1 2 66259 99909
0 22893 5 1 1 22892
0 22894 7 1 2 22889 22893
0 22895 5 1 1 22894
0 22896 7 2 2 77668 22895
0 22897 7 1 2 69143 99910
0 22898 5 1 1 22897
0 22899 7 1 2 22887 22898
0 22900 7 1 2 22885 22899
0 22901 7 1 2 22858 22900
0 22902 5 1 1 22901
0 22903 7 1 2 64389 22902
0 22904 5 1 1 22903
0 22905 7 1 2 99911 98339
0 22906 5 1 1 22905
0 22907 7 1 2 69805 95145
0 22908 5 1 1 22907
0 22909 7 1 2 86696 22908
0 22910 5 1 1 22909
0 22911 7 2 2 69806 84981
0 22912 5 1 1 99912
0 22913 7 1 2 99585 99913
0 22914 5 1 1 22913
0 22915 7 1 2 99597 22914
0 22916 7 1 2 22910 22915
0 22917 5 1 1 22916
0 22918 7 1 2 73101 22917
0 22919 5 1 1 22918
0 22920 7 1 2 91585 22919
0 22921 5 1 1 22920
0 22922 7 1 2 69505 22921
0 22923 5 2 1 22922
0 22924 7 1 2 99435 86697
0 22925 5 1 1 22924
0 22926 7 1 2 89279 22925
0 22927 5 1 1 22926
0 22928 7 1 2 69807 22927
0 22929 5 1 1 22928
0 22930 7 1 2 73905 74950
0 22931 5 4 1 22930
0 22932 7 1 2 22929 99916
0 22933 5 2 1 22932
0 22934 7 1 2 65991 99920
0 22935 5 1 1 22934
0 22936 7 1 2 99914 22935
0 22937 5 1 1 22936
0 22938 7 1 2 64090 22937
0 22939 5 1 1 22938
0 22940 7 1 2 22906 22939
0 22941 7 1 2 22904 22940
0 22942 5 1 1 22941
0 22943 7 1 2 70798 22942
0 22944 5 1 1 22943
0 22945 7 1 2 77212 99921
0 22946 5 1 1 22945
0 22947 7 1 2 99915 22946
0 22948 5 1 1 22947
0 22949 7 1 2 65791 22948
0 22950 5 1 1 22949
0 22951 7 1 2 80349 81358
0 22952 5 1 1 22951
0 22953 7 2 2 70424 97338
0 22954 5 1 1 99922
0 22955 7 1 2 85597 22954
0 22956 5 7 1 22955
0 22957 7 6 2 73458 99924
0 22958 7 1 2 68032 99931
0 22959 5 1 1 22958
0 22960 7 1 2 22952 22959
0 22961 5 1 1 22960
0 22962 7 1 2 97383 22961
0 22963 5 1 1 22962
0 22964 7 1 2 93508 95689
0 22965 5 1 1 22964
0 22966 7 2 2 78739 75074
0 22967 5 2 1 99937
0 22968 7 1 2 70425 94391
0 22969 5 1 1 22968
0 22970 7 1 2 1472 22969
0 22971 5 1 1 22970
0 22972 7 1 2 99938 22971
0 22973 5 1 1 22972
0 22974 7 1 2 22965 22973
0 22975 7 1 2 22963 22974
0 22976 5 1 1 22975
0 22977 7 1 2 70165 22976
0 22978 5 1 1 22977
0 22979 7 2 2 74851 86215
0 22980 7 1 2 76468 84130
0 22981 7 1 2 99941 22980
0 22982 5 1 1 22981
0 22983 7 1 2 22978 22982
0 22984 5 1 1 22983
0 22985 7 1 2 77335 22984
0 22986 5 1 1 22985
0 22987 7 1 2 22950 22986
0 22988 5 1 1 22987
0 22989 7 1 2 69144 22988
0 22990 5 1 1 22989
0 22991 7 1 2 74739 74169
0 22992 5 1 1 22991
0 22993 7 4 2 70166 74426
0 22994 7 1 2 74781 99943
0 22995 5 1 1 22994
0 22996 7 1 2 22992 22995
0 22997 5 1 1 22996
0 22998 7 1 2 76469 22997
0 22999 5 1 1 22998
0 23000 7 1 2 82430 80159
0 23001 5 1 1 23000
0 23002 7 1 2 22999 23001
0 23003 5 1 1 23002
0 23004 7 1 2 66529 23003
0 23005 5 1 1 23004
0 23006 7 1 2 69145 92112
0 23007 5 1 1 23006
0 23008 7 4 2 64692 74951
0 23009 5 2 1 99947
0 23010 7 1 2 83311 99951
0 23011 5 13 1 23010
0 23012 7 1 2 98301 99953
0 23013 5 1 1 23012
0 23014 7 1 2 23007 23013
0 23015 5 1 1 23014
0 23016 7 1 2 70799 23015
0 23017 5 1 1 23016
0 23018 7 1 2 23005 23017
0 23019 5 1 1 23018
0 23020 7 1 2 77336 23019
0 23021 5 1 1 23020
0 23022 7 1 2 73963 74129
0 23023 7 1 2 99768 23022
0 23024 5 1 1 23023
0 23025 7 10 2 70800 66260
0 23026 7 2 2 84351 99966
0 23027 7 1 2 77213 77868
0 23028 7 1 2 99976 23027
0 23029 5 1 1 23028
0 23030 7 1 2 23024 23029
0 23031 7 1 2 23021 23030
0 23032 5 1 1 23031
0 23033 7 1 2 80698 23032
0 23034 5 1 1 23033
0 23035 7 1 2 22990 23034
0 23036 7 1 2 22944 23035
0 23037 5 1 1 23036
0 23038 7 1 2 85271 23037
0 23039 5 1 1 23038
0 23040 7 1 2 22795 23039
0 23041 5 1 1 23040
0 23042 7 1 2 67293 23041
0 23043 5 1 1 23042
0 23044 7 1 2 76470 94315
0 23045 5 1 1 23044
0 23046 7 1 2 85359 12869
0 23047 5 2 1 23046
0 23048 7 1 2 65992 99978
0 23049 5 1 1 23048
0 23050 7 1 2 21669 23049
0 23051 5 1 1 23050
0 23052 7 1 2 76314 23051
0 23053 5 1 1 23052
0 23054 7 1 2 98672 86326
0 23055 5 1 1 23054
0 23056 7 1 2 23053 23055
0 23057 5 1 1 23056
0 23058 7 1 2 70167 23057
0 23059 5 1 1 23058
0 23060 7 1 2 99829 94611
0 23061 5 1 1 23060
0 23062 7 2 2 85272 86378
0 23063 5 1 1 99980
0 23064 7 1 2 95546 87527
0 23065 5 1 1 23064
0 23066 7 1 2 23063 23065
0 23067 5 1 1 23066
0 23068 7 2 2 68643 97384
0 23069 7 1 2 23067 99982
0 23070 5 1 1 23069
0 23071 7 1 2 23061 23070
0 23072 7 1 2 23059 23071
0 23073 5 1 1 23072
0 23074 7 1 2 71637 23073
0 23075 5 1 1 23074
0 23076 7 4 2 80077 84175
0 23077 5 1 1 99984
0 23078 7 1 2 71358 81994
0 23079 5 1 1 23078
0 23080 7 1 2 23077 23079
0 23081 5 1 1 23080
0 23082 7 1 2 69808 23081
0 23083 5 1 1 23082
0 23084 7 1 2 97357 87668
0 23085 5 1 1 23084
0 23086 7 1 2 23083 23085
0 23087 5 1 1 23086
0 23088 7 1 2 81860 23087
0 23089 5 1 1 23088
0 23090 7 1 2 99621 94310
0 23091 5 1 1 23090
0 23092 7 2 2 71359 99801
0 23093 5 1 1 99988
0 23094 7 1 2 23091 23093
0 23095 5 1 1 23094
0 23096 7 1 2 69809 23095
0 23097 5 1 1 23096
0 23098 7 2 2 64693 80294
0 23099 7 1 2 80350 79470
0 23100 7 1 2 99990 23099
0 23101 5 1 1 23100
0 23102 7 1 2 23097 23101
0 23103 7 1 2 23089 23102
0 23104 5 1 1 23103
0 23105 7 1 2 85907 23104
0 23106 5 1 1 23105
0 23107 7 1 2 99709 93437
0 23108 5 1 1 23107
0 23109 7 3 2 81861 77214
0 23110 7 1 2 85273 77920
0 23111 5 1 1 23110
0 23112 7 5 2 65077 85908
0 23113 5 1 1 99995
0 23114 7 1 2 76471 99996
0 23115 5 1 1 23114
0 23116 7 1 2 23111 23115
0 23117 5 1 1 23116
0 23118 7 1 2 99992 23117
0 23119 5 1 1 23118
0 23120 7 1 2 68377 23119
0 23121 7 1 2 23108 23120
0 23122 7 1 2 23106 23121
0 23123 7 1 2 23075 23122
0 23124 5 1 1 23123
0 23125 7 2 2 68849 93384
0 23126 7 1 2 76218 100000
0 23127 5 1 1 23126
0 23128 7 1 2 76584 93720
0 23129 5 1 1 23128
0 23130 7 1 2 23127 23129
0 23131 5 1 1 23130
0 23132 7 1 2 69506 23131
0 23133 5 1 1 23132
0 23134 7 1 2 81324 91825
0 23135 5 1 1 23134
0 23136 7 1 2 23133 23135
0 23137 5 1 1 23136
0 23138 7 1 2 81862 23137
0 23139 5 1 1 23138
0 23140 7 4 2 70168 80604
0 23141 5 3 1 100002
0 23142 7 1 2 90825 100003
0 23143 5 2 1 23142
0 23144 7 1 2 13022 100009
0 23145 5 2 1 23144
0 23146 7 1 2 97385 100011
0 23147 5 1 1 23146
0 23148 7 1 2 83846 86368
0 23149 5 1 1 23148
0 23150 7 1 2 64390 94550
0 23151 5 2 1 23150
0 23152 7 1 2 79585 100013
0 23153 5 1 1 23152
0 23154 7 1 2 23149 23153
0 23155 5 1 1 23154
0 23156 7 1 2 81720 23155
0 23157 5 1 1 23156
0 23158 7 1 2 23147 23157
0 23159 5 1 1 23158
0 23160 7 1 2 85274 23159
0 23161 5 1 1 23160
0 23162 7 1 2 81296 94619
0 23163 5 1 1 23162
0 23164 7 1 2 73459 23163
0 23165 7 1 2 23161 23164
0 23166 7 1 2 23139 23165
0 23167 5 1 1 23166
0 23168 7 1 2 23124 23167
0 23169 5 1 1 23168
0 23170 7 1 2 81863 93438
0 23171 7 1 2 87202 23170
0 23172 5 1 1 23171
0 23173 7 2 2 82007 89084
0 23174 7 1 2 95494 79052
0 23175 7 1 2 100015 23174
0 23176 5 1 1 23175
0 23177 7 1 2 68033 23176
0 23178 7 1 2 23172 23177
0 23179 7 1 2 23169 23178
0 23180 5 1 1 23179
0 23181 7 1 2 79888 83650
0 23182 5 17 1 23181
0 23183 7 1 2 85275 100017
0 23184 5 1 1 23183
0 23185 7 1 2 90715 91807
0 23186 5 1 1 23185
0 23187 7 1 2 23184 23186
0 23188 5 1 1 23187
0 23189 7 1 2 80351 23188
0 23190 5 1 1 23189
0 23191 7 2 2 68850 92762
0 23192 7 2 2 71638 76355
0 23193 7 1 2 100034 100036
0 23194 5 1 1 23193
0 23195 7 1 2 23190 23194
0 23196 5 1 1 23195
0 23197 7 1 2 70169 23196
0 23198 5 1 1 23197
0 23199 7 3 2 69810 82387
0 23200 5 1 1 100038
0 23201 7 1 2 80352 100039
0 23202 7 1 2 92222 23201
0 23203 5 1 1 23202
0 23204 7 1 2 23198 23203
0 23205 5 1 1 23204
0 23206 7 1 2 70426 23205
0 23207 5 1 1 23206
0 23208 7 1 2 13795 83443
0 23209 5 1 1 23208
0 23210 7 1 2 70170 23209
0 23211 5 1 1 23210
0 23212 7 1 2 85686 82713
0 23213 5 1 1 23212
0 23214 7 1 2 23211 23213
0 23215 5 1 1 23214
0 23216 7 1 2 90691 23215
0 23217 5 1 1 23216
0 23218 7 1 2 79900 83780
0 23219 5 8 1 23218
0 23220 7 1 2 85276 100041
0 23221 5 1 1 23220
0 23222 7 1 2 86492 85829
0 23223 7 1 2 92911 23222
0 23224 5 1 1 23223
0 23225 7 1 2 23221 23224
0 23226 5 1 1 23225
0 23227 7 1 2 70427 23226
0 23228 5 1 1 23227
0 23229 7 2 2 80927 91737
0 23230 5 1 1 100049
0 23231 7 2 2 91733 23230
0 23232 7 2 2 81721 80097
0 23233 7 4 2 73460 86346
0 23234 5 1 1 100055
0 23235 7 1 2 64694 100056
0 23236 5 1 1 23235
0 23237 7 1 2 100053 23236
0 23238 5 1 1 23237
0 23239 7 1 2 100051 23238
0 23240 5 1 1 23239
0 23241 7 1 2 85277 23240
0 23242 5 1 1 23241
0 23243 7 1 2 23228 23242
0 23244 7 1 2 23217 23243
0 23245 5 1 1 23244
0 23246 7 1 2 69507 23245
0 23247 5 1 1 23246
0 23248 7 1 2 84176 91870
0 23249 5 1 1 23248
0 23250 7 3 2 94031 74921
0 23251 5 2 1 100059
0 23252 7 1 2 94531 100060
0 23253 5 1 1 23252
0 23254 7 1 2 23249 23253
0 23255 5 1 1 23254
0 23256 7 1 2 82264 23255
0 23257 5 1 1 23256
0 23258 7 1 2 23247 23257
0 23259 7 1 2 23207 23258
0 23260 5 1 1 23259
0 23261 7 1 2 71360 23260
0 23262 5 1 1 23261
0 23263 7 2 2 71639 79811
0 23264 5 1 1 100064
0 23265 7 1 2 80850 85626
0 23266 5 1 1 23265
0 23267 7 1 2 23264 23266
0 23268 5 1 1 23267
0 23269 7 1 2 85278 23268
0 23270 5 1 1 23269
0 23271 7 2 2 63794 94063
0 23272 5 1 1 100066
0 23273 7 1 2 85909 82847
0 23274 5 1 1 23273
0 23275 7 1 2 23272 23274
0 23276 5 1 1 23275
0 23277 7 1 2 76649 23276
0 23278 5 1 1 23277
0 23279 7 1 2 23270 23278
0 23280 7 1 2 66993 84055
0 23281 5 1 1 23280
0 23282 7 1 2 100037 94396
0 23283 5 1 1 23282
0 23284 7 1 2 23281 23283
0 23285 5 1 1 23284
0 23286 7 1 2 81864 23285
0 23287 5 1 1 23286
0 23288 7 1 2 80964 89705
0 23289 5 1 1 23288
0 23290 7 1 2 94612 89068
0 23291 7 1 2 23289 23290
0 23292 5 1 1 23291
0 23293 7 1 2 23287 23292
0 23294 7 1 2 23279 23293
0 23295 5 1 1 23294
0 23296 7 1 2 66261 23295
0 23297 5 1 1 23296
0 23298 7 2 2 72053 90620
0 23299 7 1 2 95706 83965
0 23300 5 2 1 23299
0 23301 7 1 2 69811 86444
0 23302 5 1 1 23301
0 23303 7 1 2 100070 23302
0 23304 5 1 1 23303
0 23305 7 1 2 100068 23304
0 23306 5 1 1 23305
0 23307 7 1 2 86004 95066
0 23308 5 1 1 23307
0 23309 7 1 2 23306 23308
0 23310 5 1 1 23309
0 23311 7 1 2 75385 23310
0 23312 5 1 1 23311
0 23313 7 3 2 68644 76650
0 23314 5 1 1 100072
0 23315 7 1 2 85279 85736
0 23316 7 1 2 100073 23315
0 23317 5 1 1 23316
0 23318 7 1 2 23312 23317
0 23319 7 1 2 23297 23318
0 23320 5 1 1 23319
0 23321 7 1 2 69508 23320
0 23322 5 1 1 23321
0 23323 7 1 2 66994 74852
0 23324 7 1 2 99721 23323
0 23325 7 1 2 99816 23324
0 23326 5 1 1 23325
0 23327 7 1 2 73102 23326
0 23328 7 1 2 23322 23327
0 23329 7 1 2 23262 23328
0 23330 5 1 1 23329
0 23331 7 1 2 23180 23330
0 23332 5 1 1 23331
0 23333 7 1 2 23045 23332
0 23334 5 1 1 23333
0 23335 7 1 2 99382 23334
0 23336 5 1 1 23335
0 23337 7 1 2 23043 23336
0 23338 5 1 1 23337
0 23339 7 1 2 67160 23338
0 23340 5 1 1 23339
0 23341 7 1 2 85280 75515
0 23342 5 1 1 23341
0 23343 7 1 2 83500 90731
0 23344 5 1 1 23343
0 23345 7 1 2 23342 23344
0 23346 5 1 1 23345
0 23347 7 15 2 72213 67294
0 23348 7 4 2 69146 100075
0 23349 5 1 1 100090
0 23350 7 2 2 100091 95349
0 23351 5 1 1 100094
0 23352 7 1 2 23346 100095
0 23353 5 1 1 23352
0 23354 7 2 2 65993 84738
0 23355 5 3 1 100096
0 23356 7 1 2 99564 100097
0 23357 5 1 1 23356
0 23358 7 5 2 64091 77148
0 23359 5 2 1 100101
0 23360 7 1 2 70428 100102
0 23361 5 1 1 23360
0 23362 7 1 2 23357 23361
0 23363 5 1 1 23362
0 23364 7 1 2 98486 23363
0 23365 5 1 1 23364
0 23366 7 6 2 70429 72371
0 23367 7 3 2 77149 100108
0 23368 5 1 1 100114
0 23369 7 1 2 85437 100115
0 23370 5 1 1 23369
0 23371 7 4 2 84739 84337
0 23372 7 1 2 64092 97733
0 23373 7 1 2 100117 23372
0 23374 5 1 1 23373
0 23375 7 1 2 23370 23374
0 23376 7 1 2 23365 23375
0 23377 5 1 1 23376
0 23378 7 1 2 85910 23377
0 23379 5 1 1 23378
0 23380 7 4 2 85496 77150
0 23381 5 2 1 100121
0 23382 7 1 2 82431 77215
0 23383 5 1 1 23382
0 23384 7 1 2 100125 23383
0 23385 5 1 1 23384
0 23386 7 1 2 99704 23385
0 23387 5 1 1 23386
0 23388 7 1 2 23379 23387
0 23389 5 1 1 23388
0 23390 7 1 2 70171 23389
0 23391 5 1 1 23390
0 23392 7 2 2 67295 85281
0 23393 7 1 2 77216 100127
0 23394 5 1 1 23393
0 23395 7 2 2 81865 85282
0 23396 5 2 1 100129
0 23397 7 1 2 94620 100131
0 23398 5 1 1 23397
0 23399 7 1 2 23398 98286
0 23400 5 1 1 23399
0 23401 7 1 2 23394 23400
0 23402 5 1 1 23401
0 23403 7 1 2 85497 23402
0 23404 5 1 1 23403
0 23405 7 1 2 99707 99993
0 23406 5 1 1 23405
0 23407 7 1 2 23404 23406
0 23408 7 1 2 23391 23407
0 23409 5 1 1 23408
0 23410 7 1 2 67161 23409
0 23411 5 1 1 23410
0 23412 7 1 2 23353 23411
0 23413 5 1 1 23412
0 23414 7 1 2 76472 23413
0 23415 5 1 1 23414
0 23416 7 1 2 70172 98213
0 23417 7 1 2 99711 23416
0 23418 7 2 2 70801 68645
0 23419 7 13 2 69147 72214
0 23420 7 3 2 100133 100135
0 23421 5 1 1 100148
0 23422 7 1 2 99192 100149
0 23423 7 1 2 23417 23422
0 23424 5 1 1 23423
0 23425 7 1 2 23415 23424
0 23426 5 1 1 23425
0 23427 7 1 2 76315 77606
0 23428 7 1 2 23426 23427
0 23429 5 1 1 23428
0 23430 7 7 2 66995 72215
0 23431 7 1 2 99077 100151
0 23432 7 2 2 80811 23431
0 23433 7 2 2 99132 86698
0 23434 7 6 2 69148 69812
0 23435 5 1 1 100162
0 23436 7 1 2 90893 100163
0 23437 7 1 2 100160 23436
0 23438 7 1 2 100158 23437
0 23439 5 1 1 23438
0 23440 7 1 2 23429 23439
0 23441 7 1 2 23340 23440
0 23442 7 1 2 22634 23441
0 23443 5 1 1 23442
0 23444 7 54 2 90585 75666
0 23445 5 4 1 100168
0 23446 7 1 2 23443 100169
0 23447 5 1 1 23446
0 23448 7 1 2 90040 93456
0 23449 5 1 1 23448
0 23450 7 2 2 66996 99858
0 23451 7 1 2 98214 100226
0 23452 5 1 1 23451
0 23453 7 1 2 23449 23452
0 23454 5 1 1 23453
0 23455 7 1 2 68378 23454
0 23456 5 1 1 23455
0 23457 7 2 2 76473 83665
0 23458 7 1 2 86005 100228
0 23459 5 1 1 23458
0 23460 7 1 2 23456 23459
0 23461 5 1 1 23460
0 23462 7 1 2 71640 23461
0 23463 5 1 1 23462
0 23464 7 1 2 77536 93457
0 23465 5 1 1 23464
0 23466 7 1 2 23463 23465
0 23467 5 1 1 23466
0 23468 7 1 2 100170 23467
0 23469 5 1 1 23468
0 23470 7 6 2 68851 84319
0 23471 7 3 2 70677 71361
0 23472 7 1 2 71641 100236
0 23473 7 2 2 100230 23472
0 23474 7 4 2 70430 70631
0 23475 7 2 2 69813 100241
0 23476 7 1 2 76356 97716
0 23477 7 1 2 100245 23476
0 23478 7 1 2 100239 23477
0 23479 5 1 1 23478
0 23480 7 1 2 23469 23479
0 23481 5 1 1 23480
0 23482 7 1 2 70173 23481
0 23483 5 1 1 23482
0 23484 7 3 2 87699 79961
0 23485 5 1 1 100247
0 23486 7 1 2 77568 23485
0 23487 5 5 1 23486
0 23488 7 1 2 69149 100250
0 23489 5 1 1 23488
0 23490 7 3 2 74135 83322
0 23491 7 2 2 75572 100255
0 23492 5 1 1 100258
0 23493 7 1 2 23489 23492
0 23494 5 1 1 23493
0 23495 7 33 2 76805 91271
0 23496 7 1 2 99439 100260
0 23497 7 1 2 23494 23496
0 23498 5 1 1 23497
0 23499 7 1 2 23483 23498
0 23500 5 1 1 23499
0 23501 7 1 2 65792 23500
0 23502 5 1 1 23501
0 23503 7 7 2 93895 96407
0 23504 7 1 2 70431 85447
0 23505 7 1 2 100293 23504
0 23506 7 1 2 100251 23505
0 23507 5 1 1 23506
0 23508 7 1 2 23502 23507
0 23509 5 1 1 23508
0 23510 7 1 2 71062 23509
0 23511 5 1 1 23510
0 23512 7 1 2 76474 93684
0 23513 5 1 1 23512
0 23514 7 5 2 90586 85843
0 23515 7 1 2 100300 82770
0 23516 7 1 2 99610 23515
0 23517 7 1 2 23513 23516
0 23518 5 1 1 23517
0 23519 7 1 2 67296 23518
0 23520 7 1 2 23511 23519
0 23521 5 1 1 23520
0 23522 7 1 2 75573 93896
0 23523 7 3 2 94584 86524
0 23524 7 1 2 100305 95328
0 23525 7 1 2 23522 23524
0 23526 5 2 1 23525
0 23527 7 2 2 77629 77607
0 23528 5 3 1 100310
0 23529 7 3 2 75971 100311
0 23530 7 1 2 69814 100315
0 23531 5 1 1 23530
0 23532 7 1 2 99917 23531
0 23533 5 3 1 23532
0 23534 7 1 2 91821 87745
0 23535 7 1 2 91347 23534
0 23536 7 1 2 100318 23535
0 23537 5 1 1 23536
0 23538 7 1 2 100308 23537
0 23539 5 1 1 23538
0 23540 7 1 2 85498 23539
0 23541 5 1 1 23540
0 23542 7 1 2 66262 84551
0 23543 5 2 1 23542
0 23544 7 2 2 75075 77869
0 23545 5 2 1 100323
0 23546 7 1 2 100321 100325
0 23547 5 4 1 23546
0 23548 7 1 2 64695 100327
0 23549 5 1 1 23548
0 23550 7 1 2 92923 77885
0 23551 5 2 1 23550
0 23552 7 2 2 23549 100331
0 23553 5 4 1 100333
0 23554 7 9 2 70678 70802
0 23555 7 4 2 71939 100339
0 23556 7 1 2 99565 77831
0 23557 7 1 2 83883 23556
0 23558 7 1 2 100348 23557
0 23559 7 1 2 100335 23558
0 23560 5 1 1 23559
0 23561 7 1 2 23541 23560
0 23562 5 1 1 23561
0 23563 7 1 2 71063 23562
0 23564 5 1 1 23563
0 23565 7 1 2 85283 81359
0 23566 7 2 2 88892 84605
0 23567 7 1 2 93111 100352
0 23568 7 1 2 23565 23567
0 23569 5 1 1 23568
0 23570 7 1 2 72372 23569
0 23571 7 1 2 23564 23570
0 23572 5 1 1 23571
0 23573 7 1 2 67162 23572
0 23574 7 1 2 23521 23573
0 23575 5 1 1 23574
0 23576 7 1 2 85360 20675
0 23577 5 1 1 23576
0 23578 7 1 2 100171 23577
0 23579 7 1 2 100319 23578
0 23580 5 1 1 23579
0 23581 7 1 2 100309 23580
0 23582 5 1 1 23581
0 23583 7 2 2 99443 95280
0 23584 7 1 2 72216 100354
0 23585 7 1 2 23582 23584
0 23586 5 1 1 23585
0 23587 7 1 2 23575 23586
0 23588 5 1 1 23587
0 23589 7 1 2 69509 23588
0 23590 5 1 1 23589
0 23591 7 2 2 100301 82763
0 23592 7 2 2 69815 93685
0 23593 5 1 1 100358
0 23594 7 1 2 23593 86389
0 23595 7 1 2 100356 23594
0 23596 5 1 1 23595
0 23597 7 1 2 97717 83621
0 23598 7 2 2 100246 23597
0 23599 7 3 2 70679 65994
0 23600 7 1 2 73906 100362
0 23601 7 1 2 100360 23600
0 23602 7 1 2 98635 23601
0 23603 5 1 1 23602
0 23604 7 1 2 23596 23603
0 23605 5 1 1 23604
0 23606 7 1 2 71362 23605
0 23607 5 1 1 23606
0 23608 7 2 2 88893 75860
0 23609 7 3 2 66263 85284
0 23610 7 1 2 93198 100367
0 23611 7 1 2 100365 23610
0 23612 5 1 1 23611
0 23613 7 1 2 23607 23612
0 23614 5 1 1 23613
0 23615 7 1 2 85499 23614
0 23616 5 1 1 23615
0 23617 7 1 2 99550 84068
0 23618 7 1 2 100349 23617
0 23619 7 1 2 100252 23618
0 23620 5 1 1 23619
0 23621 7 1 2 99859 79812
0 23622 5 1 1 23621
0 23623 7 1 2 73461 100229
0 23624 5 1 1 23623
0 23625 7 1 2 23622 23624
0 23626 5 1 1 23625
0 23627 7 2 2 74427 76916
0 23628 7 3 2 70174 65640
0 23629 7 1 2 100372 91830
0 23630 7 1 2 100370 23629
0 23631 7 1 2 23626 23630
0 23632 5 1 1 23631
0 23633 7 1 2 23620 23632
0 23634 5 1 1 23633
0 23635 7 1 2 64391 89434
0 23636 7 1 2 23634 23635
0 23637 5 1 1 23636
0 23638 7 1 2 23616 23637
0 23639 5 1 1 23638
0 23640 7 1 2 67297 23639
0 23641 5 1 1 23640
0 23642 7 2 2 85844 76870
0 23643 7 1 2 93581 100375
0 23644 5 1 1 23643
0 23645 7 1 2 71363 100363
0 23646 7 1 2 100361 23645
0 23647 5 1 1 23646
0 23648 7 1 2 23644 23647
0 23649 5 1 1 23648
0 23650 7 8 2 70803 71642
0 23651 7 4 2 68379 100377
0 23652 7 3 2 74351 97100
0 23653 7 1 2 100385 100389
0 23654 7 1 2 23649 23653
0 23655 5 1 1 23654
0 23656 7 1 2 23641 23655
0 23657 5 1 1 23656
0 23658 7 1 2 67163 23657
0 23659 5 1 1 23658
0 23660 7 1 2 23590 23659
0 23661 5 1 1 23660
0 23662 7 1 2 82975 23661
0 23663 5 1 1 23662
0 23664 7 1 2 85361 94621
0 23665 5 1 1 23664
0 23666 7 6 2 100350 84069
0 23667 7 2 2 74536 100392
0 23668 7 1 2 98602 100398
0 23669 5 1 1 23668
0 23670 7 5 2 65641 65793
0 23671 5 1 1 100400
0 23672 7 3 2 76917 100401
0 23673 7 1 2 77608 99325
0 23674 7 1 2 100405 23673
0 23675 5 1 1 23674
0 23676 7 1 2 23669 23675
0 23677 5 1 1 23676
0 23678 7 1 2 64093 23677
0 23679 5 1 1 23678
0 23680 7 1 2 70175 88025
0 23681 7 3 2 93729 23680
0 23682 7 1 2 97963 79696
0 23683 7 1 2 100408 23682
0 23684 5 1 1 23683
0 23685 7 1 2 23679 23684
0 23686 5 1 1 23685
0 23687 7 1 2 67164 23686
0 23688 5 1 1 23687
0 23689 7 1 2 75574 100092
0 23690 7 1 2 100399 23689
0 23691 5 1 1 23690
0 23692 7 1 2 23688 23691
0 23693 5 1 1 23692
0 23694 7 1 2 76475 23693
0 23695 5 1 1 23694
0 23696 7 2 2 74389 93582
0 23697 7 2 2 66869 67165
0 23698 7 6 2 71643 67298
0 23699 7 1 2 75575 100415
0 23700 7 1 2 100413 23699
0 23701 7 1 2 100411 23700
0 23702 5 1 1 23701
0 23703 7 1 2 23695 23702
0 23704 5 1 1 23703
0 23705 7 1 2 80220 23704
0 23706 5 1 1 23705
0 23707 7 22 2 67166 72373
0 23708 7 1 2 100340 100421
0 23709 7 1 2 87864 91130
0 23710 7 1 2 23708 23709
0 23711 7 2 2 79471 93730
0 23712 7 1 2 79697 100443
0 23713 7 1 2 23710 23712
0 23714 5 1 1 23713
0 23715 7 1 2 23706 23714
0 23716 5 1 1 23715
0 23717 7 1 2 23665 23716
0 23718 5 1 1 23717
0 23719 7 1 2 83531 98806
0 23720 5 5 1 23719
0 23721 7 1 2 70432 99894
0 23722 5 1 1 23721
0 23723 7 1 2 100445 23722
0 23724 5 3 1 23723
0 23725 7 1 2 75911 84352
0 23726 7 1 2 100450 23725
0 23727 5 1 1 23726
0 23728 7 1 2 95707 93615
0 23729 7 1 2 87843 23728
0 23730 5 1 1 23729
0 23731 7 1 2 23727 23730
0 23732 5 1 1 23731
0 23733 7 1 2 85911 23732
0 23734 5 1 1 23733
0 23735 7 2 2 65078 82916
0 23736 5 3 1 100453
0 23737 7 1 2 69816 100455
0 23738 5 2 1 23737
0 23739 7 1 2 75912 100458
0 23740 5 1 1 23739
0 23741 7 1 2 64696 82917
0 23742 7 1 2 95060 23741
0 23743 5 1 1 23742
0 23744 7 1 2 23740 23743
0 23745 5 1 1 23744
0 23746 7 1 2 69150 23745
0 23747 5 1 1 23746
0 23748 7 2 2 68034 80443
0 23749 7 1 2 100256 100460
0 23750 5 1 1 23749
0 23751 7 1 2 23747 23750
0 23752 5 1 1 23751
0 23753 7 1 2 68380 23752
0 23754 5 1 1 23753
0 23755 7 2 2 74652 80353
0 23756 5 2 1 100462
0 23757 7 1 2 82741 100463
0 23758 5 1 1 23757
0 23759 7 1 2 87303 78327
0 23760 5 1 1 23759
0 23761 7 1 2 23758 23760
0 23762 5 1 1 23761
0 23763 7 1 2 66264 23762
0 23764 5 1 1 23763
0 23765 7 1 2 90101 86704
0 23766 7 1 2 93974 23765
0 23767 5 1 1 23766
0 23768 7 1 2 23764 23767
0 23769 5 1 1 23768
0 23770 7 1 2 73462 23769
0 23771 5 1 1 23770
0 23772 7 1 2 66265 90123
0 23773 5 1 1 23772
0 23774 7 1 2 23773 4059
0 23775 5 1 1 23774
0 23776 7 1 2 79838 23775
0 23777 5 2 1 23776
0 23778 7 2 2 86136 94532
0 23779 5 1 1 100468
0 23780 7 1 2 79987 100469
0 23781 5 1 1 23780
0 23782 7 1 2 100466 23781
0 23783 7 1 2 23771 23782
0 23784 5 1 1 23783
0 23785 7 1 2 69151 23784
0 23786 5 1 1 23785
0 23787 7 1 2 23754 23786
0 23788 5 1 1 23787
0 23789 7 1 2 85285 23788
0 23790 5 1 1 23789
0 23791 7 1 2 23734 23790
0 23792 5 1 1 23791
0 23793 7 1 2 67299 23792
0 23794 5 1 1 23793
0 23795 7 5 2 69817 77711
0 23796 7 1 2 99184 100470
0 23797 7 2 2 66997 74352
0 23798 7 1 2 100475 76825
0 23799 7 1 2 23796 23798
0 23800 5 1 1 23799
0 23801 7 1 2 23794 23800
0 23802 5 1 1 23801
0 23803 7 1 2 97873 23802
0 23804 5 1 1 23803
0 23805 7 2 2 83323 79249
0 23806 5 1 1 100477
0 23807 7 1 2 100478 98991
0 23808 7 1 2 100461 23807
0 23809 5 1 1 23808
0 23810 7 4 2 69510 80116
0 23811 7 1 2 99027 94835
0 23812 7 1 2 100479 23811
0 23813 7 1 2 79962 23812
0 23814 5 1 1 23813
0 23815 7 1 2 23809 23814
0 23816 5 1 1 23815
0 23817 7 1 2 68381 23816
0 23818 5 1 1 23817
0 23819 7 1 2 66731 99860
0 23820 5 1 1 23819
0 23821 7 1 2 80605 83388
0 23822 5 1 1 23821
0 23823 7 1 2 23820 23822
0 23824 5 1 1 23823
0 23825 7 1 2 73463 23824
0 23826 5 1 1 23825
0 23827 7 1 2 80606 77559
0 23828 5 1 1 23827
0 23829 7 1 2 23826 23828
0 23830 5 1 1 23829
0 23831 7 1 2 74653 23830
0 23832 5 1 1 23831
0 23833 7 1 2 74877 90132
0 23834 5 1 1 23833
0 23835 7 1 2 85605 23834
0 23836 5 1 1 23835
0 23837 7 1 2 70433 23836
0 23838 5 1 1 23837
0 23839 7 1 2 66732 87549
0 23840 5 1 1 23839
0 23841 7 1 2 23838 23840
0 23842 5 1 1 23841
0 23843 7 1 2 76219 23842
0 23844 5 1 1 23843
0 23845 7 2 2 65079 80142
0 23846 5 1 1 100483
0 23847 7 1 2 76585 83476
0 23848 7 1 2 100484 23847
0 23849 5 1 1 23848
0 23850 7 1 2 23844 23849
0 23851 7 1 2 23832 23850
0 23852 5 1 1 23851
0 23853 7 2 2 98421 77151
0 23854 7 1 2 23852 100485
0 23855 5 1 1 23854
0 23856 7 1 2 23818 23855
0 23857 5 1 1 23856
0 23858 7 1 2 69152 23857
0 23859 5 1 1 23858
0 23860 7 1 2 80812 99172
0 23861 5 1 1 23860
0 23862 7 3 2 82595 97953
0 23863 7 1 2 75913 100487
0 23864 5 1 1 23863
0 23865 7 1 2 23861 23864
0 23866 5 1 1 23865
0 23867 7 1 2 69818 23866
0 23868 5 1 1 23867
0 23869 7 1 2 99622 6758
0 23870 5 1 1 23869
0 23871 7 1 2 75276 23870
0 23872 5 1 1 23871
0 23873 7 1 2 95061 86920
0 23874 5 1 1 23873
0 23875 7 1 2 81198 23874
0 23876 7 1 2 23872 23875
0 23877 5 1 1 23876
0 23878 7 1 2 64697 23877
0 23879 5 1 1 23878
0 23880 7 1 2 65080 86921
0 23881 5 1 1 23880
0 23882 7 1 2 66530 80354
0 23883 5 2 1 23882
0 23884 7 1 2 93980 100490
0 23885 5 1 1 23884
0 23886 7 1 2 73464 23885
0 23887 5 1 1 23886
0 23888 7 1 2 23881 23887
0 23889 5 1 1 23888
0 23890 7 1 2 75914 23889
0 23891 5 1 1 23890
0 23892 7 1 2 23891 100467
0 23893 7 1 2 23879 23892
0 23894 5 1 1 23893
0 23895 7 1 2 67300 23894
0 23896 5 1 1 23895
0 23897 7 1 2 23868 23896
0 23898 5 1 1 23897
0 23899 7 4 2 95368 93557
0 23900 7 1 2 23898 100492
0 23901 5 1 1 23900
0 23902 7 1 2 23859 23901
0 23903 5 1 1 23902
0 23904 7 1 2 85286 23903
0 23905 5 1 1 23904
0 23906 7 10 2 98340 77988
0 23907 5 3 1 100496
0 23908 7 2 2 100126 100506
0 23909 5 14 1 100509
0 23910 7 8 2 67301 100511
0 23911 7 1 2 90473 100336
0 23912 5 1 1 23911
0 23913 7 2 2 82110 83472
0 23914 7 1 2 95133 100533
0 23915 5 1 1 23914
0 23916 7 2 2 23912 23915
0 23917 5 1 1 100535
0 23918 7 1 2 82918 83775
0 23919 7 1 2 99861 23918
0 23920 5 1 1 23919
0 23921 7 1 2 100536 23920
0 23922 5 1 1 23921
0 23923 7 1 2 100525 23922
0 23924 5 1 1 23923
0 23925 7 2 2 76746 99028
0 23926 7 1 2 99691 95369
0 23927 7 1 2 100537 23926
0 23928 7 1 2 100337 23927
0 23929 5 1 1 23928
0 23930 7 1 2 23924 23929
0 23931 5 1 1 23930
0 23932 7 1 2 85912 23931
0 23933 5 1 1 23932
0 23934 7 1 2 99862 93958
0 23935 5 1 1 23934
0 23936 7 6 2 73731 86540
0 23937 5 1 1 100539
0 23938 7 1 2 66531 100540
0 23939 7 1 2 81570 23938
0 23940 5 1 1 23939
0 23941 7 1 2 23935 23940
0 23942 5 1 1 23941
0 23943 7 1 2 73465 23942
0 23944 5 1 1 23943
0 23945 7 1 2 92912 81152
0 23946 5 1 1 23945
0 23947 7 1 2 93864 79191
0 23948 5 1 1 23947
0 23949 7 1 2 23946 23948
0 23950 7 1 2 23944 23949
0 23951 5 1 1 23950
0 23952 7 1 2 100390 95375
0 23953 7 1 2 23951 23952
0 23954 5 1 1 23953
0 23955 7 1 2 23933 23954
0 23956 5 1 1 23955
0 23957 7 1 2 65399 23956
0 23958 5 1 1 23957
0 23959 7 1 2 96957 97339
0 23960 5 1 1 23959
0 23961 7 3 2 69153 66532
0 23962 5 2 1 100545
0 23963 7 2 2 71818 98372
0 23964 7 1 2 100546 100550
0 23965 5 1 1 23964
0 23966 7 1 2 23960 23965
0 23967 5 1 1 23966
0 23968 7 2 2 75915 92869
0 23969 7 1 2 83966 95370
0 23970 7 1 2 100552 23969
0 23971 7 1 2 23967 23970
0 23972 5 1 1 23971
0 23973 7 1 2 71644 79472
0 23974 7 1 2 83600 23973
0 23975 7 2 2 74853 79276
0 23976 7 1 2 99591 100554
0 23977 7 1 2 23974 23976
0 23978 5 1 1 23977
0 23979 7 1 2 23972 23978
0 23980 5 1 1 23979
0 23981 7 1 2 70176 23980
0 23982 5 1 1 23981
0 23983 7 2 2 74782 98807
0 23984 7 3 2 64698 80117
0 23985 7 1 2 69511 85448
0 23986 7 2 2 100558 23985
0 23987 7 1 2 99152 100561
0 23988 7 1 2 100556 23987
0 23989 5 1 1 23988
0 23990 7 1 2 23982 23989
0 23991 5 1 1 23990
0 23992 7 1 2 85913 23991
0 23993 5 1 1 23992
0 23994 7 3 2 66998 79594
0 23995 5 1 1 100563
0 23996 7 1 2 66266 87020
0 23997 7 1 2 82048 23996
0 23998 5 1 1 23997
0 23999 7 1 2 79436 23998
0 24000 5 1 1 23999
0 24001 7 1 2 100564 24000
0 24002 5 1 1 24001
0 24003 7 1 2 99856 24002
0 24004 5 1 1 24003
0 24005 7 1 2 23995 94020
0 24006 5 1 1 24005
0 24007 7 1 2 73466 24006
0 24008 7 1 2 24004 24007
0 24009 5 1 1 24008
0 24010 7 1 2 93721 79196
0 24011 7 1 2 95409 24010
0 24012 5 1 1 24011
0 24013 7 1 2 24009 24012
0 24014 5 1 1 24013
0 24015 7 1 2 100526 24014
0 24016 5 1 1 24015
0 24017 7 3 2 70434 87997
0 24018 7 2 2 72374 87605
0 24019 7 1 2 93600 100569
0 24020 7 1 2 100566 24019
0 24021 7 1 2 100338 24020
0 24022 5 1 1 24021
0 24023 7 1 2 24016 24022
0 24024 5 1 1 24023
0 24025 7 1 2 80407 24024
0 24026 5 1 1 24025
0 24027 7 1 2 23993 24026
0 24028 7 1 2 23958 24027
0 24029 7 1 2 23905 24028
0 24030 7 1 2 23804 24029
0 24031 5 1 1 24030
0 24032 7 1 2 67167 24031
0 24033 5 1 1 24032
0 24034 7 2 2 95635 99091
0 24035 7 1 2 63795 100159
0 24036 7 1 2 100571 24035
0 24037 5 1 1 24036
0 24038 7 1 2 24033 24037
0 24039 5 1 1 24038
0 24040 7 1 2 100261 24039
0 24041 5 1 1 24040
0 24042 7 1 2 23718 24041
0 24043 7 1 2 23663 24042
0 24044 7 1 2 23447 24043
0 24045 5 1 1 24044
0 24046 7 1 2 67632 24045
0 24047 5 1 1 24046
0 24048 7 12 2 67168 72664
0 24049 7 1 2 88392 79544
0 24050 5 1 1 24049
0 24051 7 2 2 65081 86699
0 24052 5 1 1 100585
0 24053 7 1 2 71819 100586
0 24054 5 1 1 24053
0 24055 7 1 2 24050 24054
0 24056 5 1 1 24055
0 24057 7 1 2 100294 24056
0 24058 5 1 1 24057
0 24059 7 2 2 82008 99925
0 24060 5 1 1 100587
0 24061 7 2 2 65400 88472
0 24062 5 2 1 100589
0 24063 7 3 2 80499 100591
0 24064 5 3 1 100593
0 24065 7 5 2 65082 100596
0 24066 5 1 1 100599
0 24067 7 1 2 69819 100600
0 24068 5 1 1 24067
0 24069 7 1 2 24060 24068
0 24070 5 1 1 24069
0 24071 7 1 2 71364 24070
0 24072 5 1 1 24071
0 24073 7 2 2 69820 79558
0 24074 7 1 2 99926 100604
0 24075 5 1 1 24074
0 24076 7 1 2 24072 24075
0 24077 5 1 1 24076
0 24078 7 1 2 100262 24077
0 24079 5 1 1 24078
0 24080 7 2 2 64699 86685
0 24081 5 2 1 100606
0 24082 7 1 2 66267 100607
0 24083 5 1 1 24082
0 24084 7 1 2 100172 24083
0 24085 5 1 1 24084
0 24086 7 1 2 24079 24085
0 24087 5 1 1 24086
0 24088 7 1 2 85914 24087
0 24089 5 1 1 24088
0 24090 7 1 2 24058 24089
0 24091 5 1 1 24090
0 24092 7 1 2 73467 24091
0 24093 5 1 1 24092
0 24094 7 1 2 99698 97469
0 24095 5 1 1 24094
0 24096 7 1 2 97386 93819
0 24097 5 1 1 24096
0 24098 7 1 2 80295 84090
0 24099 5 1 1 24098
0 24100 7 1 2 24097 24099
0 24101 5 1 1 24100
0 24102 7 1 2 85915 24101
0 24103 5 1 1 24102
0 24104 7 2 2 85287 93809
0 24105 5 1 1 100610
0 24106 7 1 2 66268 100611
0 24107 5 1 1 24106
0 24108 7 1 2 24103 24107
0 24109 5 1 1 24108
0 24110 7 1 2 71645 24109
0 24111 5 1 1 24110
0 24112 7 2 2 85288 88393
0 24113 7 1 2 100612 78802
0 24114 5 1 1 24113
0 24115 7 1 2 72054 93829
0 24116 5 1 1 24115
0 24117 7 3 2 90709 24116
0 24118 7 2 2 97387 100614
0 24119 5 1 1 100617
0 24120 7 1 2 94421 100618
0 24121 5 1 1 24120
0 24122 7 1 2 24114 24121
0 24123 7 1 2 24111 24122
0 24124 5 1 1 24123
0 24125 7 1 2 68382 24124
0 24126 5 1 1 24125
0 24127 7 1 2 24095 24126
0 24128 5 1 1 24127
0 24129 7 1 2 100263 24128
0 24130 5 1 1 24129
0 24131 7 2 2 63796 79017
0 24132 5 2 1 100619
0 24133 7 1 2 12867 100621
0 24134 5 1 1 24133
0 24135 7 1 2 80868 95122
0 24136 5 1 1 24135
0 24137 7 1 2 24134 24136
0 24138 5 1 1 24137
0 24139 7 1 2 20464 24138
0 24140 5 1 1 24139
0 24141 7 1 2 100173 24140
0 24142 5 1 1 24141
0 24143 7 1 2 24130 24142
0 24144 7 1 2 24093 24143
0 24145 5 1 1 24144
0 24146 7 1 2 65794 24145
0 24147 5 1 1 24146
0 24148 7 1 2 100373 79602
0 24149 7 1 2 74929 24148
0 24150 7 1 2 89942 24149
0 24151 5 1 1 24150
0 24152 7 1 2 24147 24151
0 24153 5 1 1 24152
0 24154 7 1 2 68035 24153
0 24155 5 1 1 24154
0 24156 7 2 2 93210 88026
0 24157 7 1 2 89383 91878
0 24158 7 1 2 100623 24157
0 24159 5 1 1 24158
0 24160 7 2 2 89939 95816
0 24161 7 1 2 86568 84609
0 24162 7 1 2 100625 24161
0 24163 5 1 1 24162
0 24164 7 1 2 24159 24163
0 24165 5 1 1 24164
0 24166 7 1 2 65083 24165
0 24167 5 1 1 24166
0 24168 7 5 2 95718 82774
0 24169 7 1 2 19809 12847
0 24170 5 1 1 24169
0 24171 7 1 2 93810 24170
0 24172 5 1 1 24171
0 24173 7 3 2 71646 85916
0 24174 7 8 2 65401 84704
0 24175 5 4 1 100635
0 24176 7 1 2 99736 100643
0 24177 5 1 1 24176
0 24178 7 1 2 100632 24177
0 24179 5 1 1 24178
0 24180 7 1 2 94574 24179
0 24181 7 1 2 24172 24180
0 24182 5 1 1 24181
0 24183 7 1 2 100627 24182
0 24184 5 1 1 24183
0 24185 7 1 2 24167 24184
0 24186 5 1 1 24185
0 24187 7 1 2 68383 24186
0 24188 5 1 1 24187
0 24189 7 2 2 93211 100264
0 24190 7 1 2 71820 83041
0 24191 5 1 1 24190
0 24192 7 1 2 2928 24191
0 24193 5 1 1 24192
0 24194 7 1 2 80851 24193
0 24195 5 1 1 24194
0 24196 7 1 2 70435 93033
0 24197 5 1 1 24196
0 24198 7 1 2 65402 14035
0 24199 5 1 1 24198
0 24200 7 1 2 71647 89060
0 24201 7 1 2 24199 24200
0 24202 7 1 2 24197 24201
0 24203 5 1 1 24202
0 24204 7 1 2 24195 24203
0 24205 5 1 1 24204
0 24206 7 1 2 85917 24205
0 24207 5 1 1 24206
0 24208 7 1 2 24207 98784
0 24209 5 1 1 24208
0 24210 7 1 2 100647 24209
0 24211 5 1 1 24210
0 24212 7 1 2 24188 24211
0 24213 5 1 1 24212
0 24214 7 1 2 69821 24213
0 24215 5 1 1 24214
0 24216 7 1 2 93811 100648
0 24217 5 1 1 24216
0 24218 7 5 2 75667 93493
0 24219 5 1 1 100649
0 24220 7 1 2 88706 75516
0 24221 7 1 2 81602 24220
0 24222 7 1 2 100650 24221
0 24223 5 1 1 24222
0 24224 7 1 2 24217 24223
0 24225 5 1 1 24224
0 24226 7 1 2 71648 24225
0 24227 5 1 1 24226
0 24228 7 2 2 1807 99731
0 24229 5 1 1 100654
0 24230 7 1 2 73732 24229
0 24231 5 1 1 24230
0 24232 7 1 2 66733 81565
0 24233 5 1 1 24232
0 24234 7 1 2 24231 24233
0 24235 5 1 1 24234
0 24236 7 1 2 89630 92435
0 24237 7 1 2 24235 24236
0 24238 5 1 1 24237
0 24239 7 1 2 24227 24238
0 24240 5 1 1 24239
0 24241 7 1 2 85289 24240
0 24242 5 1 1 24241
0 24243 7 3 2 66870 75386
0 24244 7 1 2 68646 91307
0 24245 7 1 2 100656 24244
0 24246 5 1 1 24245
0 24247 7 1 2 100237 87910
0 24248 7 1 2 95551 24247
0 24249 5 1 1 24248
0 24250 7 1 2 24246 24249
0 24251 5 1 1 24250
0 24252 7 1 2 82414 91871
0 24253 7 1 2 24251 24252
0 24254 5 1 1 24253
0 24255 7 1 2 24242 24254
0 24256 5 1 1 24255
0 24257 7 1 2 68384 24256
0 24258 5 1 1 24257
0 24259 7 5 2 90587 84610
0 24260 7 2 2 66999 82111
0 24261 7 1 2 86327 96799
0 24262 7 1 2 100664 24261
0 24263 7 1 2 100659 24262
0 24264 5 1 1 24263
0 24265 7 1 2 24258 24264
0 24266 7 1 2 24215 24265
0 24267 5 1 1 24266
0 24268 7 1 2 73103 24267
0 24269 5 1 1 24268
0 24270 7 1 2 76316 77310
0 24271 5 1 1 24270
0 24272 7 1 2 76586 24271
0 24273 7 1 2 88845 24272
0 24274 5 1 1 24273
0 24275 7 1 2 100174 24274
0 24276 5 1 1 24275
0 24277 7 2 2 94585 75591
0 24278 7 1 2 68988 100666
0 24279 7 1 2 94541 24278
0 24280 5 1 1 24279
0 24281 7 1 2 24276 24280
0 24282 5 1 1 24281
0 24283 7 1 2 85290 24282
0 24284 5 1 1 24283
0 24285 7 6 2 93583 91959
0 24286 7 2 2 74537 87359
0 24287 5 2 1 100674
0 24288 7 1 2 76317 95112
0 24289 5 1 1 24288
0 24290 7 1 2 100676 24289
0 24291 5 1 1 24290
0 24292 7 1 2 68647 24291
0 24293 5 1 1 24292
0 24294 7 4 2 69822 75076
0 24295 5 1 1 100678
0 24296 7 1 2 81722 84214
0 24297 5 1 1 24296
0 24298 7 1 2 24295 24297
0 24299 7 1 2 24293 24298
0 24300 5 1 1 24299
0 24301 7 1 2 100668 24300
0 24302 5 1 1 24301
0 24303 7 1 2 24284 24302
0 24304 5 1 1 24303
0 24305 7 1 2 65795 24304
0 24306 5 1 1 24305
0 24307 7 1 2 24269 24306
0 24308 7 1 2 24155 24307
0 24309 5 1 1 24308
0 24310 7 1 2 69512 24309
0 24311 5 1 1 24310
0 24312 7 1 2 100320 87070
0 24313 5 1 1 24312
0 24314 7 1 2 73468 99878
0 24315 5 1 1 24314
0 24316 7 3 2 75387 99954
0 24317 5 1 1 100682
0 24318 7 1 2 68385 24317
0 24319 5 1 1 24318
0 24320 7 1 2 80607 24319
0 24321 7 1 2 24315 24320
0 24322 5 1 1 24321
0 24323 7 1 2 24313 24322
0 24324 5 1 1 24323
0 24325 7 1 2 85918 24324
0 24326 5 1 1 24325
0 24327 7 1 2 74952 82294
0 24328 5 1 1 24327
0 24329 7 2 2 68386 94264
0 24330 5 2 1 100685
0 24331 7 1 2 69823 77646
0 24332 7 1 2 100686 24331
0 24333 5 1 1 24332
0 24334 7 1 2 24328 24333
0 24335 5 1 1 24334
0 24336 7 1 2 85291 24335
0 24337 5 1 1 24336
0 24338 7 1 2 24326 24337
0 24339 5 1 1 24338
0 24340 7 1 2 68648 24339
0 24341 5 2 1 24340
0 24342 7 1 2 82371 80308
0 24343 5 1 1 24342
0 24344 7 1 2 85292 24343
0 24345 5 1 1 24344
0 24346 7 2 2 85919 88867
0 24347 5 1 1 100691
0 24348 7 1 2 68036 100692
0 24349 5 1 1 24348
0 24350 7 1 2 24345 24349
0 24351 5 1 1 24350
0 24352 7 2 2 71649 24351
0 24353 5 1 1 100693
0 24354 7 1 2 95700 86991
0 24355 5 1 1 24354
0 24356 7 1 2 24353 24355
0 24357 5 1 1 24356
0 24358 7 1 2 76476 24357
0 24359 5 1 1 24358
0 24360 7 1 2 100689 24359
0 24361 5 1 1 24360
0 24362 7 2 2 66871 24361
0 24363 7 1 2 100406 100695
0 24364 5 1 1 24363
0 24365 7 1 2 24311 24364
0 24366 5 1 1 24365
0 24367 7 1 2 71064 24366
0 24368 5 1 1 24367
0 24369 7 1 2 66269 94712
0 24370 5 1 1 24369
0 24371 7 1 2 65084 77432
0 24372 7 1 2 95222 24371
0 24373 5 1 1 24372
0 24374 7 1 2 24370 24373
0 24375 5 1 1 24374
0 24376 7 1 2 64700 24375
0 24377 5 1 1 24376
0 24378 7 1 2 94508 94127
0 24379 5 1 1 24378
0 24380 7 1 2 81723 87211
0 24381 5 1 1 24380
0 24382 7 1 2 24052 24381
0 24383 5 1 1 24382
0 24384 7 1 2 77217 24383
0 24385 5 1 1 24384
0 24386 7 1 2 24379 24385
0 24387 7 1 2 24377 24386
0 24388 5 1 1 24387
0 24389 7 1 2 73733 24388
0 24390 5 1 1 24389
0 24391 7 1 2 82519 77337
0 24392 5 1 1 24391
0 24393 7 1 2 78645 24392
0 24394 5 1 1 24393
0 24395 7 1 2 80699 89447
0 24396 5 1 1 24395
0 24397 7 1 2 24394 24396
0 24398 5 1 1 24397
0 24399 7 1 2 76220 24398
0 24400 5 1 1 24399
0 24401 7 1 2 24390 24400
0 24402 5 1 1 24401
0 24403 7 1 2 73104 24402
0 24404 5 1 1 24403
0 24405 7 1 2 86745 92163
0 24406 5 1 1 24405
0 24407 7 1 2 71365 88862
0 24408 5 1 1 24407
0 24409 7 1 2 73105 9901
0 24410 7 1 2 24408 24409
0 24411 5 1 1 24410
0 24412 7 1 2 68037 14038
0 24413 7 1 2 95142 24412
0 24414 5 1 1 24413
0 24415 7 1 2 24411 24414
0 24416 5 1 1 24415
0 24417 7 1 2 24406 24416
0 24418 5 1 1 24417
0 24419 7 1 2 77218 24418
0 24420 5 1 1 24419
0 24421 7 1 2 77219 77008
0 24422 7 1 2 86790 24421
0 24423 5 1 1 24422
0 24424 7 1 2 76686 86216
0 24425 7 1 2 81596 24424
0 24426 5 1 1 24425
0 24427 7 1 2 24423 24426
0 24428 5 1 1 24427
0 24429 7 1 2 97388 24428
0 24430 5 1 1 24429
0 24431 7 2 2 83919 94895
0 24432 5 1 1 100697
0 24433 7 1 2 77338 24432
0 24434 5 1 1 24433
0 24435 7 1 2 77339 83144
0 24436 5 1 1 24435
0 24437 7 1 2 76221 24436
0 24438 7 1 2 94748 24437
0 24439 5 1 1 24438
0 24440 7 1 2 24434 24439
0 24441 7 1 2 24430 24440
0 24442 7 1 2 24420 24441
0 24443 7 1 2 24404 24442
0 24444 5 1 1 24443
0 24445 7 1 2 85293 24444
0 24446 5 1 1 24445
0 24447 7 1 2 75077 95361
0 24448 5 1 1 24447
0 24449 7 1 2 66533 86992
0 24450 5 1 1 24449
0 24451 7 1 2 24448 24450
0 24452 5 1 1 24451
0 24453 7 1 2 65085 24452
0 24454 5 1 1 24453
0 24455 7 1 2 98369 12849
0 24456 7 1 2 86925 24455
0 24457 5 1 1 24456
0 24458 7 1 2 66270 24457
0 24459 5 1 1 24458
0 24460 7 1 2 88366 91588
0 24461 5 1 1 24460
0 24462 7 1 2 24459 24461
0 24463 7 1 2 24454 24462
0 24464 5 1 1 24463
0 24465 7 1 2 64701 24464
0 24466 5 1 1 24465
0 24467 7 1 2 86998 79215
0 24468 5 1 1 24467
0 24469 7 1 2 69513 89819
0 24470 5 1 1 24469
0 24471 7 1 2 24468 24470
0 24472 5 1 1 24471
0 24473 7 5 2 73469 92924
0 24474 7 2 2 74654 88367
0 24475 5 1 1 100704
0 24476 7 1 2 82284 24475
0 24477 5 1 1 24476
0 24478 7 1 2 100699 24477
0 24479 5 1 1 24478
0 24480 7 1 2 81866 75088
0 24481 5 1 1 24480
0 24482 7 1 2 78834 24481
0 24483 5 1 1 24482
0 24484 7 1 2 24479 24483
0 24485 7 1 2 24472 24484
0 24486 7 1 2 24466 24485
0 24487 5 1 1 24486
0 24488 7 1 2 68038 24487
0 24489 5 1 1 24488
0 24490 7 2 2 9438 83095
0 24491 5 1 1 100706
0 24492 7 1 2 71366 100707
0 24493 5 1 1 24492
0 24494 7 1 2 66271 81318
0 24495 5 3 1 24494
0 24496 7 1 2 68649 100708
0 24497 7 1 2 24493 24496
0 24498 5 1 1 24497
0 24499 7 1 2 97358 73907
0 24500 5 2 1 24499
0 24501 7 1 2 71367 95046
0 24502 5 1 1 24501
0 24503 7 1 2 84198 24502
0 24504 5 1 1 24503
0 24505 7 1 2 100711 24504
0 24506 7 1 2 24498 24505
0 24507 5 1 1 24506
0 24508 7 1 2 66734 24507
0 24509 5 1 1 24508
0 24510 7 2 2 74655 83410
0 24511 7 1 2 75078 100713
0 24512 5 1 1 24511
0 24513 7 1 2 24509 24512
0 24514 5 1 1 24513
0 24515 7 1 2 65403 24514
0 24516 5 1 1 24515
0 24517 7 1 2 93865 100679
0 24518 5 1 1 24517
0 24519 7 1 2 97389 95113
0 24520 5 1 1 24519
0 24521 7 1 2 99821 94932
0 24522 5 1 1 24521
0 24523 7 1 2 24520 24522
0 24524 5 1 1 24523
0 24525 7 1 2 68650 24524
0 24526 5 1 1 24525
0 24527 7 1 2 24518 24526
0 24528 7 1 2 24516 24527
0 24529 5 1 1 24528
0 24530 7 1 2 73106 24529
0 24531 5 1 1 24530
0 24532 7 1 2 79277 86109
0 24533 5 2 1 24532
0 24534 7 1 2 24531 100715
0 24535 7 1 2 24489 24534
0 24536 5 1 1 24535
0 24537 7 1 2 65995 24536
0 24538 5 1 1 24537
0 24539 7 1 2 87203 86981
0 24540 5 1 1 24539
0 24541 7 1 2 97390 98935
0 24542 5 1 1 24541
0 24543 7 1 2 24540 24542
0 24544 5 1 1 24543
0 24545 7 1 2 68039 24544
0 24546 5 1 1 24545
0 24547 7 2 2 85687 97826
0 24548 5 1 1 100717
0 24549 7 1 2 83283 100718
0 24550 5 1 1 24549
0 24551 7 1 2 24546 24550
0 24552 5 1 1 24551
0 24553 7 1 2 73734 24552
0 24554 5 1 1 24553
0 24555 7 2 2 76477 77870
0 24556 5 1 1 100719
0 24557 7 1 2 85737 100720
0 24558 5 1 1 24557
0 24559 7 1 2 99955 88848
0 24560 5 1 1 24559
0 24561 7 1 2 99942 90014
0 24562 5 1 1 24561
0 24563 7 1 2 24560 24562
0 24564 5 1 1 24563
0 24565 7 1 2 65086 24564
0 24566 5 1 1 24565
0 24567 7 1 2 24558 24566
0 24568 7 1 2 24554 24567
0 24569 5 1 1 24568
0 24570 7 1 2 64392 24569
0 24571 5 1 1 24570
0 24572 7 1 2 75388 24548
0 24573 5 1 1 24572
0 24574 7 1 2 73735 24573
0 24575 5 1 1 24574
0 24576 7 1 2 65087 88849
0 24577 5 1 1 24576
0 24578 7 1 2 24575 24577
0 24579 5 1 1 24578
0 24580 7 1 2 75605 76871
0 24581 7 1 2 24579 24580
0 24582 5 1 1 24581
0 24583 7 1 2 24571 24582
0 24584 7 1 2 24538 24583
0 24585 5 1 1 24584
0 24586 7 1 2 85920 24585
0 24587 5 1 1 24586
0 24588 7 1 2 24446 24587
0 24589 5 1 1 24588
0 24590 7 1 2 70804 24589
0 24591 5 1 1 24590
0 24592 7 1 2 99718 94311
0 24593 7 1 2 100555 98682
0 24594 7 1 2 24592 24593
0 24595 5 2 1 24594
0 24596 7 1 2 76478 100694
0 24597 5 1 1 24596
0 24598 7 1 2 100690 24597
0 24599 5 2 1 24598
0 24600 7 1 2 100723 93056
0 24601 5 1 1 24600
0 24602 7 1 2 100721 24601
0 24603 7 1 2 24591 24602
0 24604 5 1 1 24603
0 24605 7 1 2 100175 24604
0 24606 5 1 1 24605
0 24607 7 1 2 24368 24606
0 24608 5 1 1 24607
0 24609 7 1 2 67302 24608
0 24610 5 1 1 24609
0 24611 7 1 2 80608 99173
0 24612 5 1 1 24611
0 24613 7 3 2 81724 78954
0 24614 7 1 2 76999 98172
0 24615 7 1 2 100725 24614
0 24616 5 1 1 24615
0 24617 7 1 2 24612 24616
0 24618 5 1 1 24617
0 24619 7 1 2 66534 24618
0 24620 5 1 1 24619
0 24621 7 1 2 80609 76117
0 24622 5 1 1 24621
0 24623 7 1 2 71368 95887
0 24624 5 1 1 24623
0 24625 7 1 2 24622 24624
0 24626 5 1 1 24625
0 24627 7 1 2 75389 24626
0 24628 5 1 1 24627
0 24629 7 1 2 74953 94949
0 24630 5 1 1 24629
0 24631 7 1 2 24628 24630
0 24632 5 1 1 24631
0 24633 7 1 2 72375 24632
0 24634 5 1 1 24633
0 24635 7 1 2 24620 24634
0 24636 5 1 1 24635
0 24637 7 1 2 64702 24636
0 24638 5 1 1 24637
0 24639 7 1 2 77101 83448
0 24640 5 1 1 24639
0 24641 7 1 2 80700 79241
0 24642 5 1 1 24641
0 24643 7 1 2 85581 24642
0 24644 7 1 2 24640 24643
0 24645 5 1 1 24644
0 24646 7 1 2 65088 24645
0 24647 5 1 1 24646
0 24648 7 1 2 79216 88477
0 24649 5 1 1 24648
0 24650 7 1 2 100590 24649
0 24651 5 1 1 24650
0 24652 7 4 2 69824 82596
0 24653 5 1 1 100728
0 24654 7 1 2 66535 100729
0 24655 5 1 1 24654
0 24656 7 1 2 68040 24655
0 24657 7 1 2 24651 24656
0 24658 7 1 2 24647 24657
0 24659 5 1 1 24658
0 24660 7 3 2 88772 96450
0 24661 5 7 1 100732
0 24662 7 1 2 82295 100735
0 24663 5 1 1 24662
0 24664 7 1 2 69825 77123
0 24665 5 1 1 24664
0 24666 7 1 2 80800 24665
0 24667 5 1 1 24666
0 24668 7 1 2 80610 24667
0 24669 5 2 1 24668
0 24670 7 1 2 73107 100742
0 24671 7 1 2 24663 24670
0 24672 5 1 1 24671
0 24673 7 1 2 71369 24672
0 24674 7 1 2 24659 24673
0 24675 5 1 1 24674
0 24676 7 2 2 84080 80894
0 24677 5 2 1 100744
0 24678 7 1 2 74783 100745
0 24679 5 2 1 24678
0 24680 7 1 2 68387 100733
0 24681 5 1 1 24680
0 24682 7 1 2 73470 100006
0 24683 5 1 1 24682
0 24684 7 1 2 24683 78763
0 24685 7 1 2 24681 24684
0 24686 5 1 1 24685
0 24687 7 1 2 100748 24686
0 24688 5 1 1 24687
0 24689 7 1 2 71650 24688
0 24690 5 1 1 24689
0 24691 7 1 2 68041 96451
0 24692 7 1 2 97814 24691
0 24693 5 1 1 24692
0 24694 7 1 2 92925 87021
0 24695 7 1 2 96681 24694
0 24696 7 1 2 24693 24695
0 24697 5 1 1 24696
0 24698 7 1 2 24690 24697
0 24699 7 1 2 24675 24698
0 24700 5 1 1 24699
0 24701 7 1 2 72376 24700
0 24702 5 1 1 24701
0 24703 7 1 2 24638 24702
0 24704 5 1 1 24703
0 24705 7 1 2 77152 24704
0 24706 5 1 1 24705
0 24707 7 1 2 70177 79947
0 24708 5 1 1 24707
0 24709 7 1 2 80160 24708
0 24710 5 1 1 24709
0 24711 7 1 2 73471 24710
0 24712 5 1 1 24711
0 24713 7 1 2 24712 95903
0 24714 5 1 1 24713
0 24715 7 1 2 88394 24714
0 24716 5 1 1 24715
0 24717 7 1 2 93812 83638
0 24718 5 1 1 24717
0 24719 7 6 2 69826 80701
0 24720 5 3 1 100750
0 24721 7 3 2 73472 75972
0 24722 7 1 2 100751 100759
0 24723 7 1 2 83810 24722
0 24724 5 1 1 24723
0 24725 7 1 2 24718 24724
0 24726 5 1 1 24725
0 24727 7 1 2 71651 24726
0 24728 5 1 1 24727
0 24729 7 1 2 81645 93826
0 24730 5 1 1 24729
0 24731 7 1 2 99956 85627
0 24732 5 1 1 24731
0 24733 7 1 2 24730 24732
0 24734 7 1 2 24728 24733
0 24735 7 1 2 24716 24734
0 24736 5 1 1 24735
0 24737 7 1 2 98267 24736
0 24738 5 1 1 24737
0 24739 7 1 2 24706 24738
0 24740 5 1 1 24739
0 24741 7 1 2 85294 24740
0 24742 5 1 1 24741
0 24743 7 1 2 83127 96660
0 24744 5 1 1 24743
0 24745 7 5 2 71065 68651
0 24746 7 3 2 98609 100762
0 24747 5 1 1 100767
0 24748 7 1 2 98227 24747
0 24749 5 4 1 24748
0 24750 7 1 2 24744 100770
0 24751 5 1 1 24750
0 24752 7 2 2 68652 98173
0 24753 7 1 2 97989 100774
0 24754 5 1 1 24753
0 24755 7 1 2 100480 98196
0 24756 5 1 1 24755
0 24757 7 1 2 24754 24756
0 24758 5 1 1 24757
0 24759 7 1 2 84828 24758
0 24760 5 1 1 24759
0 24761 7 3 2 69514 74902
0 24762 7 2 2 72377 73736
0 24763 7 3 2 71066 100779
0 24764 7 1 2 100776 100781
0 24765 5 1 1 24764
0 24766 7 2 2 81603 98219
0 24767 5 1 1 100784
0 24768 7 1 2 24765 24767
0 24769 5 1 1 24768
0 24770 7 1 2 66735 24769
0 24771 5 1 1 24770
0 24772 7 1 2 100567 100782
0 24773 5 1 1 24772
0 24774 7 1 2 24771 24773
0 24775 5 1 1 24774
0 24776 7 1 2 71652 24775
0 24777 5 1 1 24776
0 24778 7 5 2 64393 99522
0 24779 7 1 2 86347 87124
0 24780 7 1 2 100786 24779
0 24781 5 1 1 24780
0 24782 7 1 2 24777 24781
0 24783 5 1 1 24782
0 24784 7 1 2 68388 24783
0 24785 5 1 1 24784
0 24786 7 1 2 24760 24785
0 24787 5 1 1 24786
0 24788 7 1 2 68042 24787
0 24789 5 1 1 24788
0 24790 7 1 2 24751 24789
0 24791 5 1 1 24790
0 24792 7 1 2 97391 24791
0 24793 5 1 1 24792
0 24794 7 1 2 84626 79298
0 24795 5 1 1 24794
0 24796 7 3 2 73908 82009
0 24797 7 1 2 99822 100791
0 24798 5 1 1 24797
0 24799 7 1 2 24795 24798
0 24800 5 1 1 24799
0 24801 7 1 2 100771 24800
0 24802 5 1 1 24801
0 24803 7 1 2 86137 98247
0 24804 5 1 1 24803
0 24805 7 1 2 82919 98268
0 24806 5 1 1 24805
0 24807 7 1 2 24804 24806
0 24808 5 1 1 24807
0 24809 7 1 2 65404 24808
0 24810 5 1 1 24809
0 24811 7 1 2 23368 98228
0 24812 5 1 1 24811
0 24813 7 1 2 80491 24812
0 24814 5 1 1 24813
0 24815 7 1 2 24810 24814
0 24816 5 1 1 24815
0 24817 7 1 2 65089 24816
0 24818 5 1 1 24817
0 24819 7 1 2 98472 94222
0 24820 5 1 1 24819
0 24821 7 1 2 24818 24820
0 24822 5 1 1 24821
0 24823 7 1 2 100680 24822
0 24824 5 1 1 24823
0 24825 7 1 2 24802 24824
0 24826 5 1 1 24825
0 24827 7 1 2 68043 24826
0 24828 5 1 1 24827
0 24829 7 1 2 83546 80552
0 24830 5 1 1 24829
0 24831 7 1 2 68389 93813
0 24832 5 2 1 24831
0 24833 7 1 2 66536 95363
0 24834 7 1 2 100794 24833
0 24835 5 1 1 24834
0 24836 7 1 2 73473 94212
0 24837 5 1 1 24836
0 24838 7 1 2 65090 93883
0 24839 5 1 1 24838
0 24840 7 1 2 71653 12218
0 24841 7 1 2 24839 24840
0 24842 7 1 2 24837 24841
0 24843 5 1 1 24842
0 24844 7 1 2 24835 24843
0 24845 5 1 1 24844
0 24846 7 1 2 24830 24845
0 24847 5 1 1 24846
0 24848 7 1 2 98269 24847
0 24849 5 1 1 24848
0 24850 7 3 2 71654 77153
0 24851 7 1 2 98186 100796
0 24852 7 1 2 88671 24851
0 24853 5 1 1 24852
0 24854 7 5 2 82112 86138
0 24855 7 1 2 98473 77520
0 24856 7 1 2 100799 24855
0 24857 5 1 1 24856
0 24858 7 1 2 24853 24857
0 24859 7 1 2 24849 24858
0 24860 5 1 1 24859
0 24861 7 1 2 83284 24860
0 24862 5 1 1 24861
0 24863 7 1 2 24828 24862
0 24864 7 1 2 24793 24863
0 24865 5 1 1 24864
0 24866 7 1 2 85921 24865
0 24867 5 1 1 24866
0 24868 7 1 2 24742 24867
0 24869 5 1 1 24868
0 24870 7 1 2 100265 24869
0 24871 5 1 1 24870
0 24872 7 11 2 63901 65642
0 24873 5 1 1 100804
0 24874 7 2 2 100805 97218
0 24875 7 1 2 71067 88676
0 24876 5 1 1 24875
0 24877 7 1 2 99918 24876
0 24878 5 1 1 24877
0 24879 7 1 2 69515 24878
0 24880 5 1 1 24879
0 24881 7 2 2 70436 77712
0 24882 7 1 2 95690 100817
0 24883 5 1 1 24882
0 24884 7 1 2 77220 24883
0 24885 5 1 1 24884
0 24886 7 1 2 69827 24885
0 24887 5 1 1 24886
0 24888 7 1 2 16722 24887
0 24889 7 1 2 24880 24888
0 24890 5 1 1 24889
0 24891 7 1 2 70178 24890
0 24892 5 1 1 24891
0 24893 7 1 2 82520 90972
0 24894 5 1 1 24893
0 24895 7 1 2 100316 24894
0 24896 5 1 1 24895
0 24897 7 1 2 77221 74889
0 24898 5 1 1 24897
0 24899 7 1 2 74954 24898
0 24900 5 1 1 24899
0 24901 7 1 2 24896 24900
0 24902 5 1 1 24901
0 24903 7 1 2 77433 24902
0 24904 5 1 1 24903
0 24905 7 3 2 68653 77154
0 24906 5 1 1 100819
0 24907 7 3 2 78018 86172
0 24908 5 1 1 100822
0 24909 7 1 2 77222 24908
0 24910 5 1 1 24909
0 24911 7 1 2 70179 77434
0 24912 7 1 2 24910 24911
0 24913 5 1 1 24912
0 24914 7 1 2 24906 24913
0 24915 5 1 1 24914
0 24916 7 1 2 95466 24915
0 24917 5 1 1 24916
0 24918 7 2 2 66272 77000
0 24919 5 1 1 100825
0 24920 7 1 2 82260 24919
0 24921 5 1 1 24920
0 24922 7 1 2 24917 24921
0 24923 7 1 2 24904 24922
0 24924 7 1 2 24892 24923
0 24925 5 1 1 24924
0 24926 7 1 2 85295 24925
0 24927 5 1 1 24926
0 24928 7 1 2 75789 87115
0 24929 5 1 1 24928
0 24930 7 1 2 70180 24929
0 24931 5 1 1 24930
0 24932 7 3 2 68390 84705
0 24933 5 1 1 100827
0 24934 7 1 2 24931 24933
0 24935 5 1 1 24934
0 24936 7 1 2 71655 24935
0 24937 5 1 1 24936
0 24938 7 2 2 68654 100828
0 24939 5 1 1 100830
0 24940 7 1 2 24937 24939
0 24941 5 1 1 24940
0 24942 7 1 2 65405 24941
0 24943 5 1 1 24942
0 24944 7 1 2 82920 81611
0 24945 5 1 1 24944
0 24946 7 1 2 24943 24945
0 24947 5 1 1 24946
0 24948 7 1 2 69828 24947
0 24949 5 1 1 24948
0 24950 7 1 2 100831 86168
0 24951 5 1 1 24950
0 24952 7 1 2 24949 24951
0 24953 5 1 1 24952
0 24954 7 1 2 82578 24953
0 24955 5 1 1 24954
0 24956 7 1 2 77569 93280
0 24957 5 1 1 24956
0 24958 7 1 2 76318 82579
0 24959 7 1 2 79940 24958
0 24960 7 1 2 95435 24959
0 24961 5 1 1 24960
0 24962 7 1 2 24957 24961
0 24963 5 1 1 24962
0 24964 7 1 2 75390 24963
0 24965 5 1 1 24964
0 24966 7 1 2 69829 91626
0 24967 5 2 1 24966
0 24968 7 1 2 71068 81283
0 24969 5 1 1 24968
0 24970 7 1 2 100832 24969
0 24971 5 1 1 24970
0 24972 7 1 2 69516 24971
0 24973 5 1 1 24972
0 24974 7 2 2 76936 91430
0 24975 5 1 1 100834
0 24976 7 1 2 24973 24975
0 24977 5 1 1 24976
0 24978 7 1 2 74784 24977
0 24979 5 1 1 24978
0 24980 7 1 2 24965 24979
0 24981 5 1 1 24980
0 24982 7 1 2 80611 24981
0 24983 5 1 1 24982
0 24984 7 1 2 68391 87148
0 24985 5 1 1 24984
0 24986 7 1 2 77621 24985
0 24987 5 1 1 24986
0 24988 7 1 2 81725 24987
0 24989 5 1 1 24988
0 24990 7 1 2 83145 75698
0 24991 5 1 1 24990
0 24992 7 1 2 71656 24991
0 24993 5 1 1 24992
0 24994 7 1 2 84200 24993
0 24995 5 1 1 24994
0 24996 7 1 2 88368 24995
0 24997 5 1 1 24996
0 24998 7 1 2 24997 92022
0 24999 7 1 2 24989 24998
0 25000 5 1 1 24999
0 25001 7 1 2 77155 25000
0 25002 5 1 1 25001
0 25003 7 1 2 24983 25002
0 25004 7 1 2 24955 25003
0 25005 5 1 1 25004
0 25006 7 1 2 85922 25005
0 25007 5 1 1 25006
0 25008 7 1 2 24927 25007
0 25009 5 1 1 25008
0 25010 7 1 2 100815 25009
0 25011 5 1 1 25010
0 25012 7 1 2 24871 25011
0 25013 5 1 1 25012
0 25014 7 1 2 70805 25013
0 25015 5 1 1 25014
0 25016 7 1 2 24610 25015
0 25017 5 1 1 25016
0 25018 7 1 2 69154 25017
0 25019 5 1 1 25018
0 25020 7 2 2 70181 99927
0 25021 5 1 1 100836
0 25022 7 5 2 73474 100837
0 25023 5 4 1 100838
0 25024 7 1 2 93839 100843
0 25025 5 3 1 25024
0 25026 7 1 2 85923 100847
0 25027 5 1 1 25026
0 25028 7 1 2 98825 25027
0 25029 5 2 1 25028
0 25030 7 1 2 64703 100850
0 25031 5 1 1 25030
0 25032 7 1 2 73475 93827
0 25033 5 1 1 25032
0 25034 7 1 2 94425 25033
0 25035 5 1 1 25034
0 25036 7 1 2 85296 25035
0 25037 5 1 1 25036
0 25038 7 1 2 25031 25037
0 25039 5 1 1 25038
0 25040 7 1 2 68044 25039
0 25041 5 1 1 25040
0 25042 7 2 2 70437 91866
0 25043 7 1 2 94397 100852
0 25044 5 1 1 25043
0 25045 7 1 2 24105 25044
0 25046 5 2 1 25045
0 25047 7 1 2 81360 100854
0 25048 5 1 1 25047
0 25049 7 1 2 25041 25048
0 25050 5 1 1 25049
0 25051 7 1 2 71370 25050
0 25052 5 1 1 25051
0 25053 7 3 2 75576 80078
0 25054 5 3 1 100856
0 25055 7 1 2 100855 100857
0 25056 5 1 1 25055
0 25057 7 1 2 25052 25056
0 25058 5 1 1 25057
0 25059 7 1 2 100266 25058
0 25060 5 1 1 25059
0 25061 7 1 2 75973 95114
0 25062 5 1 1 25061
0 25063 7 1 2 100677 25062
0 25064 5 1 1 25063
0 25065 7 1 2 68655 25064
0 25066 5 1 1 25065
0 25067 7 1 2 81726 100317
0 25068 5 1 1 25067
0 25069 7 1 2 81652 25068
0 25070 7 1 2 25066 25069
0 25071 5 1 1 25070
0 25072 7 1 2 85924 25071
0 25073 5 1 1 25072
0 25074 7 1 2 88846 100698
0 25075 5 1 1 25074
0 25076 7 1 2 85297 25075
0 25077 5 1 1 25076
0 25078 7 1 2 95547 86519
0 25079 5 1 1 25078
0 25080 7 1 2 25079 94575
0 25081 5 1 1 25080
0 25082 7 1 2 75391 25081
0 25083 5 1 1 25082
0 25084 7 1 2 25077 25083
0 25085 7 1 2 25073 25084
0 25086 5 1 1 25085
0 25087 7 1 2 100176 25086
0 25088 5 1 1 25087
0 25089 7 1 2 66273 100851
0 25090 5 1 1 25089
0 25091 7 1 2 100601 93464
0 25092 5 1 1 25091
0 25093 7 1 2 100613 89820
0 25094 5 1 1 25093
0 25095 7 1 2 25092 25094
0 25096 5 1 1 25095
0 25097 7 1 2 73476 25096
0 25098 5 1 1 25097
0 25099 7 1 2 25090 25098
0 25100 5 1 1 25099
0 25101 7 1 2 68045 25100
0 25102 5 1 1 25101
0 25103 7 1 2 94573 94539
0 25104 5 1 1 25103
0 25105 7 1 2 25102 25104
0 25106 5 1 1 25105
0 25107 7 1 2 100267 25106
0 25108 5 1 1 25107
0 25109 7 1 2 68852 85652
0 25110 5 1 1 25109
0 25111 7 1 2 75974 90710
0 25112 7 1 2 25110 25111
0 25113 5 1 1 25112
0 25114 7 1 2 68656 98789
0 25115 5 1 1 25114
0 25116 7 1 2 25113 25115
0 25117 7 1 2 70182 99979
0 25118 5 1 1 25117
0 25119 7 1 2 85362 24347
0 25120 5 1 1 25119
0 25121 7 1 2 71657 25120
0 25122 5 1 1 25121
0 25123 7 1 2 25118 25122
0 25124 7 1 2 25116 25123
0 25125 5 1 1 25124
0 25126 7 1 2 100177 25125
0 25127 5 1 1 25126
0 25128 7 1 2 91782 96647
0 25129 5 2 1 25128
0 25130 7 1 2 73477 90463
0 25131 5 1 1 25130
0 25132 7 1 2 88795 25131
0 25133 5 1 1 25132
0 25134 7 1 2 71658 25133
0 25135 5 1 1 25134
0 25136 7 1 2 83516 25135
0 25137 5 1 1 25136
0 25138 7 1 2 65406 25137
0 25139 5 2 1 25138
0 25140 7 1 2 96810 12592
0 25141 5 1 1 25140
0 25142 7 1 2 70438 25141
0 25143 5 1 1 25142
0 25144 7 1 2 96807 25143
0 25145 7 1 2 100864 25144
0 25146 5 1 1 25145
0 25147 7 1 2 71371 25146
0 25148 5 1 1 25147
0 25149 7 1 2 100862 25148
0 25150 5 1 1 25149
0 25151 7 1 2 73108 99339
0 25152 7 1 2 25150 25151
0 25153 5 1 1 25152
0 25154 7 1 2 25127 25153
0 25155 7 1 2 25108 25154
0 25156 5 1 1 25155
0 25157 7 1 2 69830 25156
0 25158 5 1 1 25157
0 25159 7 1 2 25088 25158
0 25160 7 1 2 25060 25159
0 25161 5 1 1 25160
0 25162 7 1 2 64094 25161
0 25163 5 1 1 25162
0 25164 7 2 2 70183 100242
0 25165 7 1 2 73478 92309
0 25166 7 1 2 100866 25165
0 25167 7 1 2 100240 25166
0 25168 5 1 1 25167
0 25169 7 1 2 94064 92064
0 25170 7 1 2 78169 25169
0 25171 7 1 2 100626 25170
0 25172 5 1 1 25171
0 25173 7 1 2 25168 25172
0 25174 5 1 1 25173
0 25175 7 1 2 73737 25174
0 25176 5 1 1 25175
0 25177 7 1 2 80612 77630
0 25178 5 1 1 25177
0 25179 7 1 2 1869 25178
0 25180 5 1 1 25179
0 25181 7 4 2 84320 96408
0 25182 7 1 2 25180 100868
0 25183 5 1 1 25182
0 25184 7 2 2 91308 90658
0 25185 5 1 1 100872
0 25186 7 1 2 78955 100873
0 25187 7 1 2 89789 25186
0 25188 5 1 1 25187
0 25189 7 1 2 25183 25188
0 25190 5 1 1 25189
0 25191 7 1 2 85298 25190
0 25192 5 1 1 25191
0 25193 7 1 2 25176 25192
0 25194 5 1 1 25193
0 25195 7 1 2 78740 25194
0 25196 5 1 1 25195
0 25197 7 1 2 100328 94251
0 25198 5 1 1 25197
0 25199 7 1 2 80542 76074
0 25200 5 1 1 25199
0 25201 7 1 2 79066 76158
0 25202 5 1 1 25201
0 25203 7 1 2 25200 25202
0 25204 5 1 1 25203
0 25205 7 1 2 73479 25204
0 25206 5 1 1 25205
0 25207 7 1 2 100636 85823
0 25208 5 1 1 25207
0 25209 7 1 2 25206 25208
0 25210 5 1 1 25209
0 25211 7 1 2 66537 25210
0 25212 5 1 1 25211
0 25213 7 1 2 25198 25212
0 25214 5 1 1 25213
0 25215 7 1 2 65091 25214
0 25216 5 1 1 25215
0 25217 7 2 2 74785 84131
0 25218 5 1 1 100874
0 25219 7 1 2 65407 97790
0 25220 5 1 1 25219
0 25221 7 1 2 25218 25220
0 25222 5 1 1 25221
0 25223 7 1 2 66736 25222
0 25224 5 1 1 25223
0 25225 7 1 2 85765 83130
0 25226 5 1 1 25225
0 25227 7 1 2 25224 25226
0 25228 5 1 1 25227
0 25229 7 1 2 79559 25228
0 25230 5 1 1 25229
0 25231 7 1 2 25216 25230
0 25232 5 1 1 25231
0 25233 7 5 2 64704 65643
0 25234 7 2 2 75194 78865
0 25235 7 1 2 100876 100881
0 25236 7 1 2 25232 25235
0 25237 5 1 1 25236
0 25238 7 1 2 25196 25237
0 25239 7 1 2 25163 25238
0 25240 5 1 1 25239
0 25241 7 1 2 69517 25240
0 25242 5 1 1 25241
0 25243 7 1 2 64095 93584
0 25244 7 1 2 100696 25243
0 25245 5 1 1 25244
0 25246 7 1 2 25242 25245
0 25247 5 1 1 25246
0 25248 7 1 2 71069 25247
0 25249 5 1 1 25248
0 25250 7 1 2 78124 100724
0 25251 5 1 1 25250
0 25252 7 1 2 25251 100722
0 25253 5 1 1 25252
0 25254 7 1 2 100178 25253
0 25255 5 1 1 25254
0 25256 7 1 2 25249 25255
0 25257 5 1 1 25256
0 25258 7 1 2 99444 25257
0 25259 5 1 1 25258
0 25260 7 1 2 75790 92168
0 25261 5 1 1 25260
0 25262 7 1 2 64705 25261
0 25263 5 1 1 25262
0 25264 7 1 2 76319 91297
0 25265 5 2 1 25264
0 25266 7 1 2 79293 100883
0 25267 7 1 2 25263 25266
0 25268 5 1 1 25267
0 25269 7 1 2 68392 25268
0 25270 5 1 1 25269
0 25271 7 2 2 66274 74878
0 25272 5 2 1 100885
0 25273 7 1 2 81131 100886
0 25274 5 1 1 25273
0 25275 7 1 2 25270 25274
0 25276 5 1 1 25275
0 25277 7 1 2 65996 25276
0 25278 5 1 1 25277
0 25279 7 3 2 73738 97392
0 25280 5 1 1 100889
0 25281 7 1 2 66275 91947
0 25282 5 1 1 25281
0 25283 7 1 2 25280 25282
0 25284 7 1 2 100884 25283
0 25285 5 1 1 25284
0 25286 7 1 2 82790 25285
0 25287 5 1 1 25286
0 25288 7 1 2 25278 25287
0 25289 5 1 1 25288
0 25290 7 1 2 85925 25289
0 25291 5 1 1 25290
0 25292 7 2 2 85299 82296
0 25293 5 1 1 100892
0 25294 7 1 2 100893 78043
0 25295 5 1 1 25294
0 25296 7 1 2 25291 25295
0 25297 5 1 1 25296
0 25298 7 1 2 73109 25297
0 25299 5 1 1 25298
0 25300 7 2 2 85300 75975
0 25301 5 1 1 100894
0 25302 7 1 2 92223 86852
0 25303 5 1 1 25302
0 25304 7 1 2 25301 25303
0 25305 5 1 1 25304
0 25306 7 1 2 77340 25305
0 25307 5 1 1 25306
0 25308 7 1 2 25299 25307
0 25309 5 1 1 25308
0 25310 7 1 2 82432 25309
0 25311 5 1 1 25310
0 25312 7 1 2 81501 80255
0 25313 5 1 1 25312
0 25314 7 2 2 68393 91627
0 25315 7 1 2 64706 100896
0 25316 5 1 1 25315
0 25317 7 1 2 25313 25316
0 25318 5 1 1 25317
0 25319 7 1 2 68046 25318
0 25320 5 1 1 25319
0 25321 7 1 2 76320 81502
0 25322 5 1 1 25321
0 25323 7 1 2 68394 95844
0 25324 5 1 1 25323
0 25325 7 1 2 25322 25324
0 25326 5 1 1 25325
0 25327 7 1 2 71070 25326
0 25328 5 1 1 25327
0 25329 7 1 2 25320 25328
0 25330 5 1 1 25329
0 25331 7 1 2 85926 25330
0 25332 5 1 1 25331
0 25333 7 1 2 73909 79617
0 25334 5 1 1 25333
0 25335 7 1 2 77578 25334
0 25336 5 1 1 25335
0 25337 7 1 2 85301 25336
0 25338 5 1 1 25337
0 25339 7 1 2 25332 25338
0 25340 5 1 1 25339
0 25341 7 1 2 69518 25340
0 25342 5 1 1 25341
0 25343 7 1 2 64707 83565
0 25344 5 2 1 25343
0 25345 7 1 2 83651 83556
0 25346 5 1 1 25345
0 25347 7 2 2 100898 25346
0 25348 7 1 2 85927 100900
0 25349 5 1 1 25348
0 25350 7 1 2 25293 25349
0 25351 5 1 1 25350
0 25352 7 1 2 71372 25351
0 25353 5 1 1 25352
0 25354 7 1 2 85302 82265
0 25355 5 1 1 25354
0 25356 7 1 2 25353 25355
0 25357 5 1 1 25356
0 25358 7 1 2 98939 25357
0 25359 5 1 1 25358
0 25360 7 1 2 25342 25359
0 25361 5 1 1 25360
0 25362 7 1 2 85500 25361
0 25363 5 1 1 25362
0 25364 7 1 2 77223 94419
0 25365 5 1 1 25364
0 25366 7 1 2 85928 97628
0 25367 5 1 1 25366
0 25368 7 1 2 25365 25367
0 25369 5 1 1 25368
0 25370 7 1 2 64708 25369
0 25371 5 1 1 25370
0 25372 7 1 2 91808 79106
0 25373 5 1 1 25372
0 25374 7 1 2 25371 25373
0 25375 5 1 1 25374
0 25376 7 1 2 82433 25375
0 25377 5 1 1 25376
0 25378 7 1 2 77224 86849
0 25379 5 1 1 25378
0 25380 7 4 2 77435 25379
0 25381 7 7 2 68395 85501
0 25382 7 1 2 85929 100906
0 25383 7 1 2 100902 25382
0 25384 5 1 1 25383
0 25385 7 1 2 25377 25384
0 25386 5 1 1 25385
0 25387 7 1 2 76075 25386
0 25388 5 1 1 25387
0 25389 7 1 2 25363 25388
0 25390 7 1 2 25311 25389
0 25391 5 1 1 25390
0 25392 7 1 2 100179 25391
0 25393 5 1 1 25392
0 25394 7 3 2 68047 100042
0 25395 5 2 1 100913
0 25396 7 2 2 73110 82297
0 25397 5 1 1 100918
0 25398 7 1 2 100916 25397
0 25399 5 1 1 25398
0 25400 7 1 2 71373 25399
0 25401 5 1 1 25400
0 25402 7 1 2 77609 82298
0 25403 7 1 2 78764 25402
0 25404 5 1 1 25403
0 25405 7 1 2 25401 25404
0 25406 5 1 1 25405
0 25407 7 1 2 85303 25406
0 25408 5 1 1 25407
0 25409 7 1 2 74538 99863
0 25410 5 1 1 25409
0 25411 7 1 2 24556 25410
0 25412 5 1 1 25411
0 25413 7 1 2 92224 25412
0 25414 5 1 1 25413
0 25415 7 1 2 25408 25414
0 25416 5 1 1 25415
0 25417 7 1 2 68657 100268
0 25418 7 1 2 100512 25417
0 25419 7 1 2 25416 25418
0 25420 5 1 1 25419
0 25421 7 1 2 25393 25420
0 25422 5 1 1 25421
0 25423 7 1 2 67303 25422
0 25424 5 1 1 25423
0 25425 7 1 2 71374 79729
0 25426 5 2 1 25425
0 25427 7 1 2 76039 100920
0 25428 5 2 1 25427
0 25429 7 1 2 69519 100922
0 25430 5 1 1 25429
0 25431 7 2 2 74656 80161
0 25432 5 1 1 100924
0 25433 7 2 2 69831 76023
0 25434 5 2 1 100926
0 25435 7 1 2 74539 100928
0 25436 7 1 2 6944 25435
0 25437 5 1 1 25436
0 25438 7 1 2 25432 25437
0 25439 5 1 1 25438
0 25440 7 1 2 25430 25439
0 25441 5 1 1 25440
0 25442 7 1 2 71071 25441
0 25443 5 1 1 25442
0 25444 7 4 2 69520 81132
0 25445 7 1 2 99223 100930
0 25446 5 1 1 25445
0 25447 7 2 2 69832 79730
0 25448 5 1 1 100934
0 25449 7 1 2 79423 25448
0 25450 5 1 1 25449
0 25451 7 1 2 25450 91630
0 25452 5 1 1 25451
0 25453 7 1 2 25446 25452
0 25454 7 1 2 25443 25453
0 25455 5 1 1 25454
0 25456 7 1 2 68396 25455
0 25457 5 1 1 25456
0 25458 7 1 2 69521 77580
0 25459 5 1 1 25458
0 25460 7 2 2 71072 80150
0 25461 5 1 1 100936
0 25462 7 1 2 25459 25461
0 25463 5 2 1 25462
0 25464 7 1 2 83015 100938
0 25465 5 1 1 25464
0 25466 7 1 2 25457 25465
0 25467 5 1 1 25466
0 25468 7 1 2 85930 25467
0 25469 5 1 1 25468
0 25470 7 1 2 77610 80278
0 25471 5 1 1 25470
0 25472 7 1 2 89280 77225
0 25473 5 1 1 25472
0 25474 7 1 2 25473 10508
0 25475 5 1 1 25474
0 25476 7 1 2 25471 25475
0 25477 5 1 1 25476
0 25478 7 1 2 85304 25477
0 25479 5 1 1 25478
0 25480 7 1 2 25469 25479
0 25481 5 1 1 25480
0 25482 7 1 2 99751 100180
0 25483 7 1 2 25481 25482
0 25484 5 1 1 25483
0 25485 7 1 2 25424 25484
0 25486 5 1 1 25485
0 25487 7 1 2 81867 25486
0 25488 5 1 1 25487
0 25489 7 3 2 66737 94852
0 25490 7 3 2 68853 79025
0 25491 7 1 2 100940 100943
0 25492 5 1 1 25491
0 25493 7 1 2 98785 25492
0 25494 5 1 1 25493
0 25495 7 1 2 100103 100393
0 25496 5 1 1 25495
0 25497 7 1 2 69155 100269
0 25498 7 1 2 97874 25497
0 25499 5 1 1 25498
0 25500 7 1 2 25496 25499
0 25501 5 1 1 25500
0 25502 7 1 2 25494 25501
0 25503 5 1 1 25502
0 25504 7 3 2 66738 76391
0 25505 7 2 2 77226 100946
0 25506 7 5 2 90588 87746
0 25507 5 1 1 100951
0 25508 7 1 2 82434 95999
0 25509 7 1 2 100952 25508
0 25510 7 1 2 100949 25509
0 25511 5 1 1 25510
0 25512 7 1 2 25503 25511
0 25513 5 1 1 25512
0 25514 7 1 2 71375 25513
0 25515 5 1 1 25514
0 25516 7 2 2 90716 93102
0 25517 7 4 2 65644 70806
0 25518 7 4 2 65598 100958
0 25519 7 1 2 84977 100962
0 25520 7 1 2 100956 25519
0 25521 7 1 2 100950 25520
0 25522 5 1 1 25521
0 25523 7 1 2 25515 25522
0 25524 5 1 1 25523
0 25525 7 1 2 68048 25524
0 25526 5 1 1 25525
0 25527 7 1 2 68854 89153
0 25528 7 1 2 93112 25527
0 25529 7 3 2 100877 76134
0 25530 7 1 2 100376 100966
0 25531 7 1 2 25528 25530
0 25532 5 1 1 25531
0 25533 7 1 2 25526 25532
0 25534 5 1 1 25533
0 25535 7 1 2 67304 25534
0 25536 5 1 1 25535
0 25537 7 1 2 69156 94565
0 25538 7 1 2 94669 25537
0 25539 7 3 2 70807 97101
0 25540 7 2 2 76159 86096
0 25541 7 1 2 100972 97644
0 25542 7 1 2 100969 25541
0 25543 7 1 2 25538 25542
0 25544 5 1 1 25543
0 25545 7 1 2 25536 25544
0 25546 5 1 1 25545
0 25547 7 1 2 66538 25546
0 25548 5 1 1 25547
0 25549 7 3 2 94586 94778
0 25550 7 2 2 68989 100974
0 25551 7 1 2 85305 98422
0 25552 7 1 2 86700 97555
0 25553 7 1 2 25551 25552
0 25554 7 1 2 82407 25553
0 25555 7 1 2 100977 25554
0 25556 5 1 1 25555
0 25557 7 1 2 25548 25556
0 25558 5 1 1 25557
0 25559 7 1 2 80098 25558
0 25560 5 1 1 25559
0 25561 7 3 2 65599 100402
0 25562 7 1 2 80296 99712
0 25563 7 1 2 100979 25562
0 25564 5 1 1 25563
0 25565 7 1 2 99944 100109
0 25566 7 1 2 98907 25565
0 25567 5 1 1 25566
0 25568 7 1 2 25564 25567
0 25569 5 1 1 25568
0 25570 7 1 2 77156 92207
0 25571 7 1 2 95759 25570
0 25572 7 1 2 25569 25571
0 25573 5 1 1 25572
0 25574 7 1 2 25560 25573
0 25575 7 1 2 25488 25574
0 25576 7 1 2 25259 25575
0 25577 7 1 2 25019 25576
0 25578 5 1 1 25577
0 25579 7 1 2 100573 25578
0 25580 5 1 1 25579
0 25581 7 3 2 67305 81868
0 25582 7 4 2 88379 100982
0 25583 7 1 2 70184 97875
0 25584 7 1 2 100985 25583
0 25585 5 1 1 25584
0 25586 7 1 2 84829 80852
0 25587 5 1 1 25586
0 25588 7 1 2 100756 25587
0 25589 5 1 1 25588
0 25590 7 1 2 100486 25589
0 25591 5 1 1 25590
0 25592 7 1 2 25585 25591
0 25593 5 1 1 25592
0 25594 7 1 2 76076 25593
0 25595 5 1 1 25594
0 25596 7 2 2 73111 81133
0 25597 5 1 1 100989
0 25598 7 4 2 72378 84830
0 25599 7 3 2 69522 100991
0 25600 7 1 2 95334 100995
0 25601 5 1 1 25600
0 25602 7 4 2 67306 97876
0 25603 7 1 2 81869 100998
0 25604 5 1 1 25603
0 25605 7 1 2 25601 25604
0 25606 5 1 1 25605
0 25607 7 1 2 68658 25606
0 25608 5 1 1 25607
0 25609 7 1 2 80613 100999
0 25610 5 1 1 25609
0 25611 7 1 2 25608 25610
0 25612 5 1 1 25611
0 25613 7 1 2 100990 25612
0 25614 5 1 1 25613
0 25615 7 1 2 25595 25614
0 25616 5 1 1 25615
0 25617 7 1 2 69157 25616
0 25618 5 1 1 25617
0 25619 7 10 2 71073 78125
0 25620 5 1 1 101002
0 25621 7 1 2 99133 101003
0 25622 7 1 2 100986 25621
0 25623 7 1 2 83261 25622
0 25624 5 1 1 25623
0 25625 7 1 2 25618 25624
0 25626 5 1 1 25625
0 25627 7 1 2 72665 25626
0 25628 5 1 1 25627
0 25629 7 1 2 100106 740
0 25630 5 18 1 25629
0 25631 7 1 2 98487 101012
0 25632 5 1 1 25631
0 25633 7 1 2 85449 98270
0 25634 5 1 1 25633
0 25635 7 1 2 77157 98650
0 25636 5 2 1 25635
0 25637 7 1 2 25634 101030
0 25638 7 1 2 25632 25637
0 25639 5 3 1 25638
0 25640 7 1 2 81134 85092
0 25641 7 1 2 86047 25640
0 25642 7 1 2 101032 25641
0 25643 5 1 1 25642
0 25644 7 1 2 25628 25643
0 25645 5 1 1 25644
0 25646 7 1 2 100295 25645
0 25647 5 1 1 25646
0 25648 7 1 2 98814 96088
0 25649 5 1 1 25648
0 25650 7 1 2 69523 25649
0 25651 5 1 1 25650
0 25652 7 5 2 67633 77158
0 25653 5 1 1 101035
0 25654 7 1 2 98863 25653
0 25655 5 1 1 25654
0 25656 7 1 2 25651 25655
0 25657 5 1 1 25656
0 25658 7 1 2 69158 25657
0 25659 5 1 1 25658
0 25660 7 5 2 85450 78479
0 25661 5 1 1 101040
0 25662 7 3 2 69524 101041
0 25663 5 3 1 101045
0 25664 7 1 2 25659 101048
0 25665 5 1 1 25664
0 25666 7 1 2 82307 25665
0 25667 5 1 1 25666
0 25668 7 9 2 72666 82435
0 25669 7 1 2 93814 80060
0 25670 7 1 2 101051 25669
0 25671 5 1 1 25670
0 25672 7 1 2 25667 25671
0 25673 5 1 1 25672
0 25674 7 1 2 72379 25673
0 25675 5 1 1 25674
0 25676 7 3 2 67307 80614
0 25677 7 2 2 67634 77227
0 25678 5 1 1 101063
0 25679 7 3 2 72667 80061
0 25680 5 1 1 101065
0 25681 7 1 2 25678 25680
0 25682 5 1 1 25681
0 25683 7 1 2 85502 25682
0 25684 5 1 1 25683
0 25685 7 1 2 25684 92818
0 25686 5 1 1 25685
0 25687 7 1 2 101060 25686
0 25688 5 1 1 25687
0 25689 7 1 2 25675 25688
0 25690 5 1 1 25689
0 25691 7 1 2 68049 25690
0 25692 5 1 1 25691
0 25693 7 2 2 96917 95371
0 25694 7 1 2 78409 101068
0 25695 5 1 1 25694
0 25696 7 4 2 85503 77436
0 25697 5 1 1 101070
0 25698 7 6 2 67308 87796
0 25699 7 1 2 83065 101074
0 25700 7 1 2 101071 25699
0 25701 5 1 1 25700
0 25702 7 1 2 25695 25701
0 25703 7 1 2 25692 25702
0 25704 5 1 1 25703
0 25705 7 1 2 85306 25704
0 25706 5 1 1 25705
0 25707 7 2 2 81727 96742
0 25708 5 1 1 101080
0 25709 7 1 2 97668 101081
0 25710 5 1 1 25709
0 25711 7 3 2 72380 83903
0 25712 7 3 2 70439 95262
0 25713 7 1 2 101082 101085
0 25714 5 2 1 25713
0 25715 7 1 2 25708 101088
0 25716 5 1 1 25715
0 25717 7 1 2 65796 25716
0 25718 5 1 1 25717
0 25719 7 1 2 88395 98450
0 25720 5 1 1 25719
0 25721 7 1 2 69159 25720
0 25722 7 1 2 25718 25721
0 25723 5 1 1 25722
0 25724 7 2 2 98488 84288
0 25725 7 1 2 86672 101090
0 25726 5 1 1 25725
0 25727 7 6 2 70808 96743
0 25728 5 1 1 101092
0 25729 7 1 2 81728 101093
0 25730 5 1 1 25729
0 25731 7 1 2 64096 25730
0 25732 7 1 2 25726 25731
0 25733 5 1 1 25732
0 25734 7 1 2 70185 25733
0 25735 7 1 2 25723 25734
0 25736 5 1 1 25735
0 25737 7 1 2 25710 25736
0 25738 5 1 1 25737
0 25739 7 1 2 89085 87606
0 25740 7 1 2 25738 25739
0 25741 5 1 1 25740
0 25742 7 1 2 25706 25741
0 25743 5 1 1 25742
0 25744 7 1 2 76321 25743
0 25745 5 1 1 25744
0 25746 7 1 2 98020 76937
0 25747 5 2 1 25746
0 25748 7 5 2 67309 81729
0 25749 7 1 2 75916 101100
0 25750 5 1 1 25749
0 25751 7 1 2 101098 25750
0 25752 5 1 1 25751
0 25753 7 1 2 86369 25752
0 25754 5 1 1 25753
0 25755 7 2 2 72381 76938
0 25756 7 1 2 82521 94730
0 25757 5 2 1 25756
0 25758 7 1 2 101105 101107
0 25759 5 1 1 25758
0 25760 7 1 2 25754 25759
0 25761 5 1 1 25760
0 25762 7 1 2 69833 25761
0 25763 5 1 1 25762
0 25764 7 2 2 86370 101101
0 25765 7 1 2 90918 101109
0 25766 5 1 1 25765
0 25767 7 1 2 25763 25766
0 25768 5 1 1 25767
0 25769 7 1 2 69525 25768
0 25770 5 1 1 25769
0 25771 7 1 2 71074 99864
0 25772 5 1 1 25771
0 25773 7 1 2 25772 90360
0 25774 5 2 1 25773
0 25775 7 1 2 101110 101111
0 25776 5 1 1 25775
0 25777 7 1 2 25770 25776
0 25778 5 1 1 25777
0 25779 7 1 2 67635 25778
0 25780 5 1 1 25779
0 25781 7 1 2 93774 99019
0 25782 7 1 2 80279 25781
0 25783 5 1 1 25782
0 25784 7 1 2 25780 25783
0 25785 5 1 1 25784
0 25786 7 1 2 85931 25785
0 25787 5 1 1 25786
0 25788 7 2 2 97038 95033
0 25789 7 1 2 71075 101113
0 25790 5 1 1 25789
0 25791 7 1 2 21220 25790
0 25792 5 1 1 25791
0 25793 7 1 2 92786 25792
0 25794 5 1 1 25793
0 25795 7 1 2 71076 80267
0 25796 7 1 2 99020 25795
0 25797 5 1 1 25796
0 25798 7 1 2 25794 25797
0 25799 5 1 1 25798
0 25800 7 2 2 85307 25799
0 25801 5 1 1 101115
0 25802 7 1 2 25787 25801
0 25803 5 1 1 25802
0 25804 7 1 2 65797 25803
0 25805 5 1 1 25804
0 25806 7 3 2 78753 79424
0 25807 5 15 1 101117
0 25808 7 2 2 66276 101120
0 25809 7 3 2 72382 93657
0 25810 5 1 1 101137
0 25811 7 1 2 98393 25810
0 25812 5 12 1 25811
0 25813 7 1 2 101135 101140
0 25814 5 1 1 25813
0 25815 7 2 2 71376 72383
0 25816 7 4 2 67636 101152
0 25817 7 1 2 69834 87051
0 25818 5 2 1 25817
0 25819 7 1 2 64709 80952
0 25820 5 1 1 25819
0 25821 7 1 2 101158 25820
0 25822 5 2 1 25821
0 25823 7 1 2 101154 101160
0 25824 5 1 1 25823
0 25825 7 1 2 25814 25824
0 25826 5 1 1 25825
0 25827 7 1 2 86371 25826
0 25828 5 1 1 25827
0 25829 7 4 2 77437 98021
0 25830 5 1 1 101162
0 25831 7 1 2 80274 101163
0 25832 5 1 1 25831
0 25833 7 1 2 67310 75606
0 25834 7 1 2 79473 25833
0 25835 5 1 1 25834
0 25836 7 1 2 25832 25835
0 25837 5 1 1 25836
0 25838 7 1 2 97279 25837
0 25839 5 1 1 25838
0 25840 7 1 2 25828 25839
0 25841 5 1 1 25840
0 25842 7 1 2 94613 25841
0 25843 5 1 1 25842
0 25844 7 1 2 76479 101114
0 25845 5 1 1 25844
0 25846 7 1 2 98975 99161
0 25847 5 1 1 25846
0 25848 7 1 2 25845 25847
0 25849 5 1 1 25848
0 25850 7 1 2 77228 25849
0 25851 5 1 1 25850
0 25852 7 1 2 73112 90474
0 25853 7 1 2 95179 25852
0 25854 5 1 1 25853
0 25855 7 1 2 92880 25854
0 25856 5 1 1 25855
0 25857 7 1 2 75917 93658
0 25858 7 1 2 94187 25857
0 25859 5 1 1 25858
0 25860 7 1 2 25856 25859
0 25861 5 1 1 25860
0 25862 7 1 2 72384 25861
0 25863 5 1 1 25862
0 25864 7 1 2 25851 25863
0 25865 5 1 1 25864
0 25866 7 1 2 85308 25865
0 25867 5 1 1 25866
0 25868 7 1 2 25843 25867
0 25869 5 1 1 25868
0 25870 7 1 2 70809 25869
0 25871 5 1 1 25870
0 25872 7 1 2 69160 25871
0 25873 7 1 2 25805 25872
0 25874 5 1 1 25873
0 25875 7 6 2 73113 97393
0 25876 7 1 2 93659 101166
0 25877 5 1 1 25876
0 25878 7 1 2 77438 90811
0 25879 5 1 1 25878
0 25880 7 3 2 92763 85077
0 25881 5 2 1 101172
0 25882 7 1 2 92553 101175
0 25883 7 1 2 25879 25882
0 25884 5 1 1 25883
0 25885 7 1 2 68050 25884
0 25886 5 1 1 25885
0 25887 7 1 2 25877 25886
0 25888 5 1 1 25887
0 25889 7 1 2 101102 25888
0 25890 5 1 1 25889
0 25891 7 3 2 98022 85078
0 25892 5 3 1 101177
0 25893 7 1 2 82261 101178
0 25894 5 1 1 25893
0 25895 7 1 2 25890 25894
0 25896 5 1 1 25895
0 25897 7 1 2 70810 25896
0 25898 5 1 1 25897
0 25899 7 2 2 76956 74062
0 25900 5 1 1 101183
0 25901 7 1 2 99303 101184
0 25902 5 1 1 25901
0 25903 7 1 2 25898 25902
0 25904 5 1 1 25903
0 25905 7 1 2 86372 25904
0 25906 5 1 1 25905
0 25907 7 1 2 98489 76957
0 25908 7 1 2 93077 25907
0 25909 7 1 2 101108 25908
0 25910 5 1 1 25909
0 25911 7 1 2 25906 25910
0 25912 5 1 1 25911
0 25913 7 1 2 85932 25912
0 25914 5 1 1 25913
0 25915 7 1 2 70811 101116
0 25916 5 1 1 25915
0 25917 7 1 2 64097 25916
0 25918 7 1 2 25914 25917
0 25919 5 1 1 25918
0 25920 7 1 2 25874 25919
0 25921 5 1 1 25920
0 25922 7 1 2 25745 25921
0 25923 5 1 1 25922
0 25924 7 1 2 100181 25923
0 25925 5 1 1 25924
0 25926 7 1 2 25647 25925
0 25927 5 1 1 25926
0 25928 7 1 2 67169 25927
0 25929 5 1 1 25928
0 25930 7 2 2 88894 75147
0 25931 7 3 2 75806 79636
0 25932 7 1 2 101185 101187
0 25933 5 1 1 25932
0 25934 7 2 2 97718 84070
0 25935 7 1 2 94670 101190
0 25936 5 1 1 25935
0 25937 7 1 2 100222 25936
0 25938 5 1 1 25937
0 25939 7 1 2 92159 25938
0 25940 5 1 1 25939
0 25941 7 1 2 95701 89141
0 25942 7 1 2 88904 25941
0 25943 5 1 1 25942
0 25944 7 1 2 25940 25943
0 25945 5 1 1 25944
0 25946 7 1 2 76480 25945
0 25947 5 1 1 25946
0 25948 7 1 2 25933 25947
0 25949 5 1 1 25948
0 25950 7 1 2 88316 25949
0 25951 5 1 1 25950
0 25952 7 1 2 99440 90041
0 25953 5 1 1 25952
0 25954 7 1 2 76481 95702
0 25955 5 1 1 25954
0 25956 7 1 2 25953 25955
0 25957 5 1 1 25956
0 25958 7 1 2 80444 25957
0 25959 5 1 1 25958
0 25960 7 1 2 85309 77537
0 25961 5 1 1 25960
0 25962 7 1 2 25959 25961
0 25963 5 1 1 25962
0 25964 7 1 2 100182 25963
0 25965 5 1 1 25964
0 25966 7 1 2 91272 87865
0 25967 7 1 2 84487 25966
0 25968 7 1 2 92160 86595
0 25969 7 1 2 25967 25968
0 25970 5 1 1 25969
0 25971 7 1 2 25965 25970
0 25972 7 1 2 25951 25971
0 25973 5 1 1 25972
0 25974 7 10 2 67637 100076
0 25975 7 3 2 82436 77159
0 25976 7 1 2 101192 101202
0 25977 7 1 2 25973 25976
0 25978 5 1 1 25977
0 25979 7 1 2 25929 25978
0 25980 5 1 1 25979
0 25981 7 1 2 78694 25980
0 25982 5 1 1 25981
0 25983 7 1 2 82771 100963
0 25984 7 1 2 95613 25983
0 25985 7 1 2 71077 80297
0 25986 7 1 2 100077 25985
0 25987 7 1 2 95760 25986
0 25988 7 1 2 25984 25987
0 25989 5 1 1 25988
0 25990 7 1 2 25982 25989
0 25991 7 1 2 25580 25990
0 25992 7 1 2 24047 25991
0 25993 5 1 1 25992
0 25994 7 1 2 72153 25993
0 25995 5 1 1 25994
0 25996 7 4 2 64394 81870
0 25997 5 1 1 101205
0 25998 7 1 2 19744 25997
0 25999 5 1 1 25998
0 26000 7 1 2 73910 25999
0 26001 5 1 1 26000
0 26002 7 1 2 81871 90091
0 26003 7 1 2 100687 26002
0 26004 5 1 1 26003
0 26005 7 2 2 64395 82647
0 26006 5 2 1 101209
0 26007 7 1 2 97619 101210
0 26008 5 2 1 26007
0 26009 7 1 2 98998 101213
0 26010 7 1 2 26004 26009
0 26011 5 1 1 26010
0 26012 7 1 2 70186 26011
0 26013 5 1 1 26012
0 26014 7 1 2 26001 26013
0 26015 5 1 1 26014
0 26016 7 1 2 85310 26015
0 26017 5 1 1 26016
0 26018 7 1 2 100633 95778
0 26019 5 1 1 26018
0 26020 7 1 2 81872 92979
0 26021 7 1 2 86579 26020
0 26022 5 1 1 26021
0 26023 7 1 2 26019 26022
0 26024 5 1 1 26023
0 26025 7 1 2 91131 26024
0 26026 5 1 1 26025
0 26027 7 1 2 26017 26026
0 26028 5 1 1 26027
0 26029 7 1 2 65997 26028
0 26030 5 1 1 26029
0 26031 7 2 2 96800 86982
0 26032 5 1 1 101215
0 26033 7 2 2 81873 83547
0 26034 5 1 1 101217
0 26035 7 1 2 71659 101218
0 26036 5 1 1 26035
0 26037 7 1 2 26032 26036
0 26038 5 2 1 26037
0 26039 7 2 2 73739 101219
0 26040 7 1 2 99219 101221
0 26041 5 1 1 26040
0 26042 7 1 2 26030 26041
0 26043 5 1 1 26042
0 26044 7 1 2 71377 26043
0 26045 5 1 1 26044
0 26046 7 1 2 65092 94387
0 26047 5 1 1 26046
0 26048 7 1 2 65998 2371
0 26049 5 3 1 26048
0 26050 7 1 2 81730 92735
0 26051 7 1 2 101223 26050
0 26052 7 1 2 26047 26051
0 26053 5 1 1 26052
0 26054 7 2 2 66539 83422
0 26055 5 1 1 101226
0 26056 7 1 2 80118 101227
0 26057 5 1 1 26056
0 26058 7 1 2 26053 26057
0 26059 5 1 1 26058
0 26060 7 1 2 73480 26059
0 26061 5 1 1 26060
0 26062 7 1 2 65999 99906
0 26063 5 3 1 26062
0 26064 7 1 2 71078 91524
0 26065 5 1 1 26064
0 26066 7 1 2 70440 26065
0 26067 7 1 2 101228 26066
0 26068 5 1 1 26067
0 26069 7 1 2 26061 26068
0 26070 5 1 1 26069
0 26071 7 1 2 100368 26070
0 26072 5 1 1 26071
0 26073 7 1 2 26045 26072
0 26074 5 1 1 26073
0 26075 7 1 2 69835 26074
0 26076 5 1 1 26075
0 26077 7 1 2 80813 94312
0 26078 5 2 1 26077
0 26079 7 1 2 81731 94388
0 26080 5 1 1 26079
0 26081 7 1 2 80119 83811
0 26082 7 1 2 88850 26081
0 26083 7 1 2 26080 26082
0 26084 5 1 1 26083
0 26085 7 1 2 101231 26084
0 26086 5 1 1 26085
0 26087 7 1 2 71378 26086
0 26088 5 1 1 26087
0 26089 7 1 2 76872 101222
0 26090 5 1 1 26089
0 26091 7 3 2 73481 82841
0 26092 7 5 2 78019 84081
0 26093 5 2 1 101236
0 26094 7 2 2 6815 101241
0 26095 5 1 1 101243
0 26096 7 1 2 101233 26095
0 26097 5 1 1 26096
0 26098 7 1 2 95192 87520
0 26099 5 1 1 26098
0 26100 7 1 2 26097 26099
0 26101 5 1 1 26100
0 26102 7 1 2 77439 26101
0 26103 5 1 1 26102
0 26104 7 1 2 26090 26103
0 26105 7 1 2 26088 26104
0 26106 5 1 1 26105
0 26107 7 1 2 93399 26106
0 26108 5 1 1 26107
0 26109 7 1 2 26076 26108
0 26110 5 1 1 26109
0 26111 7 1 2 67638 26110
0 26112 5 1 1 26111
0 26113 7 3 2 73911 86541
0 26114 5 1 1 101245
0 26115 7 1 2 76412 101246
0 26116 5 1 1 26115
0 26117 7 1 2 91786 79301
0 26118 5 5 1 26117
0 26119 7 2 2 80615 101248
0 26120 7 1 2 70187 101253
0 26121 5 1 1 26120
0 26122 7 1 2 26116 26121
0 26123 5 1 1 26122
0 26124 7 1 2 69836 26123
0 26125 5 1 1 26124
0 26126 7 4 2 68397 92402
0 26127 7 1 2 99782 101255
0 26128 5 2 1 26127
0 26129 7 1 2 26125 101259
0 26130 5 1 1 26129
0 26131 7 1 2 77440 26130
0 26132 5 1 1 26131
0 26133 7 1 2 80246 2275
0 26134 7 1 2 83684 26133
0 26135 5 4 1 26134
0 26136 7 1 2 66277 101261
0 26137 5 2 1 26136
0 26138 7 1 2 78784 85738
0 26139 5 1 1 26138
0 26140 7 1 2 101265 26139
0 26141 5 1 1 26140
0 26142 7 1 2 77160 26141
0 26143 5 1 1 26142
0 26144 7 1 2 26132 26143
0 26145 5 1 1 26144
0 26146 7 1 2 68659 26145
0 26147 5 1 1 26146
0 26148 7 2 2 76482 76747
0 26149 7 1 2 101216 101267
0 26150 5 1 1 26149
0 26151 7 1 2 26147 26150
0 26152 5 1 1 26151
0 26153 7 1 2 90849 26152
0 26154 5 1 1 26153
0 26155 7 1 2 26112 26154
0 26156 5 1 1 26155
0 26157 7 1 2 64098 26156
0 26158 5 1 1 26157
0 26159 7 1 2 64396 88868
0 26160 5 1 1 26159
0 26161 7 1 2 22780 26160
0 26162 5 1 1 26161
0 26163 7 1 2 79560 26162
0 26164 5 1 1 26163
0 26165 7 1 2 77981 90155
0 26166 5 1 1 26165
0 26167 7 1 2 26164 26166
0 26168 5 1 1 26167
0 26169 7 1 2 68660 26168
0 26170 5 1 1 26169
0 26171 7 1 2 83371 99989
0 26172 5 1 1 26171
0 26173 7 1 2 26170 26172
0 26174 5 1 1 26173
0 26175 7 1 2 64710 26174
0 26176 5 1 1 26175
0 26177 7 5 2 64397 79474
0 26178 5 2 1 101269
0 26179 7 1 2 99840 100700
0 26180 5 1 1 26179
0 26181 7 1 2 101274 26180
0 26182 5 1 1 26181
0 26183 7 1 2 84906 26182
0 26184 5 1 1 26183
0 26185 7 2 2 84740 92764
0 26186 5 1 1 101276
0 26187 7 1 2 83372 84978
0 26188 7 1 2 101277 26187
0 26189 5 1 1 26188
0 26190 7 1 2 26184 26189
0 26191 7 1 2 26176 26190
0 26192 5 1 1 26191
0 26193 7 1 2 66540 26192
0 26194 5 1 1 26193
0 26195 7 2 2 80079 82168
0 26196 5 1 1 101278
0 26197 7 1 2 79484 26196
0 26198 5 1 1 26197
0 26199 7 1 2 64398 26198
0 26200 5 1 1 26199
0 26201 7 6 2 64711 74151
0 26202 7 1 2 73912 101280
0 26203 5 1 1 26202
0 26204 7 1 2 26200 26203
0 26205 5 2 1 26204
0 26206 7 1 2 84907 101286
0 26207 5 1 1 26206
0 26208 7 1 2 87521 88010
0 26209 5 1 1 26208
0 26210 7 1 2 26207 26209
0 26211 5 1 1 26210
0 26212 7 1 2 65093 26211
0 26213 5 1 1 26212
0 26214 7 1 2 26194 26213
0 26215 5 1 1 26214
0 26216 7 1 2 72668 26215
0 26217 5 1 1 26216
0 26218 7 4 2 67639 81732
0 26219 7 3 2 81107 101288
0 26220 7 1 2 89742 96070
0 26221 7 1 2 101292 26220
0 26222 5 1 1 26221
0 26223 7 1 2 26217 26222
0 26224 5 1 1 26223
0 26225 7 1 2 100476 26224
0 26226 5 1 1 26225
0 26227 7 1 2 26158 26226
0 26228 5 1 1 26227
0 26229 7 1 2 68051 26228
0 26230 5 1 1 26229
0 26231 7 1 2 77441 79873
0 26232 5 2 1 26231
0 26233 7 1 2 99802 84353
0 26234 7 1 2 101295 26233
0 26235 5 1 1 26234
0 26236 7 2 2 71079 83423
0 26237 5 2 1 101297
0 26238 7 1 2 84752 101299
0 26239 5 1 1 26238
0 26240 7 1 2 94322 26239
0 26241 5 1 1 26240
0 26242 7 1 2 71080 84766
0 26243 5 1 1 26242
0 26244 7 1 2 26241 26243
0 26245 5 1 1 26244
0 26246 7 2 2 69837 101249
0 26247 5 1 1 101301
0 26248 7 1 2 100712 26247
0 26249 5 4 1 26248
0 26250 7 1 2 64099 101303
0 26251 7 1 2 26245 26250
0 26252 5 1 1 26251
0 26253 7 1 2 26235 26252
0 26254 5 1 1 26253
0 26255 7 1 2 65094 26254
0 26256 5 1 1 26255
0 26257 7 2 2 82597 80326
0 26258 7 1 2 66278 101307
0 26259 5 3 1 26258
0 26260 7 2 2 95124 77943
0 26261 7 1 2 77442 101312
0 26262 5 1 1 26261
0 26263 7 2 2 92765 84204
0 26264 5 1 1 101314
0 26265 7 1 2 26262 26264
0 26266 5 1 1 26265
0 26267 7 1 2 96648 26266
0 26268 5 1 1 26267
0 26269 7 1 2 101309 26268
0 26270 5 1 1 26269
0 26271 7 1 2 64100 68661
0 26272 7 1 2 26270 26271
0 26273 5 1 1 26272
0 26274 7 1 2 26256 26273
0 26275 5 1 1 26274
0 26276 7 1 2 73114 26275
0 26277 5 1 1 26276
0 26278 7 1 2 86448 12099
0 26279 5 1 1 26278
0 26280 7 1 2 86293 26279
0 26281 5 1 1 26280
0 26282 7 1 2 66541 92113
0 26283 7 1 2 98308 26282
0 26284 5 1 1 26283
0 26285 7 1 2 89199 26284
0 26286 5 1 1 26285
0 26287 7 1 2 65095 26286
0 26288 5 1 1 26287
0 26289 7 1 2 26281 26288
0 26290 5 1 1 26289
0 26291 7 6 2 66000 74190
0 26292 7 1 2 26290 101316
0 26293 5 1 1 26292
0 26294 7 1 2 26277 26293
0 26295 5 1 1 26294
0 26296 7 1 2 67640 26295
0 26297 5 1 1 26296
0 26298 7 3 2 76873 80020
0 26299 5 1 1 101322
0 26300 7 1 2 92821 101323
0 26301 7 1 2 88744 26300
0 26302 5 1 1 26301
0 26303 7 1 2 26297 26302
0 26304 5 1 1 26303
0 26305 7 1 2 85311 26304
0 26306 5 1 1 26305
0 26307 7 1 2 100446 100844
0 26308 5 1 1 26307
0 26309 7 2 2 73115 26308
0 26310 5 1 1 101325
0 26311 7 1 2 90475 92248
0 26312 5 1 1 26311
0 26313 7 1 2 26310 26312
0 26314 5 1 1 26313
0 26315 7 1 2 85933 26314
0 26316 5 1 1 26315
0 26317 7 1 2 73913 83137
0 26318 5 3 1 26317
0 26319 7 1 2 77689 94731
0 26320 7 2 2 101327 26319
0 26321 5 1 1 101330
0 26322 7 1 2 82748 26321
0 26323 5 1 1 26322
0 26324 7 1 2 85312 26323
0 26325 5 2 1 26324
0 26326 7 1 2 26316 101332
0 26327 5 1 1 26326
0 26328 7 1 2 64712 26327
0 26329 5 1 1 26328
0 26330 7 1 2 78328 94055
0 26331 5 2 1 26330
0 26332 7 2 2 99682 90476
0 26333 5 1 1 101336
0 26334 7 1 2 66542 101337
0 26335 5 1 1 26334
0 26336 7 1 2 101334 26335
0 26337 5 1 1 26336
0 26338 7 1 2 65408 26337
0 26339 5 1 1 26338
0 26340 7 1 2 66543 100130
0 26341 5 1 1 26340
0 26342 7 1 2 26339 26341
0 26343 5 1 1 26342
0 26344 7 1 2 73482 26343
0 26345 5 1 1 26344
0 26346 7 1 2 100067 82272
0 26347 5 1 1 26346
0 26348 7 1 2 26345 26347
0 26349 5 1 1 26348
0 26350 7 1 2 73116 26349
0 26351 5 1 1 26350
0 26352 7 1 2 26329 26351
0 26353 5 1 1 26352
0 26354 7 1 2 66279 26353
0 26355 5 1 1 26354
0 26356 7 1 2 94056 78895
0 26357 5 1 1 26356
0 26358 7 1 2 90477 94226
0 26359 5 2 1 26358
0 26360 7 1 2 94023 101338
0 26361 5 1 1 26360
0 26362 7 1 2 75079 26361
0 26363 5 1 1 26362
0 26364 7 1 2 26357 26363
0 26365 5 1 1 26364
0 26366 7 1 2 75607 26365
0 26367 5 1 1 26366
0 26368 7 1 2 66739 90670
0 26369 7 1 2 95009 26368
0 26370 5 1 1 26369
0 26371 7 1 2 76587 98683
0 26372 7 1 2 89605 26371
0 26373 5 1 1 26372
0 26374 7 1 2 26370 26373
0 26375 7 1 2 26367 26374
0 26376 5 1 1 26375
0 26377 7 1 2 65409 26376
0 26378 5 1 1 26377
0 26379 7 1 2 67641 26378
0 26380 7 1 2 26355 26379
0 26381 5 1 1 26380
0 26382 7 3 2 68398 97394
0 26383 5 1 1 101340
0 26384 7 1 2 85934 101341
0 26385 5 1 1 26384
0 26386 7 1 2 100622 26385
0 26387 5 1 1 26386
0 26388 7 1 2 73117 26387
0 26389 5 1 1 26388
0 26390 7 1 2 92225 80046
0 26391 5 1 1 26390
0 26392 7 1 2 26389 26391
0 26393 5 1 1 26392
0 26394 7 1 2 71660 26393
0 26395 5 1 1 26394
0 26396 7 1 2 74786 100620
0 26397 5 1 1 26396
0 26398 7 1 2 26395 26397
0 26399 5 1 1 26398
0 26400 7 1 2 70188 26399
0 26401 5 1 1 26400
0 26402 7 1 2 84215 89416
0 26403 5 1 1 26402
0 26404 7 1 2 26401 26403
0 26405 5 1 1 26404
0 26406 7 1 2 68662 26405
0 26407 5 1 1 26406
0 26408 7 1 2 66280 91764
0 26409 5 2 1 26408
0 26410 7 2 2 71379 79905
0 26411 5 1 1 101345
0 26412 7 1 2 101343 26411
0 26413 5 1 1 26412
0 26414 7 1 2 98684 26413
0 26415 5 1 1 26414
0 26416 7 1 2 26407 26415
0 26417 5 1 1 26416
0 26418 7 1 2 81874 26417
0 26419 5 1 1 26418
0 26420 7 2 2 71380 84552
0 26421 5 1 1 101347
0 26422 7 1 2 100859 26421
0 26423 5 2 1 26422
0 26424 7 1 2 69838 101349
0 26425 5 1 1 26424
0 26426 7 1 2 74955 83648
0 26427 5 1 1 26426
0 26428 7 1 2 26425 26427
0 26429 5 1 1 26428
0 26430 7 1 2 90478 26429
0 26431 5 1 1 26430
0 26432 7 1 2 83512 99957
0 26433 5 1 1 26432
0 26434 7 1 2 26431 26433
0 26435 5 1 1 26434
0 26436 7 1 2 65410 26435
0 26437 5 1 1 26436
0 26438 7 1 2 69839 100451
0 26439 5 1 1 26438
0 26440 7 1 2 95084 75028
0 26441 5 2 1 26440
0 26442 7 1 2 26439 101351
0 26443 5 1 1 26442
0 26444 7 1 2 76077 26443
0 26445 5 1 1 26444
0 26446 7 1 2 99948 100452
0 26447 5 1 1 26446
0 26448 7 2 2 83501 83324
0 26449 7 1 2 79067 74787
0 26450 7 1 2 101353 26449
0 26451 5 1 1 26450
0 26452 7 1 2 26447 26451
0 26453 7 1 2 26445 26452
0 26454 7 1 2 26437 26453
0 26455 5 1 1 26454
0 26456 7 1 2 85935 26455
0 26457 5 1 1 26456
0 26458 7 1 2 85739 74956
0 26459 5 1 1 26458
0 26460 7 1 2 74540 96821
0 26461 5 1 1 26460
0 26462 7 1 2 26459 26461
0 26463 5 1 1 26462
0 26464 7 1 2 69840 26463
0 26465 5 1 1 26464
0 26466 7 1 2 71381 96824
0 26467 5 1 1 26466
0 26468 7 1 2 76651 93951
0 26469 7 1 2 26467 26468
0 26470 5 1 1 26469
0 26471 7 1 2 82176 87221
0 26472 5 1 1 26471
0 26473 7 1 2 74957 26472
0 26474 5 1 1 26473
0 26475 7 1 2 75791 75653
0 26476 5 1 1 26475
0 26477 7 1 2 100730 26476
0 26478 5 1 1 26477
0 26479 7 1 2 89961 91953
0 26480 5 1 1 26479
0 26481 7 1 2 26478 26480
0 26482 5 1 1 26481
0 26483 7 1 2 75392 26482
0 26484 5 1 1 26483
0 26485 7 1 2 26474 26484
0 26486 7 1 2 26470 26485
0 26487 7 1 2 26465 26486
0 26488 5 1 1 26487
0 26489 7 1 2 85313 26488
0 26490 5 1 1 26489
0 26491 7 1 2 72669 26490
0 26492 7 1 2 26457 26491
0 26493 7 1 2 26419 26492
0 26494 5 1 1 26493
0 26495 7 1 2 101013 26494
0 26496 7 1 2 26381 26495
0 26497 5 1 1 26496
0 26498 7 1 2 26306 26497
0 26499 7 1 2 26230 26498
0 26500 5 1 1 26499
0 26501 7 1 2 72217 26500
0 26502 5 1 1 26501
0 26503 7 3 2 67170 86558
0 26504 7 2 2 63797 84525
0 26505 7 1 2 101355 101358
0 26506 7 1 2 95534 26505
0 26507 7 1 2 94146 26506
0 26508 5 1 1 26507
0 26509 7 1 2 26502 26508
0 26510 5 1 1 26509
0 26511 7 1 2 100270 26510
0 26512 5 1 1 26511
0 26513 7 3 2 81319 95039
0 26514 5 3 1 101360
0 26515 7 1 2 69841 101363
0 26516 5 1 1 26515
0 26517 7 1 2 101328 26516
0 26518 5 1 1 26517
0 26519 7 1 2 82976 26518
0 26520 5 1 1 26519
0 26521 7 1 2 26520 87862
0 26522 5 1 1 26521
0 26523 7 1 2 66001 26522
0 26524 5 1 1 26523
0 26525 7 1 2 82977 86269
0 26526 5 2 1 26525
0 26527 7 1 2 80247 101366
0 26528 5 1 1 26527
0 26529 7 2 2 73118 26528
0 26530 5 1 1 101368
0 26531 7 1 2 74541 90105
0 26532 5 3 1 26531
0 26533 7 2 2 87639 87381
0 26534 5 1 1 101373
0 26535 7 1 2 71081 101374
0 26536 5 1 1 26535
0 26537 7 1 2 101370 26536
0 26538 7 1 2 26530 26537
0 26539 5 2 1 26538
0 26540 7 5 2 64713 77443
0 26541 7 1 2 101375 101377
0 26542 5 1 1 26541
0 26543 7 1 2 78754 86733
0 26544 5 1 1 26543
0 26545 7 1 2 87083 26544
0 26546 5 1 1 26545
0 26547 7 1 2 26542 26546
0 26548 7 1 2 26524 26547
0 26549 5 1 1 26548
0 26550 7 1 2 67642 26549
0 26551 5 1 1 26550
0 26552 7 1 2 100903 93332
0 26553 5 1 1 26552
0 26554 7 2 2 76652 77444
0 26555 7 1 2 77229 432
0 26556 5 1 1 26555
0 26557 7 1 2 101382 26556
0 26558 5 1 1 26557
0 26559 7 1 2 91616 4218
0 26560 5 1 1 26559
0 26561 7 1 2 66740 26560
0 26562 7 1 2 26558 26561
0 26563 7 1 2 26553 26562
0 26564 5 1 1 26563
0 26565 7 1 2 80832 92599
0 26566 5 1 1 26565
0 26567 7 1 2 71821 26566
0 26568 5 1 1 26567
0 26569 7 1 2 72670 26568
0 26570 7 1 2 26564 26569
0 26571 5 1 1 26570
0 26572 7 1 2 26551 26571
0 26573 5 1 1 26572
0 26574 7 1 2 71382 26573
0 26575 5 1 1 26574
0 26576 7 1 2 71082 91092
0 26577 5 1 1 26576
0 26578 7 2 2 74542 80062
0 26579 7 1 2 69842 101384
0 26580 5 1 1 26579
0 26581 7 1 2 26577 26580
0 26582 5 1 1 26581
0 26583 7 1 2 95311 26582
0 26584 5 1 1 26583
0 26585 7 1 2 67643 82978
0 26586 7 1 2 2124 26585
0 26587 7 5 2 69843 74657
0 26588 5 1 1 101386
0 26589 7 1 2 26588 78057
0 26590 7 1 2 26586 26589
0 26591 5 1 1 26590
0 26592 7 1 2 26584 26591
0 26593 5 1 1 26592
0 26594 7 1 2 68399 26593
0 26595 5 1 1 26594
0 26596 7 1 2 64714 92737
0 26597 5 1 1 26596
0 26598 7 1 2 66741 92545
0 26599 7 1 2 26597 26598
0 26600 5 1 1 26599
0 26601 7 1 2 26595 26600
0 26602 5 1 1 26601
0 26603 7 1 2 68052 26602
0 26604 5 1 1 26603
0 26605 7 4 2 64715 87797
0 26606 5 5 1 101391
0 26607 7 1 2 78715 86810
0 26608 5 1 1 26607
0 26609 7 2 2 69844 91526
0 26610 5 1 1 101400
0 26611 7 1 2 26608 26610
0 26612 5 1 1 26611
0 26613 7 1 2 95312 26612
0 26614 5 1 1 26613
0 26615 7 1 2 101395 26614
0 26616 5 1 1 26615
0 26617 7 1 2 77161 26616
0 26618 5 1 1 26617
0 26619 7 1 2 26604 26618
0 26620 7 1 2 26575 26619
0 26621 5 1 1 26620
0 26622 7 1 2 65411 26621
0 26623 5 1 1 26622
0 26624 7 5 2 66281 91497
0 26625 5 1 1 101402
0 26626 7 1 2 26625 85049
0 26627 5 1 1 26626
0 26628 7 1 2 64716 26627
0 26629 5 1 1 26628
0 26630 7 1 2 86217 82193
0 26631 5 2 1 26630
0 26632 7 1 2 87679 101407
0 26633 7 1 2 26629 26632
0 26634 5 1 1 26633
0 26635 7 1 2 74543 26634
0 26636 5 1 1 26635
0 26637 7 1 2 84706 101392
0 26638 5 1 1 26637
0 26639 7 1 2 26636 26638
0 26640 5 1 1 26639
0 26641 7 1 2 68400 26640
0 26642 5 1 1 26641
0 26643 7 2 2 69845 93000
0 26644 5 1 1 101409
0 26645 7 1 2 97359 87798
0 26646 5 2 1 26645
0 26647 7 1 2 26644 101411
0 26648 5 1 1 26647
0 26649 7 1 2 83548 26648
0 26650 5 1 1 26649
0 26651 7 1 2 26642 26650
0 26652 5 1 1 26651
0 26653 7 1 2 77445 26652
0 26654 5 1 1 26653
0 26655 7 1 2 87992 1430
0 26656 7 1 2 101224 26655
0 26657 5 1 1 26656
0 26658 7 1 2 85079 26657
0 26659 5 1 1 26658
0 26660 7 1 2 75699 97679
0 26661 7 1 2 80936 26660
0 26662 5 1 1 26661
0 26663 7 1 2 26659 26662
0 26664 5 1 1 26663
0 26665 7 1 2 69846 26664
0 26666 5 1 1 26665
0 26667 7 1 2 75277 82194
0 26668 5 2 1 26667
0 26669 7 1 2 81493 101413
0 26670 5 1 1 26669
0 26671 7 1 2 92870 26670
0 26672 5 1 1 26671
0 26673 7 1 2 71383 97680
0 26674 7 1 2 94933 26673
0 26675 5 1 1 26674
0 26676 7 1 2 26672 26675
0 26677 7 1 2 26666 26676
0 26678 5 1 1 26677
0 26679 7 1 2 68053 26678
0 26680 5 1 1 26679
0 26681 7 1 2 92882 101176
0 26682 5 1 1 26681
0 26683 7 2 2 75588 83788
0 26684 7 1 2 26682 101415
0 26685 5 1 1 26684
0 26686 7 1 2 80221 92579
0 26687 5 1 1 26686
0 26688 7 1 2 94934 90762
0 26689 5 1 1 26688
0 26690 7 1 2 26687 26689
0 26691 5 1 1 26690
0 26692 7 1 2 77446 26691
0 26693 5 1 1 26692
0 26694 7 1 2 26685 26693
0 26695 7 1 2 26680 26694
0 26696 5 1 1 26695
0 26697 7 1 2 80355 26696
0 26698 5 1 1 26697
0 26699 7 1 2 97395 98960
0 26700 5 1 1 26699
0 26701 7 1 2 71384 10955
0 26702 5 1 1 26701
0 26703 7 1 2 66282 76969
0 26704 5 1 1 26703
0 26705 7 1 2 83395 26704
0 26706 7 1 2 26702 26705
0 26707 5 1 1 26706
0 26708 7 1 2 26700 26707
0 26709 5 1 1 26708
0 26710 7 1 2 67644 26709
0 26711 5 1 1 26710
0 26712 7 1 2 92546 78789
0 26713 5 1 1 26712
0 26714 7 1 2 26711 26713
0 26715 5 1 1 26714
0 26716 7 1 2 73119 26715
0 26717 5 1 1 26716
0 26718 7 1 2 81656 92024
0 26719 5 1 1 26718
0 26720 7 1 2 71083 26719
0 26721 5 1 1 26720
0 26722 7 1 2 80151 80790
0 26723 5 1 1 26722
0 26724 7 1 2 26721 26723
0 26725 5 1 1 26724
0 26726 7 1 2 81466 26725
0 26727 5 1 1 26726
0 26728 7 1 2 26717 26727
0 26729 7 1 2 26698 26728
0 26730 7 1 2 26654 26729
0 26731 5 1 1 26730
0 26732 7 1 2 70441 26731
0 26733 5 1 1 26732
0 26734 7 2 2 83601 81415
0 26735 5 1 1 101417
0 26736 7 1 2 26735 5314
0 26737 5 1 1 26736
0 26738 7 1 2 78803 26737
0 26739 5 1 1 26738
0 26740 7 1 2 71822 81379
0 26741 5 1 1 26740
0 26742 7 1 2 79930 26741
0 26743 5 1 1 26742
0 26744 7 1 2 71385 26743
0 26745 5 1 1 26744
0 26746 7 1 2 70189 100858
0 26747 5 1 1 26746
0 26748 7 1 2 81250 26747
0 26749 5 1 1 26748
0 26750 7 1 2 98956 26749
0 26751 5 1 1 26750
0 26752 7 1 2 15570 26751
0 26753 7 1 2 26745 26752
0 26754 5 1 1 26753
0 26755 7 1 2 72671 26754
0 26756 5 1 1 26755
0 26757 7 1 2 26739 26756
0 26758 5 1 1 26757
0 26759 7 1 2 69847 26758
0 26760 5 1 1 26759
0 26761 7 1 2 74544 97360
0 26762 7 1 2 101418 26761
0 26763 5 1 1 26762
0 26764 7 1 2 26760 26763
0 26765 5 1 1 26764
0 26766 7 1 2 71084 26765
0 26767 5 1 1 26766
0 26768 7 1 2 71386 81374
0 26769 5 1 1 26768
0 26770 7 1 2 100860 26769
0 26771 5 1 1 26770
0 26772 7 1 2 70190 26771
0 26773 5 2 1 26772
0 26774 7 2 2 74740 77713
0 26775 5 1 1 101421
0 26776 7 1 2 101419 26775
0 26777 5 1 1 26776
0 26778 7 1 2 69848 26777
0 26779 5 1 1 26778
0 26780 7 1 2 74958 100792
0 26781 5 1 1 26780
0 26782 7 1 2 26779 26781
0 26783 5 1 1 26782
0 26784 7 1 2 98982 26783
0 26785 5 1 1 26784
0 26786 7 1 2 71823 81642
0 26787 5 1 1 26786
0 26788 7 1 2 81637 26787
0 26789 5 1 1 26788
0 26790 7 1 2 73120 26789
0 26791 5 1 1 26790
0 26792 7 1 2 75393 100760
0 26793 5 1 1 26792
0 26794 7 1 2 81657 26793
0 26795 5 1 1 26794
0 26796 7 1 2 71824 26795
0 26797 5 1 1 26796
0 26798 7 1 2 81653 26797
0 26799 5 1 1 26798
0 26800 7 1 2 72672 26799
0 26801 5 1 1 26800
0 26802 7 1 2 26791 26801
0 26803 5 1 1 26802
0 26804 7 1 2 71085 26803
0 26805 5 1 1 26804
0 26806 7 1 2 26785 26805
0 26807 5 1 1 26806
0 26808 7 1 2 69526 26807
0 26809 5 1 1 26808
0 26810 7 1 2 26767 26809
0 26811 7 1 2 26733 26810
0 26812 7 1 2 26623 26811
0 26813 5 1 1 26812
0 26814 7 1 2 72218 26813
0 26815 5 1 1 26814
0 26816 7 2 2 77886 100574
0 26817 7 2 2 77341 81667
0 26818 7 1 2 101423 101425
0 26819 5 1 1 26818
0 26820 7 12 2 72219 67645
0 26821 7 1 2 80457 101376
0 26822 5 1 1 26821
0 26823 7 1 2 80120 78922
0 26824 5 1 1 26823
0 26825 7 1 2 77447 82079
0 26826 5 1 1 26825
0 26827 7 1 2 26824 26826
0 26828 5 1 1 26827
0 26829 7 1 2 87626 26828
0 26830 5 1 1 26829
0 26831 7 1 2 90106 87844
0 26832 5 1 1 26831
0 26833 7 1 2 2141 26832
0 26834 5 1 1 26833
0 26835 7 1 2 69527 26834
0 26836 5 1 1 26835
0 26837 7 2 2 70191 81982
0 26838 7 1 2 101439 86724
0 26839 5 1 1 26838
0 26840 7 1 2 26836 26839
0 26841 7 1 2 26830 26840
0 26842 7 1 2 26822 26841
0 26843 5 1 1 26842
0 26844 7 1 2 101427 26843
0 26845 5 1 1 26844
0 26846 7 1 2 69528 87627
0 26847 5 1 1 26846
0 26848 7 1 2 26847 95793
0 26849 5 1 1 26848
0 26850 7 1 2 82580 26849
0 26851 5 1 1 26850
0 26852 7 1 2 77230 26851
0 26853 5 1 1 26852
0 26854 7 1 2 101428 26853
0 26855 5 1 1 26854
0 26856 7 1 2 68054 86551
0 26857 5 1 1 26856
0 26858 7 5 2 67171 73483
0 26859 7 1 2 82681 83728
0 26860 7 1 2 101441 26859
0 26861 7 1 2 26857 26860
0 26862 5 1 1 26861
0 26863 7 1 2 26855 26862
0 26864 5 1 1 26863
0 26865 7 1 2 64717 26864
0 26866 5 1 1 26865
0 26867 7 1 2 64399 77669
0 26868 7 1 2 100575 93442
0 26869 7 1 2 26867 26868
0 26870 7 1 2 96896 26869
0 26871 5 1 1 26870
0 26872 7 1 2 26866 26871
0 26873 7 1 2 26845 26872
0 26874 5 1 1 26873
0 26875 7 1 2 84979 26874
0 26876 5 1 1 26875
0 26877 7 1 2 26819 26876
0 26878 7 1 2 26815 26877
0 26879 5 1 1 26878
0 26880 7 1 2 64101 26879
0 26881 5 1 1 26880
0 26882 7 2 2 66544 75508
0 26883 7 1 2 88307 101446
0 26884 5 1 1 26883
0 26885 7 1 2 64400 81604
0 26886 5 1 1 26885
0 26887 7 1 2 68055 26886
0 26888 7 1 2 26884 26887
0 26889 5 1 1 26888
0 26890 7 1 2 75782 81597
0 26891 5 2 1 26890
0 26892 7 1 2 80971 96140
0 26893 5 1 1 26892
0 26894 7 1 2 73121 26893
0 26895 7 1 2 101448 26894
0 26896 5 1 1 26895
0 26897 7 1 2 71825 26896
0 26898 7 1 2 26889 26897
0 26899 5 1 1 26898
0 26900 7 1 2 66283 79778
0 26901 5 1 1 26900
0 26902 7 1 2 77282 79767
0 26903 7 1 2 79430 26902
0 26904 5 1 1 26903
0 26905 7 1 2 26901 26904
0 26906 5 1 1 26905
0 26907 7 1 2 66742 26906
0 26908 5 1 1 26907
0 26909 7 1 2 81223 92087
0 26910 5 1 1 26909
0 26911 7 1 2 64718 26910
0 26912 5 1 1 26911
0 26913 7 1 2 1157 76058
0 26914 7 1 2 78756 26913
0 26915 5 1 1 26914
0 26916 7 1 2 64401 26915
0 26917 5 1 1 26916
0 26918 7 1 2 26912 26917
0 26919 5 1 1 26918
0 26920 7 1 2 81875 26919
0 26921 5 1 1 26920
0 26922 7 1 2 26908 26921
0 26923 7 1 2 26899 26922
0 26924 5 1 1 26923
0 26925 7 1 2 68401 26924
0 26926 5 1 1 26925
0 26927 7 1 2 90042 83291
0 26928 5 1 1 26927
0 26929 7 1 2 78597 81591
0 26930 5 3 1 26929
0 26931 7 1 2 65096 101450
0 26932 7 1 2 99958 26931
0 26933 5 1 1 26932
0 26934 7 1 2 26928 26933
0 26935 5 1 1 26934
0 26936 7 1 2 66743 26935
0 26937 5 1 1 26936
0 26938 7 1 2 101237 82080
0 26939 5 1 1 26938
0 26940 7 1 2 78841 26939
0 26941 5 1 1 26940
0 26942 7 1 2 73484 26941
0 26943 5 1 1 26942
0 26944 7 1 2 26937 26943
0 26945 7 1 2 26926 26944
0 26946 5 1 1 26945
0 26947 7 1 2 66002 26946
0 26948 5 1 1 26947
0 26949 7 2 2 71826 81605
0 26950 5 2 1 101453
0 26951 7 1 2 101455 93783
0 26952 5 2 1 26951
0 26953 7 1 2 66003 101457
0 26954 5 1 1 26953
0 26955 7 2 2 71661 101456
0 26956 5 1 1 101459
0 26957 7 1 2 101206 26956
0 26958 5 1 1 26957
0 26959 7 1 2 26954 26958
0 26960 5 1 1 26959
0 26961 7 1 2 68402 26960
0 26962 5 1 1 26961
0 26963 7 1 2 12123 26962
0 26964 5 1 1 26963
0 26965 7 1 2 99865 26964
0 26966 5 1 1 26965
0 26967 7 1 2 81571 86993
0 26968 5 1 1 26967
0 26969 7 2 2 80162 80177
0 26970 7 1 2 81733 101461
0 26971 5 1 1 26970
0 26972 7 1 2 26968 26971
0 26973 5 1 1 26972
0 26974 7 1 2 66545 26973
0 26975 5 1 1 26974
0 26976 7 1 2 99959 94010
0 26977 5 1 1 26976
0 26978 7 1 2 26975 26977
0 26979 5 1 1 26978
0 26980 7 1 2 87985 26979
0 26981 5 1 1 26980
0 26982 7 1 2 72673 26981
0 26983 7 1 2 26966 26982
0 26984 7 1 2 26948 26983
0 26985 5 1 1 26984
0 26986 7 1 2 86227 96144
0 26987 5 1 1 26986
0 26988 7 2 2 66546 26987
0 26989 5 1 1 101463
0 26990 7 1 2 26989 86917
0 26991 5 1 1 26990
0 26992 7 2 2 64719 78044
0 26993 7 1 2 26991 101465
0 26994 5 1 1 26993
0 26995 7 1 2 90112 94265
0 26996 5 2 1 26995
0 26997 7 1 2 73122 101467
0 26998 5 1 1 26997
0 26999 7 1 2 82231 86797
0 27000 7 1 2 26998 26999
0 27001 5 1 1 27000
0 27002 7 1 2 77342 27001
0 27003 5 1 1 27002
0 27004 7 1 2 26994 27003
0 27005 5 1 1 27004
0 27006 7 1 2 65097 27005
0 27007 5 1 1 27006
0 27008 7 1 2 84982 87304
0 27009 5 1 1 27008
0 27010 7 1 2 78646 27009
0 27011 5 1 1 27010
0 27012 7 1 2 78821 6602
0 27013 5 1 1 27012
0 27014 7 1 2 27011 27013
0 27015 5 1 1 27014
0 27016 7 1 2 77343 27015
0 27017 5 1 1 27016
0 27018 7 1 2 67646 27017
0 27019 7 1 2 27007 27018
0 27020 5 1 1 27019
0 27021 7 1 2 100136 27020
0 27022 7 1 2 26985 27021
0 27023 5 1 1 27022
0 27024 7 1 2 26881 27023
0 27025 5 1 1 27024
0 27026 7 1 2 85936 27025
0 27027 5 1 1 27026
0 27028 7 1 2 76222 89020
0 27029 5 1 1 27028
0 27030 7 12 2 73485 97396
0 27031 5 1 1 101469
0 27032 7 1 2 84831 101470
0 27033 5 1 1 27032
0 27034 7 1 2 27029 27033
0 27035 5 1 1 27034
0 27036 7 1 2 68663 27035
0 27037 5 1 1 27036
0 27038 7 1 2 64720 101254
0 27039 5 1 1 27038
0 27040 7 1 2 27037 27039
0 27041 5 1 1 27040
0 27042 7 1 2 97990 27041
0 27043 5 1 1 27042
0 27044 7 1 2 76588 94288
0 27045 5 1 1 27044
0 27046 7 3 2 76322 27045
0 27047 7 3 2 64102 77231
0 27048 5 1 1 101484
0 27049 7 1 2 101481 101485
0 27050 5 1 1 27049
0 27051 7 1 2 68056 27050
0 27052 7 1 2 27043 27051
0 27053 5 1 1 27052
0 27054 7 1 2 97991 83819
0 27055 5 1 1 27054
0 27056 7 1 2 82702 27055
0 27057 5 1 1 27056
0 27058 7 1 2 69849 27057
0 27059 5 1 1 27058
0 27060 7 1 2 97779 77232
0 27061 5 1 1 27060
0 27062 7 1 2 82697 27061
0 27063 5 1 1 27062
0 27064 7 4 2 69161 77233
0 27065 7 1 2 77448 77954
0 27066 5 1 1 27065
0 27067 7 1 2 101487 27066
0 27068 5 1 1 27067
0 27069 7 1 2 66284 27068
0 27070 7 1 2 27063 27069
0 27071 7 1 2 27059 27070
0 27072 5 1 1 27071
0 27073 7 1 2 64402 89031
0 27074 5 1 1 27073
0 27075 7 1 2 82703 27074
0 27076 5 1 1 27075
0 27077 7 1 2 64721 27076
0 27078 5 1 1 27077
0 27079 7 1 2 65098 86031
0 27080 5 1 1 27079
0 27081 7 2 2 69850 27080
0 27082 5 1 1 101491
0 27083 7 1 2 77344 79231
0 27084 7 1 2 101492 27083
0 27085 5 1 1 27084
0 27086 7 1 2 71387 27085
0 27087 7 1 2 27078 27086
0 27088 5 1 1 27087
0 27089 7 1 2 27072 27088
0 27090 5 1 1 27089
0 27091 7 1 2 77345 86842
0 27092 5 2 1 27091
0 27093 7 1 2 82704 101493
0 27094 5 1 1 27093
0 27095 7 1 2 71388 27094
0 27096 5 1 1 27095
0 27097 7 1 2 69162 93234
0 27098 5 1 1 27097
0 27099 7 1 2 27096 27098
0 27100 5 1 1 27099
0 27101 7 1 2 80702 27100
0 27102 5 1 1 27101
0 27103 7 6 2 66004 79278
0 27104 7 2 2 84832 75473
0 27105 5 2 1 101501
0 27106 7 2 2 71389 101502
0 27107 7 1 2 101495 101505
0 27108 5 1 1 27107
0 27109 7 1 2 27102 27108
0 27110 5 1 1 27109
0 27111 7 1 2 73486 27110
0 27112 5 1 1 27111
0 27113 7 1 2 2440 101317
0 27114 5 1 1 27113
0 27115 7 1 2 73123 27114
0 27116 7 1 2 27112 27115
0 27117 7 1 2 27090 27116
0 27118 5 1 1 27117
0 27119 7 1 2 27053 27118
0 27120 5 1 1 27119
0 27121 7 3 2 69163 77449
0 27122 5 4 1 101507
0 27123 7 7 2 68057 97397
0 27124 7 1 2 98808 101514
0 27125 5 1 1 27124
0 27126 7 1 2 73124 100471
0 27127 5 1 1 27126
0 27128 7 1 2 27125 27127
0 27129 5 1 1 27128
0 27130 7 1 2 68403 27129
0 27131 5 1 1 27130
0 27132 7 1 2 95329 95906
0 27133 5 1 1 27132
0 27134 7 1 2 27131 27133
0 27135 5 1 1 27134
0 27136 7 1 2 65099 27135
0 27137 5 1 1 27136
0 27138 7 1 2 86303 83431
0 27139 5 1 1 27138
0 27140 7 2 2 73125 27139
0 27141 7 1 2 100472 101521
0 27142 5 1 1 27141
0 27143 7 1 2 27137 27142
0 27144 5 1 1 27143
0 27145 7 1 2 101510 27144
0 27146 5 1 1 27145
0 27147 7 2 2 82670 88348
0 27148 7 1 2 81135 101523
0 27149 5 1 1 27148
0 27150 7 1 2 82705 27149
0 27151 5 1 1 27150
0 27152 7 1 2 73126 79576
0 27153 5 1 1 27152
0 27154 7 1 2 100322 27153
0 27155 5 1 1 27154
0 27156 7 1 2 27151 27155
0 27157 5 1 1 27156
0 27158 7 1 2 76483 101486
0 27159 7 1 2 95772 27158
0 27160 5 1 1 27159
0 27161 7 1 2 67647 2034
0 27162 7 1 2 27160 27161
0 27163 7 1 2 27157 27162
0 27164 7 1 2 27146 27163
0 27165 7 1 2 27120 27164
0 27166 5 1 1 27165
0 27167 7 2 2 71086 75976
0 27168 5 1 1 101525
0 27169 7 2 2 64103 101526
0 27170 5 1 1 101527
0 27171 7 1 2 79475 91132
0 27172 7 1 2 89177 27171
0 27173 5 1 1 27172
0 27174 7 1 2 27170 27173
0 27175 5 1 1 27174
0 27176 7 1 2 69851 27175
0 27177 5 1 1 27176
0 27178 7 1 2 77234 85388
0 27179 5 2 1 27178
0 27180 7 2 2 74959 93558
0 27181 5 3 1 101531
0 27182 7 1 2 101529 101533
0 27183 7 1 2 27177 27182
0 27184 5 1 1 27183
0 27185 7 1 2 71662 27184
0 27186 5 1 1 27185
0 27187 7 1 2 79994 101528
0 27188 5 1 1 27187
0 27189 7 1 2 101530 27188
0 27190 5 1 1 27189
0 27191 7 1 2 80616 27190
0 27192 5 1 1 27191
0 27193 7 1 2 64104 94266
0 27194 5 1 1 27193
0 27195 7 1 2 90873 80121
0 27196 7 1 2 98809 27195
0 27197 5 1 1 27196
0 27198 7 1 2 27194 27197
0 27199 5 1 1 27198
0 27200 7 1 2 69529 99106
0 27201 7 1 2 27199 27200
0 27202 5 1 1 27201
0 27203 7 1 2 27192 27202
0 27204 7 1 2 27186 27203
0 27205 5 1 1 27204
0 27206 7 1 2 68404 27205
0 27207 5 1 1 27206
0 27208 7 1 2 88322 97657
0 27209 5 1 1 27208
0 27210 7 2 2 64722 97780
0 27211 7 1 2 66285 101536
0 27212 5 1 1 27211
0 27213 7 1 2 77235 95895
0 27214 7 1 2 27212 27213
0 27215 5 1 1 27214
0 27216 7 1 2 27209 27215
0 27217 5 1 1 27216
0 27218 7 1 2 69164 27217
0 27219 5 1 1 27218
0 27220 7 4 2 71087 83187
0 27221 7 1 2 89663 101538
0 27222 7 1 2 99928 27221
0 27223 5 1 1 27222
0 27224 7 1 2 73127 27223
0 27225 7 1 2 27219 27224
0 27226 5 1 1 27225
0 27227 7 1 2 66286 97781
0 27228 5 2 1 27227
0 27229 7 1 2 69852 101542
0 27230 5 1 1 27229
0 27231 7 1 2 84160 83151
0 27232 5 2 1 27231
0 27233 7 1 2 77236 101544
0 27234 7 1 2 27230 27233
0 27235 5 1 1 27234
0 27236 7 1 2 82698 27235
0 27237 5 1 1 27236
0 27238 7 1 2 101296 101488
0 27239 5 1 1 27238
0 27240 7 1 2 68058 27239
0 27241 7 1 2 27237 27240
0 27242 5 1 1 27241
0 27243 7 1 2 27226 27242
0 27244 5 1 1 27243
0 27245 7 1 2 71088 101543
0 27246 5 1 1 27245
0 27247 7 1 2 64723 27246
0 27248 5 1 1 27247
0 27249 7 1 2 66005 101545
0 27250 5 1 1 27249
0 27251 7 1 2 69530 27250
0 27252 7 1 2 27248 27251
0 27253 5 1 1 27252
0 27254 7 2 2 84161 81983
0 27255 7 1 2 80895 101546
0 27256 5 1 1 27255
0 27257 7 1 2 27253 27256
0 27258 5 1 1 27257
0 27259 7 1 2 64105 27258
0 27260 5 1 1 27259
0 27261 7 1 2 69165 101270
0 27262 5 1 1 27261
0 27263 7 1 2 72674 27262
0 27264 7 1 2 27260 27263
0 27265 7 1 2 27244 27264
0 27266 7 1 2 27207 27265
0 27267 5 1 1 27266
0 27268 7 1 2 72220 27267
0 27269 7 1 2 27166 27268
0 27270 5 1 1 27269
0 27271 7 10 2 66006 84526
0 27272 7 1 2 76223 101548
0 27273 7 1 2 101424 27272
0 27274 5 1 1 27273
0 27275 7 1 2 27270 27274
0 27276 5 1 1 27275
0 27277 7 1 2 85314 27276
0 27278 5 1 1 27277
0 27279 7 1 2 69853 83673
0 27280 5 1 1 27279
0 27281 7 1 2 67172 101549
0 27282 7 1 2 27280 27281
0 27283 5 1 1 27282
0 27284 7 1 2 72221 101121
0 27285 7 1 2 80327 27284
0 27286 5 1 1 27285
0 27287 7 1 2 27283 27286
0 27288 5 1 1 27287
0 27289 7 1 2 85315 27288
0 27290 5 1 1 27289
0 27291 7 9 2 68059 77237
0 27292 5 1 1 101558
0 27293 7 1 2 69854 101559
0 27294 5 2 1 27293
0 27295 7 1 2 87118 101567
0 27296 5 1 1 27295
0 27297 7 3 2 72055 72222
0 27298 7 1 2 93701 101569
0 27299 7 1 2 27296 27298
0 27300 5 1 1 27299
0 27301 7 1 2 27290 27300
0 27302 5 1 1 27301
0 27303 7 1 2 78647 27302
0 27304 5 1 1 27303
0 27305 7 6 2 72223 68405
0 27306 7 3 2 77238 94689
0 27307 7 1 2 70442 101122
0 27308 7 1 2 101578 27307
0 27309 5 1 1 27308
0 27310 7 2 2 96000 90894
0 27311 7 1 2 81984 91068
0 27312 7 1 2 101581 27311
0 27313 5 1 1 27312
0 27314 7 1 2 27309 27313
0 27315 5 1 1 27314
0 27316 7 1 2 101572 27315
0 27317 5 1 1 27316
0 27318 7 1 2 27304 27317
0 27319 5 1 1 27318
0 27320 7 1 2 66287 27319
0 27321 5 1 1 27320
0 27322 7 3 2 68855 93605
0 27323 7 1 2 76357 81437
0 27324 7 1 2 101583 27323
0 27325 5 1 1 27324
0 27326 7 1 2 77871 83218
0 27327 7 1 2 101582 27326
0 27328 5 1 1 27327
0 27329 7 1 2 27325 27328
0 27330 5 1 1 27329
0 27331 7 1 2 71089 27330
0 27332 5 1 1 27331
0 27333 7 3 2 64724 79813
0 27334 5 3 1 101586
0 27335 7 1 2 101118 101589
0 27336 5 1 1 27335
0 27337 7 1 2 87036 79906
0 27338 7 1 2 101579 27337
0 27339 7 1 2 27336 27338
0 27340 5 1 1 27339
0 27341 7 1 2 27332 27340
0 27342 5 1 1 27341
0 27343 7 1 2 71390 27342
0 27344 5 1 1 27343
0 27345 7 2 2 75577 88349
0 27346 7 1 2 87528 93702
0 27347 7 1 2 101592 27346
0 27348 5 1 1 27347
0 27349 7 1 2 27344 27348
0 27350 5 1 1 27349
0 27351 7 1 2 72224 27350
0 27352 5 1 1 27351
0 27353 7 1 2 27321 27352
0 27354 5 1 1 27353
0 27355 7 1 2 72675 27354
0 27356 5 1 1 27355
0 27357 7 1 2 93458 82566
0 27358 5 1 1 27357
0 27359 7 2 2 100565 101511
0 27360 7 1 2 68060 101594
0 27361 5 1 1 27360
0 27362 7 1 2 27358 27361
0 27363 5 1 1 27362
0 27364 7 1 2 76484 27363
0 27365 5 1 1 27364
0 27366 7 1 2 81153 101580
0 27367 5 1 1 27366
0 27368 7 1 2 27365 27367
0 27369 5 1 1 27368
0 27370 7 1 2 78648 27369
0 27371 5 1 1 27370
0 27372 7 1 2 73914 101515
0 27373 7 1 2 101595 27372
0 27374 5 1 1 27373
0 27375 7 1 2 27371 27374
0 27376 5 1 1 27375
0 27377 7 1 2 101429 27376
0 27378 5 1 1 27377
0 27379 7 1 2 27356 27378
0 27380 5 1 1 27379
0 27381 7 1 2 90479 27380
0 27382 5 1 1 27381
0 27383 7 1 2 27278 27382
0 27384 7 1 2 27027 27383
0 27385 5 1 1 27384
0 27386 7 1 2 100183 27385
0 27387 5 1 1 27386
0 27388 7 1 2 26512 27387
0 27389 5 1 1 27388
0 27390 7 1 2 72385 27389
0 27391 5 1 1 27390
0 27392 7 1 2 65412 23917
0 27393 5 1 1 27392
0 27394 7 1 2 70192 99923
0 27395 5 1 1 27394
0 27396 7 1 2 100548 27395
0 27397 5 1 1 27396
0 27398 7 1 2 73487 27397
0 27399 5 1 1 27398
0 27400 7 1 2 100447 27399
0 27401 5 1 1 27400
0 27402 7 1 2 81154 27401
0 27403 5 1 1 27402
0 27404 7 1 2 27393 27403
0 27405 5 1 1 27404
0 27406 7 1 2 85316 27405
0 27407 5 1 1 27406
0 27408 7 1 2 65100 86802
0 27409 5 1 1 27408
0 27410 7 1 2 64725 83666
0 27411 5 1 1 27410
0 27412 7 1 2 27409 27411
0 27413 5 1 1 27412
0 27414 7 1 2 82223 94690
0 27415 7 1 2 27413 27414
0 27416 5 1 1 27415
0 27417 7 1 2 27407 27416
0 27418 5 1 1 27417
0 27419 7 1 2 100184 27418
0 27420 5 1 1 27419
0 27421 7 2 2 88027 78310
0 27422 7 2 2 66744 101596
0 27423 7 3 2 77001 83219
0 27424 7 1 2 95575 78355
0 27425 7 1 2 101600 27424
0 27426 7 1 2 101598 27425
0 27427 5 1 1 27426
0 27428 7 1 2 27420 27427
0 27429 5 1 1 27428
0 27430 7 1 2 94685 27429
0 27431 5 1 1 27430
0 27432 7 7 2 98908 97691
0 27433 5 1 1 101603
0 27434 7 1 2 65101 92015
0 27435 7 1 2 101604 27434
0 27436 5 2 1 27435
0 27437 7 2 2 76918 79448
0 27438 7 3 2 65645 93669
0 27439 7 1 2 91069 101614
0 27440 7 1 2 101612 27439
0 27441 5 2 1 27440
0 27442 7 1 2 89926 100941
0 27443 5 1 1 27442
0 27444 7 2 2 67000 90480
0 27445 7 1 2 63798 101619
0 27446 5 1 1 27445
0 27447 7 1 2 27443 27446
0 27448 5 1 1 27447
0 27449 7 2 2 73128 27448
0 27450 7 2 2 75668 91716
0 27451 7 2 2 65600 101623
0 27452 5 1 1 101625
0 27453 7 1 2 101621 101626
0 27454 5 2 1 27453
0 27455 7 1 2 10878 10916
0 27456 5 1 1 27455
0 27457 7 1 2 65413 27456
0 27458 5 1 1 27457
0 27459 7 1 2 85363 23113
0 27460 5 2 1 27459
0 27461 7 1 2 86791 101629
0 27462 5 1 1 27461
0 27463 7 1 2 27458 27462
0 27464 5 1 1 27463
0 27465 7 1 2 100185 27464
0 27466 5 1 1 27465
0 27467 7 1 2 79378 91387
0 27468 7 1 2 95231 27467
0 27469 7 1 2 84776 27468
0 27470 5 1 1 27469
0 27471 7 1 2 27466 27470
0 27472 5 1 1 27471
0 27473 7 1 2 64726 27472
0 27474 5 1 1 27473
0 27475 7 1 2 101627 27474
0 27476 5 1 1 27475
0 27477 7 1 2 73488 27476
0 27478 5 1 1 27477
0 27479 7 1 2 101617 27478
0 27480 5 1 1 27479
0 27481 7 1 2 66547 27480
0 27482 5 1 1 27481
0 27483 7 1 2 101610 27482
0 27484 5 1 1 27483
0 27485 7 1 2 66288 27484
0 27486 5 1 1 27485
0 27487 7 1 2 85317 75140
0 27488 5 1 1 27487
0 27489 7 1 2 94853 93146
0 27490 5 1 1 27489
0 27491 7 1 2 27488 27490
0 27492 5 1 1 27491
0 27493 7 1 2 66745 27492
0 27494 5 1 1 27493
0 27495 7 1 2 84573 86085
0 27496 5 1 1 27495
0 27497 7 1 2 27494 27496
0 27498 5 1 1 27497
0 27499 7 1 2 82742 27498
0 27500 5 1 1 27499
0 27501 7 1 2 83382 93919
0 27502 5 1 1 27501
0 27503 7 1 2 85318 27502
0 27504 5 1 1 27503
0 27505 7 1 2 73129 90692
0 27506 5 1 1 27505
0 27507 7 1 2 27504 27506
0 27508 5 1 1 27507
0 27509 7 1 2 66289 27508
0 27510 5 1 1 27509
0 27511 7 1 2 75625 79874
0 27512 5 1 1 27511
0 27513 7 1 2 90711 2871
0 27514 7 1 2 27512 27513
0 27515 5 1 1 27514
0 27516 7 1 2 27510 27515
0 27517 7 1 2 27500 27516
0 27518 5 1 1 27517
0 27519 7 1 2 100186 27518
0 27520 5 1 1 27519
0 27521 7 1 2 90481 78923
0 27522 5 1 1 27521
0 27523 7 3 2 73130 90464
0 27524 5 1 1 101631
0 27525 7 1 2 87573 101632
0 27526 5 1 1 27525
0 27527 7 1 2 27522 27526
0 27528 5 1 1 27527
0 27529 7 1 2 73489 27528
0 27530 5 1 1 27529
0 27531 7 2 2 82921 83789
0 27532 5 1 1 101634
0 27533 7 1 2 65102 87646
0 27534 5 2 1 27533
0 27535 7 1 2 27532 101636
0 27536 5 1 1 27535
0 27537 7 1 2 73131 27536
0 27538 5 1 1 27537
0 27539 7 2 2 27530 27538
0 27540 5 1 1 101638
0 27541 7 1 2 85937 27540
0 27542 5 1 1 27541
0 27543 7 1 2 101333 27542
0 27544 5 1 1 27543
0 27545 7 1 2 66290 27544
0 27546 5 1 1 27545
0 27547 7 1 2 100061 87369
0 27548 5 1 1 27547
0 27549 7 1 2 100062 101339
0 27550 5 1 1 27549
0 27551 7 1 2 75080 27550
0 27552 5 1 1 27551
0 27553 7 1 2 82626 80438
0 27554 5 3 1 27553
0 27555 7 1 2 94384 101640
0 27556 5 1 1 27555
0 27557 7 1 2 65414 27556
0 27558 5 1 1 27557
0 27559 7 1 2 65103 84767
0 27560 5 1 1 27559
0 27561 7 1 2 27558 27560
0 27562 5 1 1 27561
0 27563 7 1 2 85319 27562
0 27564 5 1 1 27563
0 27565 7 1 2 27552 27564
0 27566 5 1 1 27565
0 27567 7 1 2 73132 27566
0 27568 5 1 1 27567
0 27569 7 1 2 27548 27568
0 27570 7 1 2 27546 27569
0 27571 5 1 1 27570
0 27572 7 1 2 64727 27571
0 27573 5 1 1 27572
0 27574 7 1 2 85320 86439
0 27575 5 1 1 27574
0 27576 7 1 2 74788 99981
0 27577 5 1 1 27576
0 27578 7 3 2 81734 78329
0 27579 5 1 1 101643
0 27580 7 1 2 89417 101644
0 27581 5 1 1 27580
0 27582 7 1 2 100132 26333
0 27583 5 1 1 27582
0 27584 7 1 2 73133 27583
0 27585 5 1 1 27584
0 27586 7 1 2 84804 75654
0 27587 5 1 1 27586
0 27588 7 1 2 83812 93394
0 27589 7 1 2 27587 27588
0 27590 5 1 1 27589
0 27591 7 1 2 27585 27590
0 27592 5 1 1 27591
0 27593 7 1 2 66548 27592
0 27594 5 1 1 27593
0 27595 7 1 2 27581 27594
0 27596 5 1 1 27595
0 27597 7 1 2 73490 27596
0 27598 5 1 1 27597
0 27599 7 1 2 27577 27598
0 27600 5 1 1 27599
0 27601 7 1 2 66291 27600
0 27602 5 1 1 27601
0 27603 7 1 2 27575 27602
0 27604 7 1 2 27573 27603
0 27605 5 1 1 27604
0 27606 7 1 2 100271 27605
0 27607 5 1 1 27606
0 27608 7 1 2 27520 27607
0 27609 5 1 1 27608
0 27610 7 1 2 64403 27609
0 27611 5 1 1 27610
0 27612 7 1 2 27486 27611
0 27613 5 1 1 27612
0 27614 7 1 2 66007 27613
0 27615 5 1 1 27614
0 27616 7 2 2 84071 91331
0 27617 7 2 2 70680 101646
0 27618 7 1 2 84908 101648
0 27619 5 1 1 27618
0 27620 7 1 2 27452 27619
0 27621 5 1 1 27620
0 27622 7 1 2 65104 27621
0 27623 5 1 1 27622
0 27624 7 1 2 100187 86792
0 27625 5 1 1 27624
0 27626 7 1 2 27623 27625
0 27627 5 2 1 27626
0 27628 7 1 2 85321 101650
0 27629 5 1 1 27628
0 27630 7 2 2 65105 86793
0 27631 5 2 1 101652
0 27632 7 1 2 83674 101654
0 27633 5 1 1 27632
0 27634 7 2 2 85938 27633
0 27635 5 1 1 101656
0 27636 7 1 2 100188 101657
0 27637 5 1 1 27636
0 27638 7 1 2 27629 27637
0 27639 5 1 1 27638
0 27640 7 1 2 64728 27639
0 27641 5 1 1 27640
0 27642 7 1 2 101628 27641
0 27643 5 1 1 27642
0 27644 7 1 2 73491 27643
0 27645 5 1 1 27644
0 27646 7 1 2 27645 101618
0 27647 5 1 1 27646
0 27648 7 1 2 66549 27647
0 27649 5 1 1 27648
0 27650 7 1 2 27649 101611
0 27651 5 1 1 27650
0 27652 7 1 2 79893 27651
0 27653 5 1 1 27652
0 27654 7 1 2 67648 27653
0 27655 7 1 2 27615 27654
0 27656 5 1 1 27655
0 27657 7 1 2 95904 101420
0 27658 5 1 1 27657
0 27659 7 1 2 86048 27658
0 27660 5 1 1 27659
0 27661 7 2 2 68061 101635
0 27662 5 1 1 101658
0 27663 7 1 2 71391 101659
0 27664 5 1 1 27663
0 27665 7 1 2 27660 27664
0 27666 5 1 1 27665
0 27667 7 1 2 64729 27666
0 27668 5 1 1 27667
0 27669 7 1 2 71392 101639
0 27670 5 1 1 27669
0 27671 7 1 2 86049 97666
0 27672 5 1 1 27671
0 27673 7 1 2 66292 27662
0 27674 7 1 2 27672 27673
0 27675 5 1 1 27674
0 27676 7 1 2 69855 27675
0 27677 7 1 2 27670 27676
0 27678 5 1 1 27677
0 27679 7 1 2 27668 27678
0 27680 5 1 1 27679
0 27681 7 2 2 96409 95544
0 27682 7 1 2 27680 101660
0 27683 5 1 1 27682
0 27684 7 1 2 69856 101369
0 27685 5 1 1 27684
0 27686 7 1 2 94927 101371
0 27687 5 2 1 27686
0 27688 7 1 2 68062 101662
0 27689 5 1 1 27688
0 27690 7 1 2 74545 74789
0 27691 5 2 1 27690
0 27692 7 2 2 68063 88335
0 27693 5 1 1 101666
0 27694 7 1 2 101664 27693
0 27695 5 1 1 27694
0 27696 7 1 2 82979 27695
0 27697 5 2 1 27696
0 27698 7 1 2 27689 101668
0 27699 7 1 2 27685 27698
0 27700 5 1 1 27699
0 27701 7 1 2 66008 27700
0 27702 5 1 1 27701
0 27703 7 1 2 75626 100456
0 27704 5 1 1 27703
0 27705 7 1 2 71090 82743
0 27706 7 1 2 27704 27705
0 27707 5 1 1 27706
0 27708 7 1 2 101568 27707
0 27709 5 1 1 27708
0 27710 7 1 2 73492 27709
0 27711 5 1 1 27710
0 27712 7 1 2 99841 87628
0 27713 5 1 1 27712
0 27714 7 1 2 82922 92766
0 27715 5 1 1 27714
0 27716 7 1 2 27713 27715
0 27717 5 1 1 27716
0 27718 7 1 2 68064 27717
0 27719 5 1 1 27718
0 27720 7 1 2 27711 27719
0 27721 5 1 1 27720
0 27722 7 1 2 66550 27721
0 27723 5 1 1 27722
0 27724 7 1 2 91444 87640
0 27725 7 1 2 101560 27724
0 27726 5 1 1 27725
0 27727 7 1 2 27723 27726
0 27728 7 1 2 27702 27727
0 27729 5 1 1 27728
0 27730 7 1 2 66293 27729
0 27731 5 1 1 27730
0 27732 7 3 2 66551 82169
0 27733 5 1 1 101670
0 27734 7 1 2 93967 101671
0 27735 5 2 1 27734
0 27736 7 1 2 87641 101123
0 27737 5 1 1 27736
0 27738 7 1 2 74754 86891
0 27739 5 1 1 27738
0 27740 7 1 2 66552 83176
0 27741 7 1 2 27739 27740
0 27742 5 1 1 27741
0 27743 7 1 2 27737 27742
0 27744 5 1 1 27743
0 27745 7 1 2 71393 27744
0 27746 5 1 1 27745
0 27747 7 1 2 101673 27746
0 27748 5 1 1 27747
0 27749 7 1 2 65106 27748
0 27750 5 1 1 27749
0 27751 7 1 2 91589 101124
0 27752 5 1 1 27751
0 27753 7 1 2 27750 27752
0 27754 5 1 1 27753
0 27755 7 1 2 64404 27754
0 27756 5 1 1 27755
0 27757 7 5 2 70193 87336
0 27758 7 1 2 88817 101675
0 27759 5 1 1 27758
0 27760 7 2 2 81224 27759
0 27761 5 1 1 101680
0 27762 7 3 2 73134 90113
0 27763 7 1 2 75394 101682
0 27764 5 1 1 27763
0 27765 7 1 2 78774 27764
0 27766 5 1 1 27765
0 27767 7 1 2 64730 27766
0 27768 5 1 1 27767
0 27769 7 1 2 101681 27768
0 27770 5 1 1 27769
0 27771 7 1 2 71394 27770
0 27772 5 1 1 27771
0 27773 7 1 2 68065 81182
0 27774 7 1 2 12444 27773
0 27775 5 1 1 27774
0 27776 7 1 2 66553 87629
0 27777 5 2 1 27776
0 27778 7 1 2 73135 101685
0 27779 5 1 1 27778
0 27780 7 1 2 71395 27779
0 27781 7 1 2 27775 27780
0 27782 5 1 1 27781
0 27783 7 1 2 101674 27782
0 27784 5 1 1 27783
0 27785 7 1 2 65107 27784
0 27786 5 1 1 27785
0 27787 7 1 2 69531 11484
0 27788 5 1 1 27787
0 27789 7 1 2 75977 27788
0 27790 5 1 1 27789
0 27791 7 1 2 101372 27790
0 27792 5 1 1 27791
0 27793 7 1 2 69857 74132
0 27794 7 1 2 27792 27793
0 27795 5 1 1 27794
0 27796 7 1 2 27786 27795
0 27797 7 1 2 27772 27796
0 27798 5 1 1 27797
0 27799 7 1 2 66009 27798
0 27800 5 1 1 27799
0 27801 7 1 2 27756 27800
0 27802 7 1 2 27731 27801
0 27803 5 1 1 27802
0 27804 7 1 2 65415 27803
0 27805 5 1 1 27804
0 27806 7 2 2 77560 93448
0 27807 5 2 1 101687
0 27808 7 1 2 73493 101688
0 27809 5 1 1 27808
0 27810 7 1 2 76653 75046
0 27811 5 1 1 27810
0 27812 7 1 2 94928 27811
0 27813 5 2 1 27812
0 27814 7 1 2 66294 101691
0 27815 5 2 1 27814
0 27816 7 1 2 65108 101346
0 27817 5 1 1 27816
0 27818 7 1 2 90558 27817
0 27819 7 1 2 101693 27818
0 27820 5 1 1 27819
0 27821 7 1 2 65109 79878
0 27822 5 1 1 27821
0 27823 7 1 2 81630 27822
0 27824 5 1 1 27823
0 27825 7 1 2 66010 27824
0 27826 7 1 2 27820 27825
0 27827 5 1 1 27826
0 27828 7 2 2 78695 78826
0 27829 5 1 1 101695
0 27830 7 1 2 83262 87986
0 27831 7 1 2 27829 27830
0 27832 5 1 1 27831
0 27833 7 1 2 27827 27832
0 27834 5 1 1 27833
0 27835 7 1 2 86673 27834
0 27836 5 1 1 27835
0 27837 7 1 2 27809 27836
0 27838 7 1 2 27805 27837
0 27839 5 1 1 27838
0 27840 7 1 2 100189 27839
0 27841 5 1 1 27840
0 27842 7 1 2 27683 27841
0 27843 5 1 1 27842
0 27844 7 1 2 85939 27843
0 27845 5 1 1 27844
0 27846 7 1 2 83424 77239
0 27847 5 1 1 27846
0 27848 7 1 2 100098 27847
0 27849 5 3 1 27848
0 27850 7 1 2 84205 101697
0 27851 5 1 1 27850
0 27852 7 1 2 22658 94509
0 27853 5 1 1 27852
0 27854 7 1 2 101300 27853
0 27855 5 1 1 27854
0 27856 7 1 2 82224 27855
0 27857 5 1 1 27856
0 27858 7 1 2 27851 27857
0 27859 5 1 1 27858
0 27860 7 1 2 64731 27859
0 27861 5 1 1 27860
0 27862 7 1 2 101302 101698
0 27863 5 1 1 27862
0 27864 7 1 2 27861 27863
0 27865 5 1 1 27864
0 27866 7 1 2 65416 27865
0 27867 5 1 1 27866
0 27868 7 1 2 77240 101304
0 27869 5 1 1 27868
0 27870 7 1 2 82225 84406
0 27871 5 1 1 27870
0 27872 7 1 2 27869 27871
0 27873 5 1 1 27872
0 27874 7 1 2 84768 27873
0 27875 5 1 1 27874
0 27876 7 1 2 27867 27875
0 27877 5 1 1 27876
0 27878 7 1 2 65110 27877
0 27879 5 1 1 27878
0 27880 7 1 2 80356 101313
0 27881 5 1 1 27880
0 27882 7 1 2 78696 78835
0 27883 5 1 1 27882
0 27884 7 1 2 27881 27883
0 27885 5 1 1 27884
0 27886 7 1 2 70443 27885
0 27887 5 1 1 27886
0 27888 7 1 2 78836 82719
0 27889 5 1 1 27888
0 27890 7 1 2 27887 27889
0 27891 5 1 1 27890
0 27892 7 1 2 70194 27891
0 27893 5 1 1 27892
0 27894 7 1 2 81876 84216
0 27895 5 1 1 27894
0 27896 7 1 2 79941 27895
0 27897 5 1 1 27896
0 27898 7 1 2 64405 27897
0 27899 5 1 1 27898
0 27900 7 1 2 27893 27899
0 27901 5 1 1 27900
0 27902 7 1 2 66011 27901
0 27903 5 1 1 27902
0 27904 7 1 2 27879 27903
0 27905 5 1 1 27904
0 27906 7 1 2 73136 27905
0 27907 5 1 1 27906
0 27908 7 1 2 84777 86252
0 27909 5 1 1 27908
0 27910 7 1 2 101211 27909
0 27911 5 1 1 27910
0 27912 7 1 2 69858 27911
0 27913 5 1 1 27912
0 27914 7 1 2 64732 98996
0 27915 5 1 1 27914
0 27916 7 1 2 101214 27915
0 27917 5 1 1 27916
0 27918 7 1 2 70195 27917
0 27919 5 1 1 27918
0 27920 7 1 2 27913 27919
0 27921 5 1 1 27920
0 27922 7 1 2 66295 27921
0 27923 5 1 1 27922
0 27924 7 1 2 82598 78330
0 27925 5 1 1 27924
0 27926 7 1 2 101641 27925
0 27927 5 1 1 27926
0 27928 7 1 2 71396 27927
0 27929 5 1 1 27928
0 27930 7 1 2 75395 100731
0 27931 5 1 1 27930
0 27932 7 1 2 27929 27931
0 27933 5 1 1 27932
0 27934 7 1 2 65417 27933
0 27935 5 1 1 27934
0 27936 7 1 2 65418 91734
0 27937 5 1 1 27936
0 27938 7 2 2 71397 100459
0 27939 5 1 1 101700
0 27940 7 1 2 27937 101701
0 27941 5 1 1 27940
0 27942 7 1 2 27935 27941
0 27943 5 1 1 27942
0 27944 7 1 2 64406 27943
0 27945 5 1 1 27944
0 27946 7 1 2 27923 27945
0 27947 5 1 1 27946
0 27948 7 1 2 66012 27947
0 27949 5 1 1 27948
0 27950 7 1 2 68664 99807
0 27951 5 1 1 27950
0 27952 7 1 2 99804 27951
0 27953 5 4 1 27952
0 27954 7 1 2 78311 101702
0 27955 5 1 1 27954
0 27956 7 2 2 66013 101207
0 27957 5 1 1 101706
0 27958 7 1 2 27955 27957
0 27959 5 1 1 27958
0 27960 7 1 2 101250 27959
0 27961 5 1 1 27960
0 27962 7 3 2 91445 78649
0 27963 5 1 1 101708
0 27964 7 1 2 88721 101709
0 27965 7 1 2 94173 27964
0 27966 5 1 1 27965
0 27967 7 1 2 27961 27966
0 27968 7 1 2 27949 27967
0 27969 5 1 1 27968
0 27970 7 1 2 68066 27969
0 27971 5 1 1 27970
0 27972 7 4 2 66014 75396
0 27973 7 1 2 82633 101711
0 27974 7 1 2 83859 27973
0 27975 5 1 1 27974
0 27976 7 1 2 27971 27975
0 27977 7 1 2 27907 27976
0 27978 5 1 1 27977
0 27979 7 1 2 100272 27978
0 27980 5 1 1 27979
0 27981 7 2 2 64733 15252
0 27982 5 1 1 101715
0 27983 7 1 2 95784 101716
0 27984 5 8 1 27983
0 27985 7 1 2 66296 101717
0 27986 5 1 1 27985
0 27987 7 1 2 82353 79339
0 27988 5 3 1 27987
0 27989 7 1 2 71398 82372
0 27990 5 1 1 27989
0 27991 7 1 2 101725 27990
0 27992 5 1 1 27991
0 27993 7 1 2 74658 27992
0 27994 5 1 1 27993
0 27995 7 1 2 97367 95900
0 27996 7 1 2 27994 27995
0 27997 7 1 2 27986 27996
0 27998 5 1 1 27997
0 27999 7 1 2 73137 27998
0 28000 5 1 1 27999
0 28001 7 1 2 78650 76024
0 28002 5 2 1 28001
0 28003 7 1 2 82354 84132
0 28004 5 5 1 28003
0 28005 7 1 2 74755 101730
0 28006 5 1 1 28005
0 28007 7 1 2 65111 28006
0 28008 5 1 1 28007
0 28009 7 1 2 86903 101726
0 28010 7 1 2 28008 28009
0 28011 5 1 1 28010
0 28012 7 1 2 1689 28011
0 28013 5 1 1 28012
0 28014 7 1 2 101728 28013
0 28015 7 1 2 28000 28014
0 28016 5 1 1 28015
0 28017 7 1 2 77241 28016
0 28018 5 1 1 28017
0 28019 7 1 2 75978 91614
0 28020 5 1 1 28019
0 28021 7 1 2 100334 28020
0 28022 5 1 1 28021
0 28023 7 1 2 99747 28022
0 28024 5 1 1 28023
0 28025 7 1 2 78651 77450
0 28026 5 1 1 28025
0 28027 7 1 2 100448 28026
0 28028 5 1 1 28027
0 28029 7 1 2 81155 28028
0 28030 5 1 1 28029
0 28031 7 1 2 64407 79998
0 28032 5 3 1 28031
0 28033 7 1 2 28030 101735
0 28034 7 1 2 28024 28033
0 28035 7 1 2 28018 28034
0 28036 5 1 1 28035
0 28037 7 1 2 100190 28036
0 28038 5 1 1 28037
0 28039 7 1 2 27980 28038
0 28040 5 1 1 28039
0 28041 7 1 2 85322 28040
0 28042 5 1 1 28041
0 28043 7 1 2 72676 28042
0 28044 7 1 2 27845 28043
0 28045 5 1 1 28044
0 28046 7 1 2 27656 28045
0 28047 5 1 1 28046
0 28048 7 2 2 79637 89142
0 28049 7 1 2 65646 82355
0 28050 7 1 2 92511 28049
0 28051 7 1 2 101738 28050
0 28052 7 1 2 75482 28051
0 28053 7 1 2 99787 28052
0 28054 5 1 1 28053
0 28055 7 1 2 28047 28054
0 28056 5 1 1 28055
0 28057 7 1 2 64106 28056
0 28058 5 1 1 28057
0 28059 7 1 2 27431 28058
0 28060 5 1 1 28059
0 28061 7 1 2 100078 28060
0 28062 5 1 1 28061
0 28063 7 1 2 27391 28062
0 28064 5 1 1 28063
0 28065 7 1 2 65798 28064
0 28066 5 1 1 28065
0 28067 7 1 2 101516 95211
0 28068 5 1 1 28067
0 28069 7 1 2 69532 89267
0 28070 5 1 1 28069
0 28071 7 1 2 28068 28070
0 28072 5 1 1 28071
0 28073 7 1 2 98810 28072
0 28074 5 1 1 28073
0 28075 7 1 2 97799 93194
0 28076 5 1 1 28075
0 28077 7 1 2 28074 28076
0 28078 5 1 1 28077
0 28079 7 1 2 68406 28078
0 28080 5 1 1 28079
0 28081 7 1 2 73138 95263
0 28082 7 1 2 100818 28081
0 28083 7 1 2 101496 28082
0 28084 5 1 1 28083
0 28085 7 1 2 28080 28084
0 28086 5 1 1 28085
0 28087 7 1 2 65112 28086
0 28088 5 1 1 28087
0 28089 7 4 2 79476 79279
0 28090 7 1 2 82217 101740
0 28091 7 1 2 101522 28090
0 28092 5 1 1 28091
0 28093 7 1 2 28088 28092
0 28094 5 1 1 28093
0 28095 7 1 2 101605 28094
0 28096 5 1 1 28095
0 28097 7 3 2 100191 101451
0 28098 5 1 1 101744
0 28099 7 2 2 68990 66015
0 28100 7 2 2 96410 101747
0 28101 7 1 2 73915 101749
0 28102 5 1 1 28101
0 28103 7 1 2 28098 28102
0 28104 5 1 1 28103
0 28105 7 1 2 66746 28104
0 28106 5 1 1 28105
0 28107 7 2 2 73740 79693
0 28108 7 1 2 95719 101751
0 28109 7 1 2 87166 28108
0 28110 5 1 1 28109
0 28111 7 1 2 28106 28110
0 28112 5 1 1 28111
0 28113 7 1 2 64408 28112
0 28114 5 1 1 28113
0 28115 7 1 2 84964 101745
0 28116 5 1 1 28115
0 28117 7 1 2 28114 28116
0 28118 5 1 1 28117
0 28119 7 1 2 65113 28118
0 28120 5 1 1 28119
0 28121 7 3 2 70681 71827
0 28122 7 2 2 83622 101753
0 28123 7 1 2 78652 79517
0 28124 7 1 2 100867 28123
0 28125 7 1 2 101756 28124
0 28126 5 1 1 28125
0 28127 7 1 2 28120 28126
0 28128 5 1 1 28127
0 28129 7 1 2 85940 28128
0 28130 5 1 1 28129
0 28131 7 1 2 86379 97288
0 28132 5 2 1 28131
0 28133 7 1 2 101212 101758
0 28134 5 1 1 28133
0 28135 7 1 2 66016 100296
0 28136 7 1 2 28134 28135
0 28137 5 1 1 28136
0 28138 7 1 2 28130 28137
0 28139 5 1 1 28138
0 28140 7 1 2 97398 28139
0 28141 5 1 1 28140
0 28142 7 2 2 83439 84143
0 28143 5 3 1 101760
0 28144 7 1 2 83532 96554
0 28145 5 1 1 28144
0 28146 7 1 2 101762 28145
0 28147 5 5 1 28146
0 28148 7 3 2 68665 101765
0 28149 5 2 1 101770
0 28150 7 1 2 100297 101771
0 28151 5 1 1 28150
0 28152 7 3 2 65419 86270
0 28153 5 1 1 101775
0 28154 7 1 2 66747 101776
0 28155 5 1 1 28154
0 28156 7 1 2 83456 28155
0 28157 5 1 1 28156
0 28158 7 1 2 68666 28157
0 28159 5 1 1 28158
0 28160 7 2 2 26034 28159
0 28161 7 2 2 66748 83790
0 28162 5 1 1 101780
0 28163 7 1 2 86937 28162
0 28164 5 1 1 28163
0 28165 7 1 2 65420 28164
0 28166 5 1 1 28165
0 28167 7 1 2 68407 98576
0 28168 5 1 1 28167
0 28169 7 1 2 28166 28168
0 28170 7 1 2 101778 28169
0 28171 5 1 1 28170
0 28172 7 1 2 100669 28171
0 28173 5 1 1 28172
0 28174 7 1 2 28151 28173
0 28175 5 1 1 28174
0 28176 7 1 2 64734 28175
0 28177 5 1 1 28176
0 28178 7 6 2 90589 82764
0 28179 7 2 2 90659 101782
0 28180 7 1 2 83220 101788
0 28181 5 1 1 28180
0 28182 7 1 2 28177 28181
0 28183 5 1 1 28182
0 28184 7 1 2 74152 28183
0 28185 5 1 1 28184
0 28186 7 1 2 90826 93434
0 28187 5 1 1 28186
0 28188 7 2 2 65114 79477
0 28189 5 1 1 101790
0 28190 7 1 2 28187 28189
0 28191 5 1 1 28190
0 28192 7 1 2 81735 28191
0 28193 5 1 1 28192
0 28194 7 5 2 74659 89371
0 28195 5 1 1 101792
0 28196 7 1 2 74153 28195
0 28197 5 1 1 28196
0 28198 7 1 2 28193 28197
0 28199 5 1 1 28198
0 28200 7 1 2 85323 28199
0 28201 5 1 1 28200
0 28202 7 1 2 90693 99985
0 28203 7 1 2 86050 28202
0 28204 5 1 1 28203
0 28205 7 1 2 28201 28204
0 28206 5 1 1 28205
0 28207 7 1 2 100273 28206
0 28208 5 1 1 28207
0 28209 7 1 2 80256 101460
0 28210 5 1 1 28209
0 28211 7 1 2 81877 77587
0 28212 7 1 2 100670 28211
0 28213 7 1 2 28210 28212
0 28214 5 1 1 28213
0 28215 7 1 2 28208 28214
0 28216 5 1 1 28215
0 28217 7 1 2 68408 28216
0 28218 5 1 1 28217
0 28219 7 1 2 82226 101606
0 28220 5 1 1 28219
0 28221 7 1 2 100671 89224
0 28222 5 1 1 28221
0 28223 7 1 2 81878 91592
0 28224 5 1 1 28223
0 28225 7 1 2 85740 79545
0 28226 5 1 1 28225
0 28227 7 1 2 28224 28226
0 28228 5 1 1 28227
0 28229 7 1 2 100274 28228
0 28230 5 1 1 28229
0 28231 7 1 2 100223 28230
0 28232 5 1 1 28231
0 28233 7 1 2 85324 28232
0 28234 5 1 1 28233
0 28235 7 1 2 28222 28234
0 28236 5 1 1 28235
0 28237 7 1 2 66017 28236
0 28238 5 1 1 28237
0 28239 7 1 2 28220 28238
0 28240 7 1 2 28218 28239
0 28241 5 1 1 28240
0 28242 7 1 2 64409 28241
0 28243 5 1 1 28242
0 28244 7 1 2 99795 94318
0 28245 5 1 1 28244
0 28246 7 1 2 79053 91133
0 28247 7 1 2 79609 28246
0 28248 5 1 1 28247
0 28249 7 1 2 28245 28248
0 28250 5 1 1 28249
0 28251 7 1 2 101471 28250
0 28252 5 1 1 28251
0 28253 7 1 2 65115 101287
0 28254 5 1 1 28253
0 28255 7 1 2 66554 101271
0 28256 5 1 1 28255
0 28257 7 1 2 28254 28256
0 28258 5 1 1 28257
0 28259 7 1 2 73741 85325
0 28260 7 1 2 28258 28259
0 28261 5 1 1 28260
0 28262 7 1 2 28252 28261
0 28263 5 1 1 28262
0 28264 7 1 2 100275 28263
0 28265 5 1 1 28264
0 28266 7 3 2 88895 87437
0 28267 7 1 2 1417 101797
0 28268 7 1 2 94651 28267
0 28269 5 1 1 28268
0 28270 7 1 2 28265 28269
0 28271 5 1 1 28270
0 28272 7 1 2 84833 28271
0 28273 5 1 1 28272
0 28274 7 1 2 68067 28273
0 28275 7 1 2 28243 28274
0 28276 7 1 2 28185 28275
0 28277 7 1 2 28141 28276
0 28278 5 1 1 28277
0 28279 7 1 2 97399 75141
0 28280 5 1 1 28279
0 28281 7 1 2 101449 28280
0 28282 5 1 1 28281
0 28283 7 1 2 71828 28282
0 28284 5 1 1 28283
0 28285 7 1 2 92932 27939
0 28286 5 1 1 28285
0 28287 7 1 2 84133 28286
0 28288 5 1 1 28287
0 28289 7 1 2 28284 28288
0 28290 5 1 1 28289
0 28291 7 1 2 68409 28290
0 28292 5 1 1 28291
0 28293 7 1 2 91446 84707
0 28294 7 1 2 101452 28293
0 28295 5 1 1 28294
0 28296 7 1 2 28292 28295
0 28297 5 1 1 28296
0 28298 7 2 2 64410 100192
0 28299 7 1 2 28297 101800
0 28300 5 1 1 28299
0 28301 7 1 2 68410 87080
0 28302 5 1 1 28301
0 28303 7 1 2 28302 83521
0 28304 5 1 1 28303
0 28305 7 1 2 100193 28304
0 28306 5 1 1 28305
0 28307 7 2 2 71829 80099
0 28308 7 1 2 93884 101802
0 28309 5 1 1 28308
0 28310 7 1 2 99430 87566
0 28311 7 1 2 89620 28310
0 28312 5 2 1 28311
0 28313 7 1 2 28309 101804
0 28314 5 1 1 28313
0 28315 7 1 2 100194 28314
0 28316 5 1 1 28315
0 28317 7 1 2 91309 79603
0 28318 5 1 1 28317
0 28319 7 1 2 74854 83623
0 28320 7 1 2 100306 28319
0 28321 5 1 1 28320
0 28322 7 1 2 28318 28321
0 28323 5 1 1 28322
0 28324 7 1 2 81879 28323
0 28325 5 1 1 28324
0 28326 7 2 2 81736 86811
0 28327 7 1 2 100195 101806
0 28328 5 1 1 28327
0 28329 7 3 2 100243 101757
0 28330 7 1 2 101808 93535
0 28331 5 1 1 28330
0 28332 7 1 2 28328 28331
0 28333 7 1 2 28325 28332
0 28334 5 1 1 28333
0 28335 7 1 2 70196 28334
0 28336 5 1 1 28335
0 28337 7 1 2 28316 28336
0 28338 5 1 1 28337
0 28339 7 1 2 69859 28338
0 28340 5 1 1 28339
0 28341 7 1 2 28306 28340
0 28342 5 1 1 28341
0 28343 7 1 2 66297 28342
0 28344 5 1 1 28343
0 28345 7 1 2 99932 97634
0 28346 5 1 1 28345
0 28347 7 1 2 86542 97241
0 28348 5 1 1 28347
0 28349 7 1 2 28346 28348
0 28350 5 1 1 28349
0 28351 7 1 2 94587 28350
0 28352 5 1 1 28351
0 28353 7 1 2 66749 101746
0 28354 5 1 1 28353
0 28355 7 1 2 101752 101809
0 28356 5 1 1 28355
0 28357 7 1 2 28354 28356
0 28358 5 1 1 28357
0 28359 7 1 2 65116 28358
0 28360 5 1 1 28359
0 28361 7 1 2 28352 28360
0 28362 5 1 1 28361
0 28363 7 1 2 69860 28362
0 28364 5 1 1 28363
0 28365 7 1 2 64735 101458
0 28366 5 1 1 28365
0 28367 7 1 2 83425 101447
0 28368 5 1 1 28367
0 28369 7 1 2 28366 28368
0 28370 5 1 1 28369
0 28371 7 1 2 68411 28370
0 28372 5 1 1 28371
0 28373 7 2 2 82113 86320
0 28374 5 2 1 101811
0 28375 7 1 2 101813 12808
0 28376 5 1 1 28375
0 28377 7 1 2 70444 28376
0 28378 5 1 1 28377
0 28379 7 1 2 64736 93776
0 28380 5 1 1 28379
0 28381 7 1 2 82796 15505
0 28382 5 2 1 28381
0 28383 7 1 2 81880 101815
0 28384 5 1 1 28383
0 28385 7 1 2 28380 28384
0 28386 7 1 2 28378 28385
0 28387 7 1 2 28372 28386
0 28388 5 1 1 28387
0 28389 7 1 2 100196 28388
0 28390 5 1 1 28389
0 28391 7 1 2 82010 83624
0 28392 7 1 2 100307 28391
0 28393 7 1 2 87647 28392
0 28394 5 1 1 28393
0 28395 7 1 2 28390 28394
0 28396 7 1 2 28364 28395
0 28397 5 1 1 28396
0 28398 7 1 2 71399 28397
0 28399 5 1 1 28398
0 28400 7 2 2 81881 78029
0 28401 5 1 1 101817
0 28402 7 1 2 101801 101818
0 28403 5 1 1 28402
0 28404 7 1 2 28399 28403
0 28405 7 1 2 28344 28404
0 28406 5 1 1 28405
0 28407 7 1 2 66018 28406
0 28408 5 1 1 28407
0 28409 7 1 2 28300 28408
0 28410 5 1 1 28409
0 28411 7 1 2 85941 28410
0 28412 5 1 1 28411
0 28413 7 2 2 77242 100197
0 28414 7 1 2 79907 101819
0 28415 5 1 1 28414
0 28416 7 2 2 86051 91765
0 28417 5 1 1 101821
0 28418 7 1 2 91748 28417
0 28419 5 1 1 28418
0 28420 7 1 2 101661 28419
0 28421 5 1 1 28420
0 28422 7 1 2 28415 28421
0 28423 5 1 1 28422
0 28424 7 1 2 71400 28423
0 28425 5 1 1 28424
0 28426 7 1 2 101718 101820
0 28427 5 1 1 28426
0 28428 7 1 2 77451 100198
0 28429 5 1 1 28428
0 28430 7 2 2 82923 84508
0 28431 7 2 2 77162 95720
0 28432 7 1 2 101823 101825
0 28433 5 1 1 28432
0 28434 7 1 2 28429 28433
0 28435 5 1 1 28434
0 28436 7 5 2 73494 77949
0 28437 5 1 1 101827
0 28438 7 1 2 28435 101828
0 28439 5 1 1 28438
0 28440 7 1 2 28427 28439
0 28441 5 1 1 28440
0 28442 7 1 2 66298 28441
0 28443 5 1 1 28442
0 28444 7 1 2 87245 87576
0 28445 5 1 1 28444
0 28446 7 1 2 81320 28445
0 28447 5 2 1 28446
0 28448 7 1 2 91789 92070
0 28449 7 1 2 101832 28448
0 28450 5 1 1 28449
0 28451 7 1 2 28443 28450
0 28452 7 1 2 28425 28451
0 28453 5 1 1 28452
0 28454 7 1 2 85326 28453
0 28455 5 1 1 28454
0 28456 7 1 2 73139 28455
0 28457 7 1 2 28412 28456
0 28458 5 1 1 28457
0 28459 7 1 2 28278 28458
0 28460 5 1 1 28459
0 28461 7 2 2 73742 81503
0 28462 7 1 2 100298 101834
0 28463 5 1 1 28462
0 28464 7 1 2 65421 100672
0 28465 5 2 1 28464
0 28466 7 1 2 28463 101836
0 28467 5 1 1 28466
0 28468 7 1 2 66750 28467
0 28469 5 1 1 28468
0 28470 7 1 2 85830 88896
0 28471 7 1 2 87769 28470
0 28472 5 1 1 28471
0 28473 7 1 2 28469 28472
0 28474 5 1 1 28473
0 28475 7 1 2 69861 28474
0 28476 5 1 1 28475
0 28477 7 1 2 27433 28476
0 28478 5 1 1 28477
0 28479 7 1 2 101272 28478
0 28480 5 1 1 28479
0 28481 7 1 2 72677 28480
0 28482 7 1 2 28460 28481
0 28483 5 1 1 28482
0 28484 7 1 2 74808 18240
0 28485 5 1 1 28484
0 28486 7 1 2 65117 28485
0 28487 5 2 1 28486
0 28488 7 1 2 101119 2442
0 28489 5 1 1 28488
0 28490 7 1 2 73495 28489
0 28491 5 1 1 28490
0 28492 7 1 2 101838 28491
0 28493 5 1 1 28492
0 28494 7 1 2 81737 28493
0 28495 5 1 1 28494
0 28496 7 1 2 82599 79345
0 28497 5 1 1 28496
0 28498 7 1 2 64737 28497
0 28499 7 1 2 86032 28498
0 28500 5 1 1 28499
0 28501 7 1 2 28500 85761
0 28502 5 1 1 28501
0 28503 7 1 2 74660 28502
0 28504 5 1 1 28503
0 28505 7 2 2 68412 75608
0 28506 5 1 1 101840
0 28507 7 1 2 28506 2197
0 28508 7 1 2 28504 28507
0 28509 7 1 2 28495 28508
0 28510 5 1 1 28509
0 28511 7 1 2 85327 28510
0 28512 5 1 1 28511
0 28513 7 1 2 90694 101326
0 28514 5 1 1 28513
0 28515 7 1 2 28512 28514
0 28516 5 1 1 28515
0 28517 7 1 2 66299 28516
0 28518 5 1 1 28517
0 28519 7 1 2 66555 77690
0 28520 7 1 2 85590 28519
0 28521 5 1 1 28520
0 28522 7 1 2 101839 28521
0 28523 5 1 1 28522
0 28524 7 1 2 81738 28523
0 28525 5 1 1 28524
0 28526 7 1 2 65422 86228
0 28527 7 1 2 96626 28526
0 28528 5 1 1 28527
0 28529 7 1 2 78697 86229
0 28530 5 1 1 28529
0 28531 7 1 2 70445 28530
0 28532 5 1 1 28531
0 28533 7 1 2 4388 28532
0 28534 7 1 2 28528 28533
0 28535 5 1 1 28534
0 28536 7 1 2 86348 28535
0 28537 5 1 1 28536
0 28538 7 1 2 28525 28537
0 28539 5 1 1 28538
0 28540 7 1 2 93400 28539
0 28541 5 1 1 28540
0 28542 7 1 2 28518 28541
0 28543 5 1 1 28542
0 28544 7 1 2 100276 28543
0 28545 5 1 1 28544
0 28546 7 1 2 100953 94577
0 28547 5 1 1 28546
0 28548 7 2 2 75081 95941
0 28549 7 1 2 83873 91775
0 28550 7 1 2 101842 28549
0 28551 5 1 1 28550
0 28552 7 1 2 28547 28551
0 28553 5 1 1 28552
0 28554 7 1 2 73140 28553
0 28555 5 1 1 28554
0 28556 7 4 2 71940 83221
0 28557 7 2 2 83101 101844
0 28558 7 3 2 84072 90363
0 28559 5 1 1 101850
0 28560 7 1 2 66300 101851
0 28561 7 1 2 101848 28560
0 28562 5 1 1 28561
0 28563 7 1 2 28555 28562
0 28564 5 1 1 28563
0 28565 7 1 2 79839 28564
0 28566 5 1 1 28565
0 28567 7 2 2 85628 83325
0 28568 5 3 1 101853
0 28569 7 1 2 73141 101855
0 28570 5 1 1 28569
0 28571 7 1 2 93289 28570
0 28572 5 1 1 28571
0 28573 7 1 2 85328 28572
0 28574 5 1 1 28573
0 28575 7 1 2 87305 77054
0 28576 5 1 1 28575
0 28577 7 1 2 73496 28576
0 28578 5 1 1 28577
0 28579 7 1 2 86798 28578
0 28580 5 1 1 28579
0 28581 7 1 2 65118 28580
0 28582 5 1 1 28581
0 28583 7 1 2 73142 86177
0 28584 5 1 1 28583
0 28585 7 1 2 70446 28584
0 28586 5 1 1 28585
0 28587 7 1 2 93285 28586
0 28588 5 1 1 28587
0 28589 7 1 2 4519 28588
0 28590 7 1 2 28582 28589
0 28591 5 1 1 28590
0 28592 7 1 2 85942 28591
0 28593 5 1 1 28592
0 28594 7 1 2 28574 28593
0 28595 5 1 1 28594
0 28596 7 1 2 100199 28595
0 28597 5 1 1 28596
0 28598 7 1 2 28566 28597
0 28599 7 1 2 28545 28598
0 28600 5 1 1 28599
0 28601 7 1 2 77346 28600
0 28602 5 1 1 28601
0 28603 7 2 2 95721 78347
0 28604 7 1 2 87318 101858
0 28605 5 1 1 28604
0 28606 7 8 2 66872 80703
0 28607 7 1 2 93585 101860
0 28608 5 1 1 28607
0 28609 7 1 2 28605 28608
0 28610 5 1 1 28609
0 28611 7 1 2 73497 28610
0 28612 5 1 1 28611
0 28613 7 1 2 25185 28612
0 28614 5 1 1 28613
0 28615 7 1 2 85329 28614
0 28616 5 1 1 28615
0 28617 7 1 2 101798 95681
0 28618 7 1 2 101468 28617
0 28619 5 1 1 28618
0 28620 7 1 2 28616 28619
0 28621 5 1 1 28620
0 28622 7 1 2 73143 28621
0 28623 5 1 1 28622
0 28624 7 1 2 63902 85943
0 28625 7 1 2 100057 28624
0 28626 7 4 2 66556 93670
0 28627 7 1 2 95817 101868
0 28628 7 1 2 28625 28627
0 28629 5 1 1 28628
0 28630 7 1 2 28623 28629
0 28631 5 1 1 28630
0 28632 7 1 2 101466 28631
0 28633 5 1 1 28632
0 28634 7 1 2 67649 28633
0 28635 7 1 2 28602 28634
0 28636 5 1 1 28635
0 28637 7 1 2 70812 28636
0 28638 7 1 2 28483 28637
0 28639 5 1 1 28638
0 28640 7 1 2 28096 28639
0 28641 5 1 1 28640
0 28642 7 1 2 64107 28641
0 28643 5 1 1 28642
0 28644 7 1 2 100549 25021
0 28645 5 1 1 28644
0 28646 7 1 2 73498 28645
0 28647 5 1 1 28646
0 28648 7 1 2 100449 28647
0 28649 5 1 1 28648
0 28650 7 1 2 70813 28649
0 28651 5 1 1 28650
0 28652 7 1 2 69166 100839
0 28653 5 1 1 28652
0 28654 7 1 2 28651 28653
0 28655 5 1 1 28654
0 28656 7 1 2 100200 28655
0 28657 5 1 1 28656
0 28658 7 3 2 93731 96395
0 28659 7 1 2 89606 91388
0 28660 7 1 2 101872 28659
0 28661 5 1 1 28660
0 28662 7 1 2 28657 28661
0 28663 5 1 1 28662
0 28664 7 1 2 99220 82528
0 28665 7 1 2 95475 28664
0 28666 7 1 2 28663 28665
0 28667 5 1 1 28666
0 28668 7 1 2 28643 28667
0 28669 5 1 1 28668
0 28670 7 1 2 72386 28669
0 28671 5 1 1 28670
0 28672 7 1 2 96992 98447
0 28673 5 2 1 28672
0 28674 7 1 2 100201 101875
0 28675 7 1 2 93404 28674
0 28676 5 1 1 28675
0 28677 7 1 2 72056 100341
0 28678 7 1 2 96264 28677
0 28679 7 3 2 71941 87866
0 28680 7 1 2 95676 101877
0 28681 7 1 2 28678 28680
0 28682 5 1 1 28681
0 28683 7 1 2 28676 28682
0 28684 5 1 1 28683
0 28685 7 1 2 77347 28684
0 28686 5 1 1 28685
0 28687 7 2 2 97102 93771
0 28688 7 1 2 88905 81122
0 28689 7 1 2 101880 28688
0 28690 5 1 1 28689
0 28691 7 1 2 28686 28690
0 28692 5 1 1 28691
0 28693 7 1 2 84553 28692
0 28694 5 1 1 28693
0 28695 7 1 2 100342 91879
0 28696 7 1 2 74472 28695
0 28697 7 1 2 100231 98603
0 28698 7 1 2 28696 28697
0 28699 5 1 1 28698
0 28700 7 2 2 73499 91070
0 28701 7 1 2 101876 101882
0 28702 7 1 2 101789 28701
0 28703 5 1 1 28702
0 28704 7 1 2 28699 28703
0 28705 5 1 1 28704
0 28706 7 1 2 77348 28705
0 28707 5 1 1 28706
0 28708 7 1 2 71091 77670
0 28709 7 1 2 92436 28708
0 28710 7 1 2 101881 28709
0 28711 5 1 1 28710
0 28712 7 1 2 28707 28711
0 28713 5 1 1 28712
0 28714 7 1 2 97400 28713
0 28715 5 1 1 28714
0 28716 7 1 2 28694 28715
0 28717 5 1 1 28716
0 28718 7 1 2 65423 28717
0 28719 5 1 1 28718
0 28720 7 1 2 79889 101590
0 28721 5 1 1 28720
0 28722 7 1 2 76078 28721
0 28723 5 1 1 28722
0 28724 7 1 2 79410 79299
0 28725 5 2 1 28724
0 28726 7 2 2 70447 75058
0 28727 5 2 1 101886
0 28728 7 1 2 78741 101887
0 28729 5 1 1 28728
0 28730 7 1 2 101884 28729
0 28731 7 1 2 28723 28730
0 28732 5 1 1 28731
0 28733 7 1 2 77243 28732
0 28734 5 1 1 28733
0 28735 7 2 2 78653 81156
0 28736 7 1 2 71092 101890
0 28737 5 1 1 28736
0 28738 7 1 2 66019 101593
0 28739 5 1 1 28738
0 28740 7 1 2 64108 28739
0 28741 7 1 2 28737 28740
0 28742 7 1 2 28734 28741
0 28743 5 1 1 28742
0 28744 7 2 2 64411 82529
0 28745 7 1 2 101892 93282
0 28746 5 1 1 28745
0 28747 7 1 2 69167 28746
0 28748 5 1 1 28747
0 28749 7 1 2 98423 76392
0 28750 7 1 2 100954 28749
0 28751 7 1 2 28748 28750
0 28752 7 1 2 28743 28751
0 28753 5 1 1 28752
0 28754 7 1 2 28719 28753
0 28755 5 1 1 28754
0 28756 7 1 2 72678 28755
0 28757 5 1 1 28756
0 28758 7 1 2 79088 79638
0 28759 7 1 2 101186 28758
0 28760 5 1 1 28759
0 28761 7 1 2 76806 100343
0 28762 7 1 2 87911 28761
0 28763 7 1 2 93416 28762
0 28764 5 1 1 28763
0 28765 7 1 2 28760 28764
0 28766 5 1 1 28765
0 28767 7 1 2 101251 28766
0 28768 5 1 1 28767
0 28769 7 2 2 70632 100344
0 28770 7 2 2 78356 101894
0 28771 7 1 2 90950 91980
0 28772 7 1 2 101896 28771
0 28773 5 1 1 28772
0 28774 7 1 2 89276 90671
0 28775 7 1 2 100651 28774
0 28776 5 1 1 28775
0 28777 7 1 2 28773 28776
0 28778 7 1 2 28768 28777
0 28779 5 1 1 28778
0 28780 7 1 2 65424 28779
0 28781 5 1 1 28780
0 28782 7 1 2 68856 73500
0 28783 7 1 2 87912 28782
0 28784 7 1 2 95739 28783
0 28785 7 1 2 101897 28784
0 28786 5 1 1 28785
0 28787 7 1 2 28781 28786
0 28788 5 1 1 28787
0 28789 7 1 2 66020 28788
0 28790 5 1 1 28789
0 28791 7 3 2 68857 89631
0 28792 7 2 2 100964 101898
0 28793 7 1 2 79870 87945
0 28794 7 1 2 101901 28793
0 28795 5 1 1 28794
0 28796 7 1 2 28790 28795
0 28797 5 1 1 28796
0 28798 7 1 2 64412 28797
0 28799 5 1 1 28798
0 28800 7 1 2 93283 86858
0 28801 7 1 2 101902 28800
0 28802 5 1 1 28801
0 28803 7 1 2 28799 28802
0 28804 5 1 1 28803
0 28805 7 1 2 97009 28804
0 28806 5 1 1 28805
0 28807 7 1 2 28757 28806
0 28808 5 1 1 28807
0 28809 7 1 2 90482 28808
0 28810 5 1 1 28809
0 28811 7 1 2 5979 27635
0 28812 5 1 1 28811
0 28813 7 1 2 73501 94836
0 28814 7 1 2 28812 28813
0 28815 5 1 1 28814
0 28816 7 1 2 100557 93395
0 28817 5 1 1 28816
0 28818 7 1 2 28815 28817
0 28819 5 1 1 28818
0 28820 7 1 2 64738 28819
0 28821 5 1 1 28820
0 28822 7 2 2 65425 94837
0 28823 7 1 2 89154 89927
0 28824 7 1 2 101903 28823
0 28825 7 1 2 90194 28824
0 28826 5 1 1 28825
0 28827 7 1 2 28821 28826
0 28828 5 1 1 28827
0 28829 7 1 2 100202 28828
0 28830 5 1 1 28829
0 28831 7 1 2 70682 101601
0 28832 7 2 2 63799 96547
0 28833 7 1 2 96015 94995
0 28834 7 1 2 101905 28833
0 28835 7 1 2 28831 28834
0 28836 5 1 1 28835
0 28837 7 1 2 28830 28836
0 28838 5 1 1 28837
0 28839 7 2 2 66301 96744
0 28840 7 1 2 101550 101907
0 28841 7 1 2 28838 28840
0 28842 5 1 1 28841
0 28843 7 1 2 28810 28842
0 28844 7 1 2 28671 28843
0 28845 5 1 1 28844
0 28846 7 1 2 72225 28845
0 28847 5 1 1 28846
0 28848 7 2 2 77163 100454
0 28849 5 1 1 101909
0 28850 7 1 2 69862 28849
0 28851 5 1 1 28850
0 28852 7 1 2 64739 101512
0 28853 5 1 1 28852
0 28854 7 1 2 75918 28853
0 28855 7 1 2 28851 28854
0 28856 5 1 1 28855
0 28857 7 1 2 90919 101910
0 28858 5 2 1 28857
0 28859 7 1 2 87052 84354
0 28860 5 1 1 28859
0 28861 7 1 2 76079 98341
0 28862 5 1 1 28861
0 28863 7 1 2 28860 28862
0 28864 7 1 2 101911 28863
0 28865 7 1 2 28856 28864
0 28866 5 1 1 28865
0 28867 7 1 2 98691 28866
0 28868 5 1 1 28867
0 28869 7 3 2 76589 97039
0 28870 5 1 1 101913
0 28871 7 1 2 67311 89264
0 28872 5 1 1 28871
0 28873 7 1 2 28870 28872
0 28874 5 3 1 28873
0 28875 7 1 2 69168 101916
0 28876 5 1 1 28875
0 28877 7 1 2 69863 101179
0 28878 5 3 1 28877
0 28879 7 5 2 90881 90036
0 28880 7 1 2 96745 101922
0 28881 5 1 1 28880
0 28882 7 1 2 101919 28881
0 28883 5 1 1 28882
0 28884 7 1 2 100541 28883
0 28885 5 2 1 28884
0 28886 7 1 2 28876 101927
0 28887 5 1 1 28886
0 28888 7 1 2 66021 28887
0 28889 5 1 1 28888
0 28890 7 1 2 69169 98692
0 28891 7 1 2 81572 28890
0 28892 5 1 1 28891
0 28893 7 1 2 28889 28892
0 28894 5 1 1 28893
0 28895 7 1 2 64413 28894
0 28896 5 1 1 28895
0 28897 7 1 2 28868 28896
0 28898 5 1 1 28897
0 28899 7 1 2 65799 28898
0 28900 5 1 1 28899
0 28901 7 1 2 76080 100542
0 28902 5 1 1 28901
0 28903 7 1 2 3291 28902
0 28904 5 1 1 28903
0 28905 7 1 2 64740 28904
0 28906 5 1 1 28905
0 28907 7 1 2 86649 91114
0 28908 5 1 1 28907
0 28909 7 1 2 28906 28908
0 28910 5 1 1 28909
0 28911 7 1 2 28910 98718
0 28912 5 1 1 28911
0 28913 7 1 2 28900 28912
0 28914 5 1 1 28913
0 28915 7 1 2 72226 28914
0 28916 5 1 1 28915
0 28917 7 1 2 93087 97120
0 28918 5 6 1 28917
0 28919 7 1 2 101180 101929
0 28920 5 11 1 28919
0 28921 7 1 2 69864 101935
0 28922 5 2 1 28921
0 28923 7 1 2 93660 92535
0 28924 5 1 1 28923
0 28925 7 1 2 72679 27292
0 28926 7 1 2 90922 28925
0 28927 5 1 1 28926
0 28928 7 1 2 67312 28927
0 28929 7 1 2 28924 28928
0 28930 5 1 1 28929
0 28931 7 1 2 101946 28930
0 28932 5 1 1 28931
0 28933 7 1 2 100543 28932
0 28934 5 1 1 28933
0 28935 7 1 2 101164 78149
0 28936 5 1 1 28935
0 28937 7 1 2 64741 2036
0 28938 7 1 2 93469 28937
0 28939 5 1 1 28938
0 28940 7 1 2 10436 28939
0 28941 5 1 1 28940
0 28942 7 1 2 77244 28941
0 28943 5 1 1 28942
0 28944 7 2 2 77554 93516
0 28945 5 2 1 101948
0 28946 7 1 2 90874 92965
0 28947 5 1 1 28946
0 28948 7 1 2 101950 28947
0 28949 7 1 2 28943 28948
0 28950 5 1 1 28949
0 28951 7 1 2 67313 28950
0 28952 5 1 1 28951
0 28953 7 1 2 28936 28952
0 28954 7 1 2 28934 28953
0 28955 5 1 1 28954
0 28956 7 1 2 72227 28955
0 28957 5 1 1 28956
0 28958 7 1 2 76323 100457
0 28959 5 1 1 28958
0 28960 7 3 2 100576 98111
0 28961 7 1 2 99792 101952
0 28962 7 1 2 28959 28961
0 28963 5 1 1 28962
0 28964 7 1 2 28957 28963
0 28965 5 1 1 28964
0 28966 7 1 2 65800 28965
0 28967 5 1 1 28966
0 28968 7 1 2 70814 101917
0 28969 5 1 1 28968
0 28970 7 1 2 101928 28969
0 28971 5 1 1 28970
0 28972 7 1 2 66022 28971
0 28973 5 1 1 28972
0 28974 7 1 2 81573 98451
0 28975 5 1 1 28974
0 28976 7 1 2 28973 28975
0 28977 5 1 1 28976
0 28978 7 1 2 64414 28977
0 28979 5 1 1 28978
0 28980 7 3 2 64742 95335
0 28981 5 1 1 101955
0 28982 7 1 2 100544 80833
0 28983 5 1 1 28982
0 28984 7 1 2 115 28983
0 28985 5 1 1 28984
0 28986 7 1 2 69533 28985
0 28987 5 1 1 28986
0 28988 7 1 2 28981 28987
0 28989 5 1 1 28988
0 28990 7 1 2 75919 28989
0 28991 5 1 1 28990
0 28992 7 1 2 81574 77065
0 28993 5 1 1 28992
0 28994 7 1 2 101912 28993
0 28995 7 1 2 28991 28994
0 28996 5 1 1 28995
0 28997 7 1 2 98693 28996
0 28998 5 1 1 28997
0 28999 7 1 2 28979 28998
0 29000 5 1 1 28999
0 29001 7 1 2 72228 29000
0 29002 5 1 1 29001
0 29003 7 1 2 28967 29002
0 29004 5 1 1 29003
0 29005 7 1 2 64109 29004
0 29006 5 1 1 29005
0 29007 7 1 2 28916 29006
0 29008 5 1 1 29007
0 29009 7 1 2 65426 29008
0 29010 5 1 1 29009
0 29011 7 1 2 77245 81575
0 29012 5 1 1 29011
0 29013 7 1 2 90875 77452
0 29014 5 1 1 29013
0 29015 7 1 2 29012 29014
0 29016 5 1 1 29015
0 29017 7 1 2 85504 29016
0 29018 5 1 1 29017
0 29019 7 1 2 77561 100497
0 29020 5 1 1 29019
0 29021 7 1 2 29018 29020
0 29022 5 1 1 29021
0 29023 7 4 2 66751 72229
0 29024 7 1 2 29022 101958
0 29025 5 1 1 29024
0 29026 7 1 2 67173 93972
0 29027 7 1 2 96235 93423
0 29028 7 1 2 29026 29027
0 29029 5 1 1 29028
0 29030 7 1 2 29025 29029
0 29031 5 1 1 29030
0 29032 7 1 2 72680 29031
0 29033 5 1 1 29032
0 29034 7 1 2 85505 77349
0 29035 5 3 1 29034
0 29036 7 1 2 68068 85397
0 29037 5 1 1 29036
0 29038 7 1 2 101962 29037
0 29039 5 1 1 29038
0 29040 7 1 2 78150 101959
0 29041 7 1 2 29039 29040
0 29042 5 1 1 29041
0 29043 7 1 2 29033 29042
0 29044 5 1 1 29043
0 29045 7 1 2 72387 29044
0 29046 5 1 1 29045
0 29047 7 1 2 101963 3302
0 29048 5 1 1 29047
0 29049 7 2 2 73144 101960
0 29050 7 3 2 76224 96746
0 29051 5 1 1 101967
0 29052 7 1 2 101965 101968
0 29053 7 1 2 29048 29052
0 29054 5 1 1 29053
0 29055 7 1 2 29046 29054
0 29056 7 1 2 29010 29055
0 29057 5 1 1 29056
0 29058 7 1 2 100203 29057
0 29059 5 1 1 29058
0 29060 7 2 2 99770 98519
0 29061 5 1 1 101970
0 29062 7 1 2 98334 101971
0 29063 5 1 1 29062
0 29064 7 3 2 64110 80198
0 29065 7 1 2 100785 101972
0 29066 5 1 1 29065
0 29067 7 1 2 29063 29066
0 29068 5 1 1 29067
0 29069 7 1 2 79963 29068
0 29070 5 1 1 29069
0 29071 7 1 2 78822 101454
0 29072 5 1 1 29071
0 29073 7 1 2 81670 29072
0 29074 5 1 1 29073
0 29075 7 1 2 99638 101707
0 29076 7 1 2 29074 29075
0 29077 5 1 1 29076
0 29078 7 1 2 29070 29077
0 29079 5 1 1 29078
0 29080 7 1 2 67650 29079
0 29081 5 1 1 29080
0 29082 7 6 2 64111 93257
0 29083 7 1 2 100787 101975
0 29084 5 1 1 29083
0 29085 7 1 2 99771 98740
0 29086 5 1 1 29085
0 29087 7 1 2 29084 29086
0 29088 5 1 1 29087
0 29089 7 1 2 65119 29088
0 29090 5 1 1 29089
0 29091 7 2 2 96958 75104
0 29092 7 1 2 77350 80199
0 29093 7 1 2 101981 29092
0 29094 5 1 1 29093
0 29095 7 1 2 29090 29094
0 29096 5 1 1 29095
0 29097 7 1 2 86715 29096
0 29098 5 1 1 29097
0 29099 7 1 2 29081 29098
0 29100 5 1 1 29099
0 29101 7 4 2 71942 72230
0 29102 7 1 2 95722 101983
0 29103 7 1 2 29100 29102
0 29104 5 1 1 29103
0 29105 7 1 2 29059 29104
0 29106 5 1 1 29105
0 29107 7 1 2 85330 29106
0 29108 5 1 1 29107
0 29109 7 1 2 93258 88350
0 29110 7 1 2 100299 29109
0 29111 7 1 2 85064 29110
0 29112 5 1 1 29111
0 29113 7 1 2 65801 101949
0 29114 5 1 1 29113
0 29115 7 1 2 64415 10519
0 29116 5 1 1 29115
0 29117 7 1 2 29116 78452
0 29118 5 1 1 29117
0 29119 7 1 2 81157 98865
0 29120 7 1 2 29118 29119
0 29121 5 1 1 29120
0 29122 7 1 2 29114 29121
0 29123 5 1 1 29122
0 29124 7 4 2 72057 74000
0 29125 7 1 2 101624 101987
0 29126 7 1 2 29123 29125
0 29127 5 1 1 29126
0 29128 7 1 2 29112 29127
0 29129 5 1 1 29128
0 29130 7 1 2 67314 29129
0 29131 5 1 1 29130
0 29132 7 1 2 70683 74006
0 29133 7 1 2 75710 29132
0 29134 7 1 2 95232 29133
0 29135 5 1 1 29134
0 29136 7 1 2 101837 29135
0 29137 5 1 1 29136
0 29138 7 2 2 101914 29137
0 29139 5 1 1 101991
0 29140 7 1 2 101992 98705
0 29141 5 1 1 29140
0 29142 7 1 2 29131 29141
0 29143 5 1 1 29142
0 29144 7 1 2 64112 29143
0 29145 5 1 1 29144
0 29146 7 1 2 95818 101899
0 29147 7 3 2 72058 93068
0 29148 7 1 2 101993 97146
0 29149 7 1 2 29146 29148
0 29150 5 1 1 29149
0 29151 7 1 2 29139 29150
0 29152 5 1 1 29151
0 29153 7 1 2 98730 29152
0 29154 5 1 1 29153
0 29155 7 1 2 29145 29154
0 29156 5 1 1 29155
0 29157 7 1 2 72231 29156
0 29158 5 1 1 29157
0 29159 7 1 2 73145 87747
0 29160 7 1 2 100967 29159
0 29161 7 6 2 67174 98694
0 29162 7 4 2 74390 77351
0 29163 7 1 2 101994 102002
0 29164 7 1 2 101996 29163
0 29165 7 1 2 29160 29164
0 29166 5 1 1 29165
0 29167 7 1 2 29158 29166
0 29168 5 1 1 29167
0 29169 7 1 2 90483 29168
0 29170 5 1 1 29169
0 29171 7 2 2 68858 101570
0 29172 7 1 2 65427 76046
0 29173 5 2 1 29172
0 29174 7 2 2 76040 102008
0 29175 5 1 1 102010
0 29176 7 1 2 67651 100277
0 29177 7 1 2 29175 29176
0 29178 7 1 2 98741 29177
0 29179 5 1 1 29178
0 29180 7 1 2 69170 96127
0 29181 5 1 1 29180
0 29182 7 5 2 85845 93586
0 29183 7 2 2 64113 14505
0 29184 5 1 1 102017
0 29185 7 1 2 29184 93088
0 29186 7 1 2 102012 29185
0 29187 7 1 2 29181 29186
0 29188 5 1 1 29187
0 29189 7 1 2 29179 29188
0 29190 5 1 1 29189
0 29191 7 1 2 64743 29190
0 29192 5 1 1 29191
0 29193 7 2 2 93001 98742
0 29194 7 1 2 96411 79043
0 29195 7 1 2 102019 29194
0 29196 5 1 1 29195
0 29197 7 1 2 29192 29196
0 29198 5 1 1 29197
0 29199 7 1 2 72388 29198
0 29200 5 1 1 29199
0 29201 7 2 2 77570 85057
0 29202 5 1 1 102021
0 29203 7 1 2 91329 29202
0 29204 5 1 1 29203
0 29205 7 2 2 67315 29204
0 29206 7 4 2 70684 65802
0 29207 7 2 2 84321 102025
0 29208 7 1 2 79518 87962
0 29209 7 1 2 102029 29208
0 29210 7 1 2 102023 29209
0 29211 5 1 1 29210
0 29212 7 1 2 29200 29211
0 29213 5 1 1 29212
0 29214 7 1 2 65120 29213
0 29215 5 1 1 29214
0 29216 7 1 2 64416 101125
0 29217 5 1 1 29216
0 29218 7 2 2 66023 79411
0 29219 5 1 1 102031
0 29220 7 1 2 71401 29219
0 29221 7 1 2 29217 29220
0 29222 5 1 1 29221
0 29223 7 1 2 83854 99326
0 29224 7 1 2 96526 29223
0 29225 7 1 2 89947 29224
0 29226 7 1 2 100412 29225
0 29227 7 1 2 29222 29226
0 29228 5 1 1 29227
0 29229 7 1 2 29215 29228
0 29230 5 1 1 29229
0 29231 7 1 2 82924 29230
0 29232 5 1 1 29231
0 29233 7 2 2 80357 83967
0 29234 5 3 1 102033
0 29235 7 5 2 66302 98023
0 29236 7 2 2 78480 102038
0 29237 5 1 1 102043
0 29238 7 1 2 97734 93182
0 29239 5 1 1 29238
0 29240 7 1 2 29237 29239
0 29241 5 1 1 29240
0 29242 7 1 2 102034 29241
0 29243 5 1 1 29242
0 29244 7 2 2 87055 99853
0 29245 5 1 1 102045
0 29246 7 1 2 90923 102046
0 29247 5 1 1 29246
0 29248 7 1 2 96747 29247
0 29249 5 1 1 29248
0 29250 7 1 2 101920 29249
0 29251 5 1 1 29250
0 29252 7 1 2 86674 29251
0 29253 5 1 1 29252
0 29254 7 1 2 99103 98756
0 29255 5 1 1 29254
0 29256 7 1 2 29253 29255
0 29257 5 1 1 29256
0 29258 7 1 2 64417 29257
0 29259 5 1 1 29258
0 29260 7 1 2 29243 29259
0 29261 5 1 1 29260
0 29262 7 1 2 74391 29261
0 29263 5 1 1 29262
0 29264 7 11 2 67652 85506
0 29265 7 2 2 64418 102047
0 29266 5 1 1 102058
0 29267 7 1 2 90037 98457
0 29268 7 1 2 102059 29267
0 29269 5 1 1 29268
0 29270 7 1 2 29263 29269
0 29271 5 1 1 29270
0 29272 7 1 2 100204 29271
0 29273 5 1 1 29272
0 29274 7 1 2 29232 29273
0 29275 5 1 1 29274
0 29276 7 1 2 102006 29275
0 29277 5 1 1 29276
0 29278 7 1 2 29170 29277
0 29279 7 1 2 29108 29278
0 29280 5 1 1 29279
0 29281 7 1 2 73964 29280
0 29282 5 1 1 29281
0 29283 7 1 2 85364 12210
0 29284 5 2 1 29283
0 29285 7 1 2 73146 102060
0 29286 5 1 1 29285
0 29287 7 1 2 12322 29286
0 29288 5 1 1 29287
0 29289 7 1 2 82195 29288
0 29290 5 1 1 29289
0 29291 7 1 2 96539 95063
0 29292 5 1 1 29291
0 29293 7 1 2 29290 29292
0 29294 5 1 1 29293
0 29295 7 1 2 64744 29294
0 29296 5 1 1 29295
0 29297 7 1 2 82049 100895
0 29298 5 1 1 29297
0 29299 7 2 2 76081 101387
0 29300 5 1 1 102062
0 29301 7 1 2 85944 102063
0 29302 5 1 1 29301
0 29303 7 1 2 29298 29302
0 29304 5 1 1 29303
0 29305 7 1 2 72681 29304
0 29306 5 1 1 29305
0 29307 7 1 2 29296 29306
0 29308 5 1 1 29307
0 29309 7 1 2 73502 29308
0 29310 5 1 1 29309
0 29311 7 2 2 100875 81963
0 29312 5 1 1 102064
0 29313 7 1 2 99997 102065
0 29314 5 1 1 29313
0 29315 7 1 2 3236 92640
0 29316 5 1 1 29315
0 29317 7 1 2 86006 29316
0 29318 5 1 1 29317
0 29319 7 3 2 75578 93119
0 29320 7 1 2 70448 98674
0 29321 7 1 2 102066 29320
0 29322 5 1 1 29321
0 29323 7 1 2 29318 29322
0 29324 5 1 1 29323
0 29325 7 1 2 76590 29324
0 29326 5 1 1 29325
0 29327 7 1 2 29314 29326
0 29328 7 1 2 29310 29327
0 29329 5 1 1 29328
0 29330 7 1 2 64419 29329
0 29331 5 1 1 29330
0 29332 7 4 2 72682 78654
0 29333 7 1 2 93417 81123
0 29334 5 1 1 29333
0 29335 7 1 2 84574 100227
0 29336 5 1 1 29335
0 29337 7 1 2 29334 29336
0 29338 5 1 1 29337
0 29339 7 1 2 102069 29338
0 29340 5 1 1 29339
0 29341 7 1 2 29331 29340
0 29342 5 1 1 29341
0 29343 7 1 2 100205 29342
0 29344 5 1 1 29343
0 29345 7 1 2 67316 29344
0 29346 5 1 1 29345
0 29347 7 1 2 65121 75579
0 29348 7 2 2 84134 29347
0 29349 5 1 1 102073
0 29350 7 1 2 82062 29349
0 29351 5 1 1 29350
0 29352 7 1 2 76591 29351
0 29353 5 1 1 29352
0 29354 7 1 2 69865 102011
0 29355 5 1 1 29354
0 29356 7 1 2 79995 87231
0 29357 7 1 2 29355 29356
0 29358 5 1 1 29357
0 29359 7 1 2 29353 29358
0 29360 5 1 1 29359
0 29361 7 1 2 100206 29360
0 29362 5 1 1 29361
0 29363 7 1 2 66303 75647
0 29364 5 1 1 29363
0 29365 7 1 2 78966 29364
0 29366 5 1 1 29365
0 29367 7 2 2 64745 29366
0 29368 5 1 1 102075
0 29369 7 1 2 92926 87013
0 29370 5 1 1 29369
0 29371 7 1 2 29368 29370
0 29372 5 1 1 29371
0 29373 7 1 2 79925 101859
0 29374 7 1 2 29372 29373
0 29375 5 1 1 29374
0 29376 7 1 2 29362 29375
0 29377 5 1 1 29376
0 29378 7 1 2 67653 29377
0 29379 5 1 1 29378
0 29380 7 1 2 91389 95499
0 29381 7 1 2 91596 82157
0 29382 7 1 2 29380 29381
0 29383 5 1 1 29382
0 29384 7 1 2 29379 29383
0 29385 5 1 1 29384
0 29386 7 1 2 71093 29385
0 29387 5 1 1 29386
0 29388 7 1 2 70449 95384
0 29389 7 3 2 76919 100878
0 29390 7 2 2 66873 83847
0 29391 7 1 2 102077 102080
0 29392 7 1 2 29388 29391
0 29393 5 1 1 29392
0 29394 7 1 2 29387 29393
0 29395 5 1 1 29394
0 29396 7 1 2 85945 29395
0 29397 5 1 1 29396
0 29398 7 2 2 68069 93661
0 29399 7 2 2 64746 76393
0 29400 7 1 2 79068 100955
0 29401 7 1 2 102084 29400
0 29402 7 1 2 102082 29401
0 29403 5 1 1 29402
0 29404 7 1 2 79026 88028
0 29405 7 1 2 92580 29404
0 29406 7 1 2 99075 29405
0 29407 5 1 1 29406
0 29408 7 1 2 29403 29407
0 29409 5 1 1 29408
0 29410 7 1 2 75397 29409
0 29411 5 1 1 29410
0 29412 7 1 2 66557 84420
0 29413 7 1 2 91348 29412
0 29414 7 1 2 81646 84580
0 29415 7 1 2 29413 29414
0 29416 5 1 1 29415
0 29417 7 1 2 72389 29416
0 29418 7 1 2 29411 29417
0 29419 7 1 2 29397 29418
0 29420 5 1 1 29419
0 29421 7 1 2 65803 29420
0 29422 7 1 2 29346 29421
0 29423 5 1 1 29422
0 29424 7 2 2 93401 98265
0 29425 5 1 1 102086
0 29426 7 1 2 65122 102087
0 29427 5 1 1 29426
0 29428 7 2 2 77246 98137
0 29429 7 1 2 70815 74661
0 29430 7 1 2 100944 29429
0 29431 7 1 2 102088 29430
0 29432 5 1 1 29431
0 29433 7 1 2 29427 29432
0 29434 5 1 1 29433
0 29435 7 1 2 76082 29434
0 29436 5 1 1 29435
0 29437 7 4 2 66304 77872
0 29438 7 2 2 69866 98256
0 29439 5 1 1 102094
0 29440 7 1 2 93396 102095
0 29441 5 1 1 29440
0 29442 7 4 2 65428 72390
0 29443 7 2 2 71094 102096
0 29444 5 1 1 102100
0 29445 7 1 2 98284 29444
0 29446 5 1 1 29445
0 29447 7 1 2 93596 77029
0 29448 7 1 2 29446 29447
0 29449 5 1 1 29448
0 29450 7 1 2 29441 29449
0 29451 5 1 1 29450
0 29452 7 1 2 102090 29451
0 29453 5 1 1 29452
0 29454 7 2 2 77247 98024
0 29455 7 2 2 90506 102102
0 29456 7 2 2 74662 74331
0 29457 7 1 2 91804 102106
0 29458 7 1 2 102104 29457
0 29459 5 1 1 29458
0 29460 7 1 2 29453 29459
0 29461 7 1 2 29436 29460
0 29462 5 1 1 29461
0 29463 7 1 2 72683 29462
0 29464 5 1 1 29463
0 29465 7 2 2 64420 91447
0 29466 7 1 2 98685 91508
0 29467 7 1 2 102108 29466
0 29468 5 2 1 29467
0 29469 7 1 2 80259 80317
0 29470 5 1 1 29469
0 29471 7 1 2 73147 93932
0 29472 7 1 2 93235 29471
0 29473 5 1 1 29472
0 29474 7 1 2 29470 29473
0 29475 5 1 1 29474
0 29476 7 2 2 72059 29475
0 29477 7 1 2 93597 102112
0 29478 5 1 1 29477
0 29479 7 1 2 102110 29478
0 29480 5 1 1 29479
0 29481 7 1 2 97040 29480
0 29482 5 1 1 29481
0 29483 7 1 2 29464 29482
0 29484 5 1 1 29483
0 29485 7 1 2 100207 29484
0 29486 5 1 1 29485
0 29487 7 1 2 85946 78930
0 29488 5 1 1 29487
0 29489 7 1 2 65429 90725
0 29490 5 1 1 29489
0 29491 7 1 2 29488 29490
0 29492 5 1 1 29491
0 29493 7 1 2 81964 29492
0 29494 5 1 1 29493
0 29495 7 1 2 102091 98787
0 29496 5 1 1 29495
0 29497 7 1 2 29494 29496
0 29498 5 1 1 29497
0 29499 7 1 2 69867 29498
0 29500 5 1 1 29499
0 29501 7 1 2 85947 92265
0 29502 7 1 2 102076 29501
0 29503 5 1 1 29502
0 29504 7 1 2 29500 29503
0 29505 5 1 1 29504
0 29506 7 1 2 72391 29505
0 29507 5 1 1 29506
0 29508 7 1 2 90850 97121
0 29509 7 1 2 96011 29508
0 29510 5 1 1 29509
0 29511 7 1 2 29507 29510
0 29512 5 2 1 29511
0 29513 7 1 2 77352 102114
0 29514 5 1 1 29513
0 29515 7 2 2 95609 98357
0 29516 7 1 2 87314 94405
0 29517 7 1 2 102116 29516
0 29518 5 1 1 29517
0 29519 7 1 2 29514 29518
0 29520 5 1 1 29519
0 29521 7 1 2 100394 29520
0 29522 5 1 1 29521
0 29523 7 1 2 29486 29522
0 29524 5 1 1 29523
0 29525 7 1 2 73503 29524
0 29526 5 1 1 29525
0 29527 7 4 2 72060 97041
0 29528 7 2 2 91349 102118
0 29529 7 2 2 76225 87748
0 29530 7 1 2 98706 102124
0 29531 7 1 2 102122 29530
0 29532 5 1 1 29531
0 29533 7 1 2 29526 29532
0 29534 7 1 2 29423 29533
0 29535 5 1 1 29534
0 29536 7 1 2 72232 29535
0 29537 5 1 1 29536
0 29538 7 1 2 100079 90043
0 29539 5 1 1 29538
0 29540 7 6 2 72392 73504
0 29541 7 6 2 67175 73148
0 29542 7 1 2 102126 102132
0 29543 7 1 2 88323 29542
0 29544 5 2 1 29543
0 29545 7 1 2 29539 102138
0 29546 5 1 1 29545
0 29547 7 1 2 85948 29546
0 29548 5 1 1 29547
0 29549 7 1 2 87014 79880
0 29550 5 1 1 29549
0 29551 7 1 2 65430 82227
0 29552 5 1 1 29551
0 29553 7 1 2 29550 29552
0 29554 5 1 1 29553
0 29555 7 1 2 64747 29554
0 29556 5 1 1 29555
0 29557 7 1 2 77671 89813
0 29558 5 2 1 29557
0 29559 7 1 2 29556 102140
0 29560 5 1 1 29559
0 29561 7 1 2 67176 99705
0 29562 7 1 2 29560 29561
0 29563 5 1 1 29562
0 29564 7 1 2 29548 29563
0 29565 5 1 1 29564
0 29566 7 1 2 64421 29565
0 29567 5 1 1 29566
0 29568 7 3 2 97401 75398
0 29569 5 1 1 102142
0 29570 7 2 2 78790 79507
0 29571 5 1 1 102145
0 29572 7 1 2 29569 29571
0 29573 5 4 1 29572
0 29574 7 1 2 70450 102147
0 29575 5 1 1 29574
0 29576 7 1 2 74663 100681
0 29577 5 1 1 29576
0 29578 7 1 2 29575 29577
0 29579 5 1 1 29578
0 29580 7 1 2 85949 29579
0 29581 5 1 1 29580
0 29582 7 1 2 94566 83222
0 29583 5 1 1 29582
0 29584 7 1 2 73149 29583
0 29585 7 1 2 29581 29584
0 29586 5 1 1 29585
0 29587 7 1 2 68413 93343
0 29588 5 1 1 29587
0 29589 7 2 2 5102 29588
0 29590 5 1 1 102151
0 29591 7 1 2 70451 29590
0 29592 5 1 1 29591
0 29593 7 1 2 74664 101472
0 29594 5 1 1 29593
0 29595 7 1 2 29592 29594
0 29596 5 1 1 29595
0 29597 7 1 2 85950 29596
0 29598 5 1 1 29597
0 29599 7 1 2 86007 95429
0 29600 5 1 1 29599
0 29601 7 1 2 68070 29600
0 29602 7 1 2 29598 29601
0 29603 5 1 1 29602
0 29604 7 1 2 100080 29603
0 29605 7 1 2 29586 29604
0 29606 5 1 1 29605
0 29607 7 1 2 29567 29606
0 29608 5 1 1 29607
0 29609 7 1 2 100208 29608
0 29610 5 1 1 29609
0 29611 7 2 2 85951 100081
0 29612 7 1 2 77538 102153
0 29613 5 1 1 29612
0 29614 7 1 2 97103 102133
0 29615 7 1 2 95981 29614
0 29616 5 1 1 29615
0 29617 7 1 2 29613 29616
0 29618 5 1 1 29617
0 29619 7 1 2 78655 29618
0 29620 5 1 1 29619
0 29621 7 1 2 87246 102154
0 29622 7 1 2 100683 29621
0 29623 5 1 1 29622
0 29624 7 1 2 29620 29623
0 29625 5 1 1 29624
0 29626 7 1 2 100278 83292
0 29627 7 1 2 29625 29626
0 29628 5 1 1 29627
0 29629 7 1 2 29610 29628
0 29630 5 1 1 29629
0 29631 7 1 2 72684 29630
0 29632 5 1 1 29631
0 29633 7 1 2 102061 1801
0 29634 5 1 1 29633
0 29635 7 1 2 78827 93225
0 29636 5 2 1 29635
0 29637 7 1 2 94319 102155
0 29638 5 1 1 29637
0 29639 7 1 2 29634 29638
0 29640 5 1 1 29639
0 29641 7 1 2 73505 29640
0 29642 5 1 1 29641
0 29643 7 1 2 79894 93418
0 29644 5 1 1 29643
0 29645 7 1 2 90695 90938
0 29646 5 1 1 29645
0 29647 7 1 2 29644 29646
0 29648 7 1 2 29642 29647
0 29649 5 1 1 29648
0 29650 7 1 2 67317 29649
0 29651 5 1 1 29650
0 29652 7 1 2 71402 101364
0 29653 5 1 1 29652
0 29654 7 1 2 101329 29653
0 29655 5 2 1 29654
0 29656 7 1 2 69868 102157
0 29657 5 1 1 29656
0 29658 7 1 2 29657 15196
0 29659 5 3 1 29658
0 29660 7 1 2 98827 98138
0 29661 7 1 2 102159 29660
0 29662 5 1 1 29661
0 29663 7 1 2 29651 29662
0 29664 5 1 1 29663
0 29665 7 1 2 100209 29664
0 29666 5 1 1 29665
0 29667 7 1 2 78775 83798
0 29668 5 1 1 29667
0 29669 7 1 2 66305 29668
0 29670 5 1 1 29669
0 29671 7 1 2 100326 29670
0 29672 5 1 1 29671
0 29673 7 1 2 64748 29672
0 29674 5 1 1 29673
0 29675 7 1 2 100332 29674
0 29676 5 1 1 29675
0 29677 7 1 2 71943 98094
0 29678 7 1 2 91760 29677
0 29679 7 1 2 84153 29678
0 29680 7 1 2 29676 29679
0 29681 5 1 1 29680
0 29682 7 1 2 29666 29681
0 29683 5 1 1 29682
0 29684 7 1 2 101430 29683
0 29685 5 1 1 29684
0 29686 7 1 2 29632 29685
0 29687 5 1 1 29686
0 29688 7 1 2 93259 29687
0 29689 5 1 1 29688
0 29690 7 1 2 29537 29689
0 29691 5 1 1 29690
0 29692 7 1 2 64114 29691
0 29693 5 1 1 29692
0 29694 7 6 2 72233 98757
0 29695 5 2 1 102162
0 29696 7 1 2 80163 98675
0 29697 7 1 2 102163 29696
0 29698 5 1 1 29697
0 29699 7 1 2 65431 93397
0 29700 5 1 1 29699
0 29701 7 1 2 68071 29700
0 29702 5 1 1 29701
0 29703 7 1 2 67177 87882
0 29704 7 1 2 99262 29703
0 29705 7 1 2 101630 29704
0 29706 7 1 2 29702 29705
0 29707 5 1 1 29706
0 29708 7 1 2 29698 29707
0 29709 5 1 1 29708
0 29710 7 1 2 100210 29709
0 29711 5 1 1 29710
0 29712 7 4 2 91776 86503
0 29713 7 1 2 89384 101984
0 29714 7 1 2 102170 29713
0 29715 7 1 2 102024 29714
0 29716 5 1 1 29715
0 29717 7 1 2 29711 29716
0 29718 5 1 1 29717
0 29719 7 1 2 65804 29718
0 29720 5 1 1 29719
0 29721 7 1 2 100211 101918
0 29722 5 1 1 29721
0 29723 7 2 2 91761 97463
0 29724 7 1 2 87933 102174
0 29725 5 1 1 29724
0 29726 7 1 2 29722 29725
0 29727 5 1 1 29726
0 29728 7 1 2 72234 89928
0 29729 7 1 2 95618 29728
0 29730 7 1 2 29727 29729
0 29731 5 1 1 29730
0 29732 7 1 2 29720 29731
0 29733 5 1 1 29732
0 29734 7 1 2 64115 29733
0 29735 5 1 1 29734
0 29736 7 2 2 100628 84289
0 29737 7 1 2 102097 102176
0 29738 5 1 1 29737
0 29739 7 1 2 65432 98424
0 29740 5 1 1 29739
0 29741 7 1 2 97919 29740
0 29742 5 2 1 29741
0 29743 7 4 2 88897 82245
0 29744 7 1 2 76920 102180
0 29745 7 1 2 102178 29744
0 29746 5 1 1 29745
0 29747 7 1 2 29738 29746
0 29748 5 1 1 29747
0 29749 7 1 2 66306 29748
0 29750 5 1 1 29749
0 29751 7 1 2 100816 82548
0 29752 5 1 1 29751
0 29753 7 1 2 29750 29752
0 29754 5 1 1 29753
0 29755 7 1 2 64749 29754
0 29756 5 1 1 29755
0 29757 7 2 2 66874 72393
0 29758 7 1 2 82196 102184
0 29759 7 1 2 100407 29758
0 29760 5 1 1 29759
0 29761 7 1 2 29756 29760
0 29762 5 1 1 29761
0 29763 7 1 2 99998 100137
0 29764 7 1 2 29762 29763
0 29765 5 1 1 29764
0 29766 7 1 2 29735 29765
0 29767 5 1 1 29766
0 29768 7 1 2 66024 29767
0 29769 5 1 1 29768
0 29770 7 5 2 63903 74392
0 29771 7 2 2 66307 102186
0 29772 7 2 2 100082 87799
0 29773 7 2 2 65123 65647
0 29774 7 2 2 94072 102195
0 29775 7 1 2 91960 102197
0 29776 7 1 2 102193 29775
0 29777 7 1 2 102191 29776
0 29778 5 1 1 29777
0 29779 7 1 2 29769 29778
0 29780 5 1 1 29779
0 29781 7 1 2 64422 29780
0 29782 5 1 1 29781
0 29783 7 1 2 64116 102179
0 29784 5 1 1 29783
0 29785 7 2 2 69171 97964
0 29786 5 1 1 102199
0 29787 7 1 2 65433 102200
0 29788 5 1 1 29787
0 29789 7 1 2 29784 29788
0 29790 5 1 1 29789
0 29791 7 1 2 78410 29790
0 29792 5 1 1 29791
0 29793 7 1 2 97735 78541
0 29794 5 1 1 29793
0 29795 7 1 2 29792 29794
0 29796 5 1 1 29795
0 29797 7 1 2 102013 29796
0 29798 5 1 1 29797
0 29799 7 1 2 74393 99073
0 29800 7 1 2 102175 29799
0 29801 5 1 1 29800
0 29802 7 1 2 29798 29801
0 29803 5 1 1 29802
0 29804 7 1 2 102007 88747
0 29805 7 1 2 29803 29804
0 29806 5 1 1 29805
0 29807 7 1 2 29782 29806
0 29808 5 1 1 29807
0 29809 7 1 2 73965 29808
0 29810 5 1 1 29809
0 29811 7 1 2 93703 102113
0 29812 5 1 1 29811
0 29813 7 1 2 102111 29812
0 29814 5 1 1 29813
0 29815 7 1 2 98479 29814
0 29816 5 1 1 29815
0 29817 7 1 2 69172 100945
0 29818 7 2 2 102089 29817
0 29819 5 1 1 102201
0 29820 7 1 2 29425 29819
0 29821 5 1 1 29820
0 29822 7 1 2 65805 29821
0 29823 5 1 1 29822
0 29824 7 2 2 89430 82682
0 29825 7 1 2 97104 74332
0 29826 7 1 2 102203 29825
0 29827 5 1 1 29826
0 29828 7 1 2 29823 29827
0 29829 5 1 1 29828
0 29830 7 1 2 65124 29829
0 29831 5 1 1 29830
0 29832 7 1 2 92464 102202
0 29833 5 1 1 29832
0 29834 7 1 2 29831 29833
0 29835 5 1 1 29834
0 29836 7 1 2 76083 29835
0 29837 5 1 1 29836
0 29838 7 2 2 85331 91448
0 29839 5 1 1 102205
0 29840 7 1 2 97877 102206
0 29841 5 1 1 29840
0 29842 7 2 2 93704 77030
0 29843 5 1 1 102207
0 29844 7 1 2 65434 102208
0 29845 7 1 2 96129 29844
0 29846 5 1 1 29845
0 29847 7 1 2 29841 29846
0 29848 5 1 1 29847
0 29849 7 1 2 72394 29848
0 29850 5 1 1 29849
0 29851 7 1 2 29839 29843
0 29852 5 1 1 29851
0 29853 7 1 2 29852 97927
0 29854 5 1 1 29853
0 29855 7 1 2 29850 29854
0 29856 5 1 1 29855
0 29857 7 1 2 102092 29856
0 29858 5 1 1 29857
0 29859 7 1 2 92339 93705
0 29860 7 1 2 93933 29859
0 29861 7 1 2 102105 29860
0 29862 5 1 1 29861
0 29863 7 1 2 29858 29862
0 29864 7 1 2 29837 29863
0 29865 5 1 1 29864
0 29866 7 1 2 72685 29865
0 29867 5 1 1 29866
0 29868 7 1 2 29816 29867
0 29869 5 1 1 29868
0 29870 7 1 2 100212 29869
0 29871 5 1 1 29870
0 29872 7 1 2 65806 102115
0 29873 5 1 1 29872
0 29874 7 1 2 79449 84347
0 29875 7 1 2 102117 29874
0 29876 5 1 1 29875
0 29877 7 1 2 29873 29876
0 29878 5 1 1 29877
0 29879 7 1 2 77353 29878
0 29880 5 1 1 29879
0 29881 7 1 2 79168 99263
0 29882 7 1 2 93402 29881
0 29883 7 2 2 65125 93141
0 29884 7 1 2 89492 102209
0 29885 7 1 2 29882 29884
0 29886 5 1 1 29885
0 29887 7 1 2 29880 29886
0 29888 5 1 1 29887
0 29889 7 1 2 100978 29888
0 29890 5 1 1 29889
0 29891 7 1 2 29871 29890
0 29892 5 1 1 29891
0 29893 7 1 2 73506 29892
0 29894 5 1 1 29893
0 29895 7 2 2 93260 88887
0 29896 7 1 2 102211 94795
0 29897 7 1 2 102123 29896
0 29898 5 1 1 29897
0 29899 7 1 2 29894 29898
0 29900 5 1 1 29899
0 29901 7 1 2 72235 29900
0 29902 5 1 1 29901
0 29903 7 1 2 29810 29902
0 29904 7 1 2 29693 29903
0 29905 5 1 1 29904
0 29906 7 1 2 80408 29905
0 29907 5 1 1 29906
0 29908 7 1 2 87319 98271
0 29909 5 1 1 29908
0 29910 7 2 2 81882 98257
0 29911 7 1 2 73150 102213
0 29912 5 1 1 29911
0 29913 7 1 2 29909 29912
0 29914 5 1 1 29913
0 29915 7 1 2 100279 29914
0 29916 5 1 1 29915
0 29917 7 1 2 99748 78046
0 29918 5 1 1 29917
0 29919 7 1 2 77453 29918
0 29920 5 1 1 29919
0 29921 7 1 2 67318 29920
0 29922 5 1 1 29921
0 29923 7 1 2 25830 29922
0 29924 5 1 1 29923
0 29925 7 1 2 100213 29924
0 29926 5 1 1 29925
0 29927 7 1 2 29916 29926
0 29928 5 1 1 29927
0 29929 7 1 2 64750 29928
0 29930 5 1 1 29929
0 29931 7 1 2 98272 101651
0 29932 5 1 1 29931
0 29933 7 1 2 29930 29932
0 29934 5 1 1 29933
0 29935 7 1 2 65807 29934
0 29936 5 1 1 29935
0 29937 7 1 2 4533 87097
0 29938 5 1 1 29937
0 29939 7 1 2 101649 29938
0 29940 5 1 1 29939
0 29941 7 1 2 24219 29940
0 29942 5 1 1 29941
0 29943 7 2 2 98458 29942
0 29944 7 1 2 77989 102215
0 29945 5 1 1 29944
0 29946 7 1 2 29936 29945
0 29947 5 1 1 29946
0 29948 7 1 2 64117 29947
0 29949 5 1 1 29948
0 29950 7 4 2 65808 74191
0 29951 7 1 2 102216 102217
0 29952 5 1 1 29951
0 29953 7 1 2 29949 29952
0 29954 5 1 1 29953
0 29955 7 1 2 85332 29954
0 29956 5 1 1 29955
0 29957 7 1 2 64118 98490
0 29958 5 2 1 29957
0 29959 7 1 2 29786 102221
0 29960 5 7 1 29959
0 29961 7 1 2 101655 1428
0 29962 5 1 1 29961
0 29963 7 1 2 102223 29962
0 29964 5 1 1 29963
0 29965 7 1 2 97122 98152
0 29966 5 1 1 29965
0 29967 7 1 2 29964 29966
0 29968 5 1 1 29967
0 29969 7 1 2 66025 29968
0 29970 5 1 1 29969
0 29971 7 3 2 65435 98876
0 29972 7 4 2 67319 77002
0 29973 7 1 2 64119 78312
0 29974 7 1 2 102233 29973
0 29975 7 1 2 102230 29974
0 29976 5 1 1 29975
0 29977 7 1 2 29970 29976
0 29978 5 1 1 29977
0 29979 7 1 2 64423 29978
0 29980 5 1 1 29979
0 29981 7 2 2 101083 97560
0 29982 5 1 1 102237
0 29983 7 1 2 99808 102234
0 29984 5 1 1 29983
0 29985 7 1 2 29982 29984
0 29986 5 1 1 29985
0 29987 7 2 2 74394 78313
0 29988 7 1 2 29986 102239
0 29989 5 1 1 29988
0 29990 7 1 2 29980 29989
0 29991 5 1 1 29990
0 29992 7 1 2 100673 29991
0 29993 5 1 1 29992
0 29994 7 1 2 29956 29993
0 29995 5 1 1 29994
0 29996 7 1 2 67654 29995
0 29997 5 1 1 29996
0 29998 7 1 2 73743 85365
0 29999 5 1 1 29998
0 30000 7 1 2 64751 29999
0 30001 7 1 2 100615 30000
0 30002 5 1 1 30001
0 30003 7 1 2 79595 101620
0 30004 5 1 1 30003
0 30005 7 1 2 30002 30004
0 30006 5 1 1 30005
0 30007 7 1 2 97898 30006
0 30008 5 1 1 30007
0 30009 7 1 2 100970 79450
0 30010 5 1 1 30009
0 30011 7 1 2 30008 30010
0 30012 5 1 1 30011
0 30013 7 1 2 64120 30012
0 30014 5 1 1 30013
0 30015 7 2 2 84355 97965
0 30016 5 1 1 102241
0 30017 7 1 2 85333 102242
0 30018 5 1 1 30017
0 30019 7 1 2 30014 30018
0 30020 5 1 1 30019
0 30021 7 1 2 101561 30020
0 30022 5 1 1 30021
0 30023 7 1 2 101964 3084
0 30024 5 1 1 30023
0 30025 7 1 2 90696 102235
0 30026 7 1 2 87280 30025
0 30027 7 1 2 30024 30026
0 30028 5 1 1 30027
0 30029 7 1 2 30022 30028
0 30030 5 1 1 30029
0 30031 7 1 2 93587 95415
0 30032 7 1 2 30030 30031
0 30033 5 1 1 30032
0 30034 7 1 2 29997 30033
0 30035 5 1 1 30034
0 30036 7 1 2 72236 30035
0 30037 5 1 1 30036
0 30038 7 2 2 85416 91153
0 30039 7 1 2 100980 102243
0 30040 7 9 2 72686 100422
0 30041 7 1 2 102245 74324
0 30042 7 1 2 30039 30041
0 30043 7 1 2 101622 30042
0 30044 5 1 1 30043
0 30045 7 1 2 30037 30044
0 30046 5 1 1 30045
0 30047 7 1 2 79881 30046
0 30048 5 1 1 30047
0 30049 7 1 2 29907 30048
0 30050 7 1 2 29282 30049
0 30051 7 1 2 28847 30050
0 30052 7 1 2 28066 30051
0 30053 5 1 1 30052
0 30054 7 1 2 67110 30053
0 30055 5 1 1 30054
0 30056 7 27 2 7943 24873
0 30057 7 3 2 67178 102254
0 30058 7 1 2 68072 101793
0 30059 5 1 1 30058
0 30060 7 1 2 94886 30059
0 30061 5 1 1 30060
0 30062 7 1 2 73507 30061
0 30063 5 1 1 30062
0 30064 7 1 2 81739 88451
0 30065 5 1 1 30064
0 30066 7 1 2 30063 30065
0 30067 5 1 1 30066
0 30068 7 1 2 71403 30067
0 30069 5 1 1 30068
0 30070 7 1 2 73151 91752
0 30071 5 2 1 30070
0 30072 7 1 2 80445 76025
0 30073 5 1 1 30072
0 30074 7 1 2 102284 30073
0 30075 5 1 1 30074
0 30076 7 1 2 80482 30075
0 30077 5 1 1 30076
0 30078 7 1 2 30069 30077
0 30079 5 1 1 30078
0 30080 7 1 2 67655 30079
0 30081 5 1 1 30080
0 30082 7 1 2 83602 83988
0 30083 7 1 2 83210 30082
0 30084 5 2 1 30083
0 30085 7 1 2 30081 102286
0 30086 5 1 1 30085
0 30087 7 1 2 98491 30086
0 30088 5 1 1 30087
0 30089 7 1 2 99445 88707
0 30090 7 1 2 93579 30089
0 30091 5 1 1 30090
0 30092 7 2 2 74665 82925
0 30093 5 1 1 102288
0 30094 7 1 2 80972 30093
0 30095 5 2 1 30094
0 30096 7 1 2 79588 102290
0 30097 5 1 1 30096
0 30098 7 2 2 72395 94861
0 30099 5 1 1 102292
0 30100 7 1 2 97920 30099
0 30101 5 2 1 30100
0 30102 7 1 2 84290 102294
0 30103 7 1 2 30097 30102
0 30104 5 1 1 30103
0 30105 7 1 2 30091 30104
0 30106 5 1 1 30105
0 30107 7 1 2 65436 30106
0 30108 5 1 1 30107
0 30109 7 1 2 95264 97232
0 30110 5 2 1 30109
0 30111 7 1 2 19334 102296
0 30112 5 1 1 30111
0 30113 7 1 2 70816 77963
0 30114 7 1 2 30112 30113
0 30115 5 1 1 30114
0 30116 7 1 2 30108 30115
0 30117 7 1 2 30088 30116
0 30118 5 1 1 30117
0 30119 7 1 2 69173 30118
0 30120 5 1 1 30119
0 30121 7 5 2 67320 85451
0 30122 5 1 1 102298
0 30123 7 1 2 84708 88452
0 30124 5 1 1 30123
0 30125 7 1 2 88841 92919
0 30126 5 1 1 30125
0 30127 7 1 2 102291 30126
0 30128 5 1 1 30127
0 30129 7 1 2 68073 30128
0 30130 5 1 1 30129
0 30131 7 1 2 30124 30130
0 30132 5 1 1 30131
0 30133 7 1 2 65437 30132
0 30134 5 1 1 30133
0 30135 7 1 2 70197 83473
0 30136 5 2 1 30135
0 30137 7 1 2 78937 102303
0 30138 5 1 1 30137
0 30139 7 1 2 71404 30138
0 30140 5 1 1 30139
0 30141 7 1 2 76060 102285
0 30142 5 1 1 30141
0 30143 7 1 2 95176 30142
0 30144 5 1 1 30143
0 30145 7 1 2 30140 30144
0 30146 5 1 1 30145
0 30147 7 1 2 73508 30146
0 30148 5 1 1 30147
0 30149 7 1 2 30134 30148
0 30150 5 1 1 30149
0 30151 7 1 2 67656 30150
0 30152 5 1 1 30151
0 30153 7 1 2 102287 30152
0 30154 5 1 1 30153
0 30155 7 1 2 102299 30154
0 30156 5 1 1 30155
0 30157 7 1 2 30120 30156
0 30158 5 1 1 30157
0 30159 7 1 2 69869 30158
0 30160 5 1 1 30159
0 30161 7 1 2 84082 92203
0 30162 5 1 1 30161
0 30163 7 1 2 79069 90499
0 30164 5 1 1 30163
0 30165 7 1 2 71405 93786
0 30166 5 1 1 30165
0 30167 7 1 2 87078 30166
0 30168 7 1 2 30164 30167
0 30169 5 1 1 30168
0 30170 7 1 2 73152 30169
0 30171 5 1 1 30170
0 30172 7 1 2 30162 30171
0 30173 5 1 1 30172
0 30174 7 1 2 69870 30173
0 30175 5 1 1 30174
0 30176 7 2 2 76413 79731
0 30177 5 1 1 102305
0 30178 7 1 2 101676 102306
0 30179 5 1 1 30178
0 30180 7 1 2 92933 11720
0 30181 5 1 1 30180
0 30182 7 1 2 79768 30181
0 30183 5 1 1 30182
0 30184 7 1 2 79840 86187
0 30185 7 1 2 23314 30184
0 30186 5 1 1 30185
0 30187 7 1 2 84980 30186
0 30188 5 1 1 30187
0 30189 7 1 2 30183 30188
0 30190 5 1 1 30189
0 30191 7 1 2 68074 30190
0 30192 5 1 1 30191
0 30193 7 1 2 30179 30192
0 30194 7 1 2 30175 30193
0 30195 5 1 1 30194
0 30196 7 1 2 99400 30195
0 30197 5 1 1 30196
0 30198 7 3 2 80472 83839
0 30199 5 2 1 102307
0 30200 7 1 2 66308 102310
0 30201 5 1 1 30200
0 30202 7 1 2 30201 13797
0 30203 5 1 1 30202
0 30204 7 1 2 70198 30203
0 30205 5 1 1 30204
0 30206 7 1 2 68667 99817
0 30207 5 1 1 30206
0 30208 7 1 2 30205 30207
0 30209 5 1 1 30208
0 30210 7 1 2 78742 30209
0 30211 5 1 1 30210
0 30212 7 2 2 69871 86285
0 30213 5 1 1 102312
0 30214 7 1 2 77124 30213
0 30215 5 1 1 30214
0 30216 7 1 2 82317 76084
0 30217 7 1 2 30215 30216
0 30218 5 1 1 30217
0 30219 7 1 2 30211 30218
0 30220 5 1 1 30219
0 30221 7 1 2 99383 30220
0 30222 5 1 1 30221
0 30223 7 1 2 30197 30222
0 30224 5 1 1 30223
0 30225 7 1 2 67657 30224
0 30226 5 1 1 30225
0 30227 7 1 2 99401 94899
0 30228 5 1 1 30227
0 30229 7 1 2 82437 100780
0 30230 7 1 2 76085 30229
0 30231 5 1 1 30230
0 30232 7 1 2 30228 30231
0 30233 5 1 1 30232
0 30234 7 1 2 69872 30233
0 30235 5 1 1 30234
0 30236 7 2 2 82438 98025
0 30237 7 1 2 86592 102314
0 30238 5 1 1 30237
0 30239 7 1 2 30235 30238
0 30240 5 1 1 30239
0 30241 7 1 2 67658 30240
0 30242 5 1 1 30241
0 30243 7 11 2 69174 67321
0 30244 5 2 1 102316
0 30245 7 2 2 74170 102317
0 30246 7 2 2 73153 77283
0 30247 7 1 2 93089 102331
0 30248 7 1 2 102329 30247
0 30249 5 1 1 30248
0 30250 7 1 2 30242 30249
0 30251 5 1 1 30250
0 30252 7 1 2 84834 30251
0 30253 5 1 1 30252
0 30254 7 1 2 70199 100594
0 30255 5 1 1 30254
0 30256 7 1 2 30255 95185
0 30257 5 1 1 30256
0 30258 7 1 2 99420 99760
0 30259 5 1 1 30258
0 30260 7 1 2 91325 30259
0 30261 7 1 2 30257 30260
0 30262 5 1 1 30261
0 30263 7 1 2 30253 30262
0 30264 7 1 2 30226 30263
0 30265 5 1 1 30264
0 30266 7 1 2 68414 30265
0 30267 5 1 1 30266
0 30268 7 1 2 99475 85411
0 30269 7 1 2 83593 30268
0 30270 5 1 1 30269
0 30271 7 1 2 30267 30270
0 30272 7 1 2 30160 30271
0 30273 5 1 1 30272
0 30274 7 1 2 79137 30273
0 30275 5 1 1 30274
0 30276 7 1 2 99294 91703
0 30277 7 2 2 88464 30276
0 30278 7 1 2 95601 102333
0 30279 5 1 1 30278
0 30280 7 2 2 74960 79791
0 30281 7 1 2 95799 102335
0 30282 5 1 1 30281
0 30283 7 1 2 79639 94628
0 30284 5 1 1 30283
0 30285 7 1 2 30282 30284
0 30286 5 1 1 30285
0 30287 7 1 2 97042 30286
0 30288 5 1 1 30287
0 30289 7 2 2 77003 87232
0 30290 7 2 2 96748 87925
0 30291 7 1 2 78989 102339
0 30292 7 1 2 102337 30291
0 30293 5 1 1 30292
0 30294 7 1 2 30288 30293
0 30295 5 1 1 30294
0 30296 7 1 2 70817 30295
0 30297 5 1 1 30296
0 30298 7 1 2 30279 30297
0 30299 5 1 1 30298
0 30300 7 1 2 69175 30299
0 30301 5 1 1 30300
0 30302 7 1 2 102334 98106
0 30303 5 1 1 30302
0 30304 7 1 2 30301 30303
0 30305 5 1 1 30304
0 30306 7 1 2 69873 30305
0 30307 5 1 1 30306
0 30308 7 2 2 70818 101936
0 30309 5 2 1 102341
0 30310 7 2 2 74353 77901
0 30311 7 1 2 102342 102345
0 30312 5 1 1 30311
0 30313 7 1 2 30307 30312
0 30314 5 1 1 30313
0 30315 7 1 2 80704 30314
0 30316 5 1 1 30315
0 30317 7 1 2 99402 96623
0 30318 5 1 1 30317
0 30319 7 3 2 70819 99185
0 30320 5 1 1 102347
0 30321 7 1 2 73154 99551
0 30322 7 1 2 102348 30321
0 30323 5 1 1 30322
0 30324 7 1 2 30318 30323
0 30325 5 1 1 30324
0 30326 7 1 2 76324 30325
0 30327 5 1 1 30326
0 30328 7 1 2 99446 93616
0 30329 5 1 1 30328
0 30330 7 2 2 99295 92380
0 30331 5 1 1 102350
0 30332 7 6 2 70820 71830
0 30333 7 2 2 100110 102352
0 30334 5 1 1 102358
0 30335 7 1 2 76026 102359
0 30336 5 1 1 30335
0 30337 7 1 2 30331 30336
0 30338 5 1 1 30337
0 30339 7 1 2 69176 30338
0 30340 5 1 1 30339
0 30341 7 1 2 30329 30340
0 30342 7 1 2 30327 30341
0 30343 5 1 1 30342
0 30344 7 1 2 67659 30343
0 30345 5 1 1 30344
0 30346 7 1 2 97921 19957
0 30347 5 1 1 30346
0 30348 7 1 2 69177 30347
0 30349 5 1 1 30348
0 30350 7 1 2 99468 30349
0 30351 5 1 1 30350
0 30352 7 1 2 81438 90758
0 30353 7 1 2 30351 30352
0 30354 5 1 1 30353
0 30355 7 1 2 30345 30354
0 30356 5 1 1 30355
0 30357 7 1 2 78866 30356
0 30358 5 1 1 30357
0 30359 7 1 2 30316 30358
0 30360 7 1 2 30275 30359
0 30361 5 1 1 30360
0 30362 7 1 2 102281 30361
0 30363 5 1 1 30362
0 30364 7 1 2 80358 76027
0 30365 5 3 1 30364
0 30366 7 4 2 71831 79732
0 30367 5 1 1 102363
0 30368 7 1 2 76696 30367
0 30369 5 2 1 30368
0 30370 7 1 2 76325 102367
0 30371 5 1 1 30370
0 30372 7 1 2 102360 30371
0 30373 5 1 1 30372
0 30374 7 1 2 67660 30373
0 30375 5 1 1 30374
0 30376 7 4 2 68415 80409
0 30377 5 4 1 102369
0 30378 7 1 2 102373 7135
0 30379 5 2 1 30378
0 30380 7 1 2 77539 102377
0 30381 5 1 1 30380
0 30382 7 1 2 30375 30381
0 30383 5 1 1 30382
0 30384 7 1 2 70452 30383
0 30385 5 1 1 30384
0 30386 7 2 2 79027 75691
0 30387 5 1 1 102379
0 30388 7 1 2 83603 102380
0 30389 5 1 1 30388
0 30390 7 1 2 30385 30389
0 30391 5 1 1 30390
0 30392 7 1 2 72396 30391
0 30393 5 1 1 30392
0 30394 7 1 2 97043 80178
0 30395 5 2 1 30394
0 30396 7 1 2 101930 102381
0 30397 5 1 1 30396
0 30398 7 1 2 88688 30397
0 30399 5 1 1 30398
0 30400 7 1 2 30393 30399
0 30401 5 1 1 30400
0 30402 7 1 2 100214 30401
0 30403 5 1 1 30402
0 30404 7 1 2 81375 82197
0 30405 5 1 1 30404
0 30406 7 1 2 77714 92755
0 30407 5 1 1 30406
0 30408 7 1 2 30405 30407
0 30409 5 1 1 30408
0 30410 7 1 2 86052 30409
0 30411 5 1 1 30410
0 30412 7 1 2 76047 99933
0 30413 5 1 1 30412
0 30414 7 4 2 66309 80410
0 30415 5 1 1 102383
0 30416 7 1 2 86024 87027
0 30417 7 1 2 102384 30416
0 30418 5 1 1 30417
0 30419 7 1 2 30413 30418
0 30420 5 1 1 30419
0 30421 7 1 2 67661 30420
0 30422 5 1 1 30421
0 30423 7 1 2 30411 30422
0 30424 5 1 1 30423
0 30425 7 1 2 70200 30424
0 30426 5 1 1 30425
0 30427 7 1 2 82926 76028
0 30428 5 1 1 30427
0 30429 7 1 2 86904 319
0 30430 5 1 1 30429
0 30431 7 1 2 65438 88717
0 30432 7 1 2 30430 30431
0 30433 5 1 1 30432
0 30434 7 1 2 30428 30433
0 30435 5 1 1 30434
0 30436 7 1 2 97214 30435
0 30437 5 1 1 30436
0 30438 7 1 2 30426 30437
0 30439 5 1 1 30438
0 30440 7 1 2 72397 30439
0 30441 5 1 1 30440
0 30442 7 1 2 99789 101937
0 30443 5 1 1 30442
0 30444 7 1 2 66310 89178
0 30445 5 1 1 30444
0 30446 7 1 2 71406 94267
0 30447 7 1 2 98969 30446
0 30448 5 1 1 30447
0 30449 7 1 2 30445 30448
0 30450 5 1 1 30449
0 30451 7 1 2 98187 92629
0 30452 7 1 2 30450 30451
0 30453 5 1 1 30452
0 30454 7 1 2 30443 30453
0 30455 7 1 2 30441 30454
0 30456 5 1 1 30455
0 30457 7 1 2 69874 100280
0 30458 7 1 2 30456 30457
0 30459 5 1 1 30458
0 30460 7 1 2 30403 30459
0 30461 5 1 1 30460
0 30462 7 10 2 65809 72237
0 30463 7 1 2 93042 102387
0 30464 7 1 2 30461 30463
0 30465 5 1 1 30464
0 30466 7 1 2 30363 30465
0 30467 5 1 1 30466
0 30468 7 1 2 67111 30467
0 30469 5 1 1 30468
0 30470 7 3 2 99628 102255
0 30471 7 2 2 66875 102397
0 30472 7 2 2 95483 102400
0 30473 5 1 1 102402
0 30474 7 6 2 70821 67179
0 30475 7 3 2 71944 67322
0 30476 7 3 2 102404 102410
0 30477 7 1 2 95723 102413
0 30478 7 1 2 100848 30477
0 30479 5 1 1 30478
0 30480 7 1 2 30473 30479
0 30481 5 1 1 30480
0 30482 7 1 2 76086 30481
0 30483 5 1 1 30482
0 30484 7 4 2 67323 102405
0 30485 7 2 2 100806 102416
0 30486 7 3 2 86633 87002
0 30487 5 2 1 102422
0 30488 7 1 2 86113 102423
0 30489 5 2 1 30488
0 30490 7 1 2 102420 102427
0 30491 5 1 1 30490
0 30492 7 1 2 93238 102398
0 30493 7 1 2 94281 30492
0 30494 5 1 1 30493
0 30495 7 1 2 30491 30494
0 30496 5 1 1 30495
0 30497 7 1 2 77902 30496
0 30498 5 1 1 30497
0 30499 7 2 2 74790 100987
0 30500 7 3 2 70201 70685
0 30501 7 4 2 84073 102431
0 30502 7 1 2 67180 99967
0 30503 7 1 2 91880 30502
0 30504 7 1 2 102434 30503
0 30505 7 1 2 102429 30504
0 30506 5 1 1 30505
0 30507 7 1 2 30498 30506
0 30508 7 1 2 30483 30507
0 30509 5 1 1 30508
0 30510 7 1 2 67662 30509
0 30511 5 1 1 30510
0 30512 7 1 2 77112 100281
0 30513 5 1 1 30512
0 30514 7 1 2 100224 30513
0 30515 5 1 1 30514
0 30516 7 1 2 81883 30515
0 30517 5 1 1 30516
0 30518 7 5 2 83502 83152
0 30519 7 2 2 100282 102438
0 30520 5 1 1 102443
0 30521 7 1 2 30517 30520
0 30522 5 1 1 30521
0 30523 7 1 2 102417 30522
0 30524 5 1 1 30523
0 30525 7 1 2 94268 102403
0 30526 5 1 1 30525
0 30527 7 1 2 30524 30526
0 30528 5 1 1 30527
0 30529 7 1 2 68416 30528
0 30530 5 1 1 30529
0 30531 7 1 2 71663 80200
0 30532 7 1 2 86609 30531
0 30533 7 1 2 102401 30532
0 30534 5 1 1 30533
0 30535 7 1 2 30530 30534
0 30536 5 1 1 30535
0 30537 7 1 2 86716 30536
0 30538 5 1 1 30537
0 30539 7 1 2 30511 30538
0 30540 5 1 1 30539
0 30541 7 1 2 64121 30540
0 30542 5 1 1 30541
0 30543 7 7 2 66752 67324
0 30544 7 3 2 65810 102445
0 30545 5 1 1 102452
0 30546 7 2 2 70453 98425
0 30547 5 1 1 102455
0 30548 7 1 2 73744 102456
0 30549 5 1 1 30548
0 30550 7 1 2 30545 30549
0 30551 5 1 1 30550
0 30552 7 1 2 65126 30551
0 30553 5 1 1 30552
0 30554 7 3 2 70202 98426
0 30555 5 2 1 102457
0 30556 7 1 2 97922 102460
0 30557 5 1 1 30556
0 30558 7 1 2 83066 30557
0 30559 5 1 1 30558
0 30560 7 1 2 30553 30559
0 30561 5 1 1 30560
0 30562 7 1 2 71664 30561
0 30563 5 1 1 30562
0 30564 7 1 2 65127 67325
0 30565 7 1 2 79340 30564
0 30566 7 1 2 80201 30565
0 30567 5 1 1 30566
0 30568 7 1 2 30563 30567
0 30569 5 1 1 30568
0 30570 7 1 2 68417 30569
0 30571 5 1 1 30570
0 30572 7 1 2 83533 83112
0 30573 5 1 1 30572
0 30574 7 1 2 101763 30573
0 30575 5 1 1 30574
0 30576 7 1 2 98382 30575
0 30577 5 1 1 30576
0 30578 7 1 2 98427 98302
0 30579 5 1 1 30578
0 30580 7 1 2 92838 100775
0 30581 5 1 1 30580
0 30582 7 1 2 30579 30581
0 30583 5 1 1 30582
0 30584 7 1 2 84835 30583
0 30585 5 1 1 30584
0 30586 7 1 2 30577 30585
0 30587 7 1 2 30571 30586
0 30588 5 1 1 30587
0 30589 7 1 2 76087 30588
0 30590 5 1 1 30589
0 30591 7 1 2 90015 86725
0 30592 5 1 1 30591
0 30593 7 1 2 81361 101238
0 30594 5 1 1 30593
0 30595 7 1 2 30592 30594
0 30596 5 1 1 30595
0 30597 7 1 2 70203 30596
0 30598 5 1 1 30597
0 30599 7 1 2 92942 86885
0 30600 5 1 1 30599
0 30601 7 1 2 30598 30600
0 30602 5 1 1 30601
0 30603 7 1 2 98428 30602
0 30604 5 1 1 30603
0 30605 7 1 2 92839 80080
0 30606 7 1 2 102430 30605
0 30607 5 1 1 30606
0 30608 7 1 2 30604 30607
0 30609 7 1 2 30590 30608
0 30610 5 1 1 30609
0 30611 7 1 2 100283 30610
0 30612 5 1 1 30611
0 30613 7 2 2 98492 100215
0 30614 5 1 1 102462
0 30615 7 1 2 102428 102463
0 30616 5 1 1 30615
0 30617 7 1 2 67663 30616
0 30618 7 1 2 30612 30617
0 30619 5 1 1 30618
0 30620 7 4 2 69178 67181
0 30621 7 4 2 65811 100416
0 30622 5 1 1 102468
0 30623 7 1 2 91194 102435
0 30624 7 1 2 102469 30623
0 30625 5 1 1 30624
0 30626 7 1 2 30614 30625
0 30627 5 1 1 30626
0 30628 7 1 2 81884 30627
0 30629 5 1 1 30628
0 30630 7 1 2 102444 98383
0 30631 5 1 1 30630
0 30632 7 1 2 30629 30631
0 30633 5 1 1 30632
0 30634 7 1 2 74961 30633
0 30635 5 1 1 30634
0 30636 7 2 2 67326 91332
0 30637 7 2 2 101895 102472
0 30638 7 1 2 89940 75518
0 30639 7 1 2 102474 30638
0 30640 5 1 1 30639
0 30641 7 1 2 30635 30640
0 30642 5 1 1 30641
0 30643 7 1 2 68418 30642
0 30644 5 1 1 30643
0 30645 7 1 2 83067 80791
0 30646 5 1 1 30645
0 30647 7 2 2 84753 83444
0 30648 5 3 1 102476
0 30649 7 1 2 65439 102477
0 30650 5 1 1 30649
0 30651 7 1 2 70454 80524
0 30652 5 1 1 30651
0 30653 7 1 2 66558 30652
0 30654 7 1 2 30650 30653
0 30655 5 1 1 30654
0 30656 7 1 2 30646 30655
0 30657 5 1 1 30656
0 30658 7 1 2 65128 30657
0 30659 5 1 1 30658
0 30660 7 1 2 98994 30659
0 30661 5 1 1 30660
0 30662 7 3 2 73155 99153
0 30663 7 1 2 100395 102481
0 30664 7 1 2 30661 30663
0 30665 5 1 1 30664
0 30666 7 1 2 72687 30665
0 30667 7 1 2 30644 30666
0 30668 5 1 1 30667
0 30669 7 1 2 102464 30668
0 30670 7 1 2 30619 30669
0 30671 5 1 1 30670
0 30672 7 1 2 30542 30671
0 30673 5 1 1 30672
0 30674 7 1 2 69875 30673
0 30675 5 1 1 30674
0 30676 7 5 2 69179 65648
0 30677 7 3 2 102406 102484
0 30678 5 1 1 102489
0 30679 7 2 2 63904 102490
0 30680 7 2 2 85688 74962
0 30681 5 1 1 102494
0 30682 7 1 2 81885 76118
0 30683 5 1 1 30682
0 30684 7 1 2 30681 30683
0 30685 5 1 1 30684
0 30686 7 1 2 102492 30685
0 30687 5 1 1 30686
0 30688 7 1 2 76061 94282
0 30689 5 1 1 30688
0 30690 7 5 2 72238 74395
0 30691 7 2 2 102256 102496
0 30692 7 1 2 75010 94289
0 30693 5 1 1 30692
0 30694 7 1 2 102501 30693
0 30695 7 1 2 30689 30694
0 30696 5 1 1 30695
0 30697 7 1 2 30687 30696
0 30698 5 1 1 30697
0 30699 7 1 2 72398 30698
0 30700 5 1 1 30699
0 30701 7 2 2 85507 76088
0 30702 7 7 2 67182 81886
0 30703 7 2 2 67327 100807
0 30704 7 1 2 68419 102512
0 30705 7 1 2 102505 30704
0 30706 7 1 2 102503 30705
0 30707 5 1 1 30706
0 30708 7 1 2 30700 30707
0 30709 5 1 1 30708
0 30710 7 1 2 67664 30709
0 30711 5 1 1 30710
0 30712 7 3 2 73156 93090
0 30713 7 3 2 67328 85689
0 30714 7 1 2 102493 102517
0 30715 5 1 1 30714
0 30716 7 4 2 72239 102257
0 30717 7 1 2 94290 102520
0 30718 7 1 2 102224 30717
0 30719 5 1 1 30718
0 30720 7 1 2 30715 30719
0 30721 5 1 1 30720
0 30722 7 1 2 102514 30721
0 30723 5 1 1 30722
0 30724 7 1 2 30711 30723
0 30725 5 1 1 30724
0 30726 7 1 2 77903 30725
0 30727 5 1 1 30726
0 30728 7 1 2 30675 30727
0 30729 5 1 1 30728
0 30730 7 1 2 68859 30729
0 30731 5 1 1 30730
0 30732 7 2 2 78656 101938
0 30733 5 1 1 102524
0 30734 7 2 2 69876 85412
0 30735 5 1 1 102526
0 30736 7 1 2 94291 30735
0 30737 5 1 1 30736
0 30738 7 2 2 69877 93152
0 30739 5 1 1 102528
0 30740 7 1 2 3324 30739
0 30741 5 2 1 30740
0 30742 7 1 2 72399 102530
0 30743 7 1 2 30737 30742
0 30744 5 1 1 30743
0 30745 7 1 2 30733 30744
0 30746 5 1 1 30745
0 30747 7 1 2 65812 30746
0 30748 5 1 1 30747
0 30749 7 1 2 65813 101939
0 30750 5 1 1 30749
0 30751 7 2 2 99968 98358
0 30752 5 1 1 102532
0 30753 7 1 2 30750 30752
0 30754 5 3 1 30753
0 30755 7 1 2 94276 102534
0 30756 5 1 1 30755
0 30757 7 1 2 99969 98119
0 30758 5 1 1 30757
0 30759 7 1 2 30756 30758
0 30760 7 1 2 30748 30759
0 30761 5 1 1 30760
0 30762 7 1 2 64122 30761
0 30763 5 1 1 30762
0 30764 7 1 2 98651 102515
0 30765 7 1 2 94292 30764
0 30766 5 1 1 30765
0 30767 7 1 2 30763 30766
0 30768 5 1 1 30767
0 30769 7 1 2 66876 74007
0 30770 7 1 2 102521 30769
0 30771 7 1 2 30768 30770
0 30772 5 1 1 30771
0 30773 7 1 2 30731 30772
0 30774 5 1 1 30773
0 30775 7 1 2 72154 30774
0 30776 5 1 1 30775
0 30777 7 3 2 102497 97590
0 30778 5 1 1 102537
0 30779 7 1 2 71407 102538
0 30780 5 1 1 30779
0 30781 7 16 2 67112 67183
0 30782 7 3 2 70822 102540
0 30783 7 3 2 102556 97328
0 30784 5 2 1 102559
0 30785 7 2 2 70455 102560
0 30786 5 1 1 102564
0 30787 7 1 2 71832 102565
0 30788 5 1 1 30787
0 30789 7 1 2 30780 30788
0 30790 5 1 1 30789
0 30791 7 1 2 84291 30790
0 30792 5 1 1 30791
0 30793 7 1 2 80705 100312
0 30794 5 1 1 30793
0 30795 7 1 2 93291 30794
0 30796 5 2 1 30795
0 30797 7 3 2 72240 97591
0 30798 7 1 2 102568 98362
0 30799 7 1 2 102566 30798
0 30800 5 1 1 30799
0 30801 7 1 2 30792 30800
0 30802 5 1 1 30801
0 30803 7 1 2 72400 30802
0 30804 5 1 1 30803
0 30805 7 1 2 102562 30778
0 30806 5 1 1 30805
0 30807 7 1 2 75920 30806
0 30808 5 1 1 30807
0 30809 7 1 2 80706 102561
0 30810 5 1 1 30809
0 30811 7 1 2 94293 102539
0 30812 5 1 1 30811
0 30813 7 1 2 30810 30812
0 30814 5 1 1 30813
0 30815 7 1 2 75011 30814
0 30816 5 1 1 30815
0 30817 7 1 2 30808 30816
0 30818 5 1 1 30817
0 30819 7 1 2 96749 30818
0 30820 5 1 1 30819
0 30821 7 1 2 30804 30820
0 30822 5 1 1 30821
0 30823 7 1 2 78170 30822
0 30824 5 1 1 30823
0 30825 7 8 2 72155 72241
0 30826 7 2 2 77904 102571
0 30827 7 3 2 64123 93212
0 30828 7 1 2 97083 102581
0 30829 5 1 1 30828
0 30830 7 1 2 72688 102225
0 30831 7 1 2 102567 30830
0 30832 5 1 1 30831
0 30833 7 1 2 30829 30832
0 30834 5 1 1 30833
0 30835 7 1 2 102579 30834
0 30836 5 1 1 30835
0 30837 7 1 2 75278 76089
0 30838 5 2 1 30837
0 30839 7 1 2 66311 88453
0 30840 5 1 1 30839
0 30841 7 1 2 102584 30840
0 30842 5 1 1 30841
0 30843 7 1 2 66753 101052
0 30844 7 1 2 30842 30843
0 30845 5 1 1 30844
0 30846 7 2 2 85508 74963
0 30847 7 1 2 67665 11454
0 30848 7 1 2 102586 30847
0 30849 5 1 1 30848
0 30850 7 1 2 30845 30849
0 30851 5 1 1 30850
0 30852 7 1 2 67329 30851
0 30853 5 1 1 30852
0 30854 7 1 2 99384 84709
0 30855 7 1 2 92743 30854
0 30856 5 1 1 30855
0 30857 7 1 2 30853 30856
0 30858 5 1 1 30857
0 30859 7 1 2 65440 30858
0 30860 5 1 1 30859
0 30861 7 1 2 83503 101940
0 30862 5 1 1 30861
0 30863 7 1 2 67330 93183
0 30864 7 1 2 88419 30863
0 30865 5 1 1 30864
0 30866 7 1 2 30862 30865
0 30867 5 1 1 30866
0 30868 7 1 2 82439 30867
0 30869 5 1 1 30868
0 30870 7 2 2 67331 84292
0 30871 7 2 2 93213 102588
0 30872 5 2 1 102590
0 30873 7 1 2 102343 102592
0 30874 5 3 1 30873
0 30875 7 1 2 69180 102594
0 30876 5 1 1 30875
0 30877 7 2 2 99459 91467
0 30878 5 1 1 102597
0 30879 7 1 2 30876 30878
0 30880 5 3 1 30879
0 30881 7 1 2 95177 102599
0 30882 5 1 1 30881
0 30883 7 1 2 73509 30882
0 30884 7 1 2 30869 30883
0 30885 5 1 1 30884
0 30886 7 1 2 101941 93787
0 30887 5 1 1 30886
0 30888 7 1 2 72401 85413
0 30889 7 1 2 87060 30888
0 30890 5 1 1 30889
0 30891 7 1 2 30887 30890
0 30892 5 1 1 30891
0 30893 7 1 2 70823 30892
0 30894 5 1 1 30893
0 30895 7 1 2 89814 79508
0 30896 5 1 1 30895
0 30897 7 4 2 92662 30896
0 30898 5 1 1 102602
0 30899 7 1 2 96750 30898
0 30900 5 1 1 30899
0 30901 7 1 2 101181 30900
0 30902 5 1 1 30901
0 30903 7 1 2 78294 30902
0 30904 5 1 1 30903
0 30905 7 1 2 102593 30904
0 30906 5 1 1 30905
0 30907 7 1 2 84836 30906
0 30908 5 1 1 30907
0 30909 7 1 2 30894 30908
0 30910 5 1 1 30909
0 30911 7 1 2 69181 30910
0 30912 5 1 1 30911
0 30913 7 1 2 76090 90500
0 30914 5 1 1 30913
0 30915 7 1 2 10173 30914
0 30916 5 1 1 30915
0 30917 7 1 2 70456 30916
0 30918 5 1 1 30917
0 30919 7 1 2 73157 80473
0 30920 5 1 1 30919
0 30921 7 1 2 76414 30920
0 30922 7 1 2 94677 30921
0 30923 5 1 1 30922
0 30924 7 1 2 30918 30923
0 30925 5 1 1 30924
0 30926 7 1 2 67332 102048
0 30927 7 1 2 30925 30926
0 30928 5 1 1 30927
0 30929 7 1 2 84837 102598
0 30930 5 1 1 30929
0 30931 7 1 2 68420 30930
0 30932 7 1 2 30928 30931
0 30933 7 1 2 30912 30932
0 30934 5 1 1 30933
0 30935 7 1 2 30885 30934
0 30936 5 1 1 30935
0 30937 7 1 2 30860 30936
0 30938 5 1 1 30937
0 30939 7 2 2 76807 102541
0 30940 7 1 2 30938 102606
0 30941 5 1 1 30940
0 30942 7 1 2 30836 30941
0 30943 5 1 1 30942
0 30944 7 1 2 68860 30943
0 30945 5 1 1 30944
0 30946 7 1 2 30824 30945
0 30947 5 1 1 30946
0 30948 7 1 2 102258 30947
0 30949 5 1 1 30948
0 30950 7 5 2 67184 96298
0 30951 7 3 2 99552 102608
0 30952 5 1 1 102613
0 30953 7 1 2 65129 102614
0 30954 5 1 1 30953
0 30955 7 35 2 67113 72242
0 30956 7 8 2 65814 102616
0 30957 7 2 2 98147 102651
0 30958 5 1 1 102659
0 30959 7 1 2 30954 30958
0 30960 5 1 1 30959
0 30961 7 1 2 80411 30960
0 30962 5 1 1 30961
0 30963 7 8 2 74396 102617
0 30964 5 5 1 102661
0 30965 7 29 2 72156 67185
0 30966 7 9 2 70824 102674
0 30967 7 4 2 69182 74903
0 30968 7 1 2 102703 102712
0 30969 5 1 1 30968
0 30970 7 1 2 102669 30969
0 30971 5 1 1 30970
0 30972 7 2 2 82927 30971
0 30973 5 1 1 102716
0 30974 7 1 2 30962 30973
0 30975 5 1 1 30974
0 30976 7 1 2 68075 30975
0 30977 5 1 1 30976
0 30978 7 1 2 30952 102670
0 30979 5 1 1 30978
0 30980 7 1 2 30979 97795
0 30981 5 1 1 30980
0 30982 7 1 2 30977 30981
0 30983 5 1 1 30982
0 30984 7 1 2 72402 30983
0 30985 5 1 1 30984
0 30986 7 4 2 97123 102675
0 30987 7 1 2 83504 102718
0 30988 7 1 2 97669 30987
0 30989 5 1 1 30988
0 30990 7 1 2 30985 30989
0 30991 5 1 1 30990
0 30992 7 1 2 71665 30991
0 30993 5 1 1 30992
0 30994 7 1 2 68076 94944
0 30995 7 2 2 99576 80446
0 30996 7 2 2 102498 97473
0 30997 7 1 2 102722 102724
0 30998 7 1 2 30994 30997
0 30999 5 1 1 30998
0 31000 7 1 2 30993 30999
0 31001 5 1 1 31000
0 31002 7 1 2 68421 31001
0 31003 5 1 1 31002
0 31004 7 1 2 84117 96495
0 31005 5 1 1 31004
0 31006 7 1 2 102662 31005
0 31007 5 1 1 31006
0 31008 7 2 2 70825 89726
0 31009 7 4 2 70457 67186
0 31010 7 1 2 69183 102728
0 31011 7 1 2 97289 31010
0 31012 7 1 2 102726 31011
0 31013 5 1 1 31012
0 31014 7 1 2 31007 31013
0 31015 5 1 1 31014
0 31016 7 1 2 97233 31015
0 31017 5 1 1 31016
0 31018 7 1 2 31003 31017
0 31019 5 1 1 31018
0 31020 7 1 2 71408 31019
0 31021 5 1 1 31020
0 31022 7 9 2 102388 97474
0 31023 5 3 1 102732
0 31024 7 13 2 72157 67333
0 31025 7 4 2 102744 102407
0 31026 5 1 1 102757
0 31027 7 1 2 102741 31026
0 31028 5 5 1 31027
0 31029 7 1 2 64124 102761
0 31030 5 2 1 31029
0 31031 7 10 2 67334 102676
0 31032 7 1 2 85438 102768
0 31033 5 1 1 31032
0 31034 7 1 2 102766 31033
0 31035 5 3 1 31034
0 31036 7 1 2 97342 102778
0 31037 5 1 1 31036
0 31038 7 2 2 84338 92822
0 31039 7 1 2 98026 102677
0 31040 7 1 2 102781 31039
0 31041 5 1 1 31040
0 31042 7 1 2 31037 31041
0 31043 5 1 1 31042
0 31044 7 1 2 71666 31043
0 31045 5 1 1 31044
0 31046 7 2 2 98027 102618
0 31047 7 1 2 98839 80209
0 31048 7 1 2 102783 31047
0 31049 5 1 1 31048
0 31050 7 1 2 31045 31049
0 31051 5 1 1 31050
0 31052 7 1 2 71409 31051
0 31053 5 1 1 31052
0 31054 7 1 2 81566 75850
0 31055 7 1 2 102779 31054
0 31056 5 1 1 31055
0 31057 7 1 2 31053 31056
0 31058 5 1 1 31057
0 31059 7 1 2 68422 31058
0 31060 5 1 1 31059
0 31061 7 2 2 72403 74741
0 31062 7 3 2 70458 93214
0 31063 7 1 2 96866 102619
0 31064 7 1 2 102787 31063
0 31065 7 1 2 102785 31064
0 31066 5 1 1 31065
0 31067 7 1 2 31060 31066
0 31068 5 1 1 31067
0 31069 7 1 2 82980 31068
0 31070 5 1 1 31069
0 31071 7 7 2 69184 72158
0 31072 7 5 2 67187 102790
0 31073 7 1 2 97923 30547
0 31074 5 1 1 31073
0 31075 7 1 2 102797 31074
0 31076 5 1 1 31075
0 31077 7 1 2 102767 31076
0 31078 5 1 1 31077
0 31079 7 1 2 76029 80093
0 31080 7 1 2 83581 31079
0 31081 7 1 2 31078 31080
0 31082 5 1 1 31081
0 31083 7 1 2 31070 31082
0 31084 7 1 2 31021 31083
0 31085 5 1 1 31084
0 31086 7 1 2 100284 31085
0 31087 5 1 1 31086
0 31088 7 5 2 67335 68423
0 31089 7 2 2 67188 102802
0 31090 7 2 2 102807 96299
0 31091 5 1 1 102809
0 31092 7 4 2 72243 98373
0 31093 7 1 2 67114 80202
0 31094 7 1 2 102811 31093
0 31095 5 1 1 31094
0 31096 7 1 2 31091 31095
0 31097 5 1 1 31096
0 31098 7 1 2 64125 31097
0 31099 5 1 1 31098
0 31100 7 6 2 68424 98493
0 31101 7 1 2 102815 102798
0 31102 5 1 1 31101
0 31103 7 1 2 31099 31102
0 31104 5 1 1 31103
0 31105 7 1 2 70459 31104
0 31106 5 1 1 31105
0 31107 7 5 2 71833 67189
0 31108 7 2 2 77729 102821
0 31109 7 1 2 99476 102826
0 31110 5 1 1 31109
0 31111 7 1 2 31106 31110
0 31112 5 1 1 31111
0 31113 7 3 2 93588 91852
0 31114 7 1 2 31112 102828
0 31115 5 1 1 31114
0 31116 7 1 2 67666 31115
0 31117 7 1 2 31087 31116
0 31118 5 1 1 31117
0 31119 7 2 2 99566 102704
0 31120 5 1 1 102831
0 31121 7 1 2 102671 31120
0 31122 5 1 1 31121
0 31123 7 1 2 89610 93949
0 31124 5 1 1 31123
0 31125 7 1 2 31122 31124
0 31126 5 1 1 31125
0 31127 7 1 2 87700 102660
0 31128 5 2 1 31127
0 31129 7 4 2 69185 74171
0 31130 7 1 2 101442 90148
0 31131 7 1 2 102835 31130
0 31132 5 1 1 31131
0 31133 7 1 2 102833 31132
0 31134 5 1 1 31133
0 31135 7 2 2 80412 31134
0 31136 5 1 1 102839
0 31137 7 1 2 31126 31136
0 31138 5 1 1 31137
0 31139 7 1 2 76030 31138
0 31140 5 1 1 31139
0 31141 7 4 2 82440 102678
0 31142 7 1 2 101686 96817
0 31143 5 1 1 31142
0 31144 7 1 2 70460 31143
0 31145 5 1 1 31144
0 31146 7 2 2 86139 74855
0 31147 5 1 1 102845
0 31148 7 1 2 96808 31147
0 31149 7 1 2 31145 31148
0 31150 7 1 2 100865 31149
0 31151 5 1 1 31150
0 31152 7 1 2 102841 31151
0 31153 5 1 1 31152
0 31154 7 5 2 80707 80937
0 31155 7 1 2 83813 102847
0 31156 5 1 1 31155
0 31157 7 1 2 98320 31156
0 31158 5 1 1 31157
0 31159 7 1 2 102663 31158
0 31160 5 1 1 31159
0 31161 7 1 2 66312 31160
0 31162 7 1 2 31153 31161
0 31163 5 1 1 31162
0 31164 7 1 2 87642 102664
0 31165 5 1 1 31164
0 31166 7 1 2 82373 90114
0 31167 7 1 2 102832 31166
0 31168 5 1 1 31167
0 31169 7 1 2 31165 31168
0 31170 5 1 1 31169
0 31171 7 1 2 66559 31170
0 31172 5 1 1 31171
0 31173 7 2 2 71667 102842
0 31174 7 1 2 65441 102852
0 31175 5 1 1 31174
0 31176 7 1 2 102672 31175
0 31177 5 1 1 31176
0 31178 7 1 2 94011 31177
0 31179 5 1 1 31178
0 31180 7 1 2 31172 31179
0 31181 5 1 1 31180
0 31182 7 1 2 65130 31181
0 31183 5 1 1 31182
0 31184 7 1 2 65442 102834
0 31185 5 1 1 31184
0 31186 7 1 2 102840 31185
0 31187 5 1 1 31186
0 31188 7 1 2 78657 102717
0 31189 5 1 1 31188
0 31190 7 1 2 71410 31189
0 31191 7 1 2 31187 31190
0 31192 7 1 2 31183 31191
0 31193 5 1 1 31192
0 31194 7 1 2 73158 31193
0 31195 7 1 2 31163 31194
0 31196 5 1 1 31195
0 31197 7 1 2 31140 31196
0 31198 5 1 1 31197
0 31199 7 1 2 67336 31198
0 31200 5 1 1 31199
0 31201 7 9 2 67115 99629
0 31202 7 1 2 102504 102854
0 31203 7 1 2 94770 31202
0 31204 5 1 1 31203
0 31205 7 1 2 31200 31204
0 31206 5 1 1 31205
0 31207 7 1 2 100285 31206
0 31208 5 1 1 31207
0 31209 7 1 2 69186 102762
0 31210 5 1 1 31209
0 31211 7 1 2 85452 102855
0 31212 5 1 1 31211
0 31213 7 1 2 31210 31212
0 31214 5 1 1 31213
0 31215 7 1 2 85690 31214
0 31216 5 1 1 31215
0 31217 7 5 2 67337 102620
0 31218 7 1 2 88689 74397
0 31219 7 1 2 102863 31218
0 31220 5 1 1 31219
0 31221 7 1 2 31216 31220
0 31222 5 1 1 31221
0 31223 7 1 2 75012 31222
0 31224 5 1 1 31223
0 31225 7 1 2 102226 102621
0 31226 5 1 1 31225
0 31227 7 2 2 102705 102318
0 31228 5 1 1 102868
0 31229 7 1 2 31226 31228
0 31230 5 1 1 31229
0 31231 7 1 2 75921 31230
0 31232 5 1 1 31231
0 31233 7 1 2 31224 31232
0 31234 5 1 1 31233
0 31235 7 1 2 100216 31234
0 31236 5 1 1 31235
0 31237 7 1 2 72689 31236
0 31238 7 1 2 31208 31237
0 31239 5 1 1 31238
0 31240 7 1 2 68861 31239
0 31241 7 1 2 31118 31240
0 31242 5 1 1 31241
0 31243 7 1 2 30949 31242
0 31244 5 1 1 31243
0 31245 7 1 2 64752 31244
0 31246 5 1 1 31245
0 31247 7 1 2 30776 31246
0 31248 7 1 2 30469 31247
0 31249 5 1 1 31248
0 31250 7 1 2 72061 31249
0 31251 5 1 1 31250
0 31252 7 3 2 94779 96396
0 31253 7 2 2 91273 102870
0 31254 7 1 2 64753 89706
0 31255 5 2 1 31254
0 31256 7 1 2 86818 102875
0 31257 5 1 1 31256
0 31258 7 1 2 80617 31257
0 31259 5 1 1 31258
0 31260 7 1 2 88338 8842
0 31261 5 1 1 31260
0 31262 7 1 2 80708 31261
0 31263 5 1 1 31262
0 31264 7 1 2 81740 93334
0 31265 5 1 1 31264
0 31266 7 1 2 31263 31265
0 31267 7 1 2 31259 31266
0 31268 5 1 1 31267
0 31269 7 1 2 102873 31268
0 31270 5 1 1 31269
0 31271 7 3 2 73916 100004
0 31272 7 2 2 88898 79089
0 31273 7 1 2 65601 84953
0 31274 7 1 2 102880 31273
0 31275 7 1 2 102877 31274
0 31276 5 1 1 31275
0 31277 7 1 2 31270 31276
0 31278 5 1 1 31277
0 31279 7 1 2 72159 31278
0 31280 5 1 1 31279
0 31281 7 1 2 73966 83700
0 31282 5 2 1 31281
0 31283 7 1 2 86767 28437
0 31284 5 1 1 31283
0 31285 7 2 2 102882 31284
0 31286 5 1 1 102884
0 31287 7 3 2 64754 86779
0 31288 5 1 1 102886
0 31289 7 1 2 102885 31288
0 31290 5 2 1 31289
0 31291 7 4 2 67116 102259
0 31292 7 1 2 102891 102871
0 31293 7 1 2 102889 31292
0 31294 5 1 1 31293
0 31295 7 1 2 31280 31294
0 31296 5 1 1 31295
0 31297 7 1 2 71411 31296
0 31298 5 1 1 31297
0 31299 7 2 2 86780 82299
0 31300 5 1 1 102895
0 31301 7 1 2 86675 78698
0 31302 5 1 1 31301
0 31303 7 1 2 31300 31302
0 31304 5 1 1 31303
0 31305 7 1 2 102892 31304
0 31306 5 1 1 31305
0 31307 7 4 2 79841 91749
0 31308 5 9 1 102897
0 31309 7 1 2 80709 102901
0 31310 5 1 1 31309
0 31311 7 1 2 80618 94925
0 31312 5 2 1 31311
0 31313 7 1 2 100743 102910
0 31314 7 1 2 31310 31313
0 31315 5 1 1 31314
0 31316 7 1 2 98123 31315
0 31317 5 1 1 31316
0 31318 7 1 2 31306 31317
0 31319 5 1 1 31318
0 31320 7 1 2 66313 31319
0 31321 5 1 1 31320
0 31322 7 2 2 65443 102260
0 31323 7 1 2 69878 94803
0 31324 7 1 2 90092 31323
0 31325 7 1 2 102912 31324
0 31326 5 1 1 31325
0 31327 7 1 2 31321 31326
0 31328 5 1 1 31327
0 31329 7 1 2 102872 31328
0 31330 5 1 1 31329
0 31331 7 1 2 31298 31330
0 31332 5 1 1 31331
0 31333 7 1 2 63800 31332
0 31334 5 1 1 31333
0 31335 7 1 2 71412 102890
0 31336 5 1 1 31335
0 31337 7 1 2 66314 102896
0 31338 5 1 1 31337
0 31339 7 1 2 79028 82928
0 31340 5 2 1 31339
0 31341 7 1 2 101242 102914
0 31342 5 1 1 31341
0 31343 7 1 2 78699 31342
0 31344 5 1 1 31343
0 31345 7 1 2 31338 31344
0 31346 7 1 2 31336 31345
0 31347 5 1 1 31346
0 31348 7 2 2 93706 84471
0 31349 7 1 2 71945 102916
0 31350 7 1 2 102893 31349
0 31351 7 1 2 31347 31350
0 31352 5 1 1 31351
0 31353 7 1 2 67190 31352
0 31354 7 1 2 31334 31353
0 31355 5 1 1 31354
0 31356 7 3 2 89206 86449
0 31357 5 1 1 102918
0 31358 7 1 2 86304 102919
0 31359 5 2 1 31358
0 31360 7 6 2 79379 96686
0 31361 5 2 1 102923
0 31362 7 1 2 102921 102924
0 31363 5 1 1 31362
0 31364 7 8 2 102261 87272
0 31365 5 1 1 102931
0 31366 7 2 2 64755 80359
0 31367 5 2 1 102939
0 31368 7 1 2 2332 102941
0 31369 5 1 1 31368
0 31370 7 1 2 70461 31369
0 31371 5 1 1 31370
0 31372 7 1 2 90827 79197
0 31373 5 1 1 31372
0 31374 7 1 2 31371 31373
0 31375 5 1 1 31374
0 31376 7 1 2 102932 31375
0 31377 5 1 1 31376
0 31378 7 1 2 31363 31377
0 31379 5 1 1 31378
0 31380 7 1 2 71413 31379
0 31381 5 1 1 31380
0 31382 7 2 2 70462 84083
0 31383 7 2 2 94547 102943
0 31384 7 1 2 102945 102933
0 31385 5 1 1 31384
0 31386 7 1 2 31381 31385
0 31387 5 1 1 31386
0 31388 7 3 2 70633 65815
0 31389 7 2 2 71946 102947
0 31390 7 1 2 31387 102950
0 31391 5 1 1 31390
0 31392 7 4 2 70634 84488
0 31393 7 1 2 92381 102952
0 31394 7 1 2 102934 31393
0 31395 5 1 1 31394
0 31396 7 3 2 66315 92238
0 31397 7 1 2 101613 94004
0 31398 7 1 2 102956 31397
0 31399 5 1 1 31398
0 31400 7 1 2 31395 31399
0 31401 5 1 1 31400
0 31402 7 1 2 94758 31401
0 31403 5 1 1 31402
0 31404 7 1 2 95819 89639
0 31405 7 2 2 67117 78573
0 31406 7 2 2 66316 93671
0 31407 7 1 2 102959 102961
0 31408 7 1 2 31404 31407
0 31409 5 1 1 31408
0 31410 7 1 2 31403 31409
0 31411 7 1 2 31391 31410
0 31412 5 1 1 31411
0 31413 7 1 2 64126 31412
0 31414 5 1 1 31413
0 31415 7 2 2 65816 101783
0 31416 7 1 2 64756 102957
0 31417 7 1 2 102963 31416
0 31418 7 1 2 94766 31417
0 31419 5 1 1 31418
0 31420 7 1 2 31414 31419
0 31421 5 1 1 31420
0 31422 7 1 2 65131 31421
0 31423 5 1 1 31422
0 31424 7 2 2 69879 80792
0 31425 5 1 1 102965
0 31426 7 1 2 88667 102966
0 31427 5 1 1 31426
0 31428 7 1 2 68668 91738
0 31429 5 1 1 31428
0 31430 7 1 2 86646 31429
0 31431 5 1 1 31430
0 31432 7 1 2 70463 31431
0 31433 5 1 1 31432
0 31434 7 1 2 75399 86750
0 31435 5 1 1 31434
0 31436 7 1 2 31433 31435
0 31437 5 1 1 31436
0 31438 7 1 2 64757 31437
0 31439 5 1 1 31438
0 31440 7 1 2 73745 79884
0 31441 5 1 1 31440
0 31442 7 1 2 91948 83166
0 31443 5 1 1 31442
0 31444 7 1 2 78574 86169
0 31445 5 1 1 31444
0 31446 7 1 2 31443 31445
0 31447 5 1 1 31446
0 31448 7 1 2 66754 31447
0 31449 5 1 1 31448
0 31450 7 1 2 31441 31449
0 31451 7 1 2 31439 31450
0 31452 5 1 1 31451
0 31453 7 1 2 71414 31452
0 31454 5 1 1 31453
0 31455 7 1 2 31427 31454
0 31456 5 1 1 31455
0 31457 7 1 2 102935 31456
0 31458 5 1 1 31457
0 31459 7 1 2 85741 83869
0 31460 7 1 2 7979 31459
0 31461 5 1 1 31460
0 31462 7 1 2 64758 85800
0 31463 5 1 1 31462
0 31464 7 1 2 31461 31463
0 31465 5 1 1 31464
0 31466 7 1 2 102925 31465
0 31467 5 1 1 31466
0 31468 7 1 2 31458 31467
0 31469 5 1 1 31468
0 31470 7 3 2 70635 82775
0 31471 7 1 2 64127 102967
0 31472 7 1 2 31469 31471
0 31473 5 1 1 31472
0 31474 7 1 2 99774 94032
0 31475 7 2 2 77905 96278
0 31476 7 1 2 101829 102970
0 31477 7 1 2 31474 31476
0 31478 5 1 1 31477
0 31479 7 2 2 72160 93043
0 31480 7 2 2 88029 82776
0 31481 7 1 2 102972 102974
0 31482 7 1 2 102876 31481
0 31483 7 1 2 4220 31482
0 31484 5 1 1 31483
0 31485 7 1 2 31478 31484
0 31486 5 1 1 31485
0 31487 7 1 2 65444 31486
0 31488 5 1 1 31487
0 31489 7 1 2 64759 88832
0 31490 5 2 1 31489
0 31491 7 1 2 75400 94551
0 31492 7 1 2 102976 31491
0 31493 5 1 1 31492
0 31494 7 1 2 74546 84120
0 31495 5 1 1 31494
0 31496 7 1 2 76697 100491
0 31497 5 1 1 31496
0 31498 7 1 2 69880 31497
0 31499 5 1 1 31498
0 31500 7 1 2 31495 31499
0 31501 7 1 2 31493 31500
0 31502 5 1 1 31501
0 31503 7 1 2 98828 92861
0 31504 7 1 2 102975 31503
0 31505 7 1 2 31502 31504
0 31506 5 1 1 31505
0 31507 7 1 2 31488 31506
0 31508 5 1 1 31507
0 31509 7 1 2 63905 31508
0 31510 5 1 1 31509
0 31511 7 1 2 79039 102035
0 31512 5 3 1 31511
0 31513 7 2 2 65649 87273
0 31514 7 1 2 102978 102981
0 31515 5 1 1 31514
0 31516 7 4 2 67118 81887
0 31517 7 1 2 90364 102983
0 31518 5 1 1 31517
0 31519 7 1 2 31515 31518
0 31520 5 1 1 31519
0 31521 7 1 2 68425 31520
0 31522 5 1 1 31521
0 31523 7 2 2 83701 96693
0 31524 7 1 2 90717 102987
0 31525 5 1 1 31524
0 31526 7 1 2 31522 31525
0 31527 5 1 1 31526
0 31528 7 1 2 75401 31527
0 31529 5 1 1 31528
0 31530 7 1 2 102988 98844
0 31531 5 1 1 31530
0 31532 7 3 2 67119 90365
0 31533 7 1 2 85753 102989
0 31534 5 1 1 31533
0 31535 7 1 2 31531 31534
0 31536 5 1 1 31535
0 31537 7 1 2 76654 31536
0 31538 5 1 1 31537
0 31539 7 1 2 80801 8767
0 31540 5 1 1 31539
0 31541 7 1 2 88677 102982
0 31542 7 1 2 31540 31541
0 31543 5 1 1 31542
0 31544 7 1 2 31538 31543
0 31545 7 1 2 31529 31544
0 31546 5 1 1 31545
0 31547 7 3 2 84322 102951
0 31548 7 1 2 31546 102992
0 31549 5 1 1 31548
0 31550 7 1 2 31510 31549
0 31551 5 1 1 31550
0 31552 7 1 2 66317 31551
0 31553 5 1 1 31552
0 31554 7 1 2 72244 31553
0 31555 7 1 2 31473 31554
0 31556 7 1 2 31423 31555
0 31557 5 1 1 31556
0 31558 7 1 2 31355 31557
0 31559 5 1 1 31558
0 31560 7 1 2 68077 31559
0 31561 5 1 1 31560
0 31562 7 1 2 73917 77805
0 31563 5 2 1 31562
0 31564 7 4 2 100709 93755
0 31565 5 1 1 102997
0 31566 7 1 2 69881 102998
0 31567 5 1 1 31566
0 31568 7 2 2 102995 31567
0 31569 5 3 1 103001
0 31570 7 1 2 84428 103003
0 31571 5 1 1 31570
0 31572 7 1 2 85509 81174
0 31573 7 1 2 89822 31572
0 31574 5 1 1 31573
0 31575 7 1 2 31571 31574
0 31576 5 1 1 31575
0 31577 7 1 2 73746 31576
0 31578 5 1 1 31577
0 31579 7 1 2 70204 79936
0 31580 7 1 2 98153 31579
0 31581 5 1 1 31580
0 31582 7 1 2 31578 31581
0 31583 5 1 1 31582
0 31584 7 1 2 102569 31583
0 31585 5 1 1 31584
0 31586 7 1 2 71415 95581
0 31587 5 1 1 31586
0 31588 7 1 2 84201 31587
0 31589 5 1 1 31588
0 31590 7 1 2 102984 102408
0 31591 7 2 2 31589 31590
0 31592 7 1 2 97329 103006
0 31593 5 1 1 31592
0 31594 7 1 2 31585 31593
0 31595 5 1 1 31594
0 31596 7 1 2 68862 31595
0 31597 5 1 1 31596
0 31598 7 1 2 103007 94786
0 31599 5 1 1 31598
0 31600 7 1 2 31597 31599
0 31601 5 1 1 31600
0 31602 7 1 2 71947 31601
0 31603 5 1 1 31602
0 31604 7 4 2 65817 102572
0 31605 7 1 2 98148 79792
0 31606 7 1 2 103004 31605
0 31607 5 1 1 31606
0 31608 7 1 2 93617 79793
0 31609 5 1 1 31608
0 31610 7 1 2 79561 81175
0 31611 7 1 2 78867 31610
0 31612 5 1 1 31611
0 31613 7 1 2 31609 31612
0 31614 5 1 1 31613
0 31615 7 1 2 66560 31614
0 31616 5 1 1 31615
0 31617 7 1 2 862 80802
0 31618 5 1 1 31617
0 31619 7 1 2 79535 98096
0 31620 7 1 2 31618 31619
0 31621 5 1 1 31620
0 31622 7 1 2 31616 31621
0 31623 5 1 1 31622
0 31624 7 1 2 80619 31623
0 31625 5 1 1 31624
0 31626 7 1 2 98324 98097
0 31627 5 1 1 31626
0 31628 7 1 2 66877 87257
0 31629 7 1 2 87444 31628
0 31630 5 1 1 31629
0 31631 7 1 2 31627 31630
0 31632 5 1 1 31631
0 31633 7 1 2 97402 31632
0 31634 5 1 1 31633
0 31635 7 1 2 31625 31634
0 31636 7 1 2 31607 31635
0 31637 5 1 1 31636
0 31638 7 1 2 103008 31637
0 31639 5 1 1 31638
0 31640 7 7 2 67191 82441
0 31641 7 2 2 71948 84564
0 31642 7 1 2 103012 103019
0 31643 7 1 2 101482 31642
0 31644 5 1 1 31643
0 31645 7 1 2 31639 31644
0 31646 5 1 1 31645
0 31647 7 1 2 68669 31646
0 31648 5 1 1 31647
0 31649 7 1 2 31603 31648
0 31650 5 1 1 31649
0 31651 7 1 2 102262 31650
0 31652 5 1 1 31651
0 31653 7 1 2 82318 91783
0 31654 5 1 1 31653
0 31655 7 2 2 76415 87513
0 31656 5 2 1 103021
0 31657 7 1 2 99819 103023
0 31658 5 1 1 31657
0 31659 7 1 2 86943 31658
0 31660 5 1 1 31659
0 31661 7 1 2 31654 31660
0 31662 5 1 1 31661
0 31663 7 1 2 64760 31662
0 31664 5 1 1 31663
0 31665 7 1 2 100602 101473
0 31666 5 1 1 31665
0 31667 7 1 2 95067 77046
0 31668 7 1 2 86944 31667
0 31669 5 1 1 31668
0 31670 7 1 2 31666 31669
0 31671 7 1 2 31664 31670
0 31672 5 1 1 31671
0 31673 7 1 2 100217 31672
0 31674 5 1 1 31673
0 31675 7 1 2 96397 76004
0 31676 7 1 2 82228 31675
0 31677 7 1 2 101599 31676
0 31678 5 1 1 31677
0 31679 7 1 2 31674 31678
0 31680 5 1 1 31679
0 31681 7 1 2 64128 31680
0 31682 5 1 1 31681
0 31683 7 1 2 81640 100869
0 31684 5 1 1 31683
0 31685 7 1 2 94219 86945
0 31686 5 1 1 31685
0 31687 7 1 2 73510 100603
0 31688 5 1 1 31687
0 31689 7 2 2 31686 31688
0 31690 5 1 1 103025
0 31691 7 1 2 93589 93069
0 31692 7 1 2 31690 31691
0 31693 5 1 1 31692
0 31694 7 1 2 31684 31693
0 31695 5 1 1 31694
0 31696 7 1 2 69882 31695
0 31697 5 1 1 31696
0 31698 7 1 2 71416 103026
0 31699 5 1 1 31698
0 31700 7 1 2 73511 88690
0 31701 7 1 2 93815 31700
0 31702 5 1 1 31701
0 31703 7 1 2 86305 31702
0 31704 5 1 1 31703
0 31705 7 1 2 71668 31704
0 31706 5 1 1 31705
0 31707 7 1 2 85629 96801
0 31708 5 1 1 31707
0 31709 7 1 2 66318 101731
0 31710 7 1 2 31708 31709
0 31711 7 1 2 31706 31710
0 31712 5 1 1 31711
0 31713 7 1 2 100652 31712
0 31714 7 1 2 31699 31713
0 31715 5 1 1 31714
0 31716 7 1 2 76326 80917
0 31717 5 1 1 31716
0 31718 7 1 2 84202 31717
0 31719 5 1 1 31718
0 31720 7 1 2 100870 31719
0 31721 5 1 1 31720
0 31722 7 1 2 90828 75059
0 31723 7 1 2 100653 31722
0 31724 5 1 1 31723
0 31725 7 1 2 31721 31724
0 31726 5 1 1 31725
0 31727 7 1 2 81888 31726
0 31728 5 1 1 31727
0 31729 7 2 2 99558 93747
0 31730 7 2 2 76226 103027
0 31731 5 1 1 103029
0 31732 7 1 2 74136 75029
0 31733 5 1 1 31732
0 31734 7 1 2 31731 31733
0 31735 5 1 1 31734
0 31736 7 1 2 100286 31735
0 31737 5 1 1 31736
0 31738 7 1 2 31728 31737
0 31739 7 1 2 31715 31738
0 31740 7 1 2 31697 31739
0 31741 5 1 1 31740
0 31742 7 1 2 65818 31741
0 31743 5 1 1 31742
0 31744 7 1 2 31682 31743
0 31745 5 1 1 31744
0 31746 7 1 2 102622 31745
0 31747 5 1 1 31746
0 31748 7 1 2 80620 26383
0 31749 5 1 1 31748
0 31750 7 2 2 76592 80710
0 31751 5 1 1 103031
0 31752 7 1 2 75402 31751
0 31753 7 1 2 31749 31752
0 31754 5 1 1 31753
0 31755 7 1 2 97812 97547
0 31756 5 2 1 31755
0 31757 7 1 2 76485 103033
0 31758 5 1 1 31757
0 31759 7 1 2 83457 97548
0 31760 5 2 1 31759
0 31761 7 1 2 103035 92655
0 31762 5 1 1 31761
0 31763 7 1 2 31758 31762
0 31764 7 1 2 31754 31763
0 31765 5 1 1 31764
0 31766 7 1 2 102874 102679
0 31767 7 1 2 31765 31766
0 31768 5 1 1 31767
0 31769 7 1 2 31747 31768
0 31770 5 1 1 31769
0 31771 7 1 2 63801 31770
0 31772 5 1 1 31771
0 31773 7 1 2 73159 31772
0 31774 7 1 2 31652 31773
0 31775 5 1 1 31774
0 31776 7 1 2 31561 31775
0 31777 5 1 1 31776
0 31778 7 4 2 64129 70686
0 31779 7 2 2 70636 103037
0 31780 7 2 2 102652 103041
0 31781 7 1 2 79380 81504
0 31782 7 1 2 103043 31781
0 31783 5 1 1 31782
0 31784 7 2 2 82442 74033
0 31785 7 1 2 78700 102542
0 31786 7 1 2 103045 31785
0 31787 5 1 1 31786
0 31788 7 6 2 72245 73512
0 31789 7 2 2 72161 103047
0 31790 7 1 2 92840 92980
0 31791 7 1 2 93308 31790
0 31792 7 1 2 103053 31791
0 31793 5 1 1 31792
0 31794 7 1 2 31787 31793
0 31795 5 1 1 31794
0 31796 7 1 2 73747 102263
0 31797 7 1 2 31795 31796
0 31798 5 1 1 31797
0 31799 7 1 2 31783 31798
0 31800 5 1 1 31799
0 31801 7 3 2 71417 79029
0 31802 7 1 2 86402 103055
0 31803 7 1 2 31800 31802
0 31804 5 1 1 31803
0 31805 7 1 2 31777 31804
0 31806 5 1 1 31805
0 31807 7 1 2 67667 31806
0 31808 5 1 1 31807
0 31809 7 1 2 82285 102926
0 31810 5 1 1 31809
0 31811 7 1 2 86676 102936
0 31812 5 1 1 31811
0 31813 7 1 2 31810 31812
0 31814 5 1 1 31813
0 31815 7 1 2 73918 31814
0 31816 5 1 1 31815
0 31817 7 1 2 102990 87599
0 31818 7 1 2 87465 31817
0 31819 5 1 1 31818
0 31820 7 1 2 31816 31819
0 31821 5 1 1 31820
0 31822 7 1 2 102499 31821
0 31823 5 1 1 31822
0 31824 7 3 2 69187 71834
0 31825 7 1 2 68991 90366
0 31826 7 1 2 103058 31825
0 31827 7 3 2 68670 102680
0 31828 7 1 2 100386 103061
0 31829 7 1 2 31826 31828
0 31830 5 1 1 31829
0 31831 7 1 2 31823 31830
0 31832 5 1 1 31831
0 31833 7 1 2 82725 31832
0 31834 5 1 1 31833
0 31835 7 3 2 72246 73160
0 31836 7 1 2 65445 79842
0 31837 7 1 2 102991 31836
0 31838 5 1 1 31837
0 31839 7 3 2 72162 74666
0 31840 7 1 2 68863 100879
0 31841 7 1 2 103067 31840
0 31842 5 1 1 31841
0 31843 7 1 2 31838 31842
0 31844 5 1 1 31843
0 31845 7 1 2 68992 31844
0 31846 5 1 1 31845
0 31847 7 1 2 74667 96430
0 31848 7 1 2 101900 31847
0 31849 5 1 1 31848
0 31850 7 1 2 31846 31849
0 31851 5 1 1 31850
0 31852 7 1 2 85510 80413
0 31853 7 1 2 31851 31852
0 31854 5 1 1 31853
0 31855 7 4 2 68864 102264
0 31856 7 1 2 85511 103068
0 31857 7 2 2 103070 31856
0 31858 7 1 2 96001 103074
0 31859 5 1 1 31858
0 31860 7 1 2 103071 78112
0 31861 5 1 1 31860
0 31862 7 1 2 102929 31861
0 31863 5 1 1 31862
0 31864 7 2 2 85512 79843
0 31865 7 1 2 82929 103076
0 31866 7 1 2 31863 31865
0 31867 5 1 1 31866
0 31868 7 1 2 31859 31867
0 31869 7 1 2 31854 31868
0 31870 5 1 1 31869
0 31871 7 1 2 73513 31870
0 31872 5 1 1 31871
0 31873 7 3 2 96002 82930
0 31874 7 1 2 103078 103075
0 31875 5 1 1 31874
0 31876 7 1 2 31872 31875
0 31877 5 1 1 31876
0 31878 7 1 2 103064 31877
0 31879 5 1 1 31878
0 31880 7 1 2 31834 31879
0 31881 5 1 1 31880
0 31882 7 1 2 70637 31881
0 31883 5 1 1 31882
0 31884 7 1 2 63802 102706
0 31885 7 2 2 100409 31884
0 31886 5 1 1 103081
0 31887 7 3 2 70638 72247
0 31888 7 2 2 92862 103083
0 31889 7 1 2 92841 103086
0 31890 5 1 1 31889
0 31891 7 1 2 31890 102563
0 31892 5 1 1 31891
0 31893 7 1 2 68865 31892
0 31894 5 1 1 31893
0 31895 7 1 2 102557 94787
0 31896 5 1 1 31895
0 31897 7 1 2 31894 31896
0 31898 5 1 1 31897
0 31899 7 2 2 102265 31898
0 31900 5 1 1 103088
0 31901 7 1 2 70464 103089
0 31902 5 1 1 31901
0 31903 7 1 2 31886 31902
0 31904 5 1 1 31903
0 31905 7 1 2 82726 80536
0 31906 7 1 2 31904 31905
0 31907 5 1 1 31906
0 31908 7 1 2 31883 31907
0 31909 5 1 1 31908
0 31910 7 1 2 71418 31909
0 31911 5 1 1 31910
0 31912 7 1 2 101852 102615
0 31913 5 1 1 31912
0 31914 7 1 2 31900 31913
0 31915 5 1 1 31914
0 31916 7 1 2 68426 31915
0 31917 5 1 1 31916
0 31918 7 1 2 70465 103082
0 31919 5 1 1 31918
0 31920 7 1 2 31917 31919
0 31921 5 1 1 31920
0 31922 7 1 2 71669 31921
0 31923 5 1 1 31922
0 31924 7 2 2 69188 70687
0 31925 5 1 1 103090
0 31926 7 2 2 96548 103091
0 31927 7 2 2 90649 75711
0 31928 7 4 2 68427 102681
0 31929 7 1 2 103094 103096
0 31930 7 1 2 103092 31929
0 31931 5 1 1 31930
0 31932 7 1 2 31923 31931
0 31933 5 1 1 31932
0 31934 7 1 2 77540 31933
0 31935 5 1 1 31934
0 31936 7 1 2 98215 102623
0 31937 7 1 2 85513 31936
0 31938 7 1 2 79988 95724
0 31939 7 1 2 31937 31938
0 31940 7 1 2 2677 31939
0 31941 5 1 1 31940
0 31942 7 1 2 31935 31941
0 31943 5 1 1 31942
0 31944 7 1 2 82981 31943
0 31945 5 1 1 31944
0 31946 7 4 2 85691 80525
0 31947 7 1 2 75013 103100
0 31948 5 1 1 31947
0 31949 7 3 2 73161 97541
0 31950 7 1 2 73748 103104
0 31951 5 1 1 31950
0 31952 7 1 2 31948 31951
0 31953 5 1 1 31952
0 31954 7 1 2 65132 31953
0 31955 5 1 1 31954
0 31956 7 1 2 66319 94493
0 31957 5 1 1 31956
0 31958 7 1 2 31955 31957
0 31959 5 1 1 31958
0 31960 7 1 2 64761 31959
0 31961 5 1 1 31960
0 31962 7 1 2 80711 76687
0 31963 5 1 1 31962
0 31964 7 1 2 68671 101803
0 31965 5 1 1 31964
0 31966 7 1 2 31963 31965
0 31967 5 1 1 31966
0 31968 7 1 2 79989 31967
0 31969 5 1 1 31968
0 31970 7 1 2 78909 82177
0 31971 5 1 1 31970
0 31972 7 1 2 81741 83386
0 31973 7 1 2 31971 31972
0 31974 5 1 1 31973
0 31975 7 1 2 31969 31974
0 31976 5 1 1 31975
0 31977 7 1 2 66561 31976
0 31978 5 1 1 31977
0 31979 7 1 2 31961 31978
0 31980 5 1 1 31979
0 31981 7 1 2 102927 31980
0 31982 5 1 1 31981
0 31983 7 1 2 69883 94759
0 31984 5 1 1 31983
0 31985 7 1 2 102036 31984
0 31986 5 1 1 31985
0 31987 7 1 2 74668 31986
0 31988 5 1 1 31987
0 31989 7 2 2 80621 79844
0 31990 5 1 1 103107
0 31991 7 1 2 82114 103108
0 31992 5 1 1 31991
0 31993 7 1 2 73514 88437
0 31994 5 1 1 31993
0 31995 7 1 2 74904 78035
0 31996 7 1 2 31994 31995
0 31997 5 1 1 31996
0 31998 7 1 2 31992 31997
0 31999 7 1 2 31988 31998
0 32000 5 2 1 31999
0 32001 7 1 2 73162 103109
0 32002 5 1 1 32001
0 32003 7 1 2 101812 86600
0 32004 5 1 1 32003
0 32005 7 1 2 77294 93798
0 32006 5 1 1 32005
0 32007 7 2 2 73515 32006
0 32008 5 1 1 103111
0 32009 7 1 2 81321 83167
0 32010 7 1 2 97948 32009
0 32011 5 1 1 32010
0 32012 7 1 2 32008 32011
0 32013 5 1 1 32012
0 32014 7 1 2 64762 32013
0 32015 5 1 1 32014
0 32016 7 1 2 32015 16505
0 32017 5 1 1 32016
0 32018 7 1 2 68078 32017
0 32019 5 1 1 32018
0 32020 7 1 2 32004 32019
0 32021 7 1 2 32002 32020
0 32022 5 1 1 32021
0 32023 7 1 2 66320 32022
0 32024 5 1 1 32023
0 32025 7 1 2 75279 79185
0 32026 5 2 1 32025
0 32027 7 1 2 73163 80973
0 32028 5 1 1 32027
0 32029 7 1 2 103113 32028
0 32030 5 1 1 32029
0 32031 7 1 2 64763 32030
0 32032 5 1 1 32031
0 32033 7 1 2 87688 32032
0 32034 5 2 1 32033
0 32035 7 1 2 83702 103115
0 32036 5 2 1 32035
0 32037 7 4 2 65133 98976
0 32038 5 3 1 103119
0 32039 7 1 2 101830 103120
0 32040 5 1 1 32039
0 32041 7 1 2 103117 32040
0 32042 7 1 2 32024 32041
0 32043 5 1 1 32042
0 32044 7 1 2 102937 32043
0 32045 5 1 1 32044
0 32046 7 1 2 31982 32045
0 32047 5 1 1 32046
0 32048 7 1 2 85514 103084
0 32049 7 1 2 32047 32048
0 32050 5 1 1 32049
0 32051 7 1 2 31945 32050
0 32052 7 1 2 31911 32051
0 32053 5 1 1 32052
0 32054 7 1 2 71949 32053
0 32055 5 1 1 32054
0 32056 7 1 2 98793 77672
0 32057 5 1 1 32056
0 32058 7 2 2 65134 85692
0 32059 5 1 1 103126
0 32060 7 1 2 82498 76160
0 32061 7 1 2 103127 32060
0 32062 5 1 1 32061
0 32063 7 1 2 32057 32062
0 32064 5 1 1 32063
0 32065 7 1 2 71419 32064
0 32066 5 1 1 32065
0 32067 7 1 2 95101 95917
0 32068 5 1 1 32067
0 32069 7 1 2 32066 32068
0 32070 5 1 1 32069
0 32071 7 1 2 66562 32070
0 32072 5 1 1 32071
0 32073 7 1 2 82499 82931
0 32074 7 1 2 78804 32073
0 32075 7 1 2 83486 32074
0 32076 5 1 1 32075
0 32077 7 1 2 32072 32076
0 32078 5 1 1 32077
0 32079 7 1 2 69884 32078
0 32080 5 1 1 32079
0 32081 7 1 2 76048 83803
0 32082 5 1 1 32081
0 32083 7 1 2 102361 32082
0 32084 5 1 1 32083
0 32085 7 1 2 99626 32084
0 32086 5 1 1 32085
0 32087 7 1 2 99618 101517
0 32088 5 1 1 32087
0 32089 7 1 2 32086 32088
0 32090 5 1 1 32089
0 32091 7 1 2 71670 32090
0 32092 5 1 1 32091
0 32093 7 1 2 99775 96560
0 32094 7 1 2 99960 32093
0 32095 5 1 1 32094
0 32096 7 1 2 32092 32095
0 32097 5 1 1 32096
0 32098 7 1 2 68428 32097
0 32099 5 1 1 32098
0 32100 7 1 2 32080 32099
0 32101 5 1 1 32100
0 32102 7 3 2 72248 90590
0 32103 7 1 2 95921 103128
0 32104 7 1 2 32101 32103
0 32105 5 1 1 32104
0 32106 7 1 2 102389 92239
0 32107 7 1 2 93968 32106
0 32108 7 2 2 70466 90591
0 32109 7 1 2 89640 103131
0 32110 7 1 2 80108 32109
0 32111 7 1 2 32107 32110
0 32112 5 1 1 32111
0 32113 7 1 2 32105 32112
0 32114 7 1 2 32055 32113
0 32115 5 1 1 32114
0 32116 7 1 2 72690 32115
0 32117 5 1 1 32116
0 32118 7 10 2 102266 74034
0 32119 7 5 2 71950 67192
0 32120 7 1 2 100164 103143
0 32121 7 1 2 83957 32120
0 32122 7 1 2 100161 95167
0 32123 7 1 2 32121 32122
0 32124 7 1 2 103133 32123
0 32125 5 1 1 32124
0 32126 7 1 2 32117 32125
0 32127 7 1 2 31808 32126
0 32128 5 1 1 32127
0 32129 7 1 2 72404 32128
0 32130 5 1 1 32129
0 32131 7 3 2 63803 72163
0 32132 7 1 2 88396 78036
0 32133 5 1 1 32132
0 32134 7 1 2 100871 82300
0 32135 7 1 2 32133 32134
0 32136 5 2 1 32135
0 32137 7 2 2 89632 101799
0 32138 7 1 2 73749 103153
0 32139 7 1 2 87472 32138
0 32140 5 1 1 32139
0 32141 7 1 2 103151 32140
0 32142 5 1 1 32141
0 32143 7 1 2 68079 32142
0 32144 5 1 1 32143
0 32145 7 1 2 82356 83968
0 32146 5 2 1 32145
0 32147 7 2 2 69885 83703
0 32148 7 1 2 73516 103157
0 32149 5 1 1 32148
0 32150 7 1 2 103155 32149
0 32151 5 1 1 32150
0 32152 7 1 2 66563 32151
0 32153 5 1 1 32152
0 32154 7 2 2 99436 74879
0 32155 5 1 1 103159
0 32156 7 1 2 83969 103160
0 32157 5 1 1 32156
0 32158 7 1 2 32153 32157
0 32159 5 1 1 32158
0 32160 7 1 2 65135 32159
0 32161 5 1 1 32160
0 32162 7 1 2 66564 83970
0 32163 7 1 2 86932 32162
0 32164 5 1 1 32163
0 32165 7 1 2 32161 32164
0 32166 5 1 1 32165
0 32167 7 1 2 102014 32166
0 32168 5 1 1 32167
0 32169 7 1 2 32144 32168
0 32170 5 1 1 32169
0 32171 7 1 2 66321 32170
0 32172 5 1 1 32171
0 32173 7 1 2 78658 83704
0 32174 7 1 2 103154 32173
0 32175 5 1 1 32174
0 32176 7 1 2 103152 32175
0 32177 5 1 1 32176
0 32178 7 1 2 76049 32177
0 32179 5 1 1 32178
0 32180 7 1 2 100761 86033
0 32181 5 1 1 32180
0 32182 7 1 2 4770 32181
0 32183 5 1 1 32182
0 32184 7 2 2 93606 84074
0 32185 7 1 2 71671 94588
0 32186 7 1 2 103161 32185
0 32187 7 1 2 32183 32186
0 32188 5 1 1 32187
0 32189 7 1 2 32179 32188
0 32190 7 1 2 32172 32189
0 32191 5 1 1 32190
0 32192 7 1 2 67668 32191
0 32193 5 1 1 32192
0 32194 7 2 2 71951 86053
0 32195 7 1 2 100238 103162
0 32196 7 1 2 103163 32195
0 32197 5 1 1 32196
0 32198 7 5 2 65136 97403
0 32199 7 1 2 100218 83705
0 32200 7 1 2 103165 32199
0 32201 5 1 1 32200
0 32202 7 1 2 32197 32201
0 32203 5 1 1 32202
0 32204 7 1 2 73919 32203
0 32205 5 1 1 32204
0 32206 7 2 2 75783 78659
0 32207 5 1 1 103170
0 32208 7 3 2 65137 86610
0 32209 7 1 2 102881 103172
0 32210 7 1 2 103171 32209
0 32211 5 1 1 32210
0 32212 7 1 2 32205 32211
0 32213 5 1 1 32212
0 32214 7 1 2 85012 32213
0 32215 5 1 1 32214
0 32216 7 1 2 32193 32215
0 32217 5 1 1 32216
0 32218 7 1 2 70826 32217
0 32219 5 1 1 32218
0 32220 7 1 2 79173 102049
0 32221 5 1 1 32220
0 32222 7 2 2 93091 74333
0 32223 5 3 1 103175
0 32224 7 1 2 69189 103176
0 32225 5 1 1 32224
0 32226 7 1 2 32221 32225
0 32227 5 1 1 32226
0 32228 7 1 2 97930 32227
0 32229 5 1 1 32228
0 32230 7 1 2 88397 73967
0 32231 5 1 1 32230
0 32232 7 2 2 78701 32231
0 32233 7 1 2 85515 102531
0 32234 7 1 2 103180 32233
0 32235 5 1 1 32234
0 32236 7 1 2 32229 32235
0 32237 5 1 1 32236
0 32238 7 1 2 100287 32237
0 32239 5 1 1 32238
0 32240 7 1 2 95208 97264
0 32241 5 1 1 32240
0 32242 7 1 2 92188 94376
0 32243 5 1 1 32242
0 32244 7 1 2 32241 32243
0 32245 5 1 1 32244
0 32246 7 1 2 65446 32245
0 32247 5 1 1 32246
0 32248 7 1 2 87800 94393
0 32249 5 1 1 32248
0 32250 7 1 2 97785 32249
0 32251 5 1 1 32250
0 32252 7 1 2 66322 32251
0 32253 5 1 1 32252
0 32254 7 1 2 32247 32253
0 32255 5 1 1 32254
0 32256 7 1 2 64764 32255
0 32257 5 1 1 32256
0 32258 7 2 2 66323 97265
0 32259 5 1 1 103182
0 32260 7 1 2 75105 103183
0 32261 5 1 1 32260
0 32262 7 1 2 29312 32261
0 32263 5 1 1 32262
0 32264 7 1 2 66755 32263
0 32265 5 1 1 32264
0 32266 7 2 2 80526 85774
0 32267 5 1 1 103184
0 32268 7 3 2 72691 79577
0 32269 7 1 2 103185 103186
0 32270 5 1 1 32269
0 32271 7 1 2 32265 32270
0 32272 5 1 1 32271
0 32273 7 1 2 69886 32272
0 32274 5 1 1 32273
0 32275 7 1 2 32257 32274
0 32276 5 1 1 32275
0 32277 7 1 2 74428 100219
0 32278 7 1 2 32276 32277
0 32279 5 1 1 32278
0 32280 7 1 2 32239 32279
0 32281 5 1 1 32280
0 32282 7 1 2 70205 32281
0 32283 5 1 1 32282
0 32284 7 1 2 85742 75784
0 32285 5 2 1 32284
0 32286 7 1 2 76593 80360
0 32287 5 1 1 32286
0 32288 7 1 2 103189 32287
0 32289 5 1 1 32288
0 32290 7 1 2 66565 32289
0 32291 5 1 1 32290
0 32292 7 2 2 80712 97404
0 32293 5 1 1 103191
0 32294 7 1 2 83814 103192
0 32295 5 1 1 32294
0 32296 7 1 2 32291 32295
0 32297 5 1 1 32296
0 32298 7 1 2 73164 32297
0 32299 5 1 1 32298
0 32300 7 1 2 95123 89171
0 32301 5 1 1 32300
0 32302 7 1 2 78776 75067
0 32303 5 1 1 32302
0 32304 7 1 2 64765 32303
0 32305 5 1 1 32304
0 32306 7 1 2 101729 32305
0 32307 5 1 1 32306
0 32308 7 1 2 88398 32307
0 32309 5 1 1 32308
0 32310 7 1 2 32301 32309
0 32311 7 1 2 32299 32310
0 32312 5 1 1 32311
0 32313 7 1 2 100396 32312
0 32314 5 1 1 32313
0 32315 7 3 2 71672 88797
0 32316 7 2 2 63906 76486
0 32317 7 2 2 91350 103196
0 32318 7 1 2 103193 103198
0 32319 5 1 1 32318
0 32320 7 1 2 86950 95959
0 32321 7 1 2 100397 32320
0 32322 5 1 1 32321
0 32323 7 1 2 32319 32322
0 32324 5 1 1 32323
0 32325 7 1 2 85766 32324
0 32326 5 1 1 32325
0 32327 7 1 2 32314 32326
0 32328 5 1 1 32327
0 32329 7 1 2 65138 32328
0 32330 5 1 1 32329
0 32331 7 1 2 93412 89277
0 32332 5 1 1 32331
0 32333 7 1 2 93286 74334
0 32334 5 1 1 32333
0 32335 7 1 2 32332 32334
0 32336 5 1 1 32335
0 32337 7 1 2 86054 32336
0 32338 5 1 1 32337
0 32339 7 7 2 70827 73165
0 32340 7 1 2 97373 95088
0 32341 5 2 1 32340
0 32342 7 1 2 73750 83685
0 32343 7 1 2 103207 32342
0 32344 5 1 1 32343
0 32345 7 1 2 22703 32344
0 32346 5 1 1 32345
0 32347 7 1 2 66566 32346
0 32348 5 1 1 32347
0 32349 7 1 2 83068 100701
0 32350 5 1 1 32349
0 32351 7 1 2 75068 103190
0 32352 5 1 1 32351
0 32353 7 1 2 64766 32352
0 32354 5 1 1 32353
0 32355 7 1 2 32350 32354
0 32356 7 1 2 32348 32355
0 32357 5 1 1 32356
0 32358 7 1 2 103200 32357
0 32359 5 1 1 32358
0 32360 7 1 2 32338 32359
0 32361 5 1 1 32360
0 32362 7 1 2 100288 32361
0 32363 5 1 1 32362
0 32364 7 1 2 72692 32363
0 32365 7 1 2 32330 32364
0 32366 5 1 1 32365
0 32367 7 1 2 79174 92421
0 32368 5 1 1 32367
0 32369 7 2 2 77873 94822
0 32370 5 1 1 103209
0 32371 7 1 2 32368 32370
0 32372 5 1 1 32371
0 32373 7 1 2 97931 32372
0 32374 5 1 1 32373
0 32375 7 1 2 73920 83263
0 32376 5 1 1 32375
0 32377 7 1 2 83312 32376
0 32378 5 1 1 32377
0 32379 7 1 2 86055 32378
0 32380 5 1 1 32379
0 32381 7 1 2 68429 83308
0 32382 5 1 1 32381
0 32383 7 1 2 32380 32382
0 32384 5 1 1 32383
0 32385 7 1 2 65819 32384
0 32386 5 1 1 32385
0 32387 7 1 2 32374 32386
0 32388 5 1 1 32387
0 32389 7 1 2 100289 32388
0 32390 5 1 1 32389
0 32391 7 1 2 65602 100808
0 32392 7 1 2 101869 32391
0 32393 7 1 2 76784 88814
0 32394 7 1 2 32392 32393
0 32395 5 1 1 32394
0 32396 7 1 2 67669 32395
0 32397 7 1 2 32390 32396
0 32398 5 1 1 32397
0 32399 7 1 2 69190 32398
0 32400 7 1 2 32366 32399
0 32401 5 1 1 32400
0 32402 7 1 2 32283 32401
0 32403 7 1 2 32219 32402
0 32404 5 1 1 32403
0 32405 7 1 2 103148 32404
0 32406 5 1 1 32405
0 32407 7 1 2 99595 91326
0 32408 5 1 1 32407
0 32409 7 1 2 73166 101719
0 32410 5 2 1 32409
0 32411 7 1 2 68080 101856
0 32412 5 1 1 32411
0 32413 7 1 2 103211 32412
0 32414 5 1 1 32413
0 32415 7 1 2 71420 32414
0 32416 5 1 1 32415
0 32417 7 1 2 78743 94283
0 32418 5 2 1 32417
0 32419 7 1 2 76031 27982
0 32420 5 1 1 32419
0 32421 7 1 2 103213 32420
0 32422 7 1 2 32416 32421
0 32423 5 1 1 32422
0 32424 7 1 2 67670 32423
0 32425 5 1 1 32424
0 32426 7 1 2 32408 32425
0 32427 5 1 1 32426
0 32428 7 1 2 85516 32427
0 32429 5 1 1 32428
0 32430 7 1 2 66324 31286
0 32431 5 1 1 32430
0 32432 7 1 2 88860 102883
0 32433 5 2 1 32432
0 32434 7 1 2 64767 103215
0 32435 5 1 1 32434
0 32436 7 1 2 32431 32435
0 32437 5 1 1 32436
0 32438 7 1 2 73167 32437
0 32439 5 1 1 32438
0 32440 7 1 2 99431 93686
0 32441 5 1 1 32440
0 32442 7 1 2 73751 86450
0 32443 5 1 1 32442
0 32444 7 1 2 32441 32443
0 32445 5 1 1 32444
0 32446 7 1 2 86892 32445
0 32447 5 1 1 32446
0 32448 7 1 2 66325 32447
0 32449 5 1 1 32448
0 32450 7 1 2 32449 95173
0 32451 5 1 1 32450
0 32452 7 1 2 64768 32451
0 32453 5 1 1 32452
0 32454 7 3 2 70467 75922
0 32455 5 1 1 103217
0 32456 7 1 2 76091 83069
0 32457 5 1 1 32456
0 32458 7 1 2 32455 32457
0 32459 7 1 2 32453 32458
0 32460 5 1 1 32459
0 32461 7 1 2 79908 32460
0 32462 5 1 1 32461
0 32463 7 1 2 32439 32462
0 32464 5 1 1 32463
0 32465 7 1 2 101053 32464
0 32466 5 1 1 32465
0 32467 7 1 2 32429 32466
0 32468 5 1 1 32467
0 32469 7 1 2 92125 103134
0 32470 7 1 2 32468 32469
0 32471 5 1 1 32470
0 32472 7 1 2 32406 32471
0 32473 5 1 1 32472
0 32474 7 1 2 67193 32473
0 32475 5 1 1 32474
0 32476 7 1 2 89211 27579
0 32477 5 1 1 32476
0 32478 7 1 2 73517 32477
0 32479 5 2 1 32478
0 32480 7 1 2 86543 79198
0 32481 5 2 1 32480
0 32482 7 1 2 103220 103222
0 32483 5 1 1 32482
0 32484 7 1 2 75923 32483
0 32485 5 1 1 32484
0 32486 7 1 2 75014 86470
0 32487 5 2 1 32486
0 32488 7 1 2 82634 92646
0 32489 5 1 1 32488
0 32490 7 1 2 81199 32489
0 32491 7 1 2 103224 32490
0 32492 5 1 1 32491
0 32493 7 1 2 64769 32492
0 32494 5 1 1 32493
0 32495 7 1 2 82635 76092
0 32496 5 2 1 32495
0 32497 7 1 2 66326 87214
0 32498 5 1 1 32497
0 32499 7 1 2 103226 32498
0 32500 7 1 2 32494 32499
0 32501 5 1 1 32500
0 32502 7 1 2 79845 32501
0 32503 5 1 1 32502
0 32504 7 1 2 32485 32503
0 32505 5 1 1 32504
0 32506 7 1 2 102928 32505
0 32507 5 1 1 32506
0 32508 7 1 2 100608 95883
0 32509 5 1 1 32508
0 32510 7 1 2 65139 32509
0 32511 5 1 1 32510
0 32512 7 1 2 64770 100597
0 32513 5 1 1 32512
0 32514 7 1 2 32511 32513
0 32515 5 1 1 32514
0 32516 7 1 2 71421 32515
0 32517 5 1 1 32516
0 32518 7 1 2 86321 93891
0 32519 5 1 1 32518
0 32520 7 1 2 32517 32519
0 32521 5 1 1 32520
0 32522 7 1 2 73518 32521
0 32523 5 1 1 32522
0 32524 7 1 2 66327 103110
0 32525 5 1 1 32524
0 32526 7 1 2 76632 90143
0 32527 5 1 1 32526
0 32528 7 1 2 32525 32527
0 32529 7 1 2 32523 32528
0 32530 5 1 1 32529
0 32531 7 1 2 73168 32530
0 32532 5 1 1 32531
0 32533 7 1 2 75106 31565
0 32534 5 1 1 32533
0 32535 7 1 2 32534 14612
0 32536 5 1 1 32535
0 32537 7 1 2 66756 32536
0 32538 5 1 1 32537
0 32539 7 1 2 66328 103112
0 32540 5 1 1 32539
0 32541 7 1 2 32538 32540
0 32542 5 1 1 32541
0 32543 7 1 2 68081 32542
0 32544 5 1 1 32543
0 32545 7 1 2 101239 93748
0 32546 5 1 1 32545
0 32547 7 1 2 32544 32546
0 32548 5 1 1 32547
0 32549 7 1 2 64771 32548
0 32550 5 1 1 32549
0 32551 7 1 2 94128 86726
0 32552 5 1 1 32551
0 32553 7 1 2 103118 32552
0 32554 7 1 2 32550 32553
0 32555 7 1 2 32532 32554
0 32556 5 1 1 32555
0 32557 7 1 2 102938 32556
0 32558 5 1 1 32557
0 32559 7 1 2 32507 32558
0 32560 5 1 1 32559
0 32561 7 1 2 72693 32560
0 32562 5 1 1 32561
0 32563 7 1 2 31365 102930
0 32564 5 1 1 32563
0 32565 7 2 2 76227 75509
0 32566 7 3 2 87258 103228
0 32567 5 2 1 103230
0 32568 7 1 2 87801 103231
0 32569 7 1 2 32564 32568
0 32570 5 1 1 32569
0 32571 7 1 2 32562 32570
0 32572 5 1 1 32571
0 32573 7 3 2 64130 72249
0 32574 7 1 2 102968 103235
0 32575 7 1 2 32572 32574
0 32576 5 1 1 32575
0 32577 7 1 2 32475 32576
0 32578 5 1 1 32577
0 32579 7 1 2 67338 32578
0 32580 5 1 1 32579
0 32581 7 1 2 90367 102418
0 32582 7 1 2 94916 32581
0 32583 5 1 1 32582
0 32584 7 1 2 98840 99630
0 32585 7 1 2 94005 98845
0 32586 7 1 2 32584 32585
0 32587 5 1 1 32586
0 32588 7 1 2 32583 32587
0 32589 5 1 1 32588
0 32590 7 1 2 69191 32589
0 32591 5 1 1 32590
0 32592 7 3 2 66567 72250
0 32593 7 1 2 93044 102196
0 32594 7 1 2 103238 32593
0 32595 7 1 2 102816 32594
0 32596 5 1 1 32595
0 32597 7 1 2 32591 32596
0 32598 5 1 1 32597
0 32599 7 1 2 68993 32598
0 32600 5 1 1 32599
0 32601 7 1 2 103239 97093
0 32602 7 1 2 94517 32601
0 32603 7 1 2 102227 32602
0 32604 5 1 1 32603
0 32605 7 1 2 32600 32604
0 32606 5 1 1 32605
0 32607 7 1 2 76594 32606
0 32608 5 1 1 32607
0 32609 7 2 2 72251 103072
0 32610 7 1 2 88342 102228
0 32611 7 1 2 103241 32610
0 32612 5 1 1 32611
0 32613 7 1 2 32608 32612
0 32614 5 1 1 32613
0 32615 7 1 2 72694 32614
0 32616 5 1 1 32615
0 32617 7 1 2 79681 102502
0 32618 5 1 1 32617
0 32619 7 3 2 67194 68672
0 32620 7 1 2 100345 103243
0 32621 7 1 2 95576 32620
0 32622 5 1 1 32621
0 32623 7 1 2 32618 32622
0 32624 5 1 1 32623
0 32625 7 1 2 84217 32624
0 32626 5 1 1 32625
0 32627 7 3 2 71422 72252
0 32628 7 1 2 100403 103246
0 32629 7 1 2 101584 32628
0 32630 5 1 1 32629
0 32631 7 1 2 99692 90368
0 32632 7 1 2 102409 32631
0 32633 7 1 2 83932 32632
0 32634 5 1 1 32633
0 32635 7 1 2 32630 32634
0 32636 5 1 1 32635
0 32637 7 1 2 68994 32636
0 32638 5 1 1 32637
0 32639 7 2 2 102390 103038
0 32640 7 2 2 68866 71423
0 32641 7 1 2 79090 103251
0 32642 7 1 2 103249 32641
0 32643 5 1 1 32642
0 32644 7 1 2 32638 32643
0 32645 5 1 1 32644
0 32646 7 1 2 78702 32645
0 32647 5 1 1 32646
0 32648 7 1 2 32626 32647
0 32649 5 1 1 32648
0 32650 7 1 2 97044 32649
0 32651 5 1 1 32650
0 32652 7 1 2 32616 32651
0 32653 5 1 1 32652
0 32654 7 1 2 73169 32653
0 32655 5 1 1 32654
0 32656 7 2 2 83096 88339
0 32657 5 8 1 103253
0 32658 7 2 2 93215 97084
0 32659 7 1 2 103255 103263
0 32660 5 1 1 32659
0 32661 7 1 2 68082 98480
0 32662 7 1 2 102902 32661
0 32663 5 1 1 32662
0 32664 7 1 2 75280 87883
0 32665 7 1 2 102817 32664
0 32666 5 1 1 32665
0 32667 7 1 2 32663 32666
0 32668 5 1 1 32667
0 32669 7 1 2 66329 32668
0 32670 5 1 1 32669
0 32671 7 1 2 32660 32670
0 32672 5 1 1 32671
0 32673 7 1 2 64131 32672
0 32674 5 1 1 32673
0 32675 7 9 2 66330 84356
0 32676 7 3 2 66568 81416
0 32677 7 3 2 65140 72405
0 32678 7 1 2 65820 103277
0 32679 7 1 2 103274 32678
0 32680 7 1 2 103265 32679
0 32681 5 1 1 32680
0 32682 7 1 2 32674 32681
0 32683 5 1 1 32682
0 32684 7 1 2 103242 32683
0 32685 5 1 1 32684
0 32686 7 1 2 97368 101344
0 32687 5 2 1 32686
0 32688 7 3 2 70688 67195
0 32689 5 1 1 103282
0 32690 7 1 2 82443 83904
0 32691 7 1 2 103283 32690
0 32692 7 1 2 98572 32691
0 32693 7 1 2 103280 32692
0 32694 5 1 1 32693
0 32695 7 1 2 32685 32694
0 32696 7 1 2 32655 32695
0 32697 5 1 1 32696
0 32698 7 1 2 76808 32697
0 32699 5 1 1 32698
0 32700 7 3 2 99776 102399
0 32701 7 1 2 92718 103285
0 32702 5 1 1 32701
0 32703 7 2 2 72695 99296
0 32704 7 1 2 67196 100959
0 32705 7 1 2 79091 32704
0 32706 7 1 2 103288 32705
0 32707 5 1 1 32706
0 32708 7 1 2 32702 32707
0 32709 5 1 1 32708
0 32710 7 1 2 84554 32709
0 32711 5 1 1 32710
0 32712 7 1 2 97266 102421
0 32713 5 1 1 32712
0 32714 7 1 2 81449 103286
0 32715 5 1 1 32714
0 32716 7 1 2 32713 32715
0 32717 5 1 1 32716
0 32718 7 1 2 97405 32717
0 32719 5 1 1 32718
0 32720 7 1 2 32711 32719
0 32721 5 1 1 32720
0 32722 7 1 2 32721 84781
0 32723 5 1 1 32722
0 32724 7 1 2 72164 32723
0 32725 7 1 2 32699 32724
0 32726 5 1 1 32725
0 32727 7 1 2 100981 102812
0 32728 7 1 2 92590 32727
0 32729 5 1 1 32728
0 32730 7 2 2 67339 76595
0 32731 7 1 2 96412 103013
0 32732 7 1 2 103290 32731
0 32733 5 1 1 32732
0 32734 7 1 2 32729 32733
0 32735 5 1 1 32734
0 32736 7 1 2 73170 32735
0 32737 5 1 1 32736
0 32738 7 1 2 103129 84227
0 32739 7 1 2 97234 32738
0 32740 7 1 2 99983 32739
0 32741 5 1 1 32740
0 32742 7 1 2 32737 32741
0 32743 5 1 1 32742
0 32744 7 1 2 73519 32743
0 32745 5 1 1 32744
0 32746 7 9 2 67197 67340
0 32747 7 1 2 78348 103292
0 32748 7 1 2 103093 32747
0 32749 7 1 2 79964 32748
0 32750 5 1 1 32749
0 32751 7 1 2 32745 32750
0 32752 5 1 1 32751
0 32753 7 1 2 63907 32752
0 32754 5 1 1 32753
0 32755 7 1 2 77618 5077
0 32756 5 2 1 32755
0 32757 7 2 2 93732 96314
0 32758 7 1 2 102414 103303
0 32759 7 1 2 103301 32758
0 32760 5 1 1 32759
0 32761 7 1 2 32754 32760
0 32762 5 1 1 32761
0 32763 7 1 2 63804 32762
0 32764 5 1 1 32763
0 32765 7 1 2 102917 102411
0 32766 7 1 2 102282 32765
0 32767 7 1 2 103302 32766
0 32768 5 1 1 32767
0 32769 7 1 2 32764 32768
0 32770 5 1 1 32769
0 32771 7 1 2 72696 32770
0 32772 5 1 1 32771
0 32773 7 1 2 73968 95507
0 32774 7 1 2 97719 32773
0 32775 7 2 2 102283 32774
0 32776 7 1 2 94780 103305
0 32777 5 1 1 32776
0 32778 7 9 2 66331 72253
0 32779 7 1 2 66878 93239
0 32780 7 1 2 103307 32779
0 32781 7 1 2 83016 102078
0 32782 7 1 2 32780 32781
0 32783 5 1 1 32782
0 32784 7 1 2 32777 32783
0 32785 5 1 1 32784
0 32786 7 1 2 63805 32785
0 32787 5 1 1 32786
0 32788 7 3 2 65603 93707
0 32789 7 1 2 103306 103316
0 32790 5 1 1 32789
0 32791 7 1 2 32787 32790
0 32792 5 1 1 32791
0 32793 7 1 2 97045 32792
0 32794 5 1 1 32793
0 32795 7 1 2 67120 32794
0 32796 7 1 2 32772 32795
0 32797 5 1 1 32796
0 32798 7 1 2 84838 32797
0 32799 7 1 2 32726 32798
0 32800 5 1 1 32799
0 32801 7 2 2 64132 79030
0 32802 7 1 2 95648 103085
0 32803 7 1 2 103319 32802
0 32804 5 1 1 32803
0 32805 7 1 2 30786 32804
0 32806 5 1 1 32805
0 32807 7 1 2 68867 32806
0 32808 5 1 1 32807
0 32809 7 2 2 69192 67121
0 32810 7 1 2 102729 103321
0 32811 7 1 2 101906 32810
0 32812 5 1 1 32811
0 32813 7 1 2 32808 32812
0 32814 5 2 1 32813
0 32815 7 1 2 84489 103323
0 32816 5 1 1 32815
0 32817 7 1 2 78314 103149
0 32818 7 1 2 95484 32817
0 32819 7 1 2 65447 99672
0 32820 7 1 2 102962 32819
0 32821 7 1 2 32818 32820
0 32822 5 1 1 32821
0 32823 7 1 2 32816 32822
0 32824 5 1 1 32823
0 32825 7 1 2 67671 32824
0 32826 5 1 1 32825
0 32827 7 2 2 86493 76887
0 32828 7 1 2 101985 92074
0 32829 7 1 2 103325 32828
0 32830 7 1 2 98363 32829
0 32831 5 1 1 32830
0 32832 7 1 2 32826 32831
0 32833 5 1 1 32832
0 32834 7 1 2 65650 32833
0 32835 5 1 1 32834
0 32836 7 3 2 67672 81889
0 32837 7 2 2 92126 103327
0 32838 7 1 2 72254 93766
0 32839 7 1 2 100624 32838
0 32840 7 1 2 103330 32839
0 32841 5 1 1 32840
0 32842 7 1 2 32835 32841
0 32843 5 1 1 32842
0 32844 7 1 2 72406 32843
0 32845 5 1 1 32844
0 32846 7 1 2 65651 76888
0 32847 7 1 2 103009 32846
0 32848 7 2 2 68868 85417
0 32849 7 1 2 102340 103332
0 32850 7 1 2 32847 32849
0 32851 5 1 1 32850
0 32852 7 1 2 68995 32851
0 32853 7 1 2 32845 32852
0 32854 5 1 1 32853
0 32855 7 3 2 67673 94589
0 32856 7 1 2 103324 103334
0 32857 5 1 1 32856
0 32858 7 1 2 69887 22368
0 32859 5 1 1 32858
0 32860 7 1 2 64772 20623
0 32861 5 1 1 32860
0 32862 7 9 2 72255 72697
0 32863 7 1 2 103337 96290
0 32864 7 1 2 32861 32863
0 32865 7 1 2 32859 32864
0 32866 5 1 1 32865
0 32867 7 1 2 32857 32866
0 32868 5 1 1 32867
0 32869 7 1 2 71424 32868
0 32870 5 1 1 32869
0 32871 7 1 2 79138 98364
0 32872 5 1 1 32871
0 32873 7 1 2 84741 82549
0 32874 7 1 2 84782 32873
0 32875 5 1 1 32874
0 32876 7 1 2 32872 32875
0 32877 5 1 1 32876
0 32878 7 1 2 96003 103308
0 32879 7 1 2 96431 32878
0 32880 7 1 2 32877 32879
0 32881 5 1 1 32880
0 32882 7 1 2 32870 32881
0 32883 5 1 1 32882
0 32884 7 1 2 72407 32883
0 32885 5 1 1 32884
0 32886 7 4 2 64773 87926
0 32887 7 1 2 93045 102026
0 32888 7 1 2 76889 103338
0 32889 7 1 2 32887 32888
0 32890 7 1 2 103346 32889
0 32891 5 1 1 32890
0 32892 7 1 2 69888 101244
0 32893 5 1 1 32892
0 32894 7 1 2 76327 99945
0 32895 7 1 2 100609 32894
0 32896 7 1 2 32893 32895
0 32897 5 1 1 32896
0 32898 7 1 2 70828 83866
0 32899 7 1 2 84627 32898
0 32900 5 1 1 32899
0 32901 7 1 2 32897 32900
0 32902 5 1 1 32901
0 32903 7 1 2 72698 32902
0 32904 5 1 1 32903
0 32905 7 1 2 67674 74342
0 32906 7 1 2 93820 32905
0 32907 5 1 1 32906
0 32908 7 1 2 32904 32907
0 32909 5 1 1 32908
0 32910 7 3 2 88899 79640
0 32911 7 1 2 67198 103350
0 32912 7 1 2 32909 32911
0 32913 5 1 1 32912
0 32914 7 1 2 32891 32913
0 32915 5 1 1 32914
0 32916 7 1 2 102745 32915
0 32917 5 1 1 32916
0 32918 7 1 2 63908 32917
0 32919 7 1 2 32885 32918
0 32920 5 1 1 32919
0 32921 7 1 2 84555 32920
0 32922 7 1 2 32854 32921
0 32923 5 1 1 32922
0 32924 7 1 2 32800 32923
0 32925 7 1 2 32580 32924
0 32926 7 1 2 32130 32925
0 32927 5 1 1 32926
0 32928 7 1 2 67001 32927
0 32929 5 1 1 32928
0 32930 7 7 2 72408 102624
0 32931 7 1 2 102516 103353
0 32932 5 1 1 32931
0 32933 7 1 2 91468 102769
0 32934 5 1 1 32933
0 32935 7 1 2 32932 32934
0 32936 5 1 1 32935
0 32937 7 1 2 64774 100849
0 32938 5 1 1 32937
0 32939 7 1 2 65448 93866
0 32940 5 1 1 32939
0 32941 7 1 2 96900 32940
0 32942 5 1 1 32941
0 32943 7 1 2 79207 32942
0 32944 5 1 1 32943
0 32945 7 1 2 32938 32944
0 32946 5 1 1 32945
0 32947 7 4 2 85517 100290
0 32948 7 1 2 32946 103360
0 32949 5 1 1 32948
0 32950 7 2 2 90951 86504
0 32951 7 1 2 93319 98064
0 32952 7 1 2 103364 32951
0 32953 5 1 1 32952
0 32954 7 1 2 100225 32953
0 32955 5 1 1 32954
0 32956 7 1 2 85693 85518
0 32957 7 1 2 32955 32956
0 32958 5 1 1 32957
0 32959 7 1 2 32949 32958
0 32960 5 1 1 32959
0 32961 7 1 2 85952 32960
0 32962 5 1 1 32961
0 32963 7 1 2 82178 94543
0 32964 5 1 1 32963
0 32965 7 1 2 103361 32964
0 32966 5 1 1 32965
0 32967 7 1 2 100043 103362
0 32968 5 1 1 32967
0 32969 7 3 2 70206 65604
0 32970 7 2 2 79092 103366
0 32971 7 1 2 65652 92422
0 32972 7 1 2 92372 32971
0 32973 7 1 2 103369 32972
0 32974 5 1 1 32973
0 32975 7 1 2 32968 32974
0 32976 5 1 1 32975
0 32977 7 1 2 86056 32976
0 32978 5 1 1 32977
0 32979 7 1 2 32966 32978
0 32980 5 1 1 32979
0 32981 7 1 2 85334 32980
0 32982 5 1 1 32981
0 32983 7 1 2 32962 32982
0 32984 5 1 1 32983
0 32985 7 1 2 32936 32984
0 32986 5 1 1 32985
0 32987 7 1 2 32929 32986
0 32988 7 1 2 31251 32987
0 32989 5 1 1 32988
0 32990 7 1 2 81032 32989
0 32991 5 1 1 32990
0 32992 7 1 2 99693 99306
0 32993 7 1 2 92055 95501
0 32994 7 1 2 32992 32993
0 32995 5 1 1 32994
0 32996 7 1 2 76655 89445
0 32997 7 1 2 94357 32996
0 32998 5 2 1 32997
0 32999 7 2 2 91071 77021
0 33000 7 1 2 102003 103373
0 33001 7 1 2 103371 33000
0 33002 5 1 1 33001
0 33003 7 1 2 32995 33002
0 33004 5 1 1 33003
0 33005 7 1 2 79139 33004
0 33006 5 1 1 33005
0 33007 7 1 2 84255 80527
0 33008 5 1 1 33007
0 33009 7 1 2 75403 95489
0 33010 5 1 1 33009
0 33011 7 1 2 33008 33010
0 33012 5 3 1 33011
0 33013 7 2 2 76958 76845
0 33014 7 2 2 95281 78171
0 33015 7 1 2 103380 84472
0 33016 7 1 2 103378 33015
0 33017 7 1 2 103375 33016
0 33018 5 1 1 33017
0 33019 7 1 2 33006 33018
0 33020 5 1 1 33019
0 33021 7 1 2 71425 33020
0 33022 5 1 1 33021
0 33023 7 1 2 89066 95245
0 33024 5 1 1 33023
0 33025 7 1 2 66569 95106
0 33026 5 1 1 33025
0 33027 7 1 2 77939 89743
0 33028 7 1 2 83934 33027
0 33029 5 1 1 33028
0 33030 7 1 2 89664 33029
0 33031 5 1 1 33030
0 33032 7 1 2 87454 33031
0 33033 5 1 1 33032
0 33034 7 1 2 33026 33033
0 33035 7 1 2 33024 33034
0 33036 5 1 1 33035
0 33037 7 1 2 73171 33036
0 33038 5 1 1 33037
0 33039 7 1 2 33038 103233
0 33040 5 1 1 33039
0 33041 7 3 2 77248 79660
0 33042 7 1 2 33040 103382
0 33043 5 1 1 33042
0 33044 7 1 2 85607 15814
0 33045 5 1 1 33044
0 33046 7 1 2 70468 33045
0 33047 5 1 1 33046
0 33048 7 1 2 33047 85601
0 33049 5 1 1 33048
0 33050 7 1 2 64775 33049
0 33051 5 1 1 33050
0 33052 7 1 2 79217 85582
0 33053 5 1 1 33052
0 33054 7 1 2 74669 33053
0 33055 5 1 1 33054
0 33056 7 2 2 79031 82600
0 33057 5 3 1 103385
0 33058 7 1 2 33055 103387
0 33059 5 1 1 33058
0 33060 7 1 2 73172 33059
0 33061 5 1 1 33060
0 33062 7 1 2 33051 33061
0 33063 5 1 1 33062
0 33064 7 1 2 79140 33063
0 33065 5 1 1 33064
0 33066 7 1 2 78868 85815
0 33067 5 1 1 33066
0 33068 7 1 2 83484 86971
0 33069 5 3 1 33068
0 33070 7 1 2 103390 79488
0 33071 5 1 1 33070
0 33072 7 1 2 898 33071
0 33073 5 2 1 33072
0 33074 7 1 2 79846 103393
0 33075 5 1 1 33074
0 33076 7 1 2 33067 33075
0 33077 7 1 2 33065 33076
0 33078 5 1 1 33077
0 33079 7 1 2 66332 33078
0 33080 5 1 1 33079
0 33081 7 1 2 92000 103394
0 33082 5 1 1 33081
0 33083 7 1 2 77673 83815
0 33084 5 1 1 33083
0 33085 7 1 2 79847 85811
0 33086 5 1 1 33085
0 33087 7 1 2 33084 33086
0 33088 5 1 1 33087
0 33089 7 1 2 78869 33088
0 33090 5 1 1 33089
0 33091 7 1 2 85824 86403
0 33092 7 1 2 103326 33091
0 33093 5 1 1 33092
0 33094 7 1 2 85694 82744
0 33095 7 1 2 79661 33094
0 33096 5 1 1 33095
0 33097 7 1 2 33093 33096
0 33098 5 1 1 33097
0 33099 7 1 2 74670 33098
0 33100 5 1 1 33099
0 33101 7 1 2 33090 33100
0 33102 7 1 2 33082 33101
0 33103 7 1 2 33080 33102
0 33104 5 1 1 33103
0 33105 7 1 2 77354 33104
0 33106 5 1 1 33105
0 33107 7 1 2 33043 33106
0 33108 5 1 1 33107
0 33109 7 1 2 74398 74245
0 33110 7 1 2 33108 33109
0 33111 5 1 1 33110
0 33112 7 1 2 33022 33111
0 33113 5 1 1 33112
0 33114 7 1 2 67341 33113
0 33115 5 1 1 33114
0 33116 7 2 2 66333 74490
0 33117 5 1 1 103395
0 33118 7 1 2 33117 103114
0 33119 5 1 1 33118
0 33120 7 1 2 64776 33119
0 33121 5 1 1 33120
0 33122 7 1 2 33121 87689
0 33123 5 1 1 33122
0 33124 7 1 2 80414 33123
0 33125 5 1 1 33124
0 33126 7 1 2 66334 101361
0 33127 5 1 1 33126
0 33128 7 1 2 95011 33127
0 33129 5 1 1 33128
0 33130 7 1 2 64777 33129
0 33131 5 1 1 33130
0 33132 7 1 2 102141 33131
0 33133 5 2 1 33132
0 33134 7 1 2 80361 103397
0 33135 5 2 1 33134
0 33136 7 1 2 33125 103399
0 33137 5 1 1 33136
0 33138 7 1 2 70829 33137
0 33139 5 1 1 33138
0 33140 7 1 2 93216 83326
0 33141 7 1 2 95691 33140
0 33142 5 1 1 33141
0 33143 7 2 2 69889 80537
0 33144 5 1 1 103401
0 33145 7 1 2 92388 103402
0 33146 5 1 1 33145
0 33147 7 1 2 90096 74343
0 33148 5 1 1 33147
0 33149 7 1 2 33146 33148
0 33150 5 1 1 33149
0 33151 7 1 2 70207 33150
0 33152 5 1 1 33151
0 33153 7 1 2 33142 33152
0 33154 7 1 2 33139 33153
0 33155 5 1 1 33154
0 33156 7 1 2 77355 33155
0 33157 5 1 1 33156
0 33158 7 1 2 80415 103116
0 33159 5 1 1 33158
0 33160 7 1 2 103400 33159
0 33161 5 1 1 33160
0 33162 7 1 2 98520 33161
0 33163 5 1 1 33162
0 33164 7 1 2 33157 33163
0 33165 5 1 1 33164
0 33166 7 1 2 70469 33165
0 33167 5 1 1 33166
0 33168 7 2 2 83411 87233
0 33169 5 1 1 103403
0 33170 7 1 2 82982 94929
0 33171 5 1 1 33170
0 33172 7 1 2 65449 101692
0 33173 7 1 2 33171 33172
0 33174 5 1 1 33173
0 33175 7 1 2 33169 33174
0 33176 5 1 1 33175
0 33177 7 1 2 75924 33176
0 33178 5 1 1 33177
0 33179 7 2 2 96004 75281
0 33180 7 1 2 86727 103405
0 33181 5 1 1 33180
0 33182 7 1 2 33178 33181
0 33183 5 1 1 33182
0 33184 7 1 2 97878 33183
0 33185 5 1 1 33184
0 33186 7 1 2 33167 33185
0 33187 5 1 1 33186
0 33188 7 1 2 64133 33187
0 33189 5 1 1 33188
0 33190 7 1 2 69890 95051
0 33191 5 1 1 33190
0 33192 7 1 2 102037 33191
0 33193 5 1 1 33192
0 33194 7 1 2 74671 33193
0 33195 5 1 1 33194
0 33196 7 1 2 80416 103256
0 33197 5 1 1 33196
0 33198 7 1 2 82115 86160
0 33199 5 1 1 33198
0 33200 7 1 2 33197 33199
0 33201 5 1 1 33200
0 33202 7 1 2 70470 33201
0 33203 5 1 1 33202
0 33204 7 1 2 65450 101663
0 33205 5 1 1 33204
0 33206 7 1 2 33203 33205
0 33207 7 1 2 33195 33206
0 33208 5 1 1 33207
0 33209 7 1 2 73173 33208
0 33210 5 1 1 33209
0 33211 7 1 2 84118 102374
0 33212 5 1 1 33211
0 33213 7 1 2 75282 83971
0 33214 7 1 2 33212 33213
0 33215 5 1 1 33214
0 33216 7 1 2 33210 33215
0 33217 5 1 1 33216
0 33218 7 1 2 66335 33217
0 33219 5 1 1 33218
0 33220 7 5 2 66570 78315
0 33221 7 1 2 79672 88810
0 33222 5 1 1 33221
0 33223 7 1 2 66757 33222
0 33224 5 1 1 33223
0 33225 7 1 2 33224 32267
0 33226 5 1 1 33225
0 33227 7 1 2 103407 33226
0 33228 5 1 1 33227
0 33229 7 1 2 33219 33228
0 33230 5 1 1 33229
0 33231 7 1 2 98731 33230
0 33232 5 1 1 33231
0 33233 7 1 2 33189 33232
0 33234 5 1 1 33233
0 33235 7 1 2 79141 33234
0 33236 5 1 1 33235
0 33237 7 1 2 78703 95034
0 33238 5 1 1 33237
0 33239 7 1 2 77611 87285
0 33240 5 1 1 33239
0 33241 7 1 2 33238 33240
0 33242 5 1 1 33241
0 33243 7 1 2 93618 33242
0 33244 5 1 1 33243
0 33245 7 1 2 73752 101247
0 33246 5 1 1 33245
0 33247 7 2 2 80362 101234
0 33248 5 2 1 103412
0 33249 7 1 2 33246 103414
0 33250 5 2 1 33249
0 33251 7 1 2 64778 103416
0 33252 5 2 1 33251
0 33253 7 1 2 91522 86650
0 33254 5 1 1 33253
0 33255 7 1 2 103418 33254
0 33256 5 1 1 33255
0 33257 7 1 2 74964 33256
0 33258 5 1 1 33257
0 33259 7 1 2 99515 80081
0 33260 7 1 2 91954 33259
0 33261 5 1 1 33260
0 33262 7 1 2 33258 33261
0 33263 5 1 1 33262
0 33264 7 1 2 70471 33263
0 33265 5 1 1 33264
0 33266 7 1 2 77541 89035
0 33267 5 1 1 33266
0 33268 7 2 2 5641 33267
0 33269 7 1 2 65141 103420
0 33270 5 1 1 33269
0 33271 7 1 2 80164 87473
0 33272 5 1 1 33271
0 33273 7 1 2 80179 33272
0 33274 7 1 2 33270 33273
0 33275 5 2 1 33274
0 33276 7 1 2 69193 103422
0 33277 5 1 1 33276
0 33278 7 1 2 84761 92952
0 33279 7 1 2 100018 33278
0 33280 5 1 1 33279
0 33281 7 1 2 33277 33280
0 33282 7 1 2 33265 33281
0 33283 5 1 1 33282
0 33284 7 1 2 66026 33283
0 33285 5 1 1 33284
0 33286 7 1 2 33244 33285
0 33287 5 1 1 33286
0 33288 7 1 2 64424 33287
0 33289 5 1 1 33288
0 33290 7 1 2 94746 94323
0 33291 5 1 1 33290
0 33292 7 1 2 84909 100019
0 33293 5 1 1 33292
0 33294 7 1 2 33291 33293
0 33295 5 1 1 33294
0 33296 7 1 2 71426 33295
0 33297 5 1 1 33296
0 33298 7 1 2 101378 102922
0 33299 5 1 1 33298
0 33300 7 1 2 33297 33299
0 33301 5 1 1 33300
0 33302 7 1 2 65142 33301
0 33303 5 1 1 33302
0 33304 7 2 2 75089 79238
0 33305 5 4 1 103424
0 33306 7 1 2 81742 103426
0 33307 5 3 1 33306
0 33308 7 1 2 82749 103430
0 33309 5 1 1 33308
0 33310 7 1 2 101379 33309
0 33311 5 1 1 33310
0 33312 7 1 2 92779 86827
0 33313 5 1 1 33312
0 33314 7 1 2 33311 33313
0 33315 7 1 2 33303 33314
0 33316 5 1 1 33315
0 33317 7 1 2 68083 33316
0 33318 5 1 1 33317
0 33319 7 1 2 66336 85653
0 33320 5 2 1 33319
0 33321 7 1 2 103388 103433
0 33322 5 1 1 33321
0 33323 7 1 2 75404 33322
0 33324 5 1 1 33323
0 33325 7 2 2 76656 82648
0 33326 5 1 1 103435
0 33327 7 1 2 66337 103436
0 33328 5 1 1 33327
0 33329 7 1 2 33324 33328
0 33330 5 1 1 33329
0 33331 7 1 2 77454 33330
0 33332 5 1 1 33331
0 33333 7 1 2 71095 99579
0 33334 5 1 1 33333
0 33335 7 1 2 33332 33334
0 33336 5 1 1 33335
0 33337 7 1 2 73174 33336
0 33338 5 1 1 33337
0 33339 7 3 2 81890 83791
0 33340 5 1 1 103437
0 33341 7 2 2 75047 33340
0 33342 5 6 1 103440
0 33343 7 1 2 92780 103442
0 33344 5 1 1 33343
0 33345 7 1 2 101310 33344
0 33346 7 1 2 33338 33345
0 33347 7 1 2 33318 33346
0 33348 5 1 1 33347
0 33349 7 1 2 64134 33348
0 33350 5 1 1 33349
0 33351 7 1 2 33289 33350
0 33352 5 1 1 33351
0 33353 7 1 2 65821 33352
0 33354 5 1 1 33353
0 33355 7 5 2 85519 77249
0 33356 7 1 2 66338 87537
0 33357 5 1 1 33356
0 33358 7 1 2 82273 77699
0 33359 5 1 1 33358
0 33360 7 1 2 33357 33359
0 33361 5 1 1 33360
0 33362 7 1 2 64779 33361
0 33363 5 1 1 33362
0 33364 7 4 2 82601 77874
0 33365 7 1 2 95193 103453
0 33366 5 2 1 33365
0 33367 7 1 2 33363 103457
0 33368 5 1 1 33367
0 33369 7 1 2 103448 33368
0 33370 5 1 1 33369
0 33371 7 2 2 87320 100020
0 33372 5 2 1 103459
0 33373 7 1 2 92425 103460
0 33374 5 1 1 33373
0 33375 7 1 2 98707 103423
0 33376 5 1 1 33375
0 33377 7 1 2 33374 33376
0 33378 5 1 1 33377
0 33379 7 1 2 64135 33378
0 33380 5 1 1 33379
0 33381 7 1 2 33370 33380
0 33382 7 1 2 33354 33381
0 33383 5 1 1 33382
0 33384 7 1 2 78870 33383
0 33385 5 1 1 33384
0 33386 7 1 2 33236 33385
0 33387 5 1 1 33386
0 33388 7 1 2 72409 74246
0 33389 7 1 2 33387 33388
0 33390 5 1 1 33389
0 33391 7 1 2 33115 33390
0 33392 5 1 1 33391
0 33393 7 1 2 67675 33392
0 33394 5 1 1 33393
0 33395 7 1 2 74672 97406
0 33396 5 3 1 33395
0 33397 7 1 2 103463 89802
0 33398 5 1 1 33397
0 33399 7 1 2 71835 33398
0 33400 5 1 1 33399
0 33401 7 1 2 69891 88715
0 33402 5 1 1 33401
0 33403 7 1 2 97369 92169
0 33404 5 2 1 33403
0 33405 7 1 2 102478 103466
0 33406 5 1 1 33405
0 33407 7 1 2 33402 33406
0 33408 7 1 2 33400 33407
0 33409 5 1 1 33408
0 33410 7 1 2 70472 33409
0 33411 5 1 1 33410
0 33412 7 1 2 76596 80553
0 33413 7 1 2 78785 33412
0 33414 5 1 1 33413
0 33415 7 1 2 33411 33414
0 33416 5 1 1 33415
0 33417 7 1 2 97899 33416
0 33418 5 1 1 33417
0 33419 7 1 2 80363 102898
0 33420 5 2 1 33419
0 33421 7 1 2 86544 79232
0 33422 5 2 1 33421
0 33423 7 1 2 103468 103470
0 33424 5 1 1 33423
0 33425 7 1 2 95508 100111
0 33426 7 1 2 33424 33425
0 33427 5 1 1 33426
0 33428 7 1 2 33418 33427
0 33429 5 1 1 33428
0 33430 7 1 2 68084 33429
0 33431 5 1 1 33430
0 33432 7 1 2 102458 103194
0 33433 5 1 1 33432
0 33434 7 2 2 67342 93217
0 33435 7 1 2 100464 83403
0 33436 5 2 1 33435
0 33437 7 1 2 103472 103474
0 33438 5 1 1 33437
0 33439 7 1 2 33433 33438
0 33440 5 1 1 33439
0 33441 7 1 2 73175 80896
0 33442 7 1 2 33440 33441
0 33443 5 1 1 33442
0 33444 7 1 2 33431 33443
0 33445 5 1 1 33444
0 33446 7 1 2 77356 33445
0 33447 5 1 1 33446
0 33448 7 1 2 83355 92946
0 33449 5 1 1 33448
0 33450 7 1 2 88798 33449
0 33451 5 1 1 33450
0 33452 7 1 2 97361 83604
0 33453 7 1 2 86662 33452
0 33454 5 1 1 33453
0 33455 7 1 2 33451 33454
0 33456 5 1 1 33455
0 33457 7 2 2 72410 33456
0 33458 7 1 2 74063 96724
0 33459 7 1 2 103476 33458
0 33460 5 1 1 33459
0 33461 7 1 2 33447 33460
0 33462 5 1 1 33461
0 33463 7 1 2 64136 33462
0 33464 5 1 1 33463
0 33465 7 2 2 66339 74172
0 33466 7 1 2 86437 103478
0 33467 5 1 1 33466
0 33468 7 1 2 83605 102788
0 33469 5 1 1 33468
0 33470 7 1 2 33467 33469
0 33471 5 1 1 33470
0 33472 7 1 2 64780 33471
0 33473 5 1 1 33472
0 33474 7 1 2 71427 74791
0 33475 5 2 1 33474
0 33476 7 1 2 88776 103480
0 33477 5 1 1 33476
0 33478 7 1 2 69892 33477
0 33479 5 1 1 33478
0 33480 7 1 2 74965 100050
0 33481 5 1 1 33480
0 33482 7 1 2 33479 33481
0 33483 5 1 1 33482
0 33484 7 1 2 70473 33483
0 33485 5 1 1 33484
0 33486 7 1 2 83549 83327
0 33487 5 2 1 33486
0 33488 7 1 2 68430 87382
0 33489 5 1 1 33488
0 33490 7 1 2 103482 33489
0 33491 5 1 1 33490
0 33492 7 1 2 100637 33491
0 33493 5 1 1 33492
0 33494 7 1 2 33485 33493
0 33495 5 1 1 33494
0 33496 7 1 2 65822 33495
0 33497 5 1 1 33496
0 33498 7 1 2 33473 33497
0 33499 5 1 1 33498
0 33500 7 1 2 67343 33499
0 33501 5 1 1 33500
0 33502 7 2 2 83042 101677
0 33503 5 5 1 103484
0 33504 7 1 2 68085 85721
0 33505 5 1 1 33504
0 33506 7 1 2 103486 33505
0 33507 5 1 1 33506
0 33508 7 1 2 71428 33507
0 33509 5 1 1 33508
0 33510 7 1 2 85767 75030
0 33511 5 1 1 33510
0 33512 7 1 2 33509 33511
0 33513 5 1 1 33512
0 33514 7 1 2 69893 33513
0 33515 5 1 1 33514
0 33516 7 1 2 71429 102074
0 33517 5 1 1 33516
0 33518 7 1 2 33515 33517
0 33519 5 1 1 33518
0 33520 7 1 2 98429 33519
0 33521 5 1 1 33520
0 33522 7 1 2 33501 33521
0 33523 5 1 1 33522
0 33524 7 1 2 77357 33523
0 33525 5 1 1 33524
0 33526 7 1 2 98494 101891
0 33527 5 1 1 33526
0 33528 7 1 2 93413 98028
0 33529 5 1 1 33528
0 33530 7 1 2 33527 33529
0 33531 5 1 1 33530
0 33532 7 1 2 81743 33531
0 33533 5 1 1 33532
0 33534 7 1 2 74966 97966
0 33535 7 1 2 79204 33534
0 33536 7 1 2 79242 33535
0 33537 5 1 1 33536
0 33538 7 1 2 33533 33537
0 33539 5 1 1 33538
0 33540 7 1 2 65143 33539
0 33541 5 1 1 33540
0 33542 7 1 2 82602 76416
0 33543 5 5 1 33542
0 33544 7 1 2 79673 103491
0 33545 5 1 1 33544
0 33546 7 1 2 74547 33545
0 33547 5 1 1 33546
0 33548 7 1 2 66571 102495
0 33549 5 1 1 33548
0 33550 7 1 2 33547 33549
0 33551 5 1 1 33550
0 33552 7 1 2 65823 99272
0 33553 7 1 2 33551 33552
0 33554 5 1 1 33553
0 33555 7 1 2 33541 33554
0 33556 5 2 1 33555
0 33557 7 1 2 77164 103496
0 33558 5 1 1 33557
0 33559 7 1 2 64137 33558
0 33560 7 1 2 33525 33559
0 33561 5 1 1 33560
0 33562 7 1 2 77358 103497
0 33563 5 1 1 33562
0 33564 7 1 2 73520 83848
0 33565 7 1 2 93240 33564
0 33566 7 2 2 86545 77950
0 33567 7 1 2 102101 103498
0 33568 7 1 2 33565 33567
0 33569 5 1 1 33568
0 33570 7 1 2 69194 33569
0 33571 7 1 2 33563 33570
0 33572 5 1 1 33571
0 33573 7 1 2 73753 33572
0 33574 7 1 2 33561 33573
0 33575 5 1 1 33574
0 33576 7 2 2 72411 98743
0 33577 7 1 2 73176 102946
0 33578 5 1 1 33577
0 33579 7 1 2 76417 79412
0 33580 5 1 1 33579
0 33581 7 1 2 33578 33580
0 33582 5 1 1 33581
0 33583 7 1 2 68431 33582
0 33584 5 1 1 33583
0 33585 7 4 2 68086 80417
0 33586 5 1 1 103502
0 33587 7 3 2 71430 83972
0 33588 7 1 2 103503 103506
0 33589 5 1 1 33588
0 33590 7 1 2 33584 33589
0 33591 5 1 1 33590
0 33592 7 1 2 103500 33591
0 33593 5 1 1 33592
0 33594 7 1 2 100921 88777
0 33595 5 1 1 33594
0 33596 7 1 2 64781 33595
0 33597 5 1 1 33596
0 33598 7 2 2 68673 75627
0 33599 7 2 2 66340 83609
0 33600 5 1 1 103511
0 33601 7 1 2 103509 103512
0 33602 5 1 1 33601
0 33603 7 1 2 33597 33602
0 33604 5 1 1 33603
0 33605 7 1 2 68432 33604
0 33606 5 1 1 33605
0 33607 7 1 2 76487 90097
0 33608 5 1 1 33607
0 33609 7 1 2 33606 33608
0 33610 5 1 1 33609
0 33611 7 1 2 70474 33610
0 33612 5 1 1 33611
0 33613 7 1 2 83667 78030
0 33614 7 1 2 30415 33613
0 33615 5 1 1 33614
0 33616 7 1 2 33612 33615
0 33617 5 1 1 33616
0 33618 7 1 2 64138 97928
0 33619 7 1 2 33617 33618
0 33620 5 1 1 33619
0 33621 7 1 2 33593 33620
0 33622 5 1 1 33621
0 33623 7 1 2 75405 33622
0 33624 5 1 1 33623
0 33625 7 3 2 69195 82415
0 33626 7 1 2 77359 103513
0 33627 7 1 2 103477 33626
0 33628 5 1 1 33627
0 33629 7 1 2 33624 33628
0 33630 7 1 2 33575 33629
0 33631 7 1 2 33464 33630
0 33632 5 1 1 33631
0 33633 7 1 2 79142 33632
0 33634 5 1 1 33633
0 33635 7 1 2 84778 100021
0 33636 5 1 1 33635
0 33637 7 1 2 81744 79909
0 33638 5 1 1 33637
0 33639 7 1 2 82301 33638
0 33640 5 2 1 33639
0 33641 7 1 2 69196 103516
0 33642 5 1 1 33641
0 33643 7 1 2 33636 33642
0 33644 5 1 1 33643
0 33645 7 1 2 65144 33644
0 33646 5 1 1 33645
0 33647 7 1 2 69197 87474
0 33648 5 1 1 33647
0 33649 7 1 2 33648 82861
0 33650 5 1 1 33649
0 33651 7 1 2 64782 33650
0 33652 5 1 1 33651
0 33653 7 1 2 33646 33652
0 33654 5 1 1 33653
0 33655 7 1 2 77360 33654
0 33656 5 1 1 33655
0 33657 7 1 2 65145 103517
0 33658 5 1 1 33657
0 33659 7 2 2 64783 87475
0 33660 5 1 1 103518
0 33661 7 1 2 33658 33660
0 33662 5 3 1 33661
0 33663 7 1 2 77455 103520
0 33664 5 1 1 33663
0 33665 7 1 2 85654 75406
0 33666 5 1 1 33665
0 33667 7 1 2 33326 33666
0 33668 5 4 1 33667
0 33669 7 1 2 77250 103523
0 33670 5 1 1 33669
0 33671 7 1 2 103461 33670
0 33672 7 1 2 33664 33671
0 33673 5 1 1 33672
0 33674 7 1 2 64139 33673
0 33675 5 1 1 33674
0 33676 7 1 2 33656 33675
0 33677 5 1 1 33676
0 33678 7 1 2 65824 33677
0 33679 5 1 1 33678
0 33680 7 1 2 70830 103521
0 33681 5 1 1 33680
0 33682 7 1 2 103462 33681
0 33683 5 1 1 33682
0 33684 7 1 2 101551 33683
0 33685 5 1 1 33684
0 33686 7 1 2 67344 33685
0 33687 7 1 2 33679 33686
0 33688 5 1 1 33687
0 33689 7 1 2 100507 25697
0 33690 5 1 1 33689
0 33691 7 1 2 103522 33690
0 33692 5 1 1 33691
0 33693 7 1 2 75407 95708
0 33694 5 1 1 33693
0 33695 7 1 2 91927 33694
0 33696 5 1 1 33695
0 33697 7 1 2 103449 33696
0 33698 5 1 1 33697
0 33699 7 1 2 72412 33698
0 33700 7 1 2 33692 33699
0 33701 5 1 1 33700
0 33702 7 1 2 66341 33701
0 33703 7 1 2 33688 33702
0 33704 5 1 1 33703
0 33705 7 1 2 20412 102222
0 33706 5 1 1 33705
0 33707 7 1 2 79827 77251
0 33708 5 1 1 33707
0 33709 7 1 2 77456 96026
0 33710 5 1 1 33709
0 33711 7 1 2 33708 33710
0 33712 5 1 1 33711
0 33713 7 1 2 33706 33712
0 33714 5 1 1 33713
0 33715 7 1 2 82530 88751
0 33716 7 1 2 99477 33715
0 33717 5 1 1 33716
0 33718 7 1 2 33714 33717
0 33719 5 1 1 33718
0 33720 7 1 2 85743 33719
0 33721 5 1 1 33720
0 33722 7 1 2 33704 33721
0 33723 5 1 1 33722
0 33724 7 1 2 73177 33723
0 33725 5 1 1 33724
0 33726 7 2 2 68433 101562
0 33727 5 1 1 103527
0 33728 7 1 2 78660 84633
0 33729 5 1 1 33728
0 33730 7 1 2 33727 33729
0 33731 5 1 1 33730
0 33732 7 1 2 65146 33731
0 33733 5 1 1 33732
0 33734 7 1 2 101563 103427
0 33735 5 1 1 33734
0 33736 7 1 2 33733 33735
0 33737 5 1 1 33736
0 33738 7 1 2 64784 33737
0 33739 5 1 1 33738
0 33740 7 2 2 73521 77252
0 33741 7 1 2 92943 103529
0 33742 5 1 1 33741
0 33743 7 1 2 33739 33742
0 33744 5 1 1 33743
0 33745 7 1 2 81745 33744
0 33746 5 1 1 33745
0 33747 7 1 2 77361 77691
0 33748 7 1 2 93952 33747
0 33749 5 1 1 33748
0 33750 7 1 2 33746 33749
0 33751 5 1 1 33750
0 33752 7 1 2 64140 33751
0 33753 5 1 1 33752
0 33754 7 1 2 78289 103232
0 33755 5 1 1 33754
0 33756 7 1 2 33753 33755
0 33757 5 1 1 33756
0 33758 7 1 2 98495 33757
0 33759 5 1 1 33758
0 33760 7 1 2 100800 102103
0 33761 5 1 1 33760
0 33762 7 1 2 99186 77253
0 33763 7 1 2 91957 33762
0 33764 5 1 1 33763
0 33765 7 1 2 85744 77047
0 33766 7 1 2 98220 33765
0 33767 5 1 1 33766
0 33768 7 1 2 33764 33767
0 33769 5 1 1 33768
0 33770 7 1 2 65147 33769
0 33771 5 1 1 33770
0 33772 7 1 2 33761 33771
0 33773 5 1 1 33772
0 33774 7 1 2 64785 33773
0 33775 5 1 1 33774
0 33776 7 1 2 99187 77362
0 33777 7 1 2 81660 33776
0 33778 5 1 1 33777
0 33779 7 1 2 33775 33778
0 33780 5 1 1 33779
0 33781 7 1 2 85453 33780
0 33782 5 1 1 33781
0 33783 7 1 2 77457 86828
0 33784 5 1 1 33783
0 33785 7 1 2 71431 33784
0 33786 5 1 1 33785
0 33787 7 1 2 74673 103101
0 33788 5 1 1 33787
0 33789 7 1 2 23779 103492
0 33790 7 1 2 33788 33789
0 33791 5 1 1 33790
0 33792 7 1 2 64786 33791
0 33793 5 1 1 33792
0 33794 7 1 2 33786 33793
0 33795 5 1 1 33794
0 33796 7 1 2 68087 101489
0 33797 7 1 2 33795 33796
0 33798 5 1 1 33797
0 33799 7 1 2 74137 80458
0 33800 5 1 1 33799
0 33801 7 1 2 25620 33800
0 33802 5 1 1 33801
0 33803 7 1 2 103376 33802
0 33804 5 1 1 33803
0 33805 7 1 2 77458 103030
0 33806 5 1 1 33805
0 33807 7 2 2 64141 78005
0 33808 5 1 1 103531
0 33809 7 1 2 78290 91924
0 33810 5 1 1 33809
0 33811 7 1 2 33808 33810
0 33812 7 1 2 33806 33811
0 33813 7 1 2 33804 33812
0 33814 7 1 2 33798 33813
0 33815 5 1 1 33814
0 33816 7 1 2 72413 33815
0 33817 5 1 1 33816
0 33818 7 1 2 77459 91766
0 33819 5 1 1 33818
0 33820 7 1 2 101564 33819
0 33821 5 1 1 33820
0 33822 7 1 2 101275 33821
0 33823 5 1 1 33822
0 33824 7 1 2 81891 33823
0 33825 5 1 1 33824
0 33826 7 1 2 84910 101565
0 33827 7 1 2 102899 33826
0 33828 5 1 1 33827
0 33829 7 1 2 33825 33828
0 33830 5 1 1 33829
0 33831 7 1 2 96959 33830
0 33832 5 1 1 33831
0 33833 7 1 2 33817 33832
0 33834 5 1 1 33833
0 33835 7 1 2 65825 33834
0 33836 5 1 1 33835
0 33837 7 1 2 33782 33836
0 33838 7 1 2 33759 33837
0 33839 7 1 2 33725 33838
0 33840 5 1 1 33839
0 33841 7 1 2 78871 33840
0 33842 5 1 1 33841
0 33843 7 1 2 33634 33842
0 33844 5 1 1 33843
0 33845 7 1 2 96392 33844
0 33846 5 1 1 33845
0 33847 7 2 2 64787 80248
0 33848 5 2 1 103533
0 33849 7 1 2 87383 103534
0 33850 5 2 1 33849
0 33851 7 1 2 99854 103537
0 33852 5 1 1 33851
0 33853 7 1 2 77254 33852
0 33854 5 1 1 33853
0 33855 7 1 2 101736 33854
0 33856 5 1 1 33855
0 33857 7 1 2 72414 78366
0 33858 7 1 2 95649 33857
0 33859 7 1 2 33856 33858
0 33860 5 1 1 33859
0 33861 7 3 2 98758 76846
0 33862 7 1 2 70831 103539
0 33863 7 1 2 78006 33862
0 33864 5 1 1 33863
0 33865 7 3 2 97105 91486
0 33866 7 1 2 75925 97863
0 33867 7 1 2 103542 33866
0 33868 5 1 1 33867
0 33869 7 1 2 33864 33868
0 33870 5 1 1 33869
0 33871 7 1 2 80938 33870
0 33872 5 1 1 33871
0 33873 7 2 2 99447 84293
0 33874 7 1 2 76939 103379
0 33875 7 1 2 103545 33874
0 33876 5 1 1 33875
0 33877 7 1 2 33872 33876
0 33878 7 1 2 33860 33877
0 33879 5 1 1 33878
0 33880 7 1 2 78872 33879
0 33881 5 1 1 33880
0 33882 7 2 2 91881 76847
0 33883 7 1 2 70639 99448
0 33884 7 1 2 89086 33883
0 33885 7 1 2 103547 33884
0 33886 7 1 2 95626 33885
0 33887 5 1 1 33886
0 33888 7 1 2 33881 33887
0 33889 5 1 1 33888
0 33890 7 1 2 69198 33889
0 33891 5 1 1 33890
0 33892 7 2 2 73178 91767
0 33893 5 1 1 103549
0 33894 7 1 2 66342 103550
0 33895 5 1 1 33894
0 33896 7 1 2 103538 33895
0 33897 5 1 1 33896
0 33898 7 1 2 77255 33897
0 33899 5 1 1 33898
0 33900 7 1 2 101737 33899
0 33901 5 1 1 33900
0 33902 7 1 2 70832 33901
0 33903 5 1 1 33902
0 33904 7 1 2 65826 81192
0 33905 7 1 2 80280 33904
0 33906 5 1 1 33905
0 33907 7 1 2 33903 33906
0 33908 5 1 1 33907
0 33909 7 1 2 78172 92557
0 33910 7 1 2 103543 33909
0 33911 7 1 2 33908 33910
0 33912 5 1 1 33911
0 33913 7 1 2 33891 33912
0 33914 5 1 1 33913
0 33915 7 1 2 70475 33914
0 33916 5 1 1 33915
0 33917 7 1 2 67676 102152
0 33918 5 1 1 33917
0 33919 7 2 2 72699 6579
0 33920 5 1 1 103551
0 33921 7 1 2 73179 33920
0 33922 7 1 2 33918 33921
0 33923 5 1 1 33922
0 33924 7 1 2 83093 96043
0 33925 5 1 1 33924
0 33926 7 1 2 99949 81555
0 33927 5 1 1 33926
0 33928 7 1 2 33925 33927
0 33929 7 1 2 33923 33928
0 33930 5 1 1 33929
0 33931 7 1 2 97891 33930
0 33932 5 1 1 33931
0 33933 7 1 2 73180 86271
0 33934 7 1 2 94686 102351
0 33935 7 1 2 33933 33934
0 33936 5 1 1 33935
0 33937 7 1 2 33932 33936
0 33938 5 1 1 33937
0 33939 7 1 2 64142 33938
0 33940 5 1 1 33939
0 33941 7 3 2 67677 79990
0 33942 5 1 1 103553
0 33943 7 2 2 66572 103554
0 33944 5 2 1 103556
0 33945 7 1 2 65148 103557
0 33946 5 1 1 33945
0 33947 7 1 2 81136 87900
0 33948 5 1 1 33947
0 33949 7 1 2 33946 33948
0 33950 5 1 1 33949
0 33951 7 1 2 68434 33950
0 33952 5 1 1 33951
0 33953 7 1 2 93002 103257
0 33954 5 1 1 33953
0 33955 7 1 2 33952 33954
0 33956 5 1 1 33955
0 33957 7 1 2 33956 97971
0 33958 5 1 1 33957
0 33959 7 1 2 33940 33958
0 33960 5 1 1 33959
0 33961 7 1 2 65451 33960
0 33962 5 1 1 33961
0 33963 7 6 2 71673 72415
0 33964 7 2 2 71432 103560
0 33965 7 2 2 95385 103566
0 33966 5 1 1 103568
0 33967 7 2 2 93261 79280
0 33968 7 1 2 96867 103570
0 33969 7 1 2 103569 33968
0 33970 5 1 1 33969
0 33971 7 1 2 33962 33970
0 33972 5 1 1 33971
0 33973 7 1 2 79143 74247
0 33974 7 1 2 33972 33973
0 33975 5 1 1 33974
0 33976 7 1 2 33916 33975
0 33977 5 1 1 33976
0 33978 7 1 2 82983 33977
0 33979 5 1 1 33978
0 33980 7 1 2 33846 33979
0 33981 7 1 2 33394 33980
0 33982 5 1 1 33981
0 33983 7 1 2 72256 33982
0 33984 5 1 1 33983
0 33985 7 4 2 75926 82134
0 33986 5 3 1 103572
0 33987 7 1 2 95018 103576
0 33988 5 1 1 33987
0 33989 7 1 2 84742 33988
0 33990 5 1 1 33989
0 33991 7 1 2 87015 77048
0 33992 5 2 1 33991
0 33993 7 1 2 69894 103579
0 33994 5 2 1 33993
0 33995 7 1 2 103580 102603
0 33996 5 1 1 33995
0 33997 7 3 2 103581 33996
0 33998 7 1 2 73754 95265
0 33999 7 1 2 103583 33998
0 34000 5 1 1 33999
0 34001 7 1 2 33990 34000
0 34002 5 1 1 34001
0 34003 7 1 2 65452 34002
0 34004 5 1 1 34003
0 34005 7 1 2 85050 101408
0 34006 5 1 1 34005
0 34007 7 1 2 79848 34006
0 34008 5 1 1 34007
0 34009 7 1 2 75015 96031
0 34010 7 1 2 96027 34009
0 34011 5 1 1 34010
0 34012 7 1 2 34008 34011
0 34013 5 1 1 34012
0 34014 7 1 2 83102 34013
0 34015 5 1 1 34014
0 34016 7 1 2 34004 34015
0 34017 5 1 1 34016
0 34018 7 1 2 98430 34017
0 34019 5 1 1 34018
0 34020 7 1 2 84791 94896
0 34021 5 1 1 34020
0 34022 7 1 2 83426 83668
0 34023 5 1 1 34022
0 34024 7 1 2 34021 34023
0 34025 5 1 1 34024
0 34026 7 1 2 65827 98550
0 34027 7 1 2 86721 34026
0 34028 7 1 2 34025 34027
0 34029 5 1 1 34028
0 34030 7 1 2 34019 34029
0 34031 5 1 1 34030
0 34032 7 1 2 68435 34031
0 34033 5 1 1 34032
0 34034 7 1 2 64788 75979
0 34035 7 1 2 102210 34034
0 34036 7 3 2 67678 98551
0 34037 7 1 2 103586 88718
0 34038 7 1 2 34035 34037
0 34039 5 1 1 34038
0 34040 7 2 2 80622 98452
0 34041 5 1 1 103589
0 34042 7 1 2 82116 92092
0 34043 7 1 2 103590 34042
0 34044 5 1 1 34043
0 34045 7 1 2 34039 34044
0 34046 7 1 2 34033 34045
0 34047 5 1 1 34046
0 34048 7 1 2 77165 34047
0 34049 5 1 1 34048
0 34050 7 1 2 79814 94897
0 34051 5 1 1 34050
0 34052 7 1 2 102009 34051
0 34053 5 1 1 34052
0 34054 7 1 2 66758 34053
0 34055 5 1 1 34054
0 34056 7 1 2 85995 96890
0 34057 5 1 1 34056
0 34058 7 1 2 34055 34057
0 34059 5 1 1 34058
0 34060 7 2 2 103587 34059
0 34061 7 1 2 78316 98708
0 34062 7 1 2 103591 34061
0 34063 5 1 1 34062
0 34064 7 1 2 34049 34063
0 34065 5 1 1 34064
0 34066 7 1 2 69199 34065
0 34067 5 1 1 34066
0 34068 7 1 2 98496 77166
0 34069 5 1 1 34068
0 34070 7 2 2 97736 77990
0 34071 5 3 1 103593
0 34072 7 1 2 34069 103595
0 34073 5 2 1 34072
0 34074 7 1 2 69200 103598
0 34075 5 1 1 34074
0 34076 7 1 2 99460 77167
0 34077 5 2 1 34076
0 34078 7 2 2 34075 103600
0 34079 5 4 1 103602
0 34080 7 2 2 93003 103604
0 34081 5 1 1 103608
0 34082 7 1 2 73522 103609
0 34083 5 1 1 34082
0 34084 7 2 2 75785 85013
0 34085 5 1 1 103610
0 34086 7 1 2 99385 77168
0 34087 7 1 2 103611 34086
0 34088 5 1 1 34087
0 34089 7 1 2 34083 34088
0 34090 5 1 1 34089
0 34091 7 1 2 74674 34090
0 34092 5 1 1 34091
0 34093 7 1 2 75283 93004
0 34094 5 1 1 34093
0 34095 7 1 2 76785 90932
0 34096 5 1 1 34095
0 34097 7 1 2 34094 34096
0 34098 5 1 1 34097
0 34099 7 1 2 100527 34098
0 34100 5 1 1 34099
0 34101 7 1 2 70208 75016
0 34102 7 1 2 77612 34101
0 34103 5 1 1 34102
0 34104 7 1 2 21689 34103
0 34105 5 1 1 34104
0 34106 7 1 2 83989 34105
0 34107 5 1 1 34106
0 34108 7 1 2 89815 87802
0 34109 5 1 1 34108
0 34110 7 1 2 34107 34109
0 34111 5 1 1 34110
0 34112 7 5 2 72416 95636
0 34113 7 5 2 95336 103612
0 34114 7 1 2 34111 103617
0 34115 5 1 1 34114
0 34116 7 1 2 34100 34115
0 34117 7 1 2 34092 34116
0 34118 5 1 1 34117
0 34119 7 1 2 81746 34118
0 34120 5 1 1 34119
0 34121 7 1 2 93005 93749
0 34122 5 1 1 34121
0 34123 7 4 2 72700 74792
0 34124 7 1 2 84084 103622
0 34125 7 1 2 79490 34124
0 34126 5 1 1 34125
0 34127 7 1 2 34122 34126
0 34128 5 1 1 34127
0 34129 7 1 2 103605 34128
0 34130 5 1 1 34129
0 34131 7 1 2 97124 99318
0 34132 5 1 1 34131
0 34133 7 1 2 70833 102039
0 34134 5 1 1 34133
0 34135 7 1 2 34132 34134
0 34136 5 1 1 34135
0 34137 7 1 2 77169 34136
0 34138 5 1 1 34137
0 34139 7 2 2 64425 99134
0 34140 7 1 2 82388 97125
0 34141 7 1 2 103626 34140
0 34142 5 1 1 34141
0 34143 7 1 2 34138 34142
0 34144 5 1 1 34143
0 34145 7 1 2 69201 34144
0 34146 5 1 1 34145
0 34147 7 1 2 100797 83349
0 34148 7 1 2 102300 34147
0 34149 5 1 1 34148
0 34150 7 1 2 34146 34149
0 34151 5 1 1 34150
0 34152 7 1 2 82117 98985
0 34153 7 1 2 34151 34152
0 34154 5 1 1 34153
0 34155 7 1 2 34130 34154
0 34156 7 1 2 34120 34155
0 34157 7 1 2 73921 102535
0 34158 5 1 1 34157
0 34159 7 1 2 98431 92581
0 34160 7 1 2 100923 34159
0 34161 5 1 1 34160
0 34162 7 1 2 34158 34161
0 34163 5 1 1 34162
0 34164 7 1 2 70209 34163
0 34165 5 1 1 34164
0 34166 7 1 2 76161 75060
0 34167 5 1 1 34166
0 34168 7 2 2 73969 78704
0 34169 7 1 2 75637 76050
0 34170 7 1 2 103628 34169
0 34171 5 1 1 34170
0 34172 7 1 2 34167 34171
0 34173 5 1 1 34172
0 34174 7 1 2 98453 34173
0 34175 5 1 1 34174
0 34176 7 1 2 34165 34175
0 34177 5 1 1 34176
0 34178 7 1 2 77170 34177
0 34179 5 1 1 34178
0 34180 7 1 2 91134 97636
0 34181 7 1 2 102595 34180
0 34182 5 1 1 34181
0 34183 7 1 2 69202 34182
0 34184 7 1 2 34179 34183
0 34185 5 1 1 34184
0 34186 7 1 2 77171 102596
0 34187 5 1 1 34186
0 34188 7 1 2 99304 98709
0 34189 5 1 1 34188
0 34190 7 1 2 34187 34189
0 34191 5 1 1 34190
0 34192 7 1 2 81309 34191
0 34193 5 1 1 34192
0 34194 7 1 2 64143 34193
0 34195 5 1 1 34194
0 34196 7 1 2 81892 34195
0 34197 7 1 2 34185 34196
0 34198 5 1 1 34197
0 34199 7 4 2 82246 102127
0 34200 7 1 2 101203 103630
0 34201 5 1 1 34200
0 34202 7 2 2 101033 92955
0 34203 5 1 1 103634
0 34204 7 1 2 34201 34203
0 34205 5 1 1 34204
0 34206 7 1 2 75408 34205
0 34207 5 1 1 34206
0 34208 7 1 2 74548 90990
0 34209 7 1 2 101034 34208
0 34210 5 1 1 34209
0 34211 7 1 2 34207 34210
0 34212 5 1 1 34211
0 34213 7 1 2 80623 34212
0 34214 5 1 1 34213
0 34215 7 1 2 74549 103635
0 34216 5 1 1 34215
0 34217 7 1 2 34214 34216
0 34218 5 1 1 34217
0 34219 7 1 2 71433 34218
0 34220 5 1 1 34219
0 34221 7 1 2 34198 34220
0 34222 7 1 2 34156 34221
0 34223 5 1 1 34222
0 34224 7 1 2 69895 34223
0 34225 5 1 1 34224
0 34226 7 1 2 100562 103592
0 34227 5 1 1 34226
0 34228 7 1 2 64789 94194
0 34229 5 1 1 34228
0 34230 7 1 2 68436 94171
0 34231 5 1 1 34230
0 34232 7 1 2 34229 34231
0 34233 5 1 1 34232
0 34234 7 1 2 100528 34233
0 34235 5 1 1 34234
0 34236 7 1 2 83573 97607
0 34237 5 2 1 34236
0 34238 7 5 2 69203 74335
0 34239 7 1 2 98248 103638
0 34240 7 1 2 103636 34239
0 34241 5 1 1 34240
0 34242 7 1 2 34235 34241
0 34243 5 1 1 34242
0 34244 7 1 2 93006 34243
0 34245 5 1 1 34244
0 34246 7 1 2 34227 34245
0 34247 7 1 2 34225 34246
0 34248 7 1 2 34067 34247
0 34249 5 1 1 34248
0 34250 7 1 2 76848 34249
0 34251 5 1 1 34250
0 34252 7 2 2 73755 103631
0 34253 7 1 2 74922 96236
0 34254 7 3 2 66573 84598
0 34255 7 1 2 93424 103645
0 34256 7 1 2 34253 34255
0 34257 7 1 2 103643 34256
0 34258 5 1 1 34257
0 34259 7 1 2 34251 34258
0 34260 5 1 1 34259
0 34261 7 1 2 79144 34260
0 34262 5 1 1 34261
0 34263 7 2 2 75409 92767
0 34264 5 1 1 103648
0 34265 7 1 2 87247 103649
0 34266 5 3 1 34265
0 34267 7 2 2 64790 80869
0 34268 5 3 1 103653
0 34269 7 1 2 23846 103655
0 34270 5 1 1 34269
0 34271 7 2 2 73181 34270
0 34272 5 1 1 103658
0 34273 7 1 2 71096 103659
0 34274 5 1 1 34273
0 34275 7 1 2 103650 34274
0 34276 5 1 1 34275
0 34277 7 1 2 71836 34276
0 34278 5 1 1 34277
0 34279 7 1 2 75609 94510
0 34280 5 1 1 34279
0 34281 7 1 2 103651 34280
0 34282 5 1 1 34281
0 34283 7 1 2 68674 34282
0 34284 5 1 1 34283
0 34285 7 1 2 34278 34284
0 34286 5 1 1 34285
0 34287 7 1 2 67679 34286
0 34288 5 1 1 34287
0 34289 7 1 2 68675 101781
0 34290 5 1 1 34289
0 34291 7 1 2 86515 34290
0 34292 5 1 1 34291
0 34293 7 1 2 77460 92665
0 34294 7 1 2 34292 34293
0 34295 5 1 1 34294
0 34296 7 1 2 34288 34295
0 34297 5 1 1 34296
0 34298 7 1 2 70476 34297
0 34299 5 1 1 34298
0 34300 7 1 2 81149 97215
0 34301 5 1 1 34300
0 34302 7 1 2 101396 9172
0 34303 5 1 1 34302
0 34304 7 1 2 94324 34303
0 34305 5 1 1 34304
0 34306 7 3 2 69896 78435
0 34307 5 2 1 103660
0 34308 7 1 2 80939 103661
0 34309 5 1 1 34308
0 34310 7 1 2 34305 34309
0 34311 5 1 1 34310
0 34312 7 1 2 80364 34311
0 34313 5 1 1 34312
0 34314 7 1 2 34301 34313
0 34315 7 1 2 34299 34314
0 34316 5 1 1 34315
0 34317 7 1 2 67345 34316
0 34318 5 1 1 34317
0 34319 7 6 2 77172 97046
0 34320 5 3 1 103665
0 34321 7 2 2 69897 103666
0 34322 7 1 2 101833 103674
0 34323 5 1 1 34322
0 34324 7 1 2 34318 34323
0 34325 5 1 1 34324
0 34326 7 1 2 65828 34325
0 34327 5 1 1 34326
0 34328 7 2 2 79849 92582
0 34329 7 1 2 101103 103676
0 34330 5 1 1 34329
0 34331 7 1 2 80897 98517
0 34332 5 1 1 34331
0 34333 7 1 2 34330 34332
0 34334 5 1 1 34333
0 34335 7 1 2 99796 34334
0 34336 5 1 1 34335
0 34337 7 1 2 79281 14793
0 34338 5 1 1 34337
0 34339 7 1 2 82170 101712
0 34340 5 1 1 34339
0 34341 7 1 2 34338 34340
0 34342 5 1 1 34341
0 34343 7 1 2 71837 34342
0 34344 5 1 1 34343
0 34345 7 1 2 26186 34344
0 34346 5 1 1 34345
0 34347 7 1 2 70477 34346
0 34348 5 1 1 34347
0 34349 7 1 2 85593 92768
0 34350 5 1 1 34349
0 34351 7 1 2 34348 34350
0 34352 5 1 1 34351
0 34353 7 1 2 97047 34352
0 34354 5 1 1 34353
0 34355 7 1 2 34336 34354
0 34356 5 1 1 34355
0 34357 7 1 2 70834 34356
0 34358 5 1 1 34357
0 34359 7 1 2 69898 88759
0 34360 5 1 1 34359
0 34361 7 1 2 102911 34360
0 34362 5 1 1 34361
0 34363 7 1 2 77461 34362
0 34364 5 1 1 34363
0 34365 7 1 2 80898 101298
0 34366 5 1 1 34365
0 34367 7 1 2 34364 34366
0 34368 5 1 1 34367
0 34369 7 1 2 72701 34368
0 34370 5 1 1 34369
0 34371 7 1 2 85745 78481
0 34372 7 1 2 94910 34371
0 34373 5 1 1 34372
0 34374 7 1 2 34370 34373
0 34375 5 1 1 34374
0 34376 7 1 2 98497 34375
0 34377 5 1 1 34376
0 34378 7 1 2 86253 86034
0 34379 5 1 1 34378
0 34380 7 1 2 18985 98252
0 34381 5 2 1 34380
0 34382 7 1 2 67680 92382
0 34383 7 1 2 103678 34382
0 34384 7 1 2 34379 34383
0 34385 5 1 1 34384
0 34386 7 1 2 34377 34385
0 34387 7 1 2 34358 34386
0 34388 5 1 1 34387
0 34389 7 1 2 68088 34388
0 34390 5 1 1 34389
0 34391 7 1 2 88760 83792
0 34392 5 1 1 34391
0 34393 7 1 2 80805 34392
0 34394 5 3 1 34393
0 34395 7 2 2 69899 98432
0 34396 7 1 2 97681 103683
0 34397 7 1 2 103680 34396
0 34398 5 1 1 34397
0 34399 7 1 2 69204 34398
0 34400 7 1 2 34390 34399
0 34401 7 1 2 34327 34400
0 34402 5 1 1 34401
0 34403 7 1 2 86057 81193
0 34404 5 1 1 34403
0 34405 7 1 2 101362 34404
0 34406 5 2 1 34405
0 34407 7 1 2 103675 103685
0 34408 5 1 1 34407
0 34409 7 1 2 67681 34272
0 34410 5 1 1 34409
0 34411 7 1 2 68089 94552
0 34412 7 1 2 103535 34411
0 34413 5 1 1 34412
0 34414 7 1 2 72702 103483
0 34415 7 1 2 34413 34414
0 34416 5 1 1 34415
0 34417 7 1 2 71097 34416
0 34418 7 1 2 34410 34417
0 34419 5 1 1 34418
0 34420 7 1 2 78446 98566
0 34421 5 1 1 34420
0 34422 7 1 2 74550 34421
0 34423 5 1 1 34422
0 34424 7 1 2 93202 34423
0 34425 5 1 1 34424
0 34426 7 1 2 69900 34425
0 34427 5 1 1 34426
0 34428 7 4 2 69534 85014
0 34429 5 2 1 103687
0 34430 7 1 2 64791 103688
0 34431 5 1 1 34430
0 34432 7 1 2 103663 34431
0 34433 5 1 1 34432
0 34434 7 1 2 80230 34433
0 34435 5 1 1 34434
0 34436 7 1 2 34427 34435
0 34437 7 1 2 34419 34436
0 34438 5 1 1 34437
0 34439 7 1 2 71838 34438
0 34440 5 1 1 34439
0 34441 7 2 2 81194 92666
0 34442 5 1 1 103693
0 34443 7 1 2 101397 34442
0 34444 5 2 1 34443
0 34445 7 1 2 94511 103695
0 34446 5 1 1 34445
0 34447 7 3 2 67682 92769
0 34448 7 1 2 81195 103697
0 34449 5 1 1 34448
0 34450 7 1 2 34446 34449
0 34451 5 1 1 34450
0 34452 7 1 2 68676 34451
0 34453 5 1 1 34452
0 34454 7 1 2 70478 34453
0 34455 7 1 2 34440 34454
0 34456 5 1 1 34455
0 34457 7 1 2 64792 90124
0 34458 5 1 1 34457
0 34459 7 1 2 96897 88459
0 34460 5 1 1 34459
0 34461 7 1 2 34458 34460
0 34462 5 1 1 34461
0 34463 7 1 2 67683 34462
0 34464 5 1 1 34463
0 34465 7 1 2 80365 103694
0 34466 5 1 1 34465
0 34467 7 1 2 34464 34466
0 34468 5 1 1 34467
0 34469 7 1 2 71098 34468
0 34470 5 1 1 34469
0 34471 7 4 2 69535 71839
0 34472 7 1 2 68677 103700
0 34473 7 1 2 103696 34472
0 34474 5 1 1 34473
0 34475 7 1 2 65453 34474
0 34476 7 1 2 34470 34475
0 34477 5 1 1 34476
0 34478 7 1 2 34456 34477
0 34479 5 1 1 34478
0 34480 7 1 2 103698 103377
0 34481 5 1 1 34480
0 34482 7 1 2 34479 34481
0 34483 5 1 1 34482
0 34484 7 1 2 67346 34483
0 34485 5 1 1 34484
0 34486 7 1 2 34408 34485
0 34487 5 1 1 34486
0 34488 7 1 2 70835 34487
0 34489 5 1 1 34488
0 34490 7 2 2 74064 98759
0 34491 5 2 1 103704
0 34492 7 1 2 76959 103705
0 34493 7 1 2 103686 34492
0 34494 5 1 1 34493
0 34495 7 1 2 64144 34494
0 34496 7 1 2 34489 34495
0 34497 5 1 1 34496
0 34498 7 1 2 71434 34497
0 34499 7 1 2 34402 34498
0 34500 5 1 1 34499
0 34501 7 1 2 90769 89242
0 34502 5 1 1 34501
0 34503 7 1 2 77256 34502
0 34504 5 1 1 34503
0 34505 7 1 2 82567 93092
0 34506 5 2 1 34505
0 34507 7 1 2 34504 103708
0 34508 5 1 1 34507
0 34509 7 1 2 67347 34508
0 34510 5 1 1 34509
0 34511 7 1 2 97464 97561
0 34512 5 1 1 34511
0 34513 7 1 2 34510 34512
0 34514 5 1 1 34513
0 34515 7 1 2 64793 34514
0 34516 5 1 1 34515
0 34517 7 1 2 95212 97126
0 34518 5 1 1 34517
0 34519 7 1 2 34516 34518
0 34520 5 1 1 34519
0 34521 7 1 2 78661 34520
0 34522 5 1 1 34521
0 34523 7 3 2 100788 98657
0 34524 5 1 1 103710
0 34525 7 1 2 29245 103711
0 34526 5 1 1 34525
0 34527 7 1 2 34522 34526
0 34528 5 1 1 34527
0 34529 7 1 2 80870 34528
0 34530 5 1 1 34529
0 34531 7 1 2 80231 86182
0 34532 5 2 1 34531
0 34533 7 1 2 2482 80803
0 34534 5 1 1 34533
0 34535 7 1 2 80624 34534
0 34536 5 1 1 34535
0 34537 7 1 2 76657 88761
0 34538 5 1 1 34537
0 34539 7 1 2 34536 34538
0 34540 7 1 2 103713 34539
0 34541 5 1 1 34540
0 34542 7 1 2 98406 34541
0 34543 5 1 1 34542
0 34544 7 3 2 67684 98610
0 34545 5 1 1 103715
0 34546 7 1 2 71840 94937
0 34547 5 1 1 34546
0 34548 7 1 2 88762 91768
0 34549 5 1 1 34548
0 34550 7 1 2 3038 34549
0 34551 7 1 2 34547 34550
0 34552 5 1 1 34551
0 34553 7 1 2 103716 34552
0 34554 5 1 1 34553
0 34555 7 1 2 34543 34554
0 34556 5 1 1 34555
0 34557 7 1 2 66343 34556
0 34558 5 1 1 34557
0 34559 7 1 2 80232 98287
0 34560 5 1 1 34559
0 34561 7 1 2 29439 34560
0 34562 5 1 1 34561
0 34563 7 1 2 86835 34562
0 34564 5 1 1 34563
0 34565 7 1 2 34558 34564
0 34566 5 1 1 34565
0 34567 7 1 2 73182 34566
0 34568 5 1 1 34567
0 34569 7 1 2 2002 89243
0 34570 5 1 1 34569
0 34571 7 1 2 98273 34570
0 34572 5 1 1 34571
0 34573 7 2 2 69536 77521
0 34574 7 1 2 99188 85015
0 34575 7 1 2 103718 34574
0 34576 5 1 1 34575
0 34577 7 1 2 34572 34576
0 34578 5 1 1 34577
0 34579 7 1 2 64794 34578
0 34580 5 1 1 34579
0 34581 7 1 2 88763 81196
0 34582 5 1 1 34581
0 34583 7 1 2 34582 80806
0 34584 5 1 1 34583
0 34585 7 1 2 98234 81467
0 34586 7 1 2 34584 34585
0 34587 5 1 1 34586
0 34588 7 1 2 34580 34587
0 34589 7 1 2 34568 34588
0 34590 7 1 2 34530 34589
0 34591 5 1 1 34590
0 34592 7 1 2 82444 34591
0 34593 5 1 1 34592
0 34594 7 1 2 95330 93162
0 34595 5 1 1 34594
0 34596 7 2 2 68437 75107
0 34597 7 1 2 84710 103720
0 34598 5 1 1 34597
0 34599 7 1 2 100746 34598
0 34600 5 1 1 34599
0 34601 7 1 2 73183 34600
0 34602 5 1 1 34601
0 34603 7 1 2 64795 100644
0 34604 7 1 2 83432 34603
0 34605 5 1 1 34604
0 34606 7 1 2 68090 86178
0 34607 7 1 2 22912 34606
0 34608 7 1 2 34605 34607
0 34609 5 1 1 34608
0 34610 7 1 2 34602 34609
0 34611 5 1 1 34610
0 34612 7 1 2 67685 34611
0 34613 5 1 1 34612
0 34614 7 1 2 34595 34613
0 34615 5 1 1 34614
0 34616 7 1 2 99403 34615
0 34617 5 1 1 34616
0 34618 7 1 2 95386 103079
0 34619 5 1 1 34618
0 34620 7 1 2 80625 101410
0 34621 5 1 1 34620
0 34622 7 1 2 34619 34621
0 34623 5 1 1 34622
0 34624 7 1 2 99386 34623
0 34625 5 1 1 34624
0 34626 7 1 2 34617 34625
0 34627 5 1 1 34626
0 34628 7 1 2 71099 34627
0 34629 5 1 1 34628
0 34630 7 1 2 103080 103528
0 34631 5 1 1 34630
0 34632 7 1 2 99847 87167
0 34633 5 1 1 34632
0 34634 7 1 2 34631 34633
0 34635 5 1 1 34634
0 34636 7 1 2 96751 34635
0 34637 5 1 1 34636
0 34638 7 2 2 98029 95266
0 34639 7 1 2 70479 81325
0 34640 7 1 2 103722 34639
0 34641 5 1 1 34640
0 34642 7 1 2 34637 34641
0 34643 5 1 1 34642
0 34644 7 1 2 82445 34643
0 34645 5 1 1 34644
0 34646 7 1 2 34629 34645
0 34647 5 1 1 34646
0 34648 7 1 2 74675 34647
0 34649 5 1 1 34648
0 34650 7 1 2 80233 82198
0 34651 5 1 1 34650
0 34652 7 1 2 103691 34651
0 34653 5 1 1 34652
0 34654 7 1 2 64796 34653
0 34655 5 1 1 34654
0 34656 7 1 2 81468 103536
0 34657 5 1 1 34656
0 34658 7 1 2 69901 101403
0 34659 5 1 1 34658
0 34660 7 1 2 34657 34659
0 34661 5 1 1 34660
0 34662 7 1 2 73184 34661
0 34663 5 1 1 34662
0 34664 7 1 2 34655 34663
0 34665 5 1 1 34664
0 34666 7 1 2 80626 34665
0 34667 5 1 1 34666
0 34668 7 1 2 64426 95040
0 34669 5 1 1 34668
0 34670 7 1 2 83938 34669
0 34671 5 1 1 34670
0 34672 7 1 2 34667 34671
0 34673 5 1 1 34672
0 34674 7 1 2 71100 34673
0 34675 5 1 1 34674
0 34676 7 1 2 78411 87540
0 34677 5 1 1 34676
0 34678 7 1 2 87098 5296
0 34679 5 1 1 34678
0 34680 7 1 2 75628 82199
0 34681 7 1 2 34679 34680
0 34682 5 1 1 34681
0 34683 7 1 2 34677 34682
0 34684 5 1 1 34683
0 34685 7 1 2 69537 34684
0 34686 5 1 1 34685
0 34687 7 3 2 67686 76874
0 34688 5 1 1 103724
0 34689 7 1 2 69902 103725
0 34690 7 1 2 88729 34689
0 34691 5 1 1 34690
0 34692 7 1 2 34686 34691
0 34693 5 1 1 34692
0 34694 7 1 2 68678 34693
0 34695 5 1 1 34694
0 34696 7 1 2 68091 85630
0 34697 5 2 1 34696
0 34698 7 1 2 98666 103727
0 34699 5 1 1 34698
0 34700 7 1 2 34699 92875
0 34701 5 1 1 34700
0 34702 7 1 2 92554 92197
0 34703 5 1 1 34702
0 34704 7 1 2 77462 34703
0 34705 7 1 2 103681 34704
0 34706 5 1 1 34705
0 34707 7 1 2 34701 34706
0 34708 7 1 2 34695 34707
0 34709 7 1 2 34675 34708
0 34710 5 1 1 34709
0 34711 7 1 2 99404 34710
0 34712 5 1 1 34711
0 34713 7 1 2 34649 34712
0 34714 7 1 2 34593 34713
0 34715 7 1 2 34500 34714
0 34716 5 1 1 34715
0 34717 7 1 2 76849 34716
0 34718 5 1 1 34717
0 34719 7 4 2 68092 96752
0 34720 7 2 2 73756 78317
0 34721 5 1 1 103733
0 34722 7 1 2 71101 34721
0 34723 5 1 1 34722
0 34724 7 1 2 103729 34723
0 34725 5 1 1 34724
0 34726 7 1 2 101947 34725
0 34727 5 1 1 34726
0 34728 7 1 2 80627 34727
0 34729 5 1 1 34728
0 34730 7 1 2 77588 101075
0 34731 7 1 2 89056 34730
0 34732 5 1 1 34731
0 34733 7 1 2 34729 34732
0 34734 5 1 1 34733
0 34735 7 1 2 64427 34734
0 34736 5 1 1 34735
0 34737 7 1 2 66344 78457
0 34738 7 1 2 95031 34737
0 34739 5 1 1 34738
0 34740 7 1 2 66027 79769
0 34741 7 1 2 93163 34740
0 34742 5 1 1 34741
0 34743 7 1 2 34739 34742
0 34744 5 1 1 34743
0 34745 7 1 2 67348 34744
0 34746 5 1 1 34745
0 34747 7 2 2 71102 79770
0 34748 7 1 2 103723 103735
0 34749 5 1 1 34748
0 34750 7 1 2 34746 34749
0 34751 5 1 1 34750
0 34752 7 1 2 89257 34751
0 34753 5 1 1 34752
0 34754 7 1 2 34736 34753
0 34755 5 1 1 34754
0 34756 7 1 2 70836 34755
0 34757 5 1 1 34756
0 34758 7 2 2 84162 101076
0 34759 7 1 2 83973 74065
0 34760 7 1 2 103737 34759
0 34761 5 1 1 34760
0 34762 7 1 2 34757 34761
0 34763 5 1 1 34762
0 34764 7 1 2 69205 34763
0 34765 5 1 1 34764
0 34766 7 2 2 70837 85418
0 34767 7 1 2 77522 103739
0 34768 7 1 2 103738 34767
0 34769 5 1 1 34768
0 34770 7 1 2 34765 34769
0 34771 5 1 1 34770
0 34772 7 1 2 76850 34771
0 34773 5 1 1 34772
0 34774 7 4 2 82319 98963
0 34775 7 2 2 101552 96161
0 34776 7 1 2 103745 74248
0 34777 7 1 2 103741 34776
0 34778 5 1 1 34777
0 34779 7 1 2 34773 34778
0 34780 5 1 1 34779
0 34781 7 1 2 73970 34780
0 34782 5 1 1 34781
0 34783 7 4 2 85520 98940
0 34784 7 1 2 86058 103747
0 34785 5 1 1 34784
0 34786 7 1 2 100508 34785
0 34787 5 1 1 34786
0 34788 7 1 2 66574 34787
0 34789 5 1 1 34788
0 34790 7 1 2 744 34789
0 34791 5 1 1 34790
0 34792 7 1 2 65149 34791
0 34793 5 1 1 34792
0 34794 7 1 2 100498 94732
0 34795 5 1 1 34794
0 34796 7 3 2 73523 88764
0 34797 7 1 2 103748 103751
0 34798 5 1 1 34797
0 34799 7 1 2 34795 34798
0 34800 5 1 1 34799
0 34801 7 1 2 74676 34800
0 34802 5 1 1 34801
0 34803 7 2 2 69206 81108
0 34804 5 1 1 103754
0 34805 7 1 2 77991 103755
0 34806 7 1 2 86794 34805
0 34807 5 1 1 34806
0 34808 7 1 2 34802 34807
0 34809 7 1 2 34793 34808
0 34810 5 1 1 34809
0 34811 7 1 2 103540 34810
0 34812 5 1 1 34811
0 34813 7 4 2 67122 98760
0 34814 7 2 2 69207 95619
0 34815 7 2 2 103756 103760
0 34816 5 1 1 103762
0 34817 7 1 2 73757 103763
0 34818 5 1 1 34817
0 34819 7 1 2 101976 103544
0 34820 5 1 1 34819
0 34821 7 1 2 34818 34820
0 34822 5 1 1 34821
0 34823 7 1 2 64428 34822
0 34824 5 1 1 34823
0 34825 7 2 2 73758 82446
0 34826 7 3 2 67349 76851
0 34827 7 1 2 78458 103766
0 34828 7 1 2 103764 34827
0 34829 5 1 1 34828
0 34830 7 1 2 34824 34829
0 34831 5 2 1 34830
0 34832 7 1 2 83669 89195
0 34833 7 1 2 103769 34832
0 34834 5 1 1 34833
0 34835 7 1 2 34812 34834
0 34836 5 1 1 34835
0 34837 7 1 2 76597 34836
0 34838 5 1 1 34837
0 34839 7 1 2 100726 103770
0 34840 5 1 1 34839
0 34841 7 1 2 100499 91498
0 34842 7 1 2 103767 34841
0 34843 5 1 1 34842
0 34844 7 1 2 34840 34843
0 34845 5 1 1 34844
0 34846 7 1 2 64797 34845
0 34847 5 1 1 34846
0 34848 7 1 2 71435 87286
0 34849 5 1 1 34848
0 34850 7 1 2 103541 78300
0 34851 7 1 2 34849 34850
0 34852 5 1 1 34851
0 34853 7 1 2 34847 34852
0 34854 5 1 1 34853
0 34855 7 1 2 87037 34854
0 34856 5 1 1 34855
0 34857 7 2 2 96265 96018
0 34858 7 1 2 102212 94891
0 34859 7 1 2 103771 34858
0 34860 5 1 1 34859
0 34861 7 1 2 34856 34860
0 34862 7 1 2 34838 34861
0 34863 7 1 2 34782 34862
0 34864 7 1 2 34718 34863
0 34865 5 1 1 34864
0 34866 7 1 2 78873 34865
0 34867 5 1 1 34866
0 34868 7 1 2 34262 34867
0 34869 5 1 1 34868
0 34870 7 1 2 67199 34869
0 34871 5 1 1 34870
0 34872 7 2 2 72257 98695
0 34873 7 1 2 74249 78137
0 34874 7 1 2 103773 34873
0 34875 5 2 1 34874
0 34876 7 3 2 100152 95650
0 34877 7 1 2 99994 103777
0 34878 5 1 1 34877
0 34879 7 2 2 77173 95620
0 34880 7 1 2 80366 102543
0 34881 7 1 2 103780 34880
0 34882 5 1 1 34881
0 34883 7 1 2 34878 34882
0 34884 5 1 1 34883
0 34885 7 1 2 64145 34884
0 34886 5 1 1 34885
0 34887 7 1 2 84839 77066
0 34888 5 1 1 34887
0 34889 7 1 2 71841 92815
0 34890 5 1 1 34889
0 34891 7 1 2 34888 34890
0 34892 5 1 1 34891
0 34893 7 3 2 76852 102465
0 34894 7 1 2 68679 103782
0 34895 7 1 2 34892 34894
0 34896 5 1 1 34895
0 34897 7 1 2 34886 34896
0 34898 5 1 1 34897
0 34899 7 1 2 67687 34898
0 34900 5 1 1 34899
0 34901 7 3 2 67002 102573
0 34902 7 2 2 101973 103785
0 34903 5 1 1 103788
0 34904 7 3 2 67200 76853
0 34905 7 2 2 84840 103790
0 34906 7 1 2 82447 103793
0 34907 5 1 1 34906
0 34908 7 1 2 34903 34907
0 34909 5 1 1 34908
0 34910 7 1 2 101066 34909
0 34911 5 1 1 34910
0 34912 7 1 2 34900 34911
0 34913 5 1 1 34912
0 34914 7 1 2 72417 34913
0 34915 5 1 1 34914
0 34916 7 2 2 66028 95267
0 34917 5 2 1 103795
0 34918 7 1 2 84841 92966
0 34919 5 1 1 34918
0 34920 7 1 2 103797 34919
0 34921 5 1 1 34920
0 34922 7 1 2 85521 34921
0 34923 5 1 1 34922
0 34924 7 1 2 95268 78138
0 34925 5 1 1 34924
0 34926 7 1 2 34923 34925
0 34927 5 1 1 34926
0 34928 7 1 2 67201 34927
0 34929 5 1 1 34928
0 34930 7 4 2 95350 100138
0 34931 5 1 1 103799
0 34932 7 1 2 95269 103800
0 34933 5 1 1 34932
0 34934 7 1 2 34929 34933
0 34935 5 1 1 34934
0 34936 7 1 2 79054 97437
0 34937 7 1 2 34935 34936
0 34938 5 1 1 34937
0 34939 7 1 2 34915 34938
0 34940 5 1 1 34939
0 34941 7 1 2 75580 34940
0 34942 5 1 1 34941
0 34943 7 1 2 103775 34942
0 34944 5 1 1 34943
0 34945 7 1 2 75410 34944
0 34946 5 1 1 34945
0 34947 7 1 2 99478 103794
0 34948 5 1 1 34947
0 34949 7 1 2 72418 103789
0 34950 5 1 1 34949
0 34951 7 1 2 34948 34950
0 34952 5 1 1 34951
0 34953 7 1 2 68680 34952
0 34954 5 1 1 34953
0 34955 7 2 2 103786 97568
0 34956 7 1 2 77692 103803
0 34957 5 1 1 34956
0 34958 7 1 2 34954 34957
0 34959 5 1 1 34958
0 34960 7 1 2 92547 34959
0 34961 5 1 1 34960
0 34962 7 1 2 34946 34961
0 34963 5 1 1 34962
0 34964 7 1 2 78874 34963
0 34965 5 1 1 34964
0 34966 7 1 2 92967 103804
0 34967 5 1 1 34966
0 34968 7 1 2 85522 103679
0 34969 5 1 1 34968
0 34970 7 1 2 97900 101004
0 34971 5 1 1 34970
0 34972 7 1 2 34969 34971
0 34973 5 1 1 34972
0 34974 7 1 2 67202 34973
0 34975 5 1 1 34974
0 34976 7 1 2 23351 34975
0 34977 5 1 1 34976
0 34978 7 1 2 67688 76854
0 34979 7 1 2 34977 34978
0 34980 5 1 1 34979
0 34981 7 1 2 34967 34980
0 34982 5 1 1 34981
0 34983 7 1 2 87831 34982
0 34984 5 1 1 34983
0 34985 7 1 2 34984 103776
0 34986 5 1 1 34985
0 34987 7 2 2 98216 77906
0 34988 7 1 2 34986 103805
0 34989 5 1 1 34988
0 34990 7 2 2 74491 89900
0 34991 7 1 2 100083 82791
0 34992 7 1 2 96527 86090
0 34993 7 1 2 34991 34992
0 34994 7 1 2 95560 34993
0 34995 7 1 2 103807 34994
0 34996 5 1 1 34995
0 34997 7 1 2 34989 34996
0 34998 5 1 1 34997
0 34999 7 1 2 82984 34998
0 35000 5 1 1 34999
0 35001 7 1 2 71952 94012
0 35002 7 2 2 84505 35001
0 35003 7 1 2 97879 103809
0 35004 5 1 1 35003
0 35005 7 1 2 80528 78875
0 35006 7 1 2 92540 35005
0 35007 5 1 1 35006
0 35008 7 1 2 35004 35007
0 35009 5 1 1 35008
0 35010 7 1 2 98030 35009
0 35011 5 1 1 35010
0 35012 7 3 2 78990 88351
0 35013 7 2 2 73185 97901
0 35014 7 1 2 79519 103814
0 35015 7 1 2 103811 35014
0 35016 7 1 2 84121 35015
0 35017 5 1 1 35016
0 35018 7 1 2 35011 35017
0 35019 5 1 1 35018
0 35020 7 1 2 103787 35019
0 35021 5 1 1 35020
0 35022 7 1 2 84770 83686
0 35023 7 3 2 87574 35022
0 35024 5 1 1 103816
0 35025 7 2 2 77463 103817
0 35026 7 3 2 84473 102544
0 35027 7 6 2 78173 95740
0 35028 7 1 2 67350 103824
0 35029 7 1 2 103821 35028
0 35030 7 1 2 103819 35029
0 35031 5 1 1 35030
0 35032 7 1 2 35021 35031
0 35033 5 1 1 35032
0 35034 7 1 2 64146 35033
0 35035 5 1 1 35034
0 35036 7 3 2 102545 99283
0 35037 7 1 2 98498 103830
0 35038 7 1 2 103820 35037
0 35039 5 1 1 35038
0 35040 7 1 2 83293 79145
0 35041 7 3 2 72419 82932
0 35042 7 1 2 103833 103010
0 35043 7 1 2 96136 35042
0 35044 7 1 2 35040 35043
0 35045 5 1 1 35044
0 35046 7 1 2 35039 35045
0 35047 5 1 1 35046
0 35048 7 1 2 95569 35047
0 35049 5 1 1 35048
0 35050 7 1 2 35035 35049
0 35051 5 1 1 35050
0 35052 7 1 2 72703 35051
0 35053 5 1 1 35052
0 35054 7 1 2 80529 102546
0 35055 7 1 2 103781 35054
0 35056 5 1 1 35055
0 35057 7 1 2 82649 77257
0 35058 7 1 2 103778 35057
0 35059 5 1 1 35058
0 35060 7 1 2 35056 35059
0 35061 5 1 1 35060
0 35062 7 1 2 64147 35061
0 35063 5 1 1 35062
0 35064 7 1 2 77067 103818
0 35065 5 1 1 35064
0 35066 7 1 2 80530 98521
0 35067 5 1 1 35066
0 35068 7 1 2 35065 35067
0 35069 5 1 1 35068
0 35070 7 1 2 35069 103783
0 35071 5 1 1 35070
0 35072 7 1 2 35063 35071
0 35073 5 1 1 35072
0 35074 7 1 2 72420 35073
0 35075 5 1 1 35074
0 35076 7 2 2 69208 93262
0 35077 5 1 1 103836
0 35078 7 1 2 97867 102018
0 35079 5 1 1 35078
0 35080 7 1 2 35077 35079
0 35081 5 1 1 35080
0 35082 7 1 2 67203 35081
0 35083 5 1 1 35082
0 35084 7 1 2 35083 34931
0 35085 5 1 1 35084
0 35086 7 1 2 67351 91836
0 35087 7 1 2 35085 35086
0 35088 5 1 1 35087
0 35089 7 1 2 35075 35088
0 35090 5 1 1 35089
0 35091 7 1 2 68093 95411
0 35092 7 1 2 35090 35091
0 35093 5 1 1 35092
0 35094 7 1 2 35053 35093
0 35095 5 1 1 35094
0 35096 7 1 2 74551 35095
0 35097 5 1 1 35096
0 35098 7 1 2 35000 35097
0 35099 7 1 2 34965 35098
0 35100 5 1 1 35099
0 35101 7 1 2 76328 35100
0 35102 5 1 1 35101
0 35103 7 1 2 64429 79509
0 35104 5 1 1 35103
0 35105 7 1 2 64798 35104
0 35106 5 1 1 35105
0 35107 7 1 2 78805 79233
0 35108 5 2 1 35107
0 35109 7 1 2 35106 103838
0 35110 5 1 1 35109
0 35111 7 1 2 102050 35110
0 35112 5 1 1 35111
0 35113 7 1 2 35112 10360
0 35114 5 1 1 35113
0 35115 7 1 2 71103 35114
0 35116 5 1 1 35115
0 35117 7 1 2 85080 80021
0 35118 7 1 2 85523 35117
0 35119 7 1 2 93756 35118
0 35120 5 1 1 35119
0 35121 7 1 2 35116 35120
0 35122 5 1 1 35121
0 35123 7 1 2 103768 35122
0 35124 5 1 1 35123
0 35125 7 3 2 98696 92410
0 35126 7 1 2 92863 85835
0 35127 7 1 2 103840 35126
0 35128 5 1 1 35127
0 35129 7 1 2 34816 35128
0 35130 5 1 1 35129
0 35131 7 1 2 79850 77363
0 35132 7 1 2 35130 35131
0 35133 5 1 1 35132
0 35134 7 1 2 35124 35133
0 35135 5 1 1 35134
0 35136 7 1 2 73186 35135
0 35137 5 1 1 35136
0 35138 7 1 2 98197 93370
0 35139 5 1 1 35138
0 35140 7 4 2 97737 84941
0 35141 5 2 1 103843
0 35142 7 1 2 35139 103847
0 35143 5 1 1 35142
0 35144 7 1 2 70838 35143
0 35145 5 1 1 35144
0 35146 7 1 2 77258 75048
0 35147 5 1 1 35146
0 35148 7 1 2 98499 92968
0 35149 7 1 2 35147 35148
0 35150 5 1 1 35149
0 35151 7 1 2 35145 35150
0 35152 5 1 1 35151
0 35153 7 1 2 69903 35152
0 35154 5 1 1 35153
0 35155 7 2 2 71104 86272
0 35156 5 1 1 103849
0 35157 7 1 2 98500 81469
0 35158 7 1 2 103850 35157
0 35159 5 1 1 35158
0 35160 7 1 2 35154 35159
0 35161 5 1 1 35160
0 35162 7 1 2 69209 35161
0 35163 5 1 1 35162
0 35164 7 3 2 85454 96753
0 35165 5 1 1 103851
0 35166 7 4 2 71105 73922
0 35167 7 1 2 81137 103854
0 35168 5 1 1 35167
0 35169 7 1 2 64799 35156
0 35170 5 1 1 35169
0 35171 7 1 2 66029 75049
0 35172 5 2 1 35171
0 35173 7 1 2 69538 103858
0 35174 7 1 2 35170 35173
0 35175 5 1 1 35174
0 35176 7 1 2 35168 35175
0 35177 5 1 1 35176
0 35178 7 1 2 103852 35177
0 35179 5 1 1 35178
0 35180 7 1 2 35163 35179
0 35181 5 1 1 35180
0 35182 7 1 2 75980 35181
0 35183 5 1 1 35182
0 35184 7 3 2 99752 78482
0 35185 5 1 1 103860
0 35186 7 1 2 75581 92001
0 35187 7 1 2 103861 35186
0 35188 5 1 1 35187
0 35189 7 1 2 35183 35188
0 35190 5 1 1 35189
0 35191 7 1 2 76855 35190
0 35192 5 1 1 35191
0 35193 7 1 2 35137 35192
0 35194 5 1 1 35193
0 35195 7 1 2 67204 35194
0 35196 5 1 1 35195
0 35197 7 1 2 77464 102533
0 35198 5 1 1 35197
0 35199 7 4 2 66030 98761
0 35200 7 1 2 95524 103863
0 35201 5 1 1 35200
0 35202 7 1 2 35198 35201
0 35203 5 1 1 35202
0 35204 7 1 2 79851 35203
0 35205 5 1 1 35204
0 35206 7 1 2 99154 96095
0 35207 5 1 1 35206
0 35208 7 1 2 35205 35207
0 35209 5 1 1 35208
0 35210 7 1 2 64148 35209
0 35211 5 1 1 35210
0 35212 7 1 2 96124 9574
0 35213 5 1 1 35212
0 35214 7 3 2 66345 98697
0 35215 7 1 2 79852 93377
0 35216 7 1 2 103867 35215
0 35217 7 1 2 35213 35216
0 35218 5 1 1 35217
0 35219 7 1 2 35211 35218
0 35220 5 1 1 35219
0 35221 7 2 2 100153 74222
0 35222 7 1 2 73524 103870
0 35223 7 1 2 35220 35222
0 35224 5 1 1 35223
0 35225 7 1 2 35196 35224
0 35226 5 1 1 35225
0 35227 7 1 2 78876 35226
0 35228 5 1 1 35227
0 35229 7 1 2 100559 97981
0 35230 5 1 1 35229
0 35231 7 1 2 73759 93517
0 35232 5 1 1 35231
0 35233 7 1 2 35230 35232
0 35234 5 1 1 35233
0 35235 7 1 2 75927 35234
0 35236 5 1 1 35235
0 35237 7 1 2 86349 82135
0 35238 5 1 1 35237
0 35239 7 1 2 85051 35238
0 35240 5 1 1 35239
0 35241 7 1 2 73971 35240
0 35242 5 1 1 35241
0 35243 7 1 2 91499 92988
0 35244 5 1 1 35243
0 35245 7 1 2 91462 35244
0 35246 7 1 2 35242 35245
0 35247 5 1 1 35246
0 35248 7 1 2 77364 35247
0 35249 5 1 1 35248
0 35250 7 1 2 35236 35249
0 35251 5 1 1 35250
0 35252 7 1 2 67352 35251
0 35253 5 1 1 35252
0 35254 7 1 2 90882 90237
0 35255 5 1 1 35254
0 35256 7 1 2 92002 91469
0 35257 5 1 1 35256
0 35258 7 1 2 35255 35257
0 35259 5 1 1 35258
0 35260 7 1 2 73525 98235
0 35261 7 1 2 35259 35260
0 35262 5 1 1 35261
0 35263 7 1 2 35253 35262
0 35264 5 1 1 35263
0 35265 7 1 2 72258 35264
0 35266 5 1 1 35265
0 35267 7 2 2 100577 92523
0 35268 5 1 1 103872
0 35269 7 1 2 98112 94332
0 35270 7 1 2 103873 35269
0 35271 5 1 1 35270
0 35272 7 1 2 35266 35271
0 35273 5 1 1 35272
0 35274 7 1 2 74399 35273
0 35275 5 1 1 35274
0 35276 7 2 2 65150 77068
0 35277 7 3 2 69210 84457
0 35278 7 1 2 103876 103309
0 35279 7 1 2 103874 35278
0 35280 7 1 2 98120 35279
0 35281 5 1 1 35280
0 35282 7 1 2 35275 35281
0 35283 5 1 1 35282
0 35284 7 1 2 76905 35283
0 35285 5 1 1 35284
0 35286 7 1 2 17918 101931
0 35287 5 2 1 35286
0 35288 7 1 2 77365 103879
0 35289 5 1 1 35288
0 35290 7 1 2 76875 98359
0 35291 5 1 1 35290
0 35292 7 1 2 35289 35291
0 35293 5 1 1 35292
0 35294 7 5 2 66879 72259
0 35295 7 9 2 75823 103881
0 35296 7 1 2 35293 103886
0 35297 5 1 1 35296
0 35298 7 2 2 67205 99084
0 35299 7 1 2 103895 99286
0 35300 5 1 1 35299
0 35301 7 1 2 35297 35300
0 35302 5 1 1 35301
0 35303 7 1 2 75284 35302
0 35304 5 1 1 35303
0 35305 7 5 2 67003 67206
0 35306 7 2 2 97438 103897
0 35307 7 1 2 71953 92164
0 35308 7 1 2 103902 35307
0 35309 7 1 2 102083 35308
0 35310 5 1 1 35309
0 35311 7 1 2 35304 35310
0 35312 5 1 1 35311
0 35313 7 1 2 73526 35312
0 35314 5 1 1 35313
0 35315 7 1 2 65151 84206
0 35316 5 1 1 35315
0 35317 7 1 2 1005 35316
0 35318 5 1 1 35317
0 35319 7 7 2 71106 67353
0 35320 7 1 2 103144 103904
0 35321 7 1 2 92212 35320
0 35322 7 1 2 35318 35321
0 35323 5 1 1 35322
0 35324 7 1 2 35314 35323
0 35325 5 1 1 35324
0 35326 7 1 2 64800 35325
0 35327 5 1 1 35326
0 35328 7 2 2 77840 103293
0 35329 7 1 2 102067 77814
0 35330 5 1 1 35329
0 35331 7 1 2 77600 103726
0 35332 5 1 1 35331
0 35333 7 1 2 35330 35332
0 35334 5 1 1 35333
0 35335 7 1 2 69539 35334
0 35336 5 1 1 35335
0 35337 7 1 2 83138 78496
0 35338 7 1 2 4940 1229
0 35339 7 1 2 35337 35338
0 35340 7 1 2 95894 35339
0 35341 5 1 1 35340
0 35342 7 1 2 35336 35341
0 35343 5 1 1 35342
0 35344 7 1 2 103911 35343
0 35345 5 1 1 35344
0 35346 7 1 2 35327 35345
0 35347 5 1 1 35346
0 35348 7 1 2 85524 35347
0 35349 5 1 1 35348
0 35350 7 1 2 76598 84242
0 35351 5 1 1 35350
0 35352 7 1 2 11984 35351
0 35353 5 1 1 35352
0 35354 7 1 2 81529 35353
0 35355 5 1 1 35354
0 35356 7 1 2 95134 102068
0 35357 5 1 1 35356
0 35358 7 1 2 35355 35357
0 35359 5 1 1 35358
0 35360 7 2 2 96398 103903
0 35361 7 1 2 98342 103913
0 35362 7 1 2 35359 35361
0 35363 5 1 1 35362
0 35364 7 1 2 35349 35363
0 35365 7 1 2 35285 35364
0 35366 5 1 1 35365
0 35367 7 1 2 74035 35366
0 35368 5 1 1 35367
0 35369 7 3 2 71107 97407
0 35370 7 1 2 78295 103831
0 35371 7 1 2 103915 35370
0 35372 5 1 1 35371
0 35373 7 1 2 70640 93263
0 35374 7 2 2 91970 35373
0 35375 7 1 2 68869 84458
0 35376 7 1 2 103054 35375
0 35377 7 1 2 103918 35376
0 35378 5 1 1 35377
0 35379 7 1 2 35372 35378
0 35380 5 1 1 35379
0 35381 7 1 2 67689 35380
0 35382 5 1 1 35381
0 35383 7 1 2 78991 103339
0 35384 7 1 2 84271 35383
0 35385 7 1 2 101845 103571
0 35386 7 1 2 35384 35385
0 35387 5 1 1 35386
0 35388 7 1 2 35382 35387
0 35389 5 1 1 35388
0 35390 7 1 2 68094 35389
0 35391 5 1 1 35390
0 35392 7 1 2 95529 103871
0 35393 5 1 1 35392
0 35394 7 1 2 77674 99092
0 35395 7 1 2 103791 35394
0 35396 5 1 1 35395
0 35397 7 1 2 35393 35396
0 35398 5 1 1 35397
0 35399 7 1 2 95412 35398
0 35400 5 1 1 35399
0 35401 7 1 2 35391 35400
0 35402 5 1 1 35401
0 35403 7 1 2 64149 35402
0 35404 5 1 1 35403
0 35405 7 2 2 79662 103784
0 35406 7 1 2 68095 100890
0 35407 5 1 1 35406
0 35408 7 1 2 99939 35407
0 35409 5 1 1 35408
0 35410 7 1 2 74066 35409
0 35411 5 1 1 35410
0 35412 7 1 2 88725 75657
0 35413 5 1 1 35412
0 35414 7 1 2 98710 35413
0 35415 5 1 1 35414
0 35416 7 1 2 35411 35415
0 35417 5 1 1 35416
0 35418 7 1 2 67690 35417
0 35419 5 1 1 35418
0 35420 7 1 2 75928 92583
0 35421 7 1 2 101956 35420
0 35422 5 1 1 35421
0 35423 7 1 2 35419 35422
0 35424 5 1 1 35423
0 35425 7 1 2 103920 35424
0 35426 5 1 1 35425
0 35427 7 1 2 35404 35426
0 35428 5 1 1 35427
0 35429 7 1 2 67354 35428
0 35430 5 1 1 35429
0 35431 7 3 2 70839 72260
0 35432 7 1 2 69211 103922
0 35433 5 1 1 35432
0 35434 7 9 2 65829 67207
0 35435 7 10 2 64150 103925
0 35436 5 2 1 103934
0 35437 7 1 2 35433 103944
0 35438 5 19 1 35437
0 35439 7 1 2 77366 103946
0 35440 5 1 1 35439
0 35441 7 1 2 72261 101072
0 35442 5 1 1 35441
0 35443 7 1 2 35440 35442
0 35444 5 1 1 35443
0 35445 7 2 2 73760 35444
0 35446 7 1 2 97310 92075
0 35447 7 1 2 103965 35446
0 35448 5 1 1 35447
0 35449 7 2 2 71436 76856
0 35450 7 1 2 71108 82448
0 35451 7 1 2 84294 101443
0 35452 7 1 2 35450 35451
0 35453 7 1 2 103967 35452
0 35454 5 1 1 35453
0 35455 7 1 2 35448 35454
0 35456 5 1 1 35455
0 35457 7 1 2 97219 79451
0 35458 7 1 2 35456 35457
0 35459 5 1 1 35458
0 35460 7 1 2 35430 35459
0 35461 5 1 1 35460
0 35462 7 1 2 74677 35461
0 35463 5 1 1 35462
0 35464 7 1 2 95351 103832
0 35465 5 1 1 35464
0 35466 7 6 2 72262 68096
0 35467 7 1 2 72165 79107
0 35468 7 1 2 103969 35467
0 35469 7 1 2 103919 35468
0 35470 5 1 1 35469
0 35471 7 1 2 35465 35470
0 35472 5 1 1 35471
0 35473 7 1 2 64151 35472
0 35474 5 1 1 35473
0 35475 7 2 2 75929 77069
0 35476 5 2 1 103975
0 35477 7 1 2 9987 103977
0 35478 5 1 1 35477
0 35479 7 1 2 103921 35478
0 35480 5 1 1 35479
0 35481 7 1 2 35474 35480
0 35482 5 1 1 35481
0 35483 7 1 2 67355 35482
0 35484 5 1 1 35483
0 35485 7 3 2 76857 98901
0 35486 7 1 2 100423 103979
0 35487 7 1 2 95599 35486
0 35488 5 1 1 35487
0 35489 7 1 2 35484 35488
0 35490 5 1 1 35489
0 35491 7 1 2 72704 35490
0 35492 5 1 1 35491
0 35493 7 1 2 78436 84474
0 35494 7 1 2 102466 35493
0 35495 7 1 2 98031 94567
0 35496 7 1 2 79353 35495
0 35497 7 1 2 35494 35496
0 35498 5 1 1 35497
0 35499 7 1 2 35492 35498
0 35500 5 1 1 35499
0 35501 7 1 2 102903 35500
0 35502 5 1 1 35501
0 35503 7 1 2 100424 93708
0 35504 7 1 2 103548 35503
0 35505 7 2 2 83188 87867
0 35506 7 2 2 70840 76940
0 35507 7 1 2 103982 103984
0 35508 7 1 2 97435 35507
0 35509 7 1 2 35504 35508
0 35510 5 1 1 35509
0 35511 7 1 2 35502 35510
0 35512 7 1 2 35463 35511
0 35513 7 1 2 35368 35512
0 35514 7 1 2 35228 35513
0 35515 7 1 2 68438 101383
0 35516 5 1 1 35515
0 35517 7 1 2 77259 35516
0 35518 5 1 1 35517
0 35519 7 1 2 103822 35518
0 35520 5 1 1 35519
0 35521 7 1 2 103011 79677
0 35522 7 1 2 98637 35521
0 35523 5 1 1 35522
0 35524 7 1 2 35520 35523
0 35525 5 1 1 35524
0 35526 7 1 2 69212 35525
0 35527 5 1 1 35526
0 35528 7 1 2 92383 103855
0 35529 5 1 1 35528
0 35530 7 1 2 10321 35529
0 35531 5 2 1 35530
0 35532 7 1 2 65152 103986
0 35533 5 1 1 35532
0 35534 7 1 2 73972 97880
0 35535 5 1 1 35534
0 35536 7 1 2 35533 35535
0 35537 5 1 1 35536
0 35538 7 1 2 35537 103087
0 35539 5 1 1 35538
0 35540 7 1 2 35527 35539
0 35541 5 1 1 35540
0 35542 7 1 2 63806 35541
0 35543 5 1 1 35542
0 35544 7 1 2 73973 98744
0 35545 5 1 1 35544
0 35546 7 1 2 64152 103987
0 35547 5 1 1 35546
0 35548 7 1 2 98736 35547
0 35549 5 1 1 35548
0 35550 7 1 2 65153 35549
0 35551 5 1 1 35550
0 35552 7 1 2 35545 35551
0 35553 5 1 1 35552
0 35554 7 1 2 74001 102574
0 35555 7 1 2 35553 35554
0 35556 5 1 1 35555
0 35557 7 1 2 35543 35556
0 35558 5 1 1 35557
0 35559 7 1 2 72421 35558
0 35560 5 1 1 35559
0 35561 7 1 2 101073 91742
0 35562 5 1 1 35561
0 35563 7 1 2 100510 35562
0 35564 5 1 1 35563
0 35565 7 4 2 67356 102547
0 35566 7 1 2 79641 103988
0 35567 7 1 2 35564 35566
0 35568 5 1 1 35567
0 35569 7 1 2 35560 35568
0 35570 5 1 1 35569
0 35571 7 1 2 66880 35570
0 35572 5 1 1 35571
0 35573 7 2 2 67208 78992
0 35574 7 1 2 103992 92127
0 35575 7 1 2 103404 35574
0 35576 7 1 2 103606 35575
0 35577 5 1 1 35576
0 35578 7 1 2 35572 35577
0 35579 5 1 1 35578
0 35580 7 1 2 72062 35579
0 35581 5 1 1 35580
0 35582 7 2 2 72263 95604
0 35583 7 2 2 64801 102746
0 35584 7 1 2 103996 95606
0 35585 7 1 2 103994 35584
0 35586 5 1 1 35585
0 35587 7 4 2 99479 77465
0 35588 5 1 1 103998
0 35589 7 2 2 84056 77907
0 35590 7 1 2 103792 104002
0 35591 7 1 2 103999 35590
0 35592 5 1 1 35591
0 35593 7 1 2 35586 35592
0 35594 5 1 1 35593
0 35595 7 1 2 75411 35594
0 35596 5 1 1 35595
0 35597 7 2 2 73527 103069
0 35598 7 1 2 99631 97640
0 35599 7 1 2 104004 35598
0 35600 5 1 1 35599
0 35601 7 1 2 87438 103989
0 35602 7 1 2 103856 35601
0 35603 5 1 1 35602
0 35604 7 1 2 35600 35603
0 35605 5 1 1 35604
0 35606 7 1 2 68870 35605
0 35607 5 1 1 35606
0 35608 7 1 2 86505 98795
0 35609 7 1 2 98201 35608
0 35610 7 1 2 102808 35609
0 35611 5 1 1 35610
0 35612 7 1 2 35607 35611
0 35613 5 1 1 35612
0 35614 7 1 2 85525 35613
0 35615 5 1 1 35614
0 35616 7 2 2 99632 78139
0 35617 7 1 2 78993 104005
0 35618 7 1 2 104006 35617
0 35619 5 1 1 35618
0 35620 7 1 2 35615 35619
0 35621 5 1 1 35620
0 35622 7 1 2 69904 35621
0 35623 5 1 1 35622
0 35624 7 1 2 75285 97738
0 35625 7 1 2 77730 35624
0 35626 7 1 2 103995 35625
0 35627 5 1 1 35626
0 35628 7 1 2 35623 35627
0 35629 5 1 1 35628
0 35630 7 1 2 75752 35629
0 35631 5 1 1 35630
0 35632 7 1 2 35596 35631
0 35633 7 1 2 35581 35632
0 35634 5 1 1 35633
0 35635 7 1 2 93007 35634
0 35636 5 1 1 35635
0 35637 7 1 2 64802 103428
0 35638 5 2 1 35637
0 35639 7 1 2 73528 87550
0 35640 5 1 1 35639
0 35641 7 1 2 104008 35640
0 35642 5 1 1 35641
0 35643 7 1 2 75629 95292
0 35644 7 1 2 35642 35643
0 35645 5 1 1 35644
0 35646 7 1 2 79302 82179
0 35647 5 2 1 35646
0 35648 7 1 2 86350 85016
0 35649 7 1 2 104010 35648
0 35650 5 1 1 35649
0 35651 7 1 2 35645 35650
0 35652 5 1 1 35651
0 35653 7 1 2 85979 35652
0 35654 5 1 1 35653
0 35655 7 3 2 71674 81417
0 35656 5 1 1 104012
0 35657 7 1 2 99848 104013
0 35658 5 2 1 35657
0 35659 7 2 2 64803 93008
0 35660 7 1 2 78662 104017
0 35661 5 1 1 35660
0 35662 7 1 2 104015 35661
0 35663 5 1 1 35662
0 35664 7 2 2 65154 85986
0 35665 7 1 2 35663 104019
0 35666 5 1 1 35665
0 35667 7 1 2 35654 35666
0 35668 5 1 1 35667
0 35669 7 1 2 85526 35668
0 35670 5 1 1 35669
0 35671 7 1 2 100259 82550
0 35672 7 1 2 104020 35671
0 35673 5 1 1 35672
0 35674 7 1 2 35670 35673
0 35675 5 1 1 35674
0 35676 7 1 2 72422 35675
0 35677 5 1 1 35676
0 35678 7 1 2 95464 91500
0 35679 5 1 1 35678
0 35680 7 1 2 74742 103187
0 35681 5 1 1 35680
0 35682 7 1 2 35679 35681
0 35683 5 1 1 35682
0 35684 7 1 2 64804 35683
0 35685 5 1 1 35684
0 35686 7 1 2 104016 35685
0 35687 5 1 1 35686
0 35688 7 1 2 65155 35687
0 35689 5 1 1 35688
0 35690 7 2 2 82229 101393
0 35691 7 1 2 73761 104021
0 35692 5 1 1 35691
0 35693 7 1 2 35689 35692
0 35694 5 1 1 35693
0 35695 7 1 2 85987 35694
0 35696 5 1 1 35695
0 35697 7 2 2 76228 79642
0 35698 7 1 2 97303 104023
0 35699 7 1 2 93761 35698
0 35700 5 1 1 35699
0 35701 7 1 2 35696 35700
0 35702 5 1 1 35701
0 35703 7 1 2 97696 35702
0 35704 5 1 1 35703
0 35705 7 1 2 35677 35704
0 35706 5 1 1 35705
0 35707 7 1 2 102575 35706
0 35708 5 1 1 35707
0 35709 7 1 2 90770 9909
0 35710 5 1 1 35709
0 35711 7 1 2 75286 35710
0 35712 5 1 1 35711
0 35713 7 1 2 87234 93009
0 35714 5 1 1 35713
0 35715 7 1 2 35712 35714
0 35716 5 1 1 35715
0 35717 7 2 2 74354 95621
0 35718 7 1 2 94073 104025
0 35719 7 1 2 103990 35718
0 35720 7 1 2 35716 35719
0 35721 5 1 1 35720
0 35722 7 1 2 35708 35721
0 35723 5 1 1 35722
0 35724 7 1 2 66881 35723
0 35725 5 1 1 35724
0 35726 7 1 2 103991 102836
0 35727 7 1 2 103347 35726
0 35728 7 1 2 97267 83203
0 35729 7 1 2 35727 35728
0 35730 5 1 1 35729
0 35731 7 1 2 35725 35730
0 35732 5 1 1 35731
0 35733 7 1 2 77260 35732
0 35734 5 1 1 35733
0 35735 7 2 2 102576 74036
0 35736 7 2 2 97902 78575
0 35737 5 1 1 104029
0 35738 7 1 2 64805 98433
0 35739 5 1 1 35738
0 35740 7 1 2 35737 35739
0 35741 5 1 1 35740
0 35742 7 1 2 64153 35741
0 35743 5 1 1 35742
0 35744 7 1 2 30016 35743
0 35745 5 1 1 35744
0 35746 7 1 2 104027 35745
0 35747 5 1 1 35746
0 35748 7 1 2 74355 98174
0 35749 7 1 2 103823 35748
0 35750 5 1 1 35749
0 35751 7 1 2 35747 35750
0 35752 5 1 1 35751
0 35753 7 1 2 72063 35752
0 35754 5 1 1 35753
0 35755 7 1 2 67357 74927
0 35756 7 1 2 93767 35755
0 35757 7 1 2 103779 35756
0 35758 5 1 1 35757
0 35759 7 1 2 35754 35758
0 35760 5 1 1 35759
0 35761 7 1 2 74678 35760
0 35762 5 1 1 35761
0 35763 7 1 2 79853 102577
0 35764 7 1 2 85988 35763
0 35765 7 1 2 99007 35764
0 35766 5 1 1 35765
0 35767 7 1 2 35762 35766
0 35768 5 1 1 35767
0 35769 7 1 2 77367 35768
0 35770 5 1 1 35769
0 35771 7 1 2 95597 102558
0 35772 5 1 1 35771
0 35773 7 1 2 73974 74400
0 35774 7 1 2 104028 35773
0 35775 5 1 1 35774
0 35776 7 1 2 35772 35775
0 35777 5 1 1 35776
0 35778 7 1 2 100570 80022
0 35779 7 1 2 35777 35778
0 35780 5 1 1 35779
0 35781 7 1 2 35770 35780
0 35782 5 1 1 35781
0 35783 7 1 2 67691 35782
0 35784 5 1 1 35783
0 35785 7 2 2 78318 94642
0 35786 7 2 2 102128 91487
0 35787 7 1 2 104033 82822
0 35788 7 1 2 104031 35787
0 35789 7 1 2 103966 35788
0 35790 5 1 1 35789
0 35791 7 1 2 35784 35790
0 35792 5 1 1 35791
0 35793 7 1 2 66882 35792
0 35794 5 1 1 35793
0 35795 7 2 2 75753 98762
0 35796 7 2 2 101444 84565
0 35797 7 1 2 100513 104037
0 35798 5 1 1 35797
0 35799 7 2 2 80318 102391
0 35800 7 1 2 82792 86506
0 35801 7 1 2 102973 35800
0 35802 7 1 2 104039 35801
0 35803 5 1 1 35802
0 35804 7 1 2 35798 35803
0 35805 5 1 1 35804
0 35806 7 1 2 64806 35805
0 35807 5 1 1 35806
0 35808 7 2 2 94838 92823
0 35809 7 1 2 77368 104041
0 35810 7 1 2 104038 35809
0 35811 5 1 1 35810
0 35812 7 1 2 35807 35811
0 35813 5 1 1 35812
0 35814 7 1 2 104035 35813
0 35815 5 1 1 35814
0 35816 7 1 2 35794 35815
0 35817 5 1 1 35816
0 35818 7 1 2 75017 35817
0 35819 5 1 1 35818
0 35820 7 1 2 35734 35819
0 35821 7 1 2 35636 35820
0 35822 7 1 2 35514 35821
0 35823 5 1 1 35822
0 35824 7 1 2 80713 35823
0 35825 5 1 1 35824
0 35826 7 1 2 35102 35825
0 35827 7 1 2 34871 35826
0 35828 7 1 2 70210 79055
0 35829 7 1 2 94137 35828
0 35830 5 1 1 35829
0 35831 7 1 2 86576 35830
0 35832 5 1 1 35831
0 35833 7 1 2 63807 35832
0 35834 5 1 1 35833
0 35835 7 1 2 90732 94403
0 35836 5 1 1 35835
0 35837 7 1 2 35834 35836
0 35838 5 1 1 35837
0 35839 7 1 2 73529 35838
0 35840 5 1 1 35839
0 35841 7 1 2 74823 85980
0 35842 5 1 1 35841
0 35843 7 1 2 35840 35842
0 35844 5 1 1 35843
0 35845 7 1 2 66031 35844
0 35846 5 1 1 35845
0 35847 7 1 2 83373 77951
0 35848 5 2 1 35847
0 35849 7 1 2 98641 104043
0 35850 5 1 1 35849
0 35851 7 1 2 86569 79643
0 35852 7 1 2 35850 35851
0 35853 5 1 1 35852
0 35854 7 1 2 35846 35853
0 35855 5 1 1 35854
0 35856 7 1 2 84842 35855
0 35857 5 1 1 35856
0 35858 7 1 2 93821 100022
0 35859 5 1 1 35858
0 35860 7 1 2 69905 87476
0 35861 5 1 1 35860
0 35862 7 1 2 35861 103156
0 35863 5 1 1 35862
0 35864 7 1 2 86351 35863
0 35865 5 1 1 35864
0 35866 7 2 2 35859 35865
0 35867 5 1 1 104045
0 35868 7 1 2 64430 101720
0 35869 5 2 1 35868
0 35870 7 1 2 99991 87158
0 35871 5 1 1 35870
0 35872 7 1 2 104047 35871
0 35873 5 1 1 35872
0 35874 7 1 2 66032 35873
0 35875 5 1 1 35874
0 35876 7 1 2 104046 35875
0 35877 5 1 1 35876
0 35878 7 1 2 85989 35877
0 35879 5 1 1 35878
0 35880 7 1 2 81893 100044
0 35881 5 1 1 35880
0 35882 7 1 2 69906 87287
0 35883 5 3 1 35882
0 35884 7 2 2 68439 104049
0 35885 5 3 1 104052
0 35886 7 1 2 73530 101645
0 35887 5 1 1 35886
0 35888 7 1 2 104054 35887
0 35889 7 1 2 35881 35888
0 35890 5 1 1 35889
0 35891 7 1 2 85981 35890
0 35892 5 1 1 35891
0 35893 7 1 2 35879 35892
0 35894 5 1 1 35893
0 35895 7 1 2 77261 35894
0 35896 5 1 1 35895
0 35897 7 1 2 35857 35896
0 35898 5 1 1 35897
0 35899 7 1 2 64154 35898
0 35900 5 1 1 35899
0 35901 7 1 2 64431 89431
0 35902 7 1 2 76135 35901
0 35903 7 1 2 100665 103499
0 35904 7 1 2 35902 35903
0 35905 5 1 1 35904
0 35906 7 1 2 35900 35905
0 35907 5 1 1 35906
0 35908 7 1 2 65830 35907
0 35909 5 1 1 35908
0 35910 7 8 2 73531 84843
0 35911 7 4 2 65605 84575
0 35912 7 1 2 64807 104065
0 35913 7 2 2 104057 35912
0 35914 7 1 2 86570 80319
0 35915 7 1 2 93390 35914
0 35916 7 1 2 104069 35915
0 35917 5 1 1 35916
0 35918 7 1 2 35909 35917
0 35919 5 1 1 35918
0 35920 7 1 2 99327 35919
0 35921 5 1 1 35920
0 35922 7 1 2 64432 35867
0 35923 5 1 1 35922
0 35924 7 1 2 24066 95884
0 35925 5 1 1 35924
0 35926 7 1 2 73532 35925
0 35927 5 2 1 35926
0 35928 7 1 2 69540 86286
0 35929 7 1 2 104071 35928
0 35930 5 1 1 35929
0 35931 7 1 2 69907 35930
0 35932 5 1 1 35931
0 35933 7 1 2 64808 93834
0 35934 5 1 1 35933
0 35935 7 1 2 64433 94269
0 35936 5 1 1 35935
0 35937 7 1 2 35934 35936
0 35938 5 1 1 35937
0 35939 7 1 2 68440 35938
0 35940 5 1 1 35939
0 35941 7 1 2 71675 94207
0 35942 5 1 1 35941
0 35943 7 1 2 82011 99934
0 35944 5 3 1 35943
0 35945 7 1 2 35942 104073
0 35946 7 1 2 35940 35945
0 35947 7 1 2 35932 35946
0 35948 5 1 1 35947
0 35949 7 1 2 66033 35948
0 35950 5 1 1 35949
0 35951 7 1 2 35923 35950
0 35952 5 1 1 35951
0 35953 7 1 2 85439 35952
0 35954 5 1 1 35953
0 35955 7 1 2 104072 102313
0 35956 5 1 1 35955
0 35957 7 1 2 64809 93840
0 35958 5 1 1 35957
0 35959 7 1 2 77262 35958
0 35960 7 1 2 35956 35959
0 35961 5 1 1 35960
0 35962 7 1 2 81109 100588
0 35963 5 1 1 35962
0 35964 7 1 2 100688 101537
0 35965 5 1 1 35964
0 35966 7 1 2 77369 35965
0 35967 5 1 1 35966
0 35968 7 1 2 35963 35967
0 35969 7 1 2 35961 35968
0 35970 5 1 1 35969
0 35971 7 1 2 70841 35970
0 35972 5 1 1 35971
0 35973 7 1 2 86059 92569
0 35974 7 1 2 100904 35973
0 35975 5 1 1 35974
0 35976 7 1 2 25900 35975
0 35977 7 1 2 35972 35976
0 35978 5 1 1 35977
0 35979 7 1 2 64155 35978
0 35980 5 1 1 35979
0 35981 7 1 2 35954 35980
0 35982 5 1 1 35981
0 35983 7 1 2 35982 86203
0 35984 5 1 1 35983
0 35985 7 2 2 88399 103383
0 35986 5 1 1 104076
0 35987 7 1 2 70842 104077
0 35988 5 1 1 35987
0 35989 7 2 2 78994 84449
0 35990 7 1 2 90701 104078
0 35991 7 1 2 97881 35990
0 35992 5 1 1 35991
0 35993 7 1 2 35988 35992
0 35994 5 1 1 35993
0 35995 7 1 2 64156 35994
0 35996 5 1 1 35995
0 35997 7 2 2 71842 100244
0 35998 7 1 2 82389 79108
0 35999 7 1 2 91195 35998
0 36000 7 1 2 104080 35999
0 36001 5 1 1 36000
0 36002 7 1 2 35986 36001
0 36003 5 1 1 36002
0 36004 7 1 2 85440 36003
0 36005 5 1 1 36004
0 36006 7 1 2 35996 36005
0 36007 5 1 1 36006
0 36008 7 1 2 70211 36007
0 36009 5 1 1 36008
0 36010 7 1 2 88400 104003
0 36011 7 1 2 103450 36010
0 36012 5 1 1 36011
0 36013 7 1 2 36009 36012
0 36014 5 1 1 36013
0 36015 7 1 2 73533 36014
0 36016 5 1 1 36015
0 36017 7 2 2 78995 91196
0 36018 7 1 2 101497 104082
0 36019 5 1 1 36018
0 36020 7 2 2 79663 103530
0 36021 5 1 1 104084
0 36022 7 1 2 36019 36021
0 36023 5 1 1 36022
0 36024 7 1 2 85527 36023
0 36025 5 1 1 36024
0 36026 7 2 2 90718 94233
0 36027 7 1 2 84502 91197
0 36028 7 1 2 104086 36027
0 36029 5 1 1 36028
0 36030 7 1 2 36025 36029
0 36031 5 1 1 36030
0 36032 7 1 2 80628 36031
0 36033 5 1 1 36032
0 36034 7 1 2 97670 104085
0 36035 5 1 1 36034
0 36036 7 1 2 36033 36035
0 36037 5 1 1 36036
0 36038 7 1 2 89216 36037
0 36039 5 1 1 36038
0 36040 7 1 2 79664 103451
0 36041 7 1 2 27082 36040
0 36042 5 1 1 36041
0 36043 7 1 2 76658 79146
0 36044 7 1 2 95203 36043
0 36045 7 1 2 98745 36044
0 36046 5 1 1 36045
0 36047 7 1 2 36042 36046
0 36048 5 1 1 36047
0 36049 7 1 2 68441 36048
0 36050 5 1 1 36049
0 36051 7 1 2 86060 103384
0 36052 7 1 2 103077 36051
0 36053 5 1 1 36052
0 36054 7 1 2 36050 36053
0 36055 7 1 2 36039 36054
0 36056 7 1 2 36016 36055
0 36057 5 1 1 36056
0 36058 7 1 2 67004 36057
0 36059 5 1 1 36058
0 36060 7 1 2 35984 36059
0 36061 5 1 1 36060
0 36062 7 1 2 72423 36061
0 36063 5 1 1 36062
0 36064 7 1 2 95198 86754
0 36065 5 1 1 36064
0 36066 7 1 2 69908 36065
0 36067 5 1 1 36066
0 36068 7 1 2 71843 80903
0 36069 7 1 2 78041 36068
0 36070 5 2 1 36069
0 36071 7 1 2 36067 104088
0 36072 5 2 1 36071
0 36073 7 2 2 95607 104090
0 36074 7 1 2 104092 96346
0 36075 5 1 1 36074
0 36076 7 1 2 85631 86204
0 36077 5 1 1 36076
0 36078 7 1 2 104091 86166
0 36079 5 1 1 36078
0 36080 7 1 2 36077 36079
0 36081 5 1 1 36080
0 36082 7 1 2 98522 36081
0 36083 5 1 1 36082
0 36084 7 1 2 36075 36083
0 36085 5 1 1 36084
0 36086 7 1 2 64157 36085
0 36087 5 1 1 36086
0 36088 7 1 2 85441 92479
0 36089 7 1 2 104093 36088
0 36090 5 1 1 36089
0 36091 7 1 2 36087 36090
0 36092 5 1 1 36091
0 36093 7 1 2 72424 36092
0 36094 5 1 1 36093
0 36095 7 1 2 99713 102948
0 36096 7 1 2 101553 36095
0 36097 7 1 2 75793 86099
0 36098 7 1 2 36096 36097
0 36099 5 1 1 36098
0 36100 7 1 2 36094 36099
0 36101 5 1 1 36100
0 36102 7 1 2 75412 36101
0 36103 5 1 1 36102
0 36104 7 1 2 36063 36103
0 36105 7 1 2 35921 36104
0 36106 5 1 1 36105
0 36107 7 1 2 72705 36106
0 36108 5 1 1 36107
0 36109 7 1 2 98746 103810
0 36110 5 1 1 36109
0 36111 7 1 2 85372 85399
0 36112 5 1 1 36111
0 36113 7 1 2 36110 36112
0 36114 5 1 1 36113
0 36115 7 1 2 79854 36114
0 36116 5 1 1 36115
0 36117 7 1 2 104055 103221
0 36118 5 1 1 36117
0 36119 7 1 2 77466 36118
0 36120 5 1 1 36119
0 36121 7 2 2 69909 98306
0 36122 5 1 1 104094
0 36123 7 1 2 36120 36122
0 36124 5 1 1 36123
0 36125 7 1 2 64158 36124
0 36126 5 1 1 36125
0 36127 7 1 2 64810 99905
0 36128 5 3 1 36127
0 36129 7 1 2 69910 103417
0 36130 5 1 1 36129
0 36131 7 1 2 104096 36130
0 36132 5 1 1 36131
0 36133 7 1 2 70480 36132
0 36134 5 1 1 36133
0 36135 7 5 2 91449 73923
0 36136 5 1 1 104099
0 36137 7 1 2 84762 104100
0 36138 5 1 1 36137
0 36139 7 1 2 36134 36138
0 36140 5 1 1 36139
0 36141 7 1 2 77370 36140
0 36142 5 1 1 36141
0 36143 7 1 2 36126 36142
0 36144 5 1 1 36143
0 36145 7 1 2 65831 36144
0 36146 5 1 1 36145
0 36147 7 1 2 101554 104095
0 36148 5 1 1 36147
0 36149 7 1 2 36146 36148
0 36150 5 1 1 36149
0 36151 7 1 2 78877 36150
0 36152 5 1 1 36151
0 36153 7 1 2 36116 36152
0 36154 5 1 1 36153
0 36155 7 1 2 67005 36154
0 36156 5 1 1 36155
0 36157 7 1 2 76633 85575
0 36158 7 1 2 98747 36157
0 36159 5 1 1 36158
0 36160 7 2 2 74067 90664
0 36161 7 1 2 93607 87439
0 36162 7 1 2 104104 36161
0 36163 5 1 1 36162
0 36164 7 1 2 36159 36163
0 36165 5 1 1 36164
0 36166 7 1 2 68871 36165
0 36167 5 1 1 36166
0 36168 7 1 2 99728 74008
0 36169 7 1 2 104105 36168
0 36170 5 1 1 36169
0 36171 7 1 2 36167 36170
0 36172 5 1 1 36171
0 36173 7 1 2 94760 36172
0 36174 5 1 1 36173
0 36175 7 1 2 71109 93836
0 36176 5 1 1 36175
0 36177 7 1 2 77467 100840
0 36178 5 1 1 36177
0 36179 7 1 2 64811 36178
0 36180 7 1 2 36176 36179
0 36181 5 1 1 36180
0 36182 7 1 2 74679 98315
0 36183 5 1 1 36182
0 36184 7 1 2 69911 36183
0 36185 7 1 2 89033 36184
0 36186 5 1 1 36185
0 36187 7 1 2 74037 78528
0 36188 7 1 2 36186 36187
0 36189 7 1 2 36181 36188
0 36190 5 1 1 36189
0 36191 7 1 2 36174 36190
0 36192 7 1 2 36156 36191
0 36193 5 1 1 36192
0 36194 7 1 2 97048 36193
0 36195 5 1 1 36194
0 36196 7 1 2 36108 36195
0 36197 5 1 1 36196
0 36198 7 1 2 102578 36197
0 36199 5 1 1 36198
0 36200 7 1 2 68442 93788
0 36201 5 1 1 36200
0 36202 7 1 2 87353 36201
0 36203 5 1 1 36202
0 36204 7 1 2 69912 36203
0 36205 5 1 1 36204
0 36206 7 1 2 77113 88869
0 36207 5 1 1 36206
0 36208 7 1 2 36205 36207
0 36209 5 1 1 36208
0 36210 7 1 2 103618 36209
0 36211 5 1 1 36210
0 36212 7 1 2 69913 86965
0 36213 5 1 1 36212
0 36214 7 2 2 68681 100675
0 36215 5 1 1 104106
0 36216 7 1 2 36213 36215
0 36217 5 1 1 36216
0 36218 7 1 2 100529 36217
0 36219 5 1 1 36218
0 36220 7 1 2 36211 36219
0 36221 5 1 1 36220
0 36222 7 1 2 72706 36221
0 36223 5 1 1 36222
0 36224 7 1 2 67692 94360
0 36225 5 1 1 36224
0 36226 7 1 2 98299 36225
0 36227 5 1 1 36226
0 36228 7 1 2 103607 36227
0 36229 5 1 1 36228
0 36230 7 1 2 74173 97769
0 36231 7 1 2 103613 36230
0 36232 7 1 2 95161 36231
0 36233 5 1 1 36232
0 36234 7 1 2 36229 36233
0 36235 5 1 1 36234
0 36236 7 1 2 64812 36235
0 36237 5 1 1 36236
0 36238 7 1 2 36223 36237
0 36239 5 1 1 36238
0 36240 7 1 2 83884 36239
0 36241 5 1 1 36240
0 36242 7 1 2 69541 101229
0 36243 5 1 1 36242
0 36244 7 1 2 88824 101440
0 36245 5 1 1 36244
0 36246 7 1 2 36243 36245
0 36247 5 1 1 36246
0 36248 7 1 2 72425 36247
0 36249 5 1 1 36248
0 36250 7 1 2 98229 36249
0 36251 5 1 1 36250
0 36252 7 1 2 70481 36251
0 36253 5 1 1 36252
0 36254 7 1 2 82842 77974
0 36255 7 1 2 100488 36254
0 36256 5 1 1 36255
0 36257 7 1 2 36253 36256
0 36258 5 1 1 36257
0 36259 7 1 2 69914 36258
0 36260 5 1 1 36259
0 36261 7 1 2 83776 83831
0 36262 5 1 1 36261
0 36263 7 1 2 100116 91729
0 36264 7 1 2 36262 36263
0 36265 5 1 1 36264
0 36266 7 1 2 36260 36265
0 36267 5 1 1 36266
0 36268 7 1 2 72707 36267
0 36269 5 1 1 36268
0 36270 7 1 2 64813 99002
0 36271 5 1 1 36270
0 36272 7 1 2 95068 86807
0 36273 5 1 1 36272
0 36274 7 1 2 36271 36273
0 36275 5 1 1 36274
0 36276 7 1 2 77468 36275
0 36277 5 1 1 36276
0 36278 7 1 2 69915 94159
0 36279 5 1 1 36278
0 36280 7 1 2 36277 36279
0 36281 5 1 1 36280
0 36282 7 1 2 70212 36281
0 36283 5 1 1 36282
0 36284 7 1 2 80328 94379
0 36285 5 1 1 36284
0 36286 7 1 2 36283 36285
0 36287 5 1 1 36286
0 36288 7 1 2 97049 36287
0 36289 5 1 1 36288
0 36290 7 1 2 36269 36289
0 36291 5 1 1 36290
0 36292 7 1 2 82449 36291
0 36293 5 1 1 36292
0 36294 7 2 2 98434 95282
0 36295 7 1 2 75510 89247
0 36296 5 1 1 36295
0 36297 7 1 2 81494 36296
0 36298 5 1 1 36297
0 36299 7 1 2 104108 36298
0 36300 5 1 1 36299
0 36301 7 1 2 71110 83645
0 36302 5 1 1 36301
0 36303 7 1 2 64434 36302
0 36304 5 1 1 36303
0 36305 7 1 2 86254 77975
0 36306 5 1 1 36305
0 36307 7 1 2 36304 36306
0 36308 5 1 1 36307
0 36309 7 1 2 101054 36308
0 36310 5 1 1 36309
0 36311 7 1 2 85528 92351
0 36312 7 1 2 82396 36311
0 36313 5 1 1 36312
0 36314 7 4 2 69542 85529
0 36315 7 1 2 78412 104110
0 36316 5 2 1 36315
0 36317 7 1 2 36313 104114
0 36318 7 1 2 36310 36317
0 36319 5 1 1 36318
0 36320 7 1 2 67358 36319
0 36321 5 1 1 36320
0 36322 7 1 2 36300 36321
0 36323 5 1 1 36322
0 36324 7 1 2 69916 36323
0 36325 5 1 1 36324
0 36326 7 2 2 64814 75511
0 36327 7 1 2 82218 104116
0 36328 5 1 1 36327
0 36329 7 3 2 75413 81470
0 36330 5 1 1 104118
0 36331 7 1 2 36328 36330
0 36332 5 1 1 36331
0 36333 7 1 2 99753 76621
0 36334 7 1 2 36332 36333
0 36335 5 1 1 36334
0 36336 7 1 2 36325 36335
0 36337 5 1 1 36336
0 36338 7 1 2 82985 36337
0 36339 5 1 1 36338
0 36340 7 1 2 92770 95582
0 36341 5 1 1 36340
0 36342 7 1 2 101380 104058
0 36343 5 1 1 36342
0 36344 7 1 2 36341 36343
0 36345 5 1 1 36344
0 36346 7 1 2 80853 36345
0 36347 5 1 1 36346
0 36348 7 1 2 89607 84697
0 36349 5 1 1 36348
0 36350 7 1 2 36347 36349
0 36351 5 1 1 36350
0 36352 7 1 2 67693 36351
0 36353 5 1 1 36352
0 36354 7 1 2 80899 92548
0 36355 5 1 1 36354
0 36356 7 1 2 36353 36355
0 36357 5 1 1 36356
0 36358 7 1 2 99405 36357
0 36359 5 1 1 36358
0 36360 7 2 2 77263 96754
0 36361 5 1 1 104121
0 36362 7 1 2 98402 36361
0 36363 5 10 1 36362
0 36364 7 1 2 79885 104123
0 36365 5 1 1 36364
0 36366 7 1 2 101256 98398
0 36367 5 1 1 36366
0 36368 7 1 2 36365 36367
0 36369 5 1 1 36368
0 36370 7 1 2 99604 36369
0 36371 5 1 1 36370
0 36372 7 2 2 98175 92266
0 36373 7 1 2 84276 104133
0 36374 5 1 1 36373
0 36375 7 1 2 36371 36374
0 36376 5 1 1 36375
0 36377 7 1 2 69213 36376
0 36378 5 1 1 36377
0 36379 7 2 2 85455 80834
0 36380 7 1 2 104134 104135
0 36381 5 1 1 36380
0 36382 7 1 2 36378 36381
0 36383 5 1 1 36382
0 36384 7 1 2 80418 36383
0 36385 5 1 1 36384
0 36386 7 1 2 88473 81398
0 36387 7 1 2 84698 36386
0 36388 7 1 2 99406 36387
0 36389 5 1 1 36388
0 36390 7 1 2 36385 36389
0 36391 5 1 1 36390
0 36392 7 1 2 65156 36391
0 36393 5 1 1 36392
0 36394 7 1 2 36359 36393
0 36395 7 1 2 36339 36394
0 36396 7 1 2 36293 36395
0 36397 5 1 1 36396
0 36398 7 1 2 83204 36397
0 36399 5 1 1 36398
0 36400 7 1 2 36241 36399
0 36401 5 1 1 36400
0 36402 7 1 2 71954 36401
0 36403 5 1 1 36402
0 36404 7 1 2 83028 97686
0 36405 5 1 1 36404
0 36406 7 1 2 78483 97833
0 36407 5 1 1 36406
0 36408 7 1 2 36405 36407
0 36409 5 1 1 36408
0 36410 7 1 2 72426 36409
0 36411 5 1 1 36410
0 36412 7 1 2 104122 97834
0 36413 5 1 1 36412
0 36414 7 1 2 69917 36413
0 36415 7 1 2 36411 36414
0 36416 5 1 1 36415
0 36417 7 1 2 75414 101141
0 36418 5 1 1 36417
0 36419 7 6 2 72427 90862
0 36420 7 1 2 68443 104137
0 36421 5 1 1 36420
0 36422 7 1 2 36418 36421
0 36423 5 1 1 36422
0 36424 7 1 2 80714 36423
0 36425 5 1 1 36424
0 36426 7 1 2 88765 101142
0 36427 5 1 1 36426
0 36428 7 1 2 80629 89707
0 36429 7 1 2 104124 36428
0 36430 5 1 1 36429
0 36431 7 1 2 64815 36430
0 36432 7 1 2 36427 36431
0 36433 7 1 2 36425 36432
0 36434 5 1 1 36433
0 36435 7 1 2 36416 36434
0 36436 5 1 1 36435
0 36437 7 2 2 77284 87360
0 36438 5 1 1 104143
0 36439 7 1 2 83079 94270
0 36440 5 1 1 36439
0 36441 7 1 2 68444 36440
0 36442 5 2 1 36441
0 36443 7 1 2 70482 91739
0 36444 7 1 2 83828 36443
0 36445 5 1 1 36444
0 36446 7 1 2 104145 36445
0 36447 5 2 1 36446
0 36448 7 1 2 65157 104147
0 36449 5 1 1 36448
0 36450 7 1 2 36438 36449
0 36451 5 1 1 36450
0 36452 7 1 2 104125 36451
0 36453 5 1 1 36452
0 36454 7 1 2 98258 86836
0 36455 5 1 1 36454
0 36456 7 1 2 82450 36455
0 36457 7 1 2 36453 36456
0 36458 7 1 2 36436 36457
0 36459 5 1 1 36458
0 36460 7 1 2 75415 78031
0 36461 5 2 1 36460
0 36462 7 1 2 77264 104149
0 36463 5 1 1 36462
0 36464 7 1 2 92969 36463
0 36465 5 1 1 36464
0 36466 7 1 2 78484 95800
0 36467 5 1 1 36466
0 36468 7 1 2 36465 36467
0 36469 5 1 1 36468
0 36470 7 1 2 80630 36469
0 36471 5 1 1 36470
0 36472 7 1 2 82603 91501
0 36473 7 1 2 84699 36472
0 36474 5 1 1 36473
0 36475 7 1 2 36471 36474
0 36476 5 1 1 36475
0 36477 7 1 2 67359 36476
0 36478 5 1 1 36477
0 36479 7 1 2 82500 36478
0 36480 5 1 1 36479
0 36481 7 1 2 74429 99284
0 36482 7 1 2 36480 36481
0 36483 7 1 2 36459 36482
0 36484 5 1 1 36483
0 36485 7 1 2 36403 36484
0 36486 5 1 1 36485
0 36487 7 1 2 102548 36486
0 36488 5 1 1 36487
0 36489 7 1 2 36199 36488
0 36490 5 1 1 36489
0 36491 7 1 2 76093 36490
0 36492 5 1 1 36491
0 36493 7 10 2 75754 102549
0 36494 7 2 2 64435 86850
0 36495 5 2 1 104161
0 36496 7 1 2 82986 104163
0 36497 5 1 1 36496
0 36498 7 2 2 80854 86173
0 36499 5 1 1 104165
0 36500 7 1 2 36497 36499
0 36501 5 1 1 36500
0 36502 7 1 2 72708 36501
0 36503 5 1 1 36502
0 36504 7 1 2 82136 102289
0 36505 5 1 1 36504
0 36506 7 1 2 36503 36505
0 36507 5 1 1 36506
0 36508 7 1 2 65454 36507
0 36509 5 1 1 36508
0 36510 7 1 2 69543 77102
0 36511 5 1 1 36510
0 36512 7 1 2 69918 99885
0 36513 5 1 1 36512
0 36514 7 1 2 36511 36513
0 36515 5 1 1 36514
0 36516 7 1 2 98658 36515
0 36517 5 1 1 36516
0 36518 7 1 2 92267 90457
0 36519 5 1 1 36518
0 36520 7 1 2 36517 36519
0 36521 7 1 2 36509 36520
0 36522 5 1 1 36521
0 36523 7 1 2 73534 36522
0 36524 5 1 1 36523
0 36525 7 1 2 65455 104044
0 36526 5 1 1 36525
0 36527 7 1 2 82933 36526
0 36528 5 1 1 36527
0 36529 7 1 2 69919 100592
0 36530 5 1 1 36529
0 36531 7 1 2 69544 36530
0 36532 7 1 2 36528 36531
0 36533 5 1 1 36532
0 36534 7 1 2 69920 4635
0 36535 5 1 1 36534
0 36536 7 1 2 64436 74880
0 36537 5 1 1 36536
0 36538 7 1 2 36535 36537
0 36539 5 1 1 36538
0 36540 7 1 2 99887 36539
0 36541 5 1 1 36540
0 36542 7 1 2 70483 3073
0 36543 7 1 2 36541 36542
0 36544 5 1 1 36543
0 36545 7 1 2 36533 36544
0 36546 5 1 1 36545
0 36547 7 1 2 72709 36546
0 36548 5 1 1 36547
0 36549 7 1 2 36524 36548
0 36550 5 1 1 36549
0 36551 7 1 2 71437 36550
0 36552 5 1 1 36551
0 36553 7 3 2 95248 77295
0 36554 7 1 2 70213 104167
0 36555 5 1 1 36554
0 36556 7 1 2 83588 36555
0 36557 5 1 1 36556
0 36558 7 1 2 83043 36557
0 36559 5 1 1 36558
0 36560 7 1 2 22356 102915
0 36561 5 1 1 36560
0 36562 7 1 2 86273 36561
0 36563 5 1 1 36562
0 36564 7 1 2 92913 75061
0 36565 5 1 1 36564
0 36566 7 1 2 22166 3703
0 36567 5 1 1 36566
0 36568 7 1 2 70484 36567
0 36569 5 1 1 36568
0 36570 7 1 2 36565 36569
0 36571 7 1 2 36563 36570
0 36572 7 1 2 36559 36571
0 36573 5 1 1 36572
0 36574 7 1 2 81471 36573
0 36575 5 1 1 36574
0 36576 7 1 2 99532 93985
0 36577 5 1 1 36576
0 36578 7 1 2 68445 36577
0 36579 5 1 1 36578
0 36580 7 1 2 71676 94952
0 36581 5 1 1 36580
0 36582 7 1 2 36579 36581
0 36583 5 1 1 36582
0 36584 7 1 2 83939 36583
0 36585 5 1 1 36584
0 36586 7 1 2 36575 36585
0 36587 7 1 2 36552 36586
0 36588 5 1 1 36587
0 36589 7 1 2 68097 36588
0 36590 5 1 1 36589
0 36591 7 1 2 64816 5644
0 36592 5 2 1 36591
0 36593 7 1 2 99723 104059
0 36594 5 1 1 36593
0 36595 7 1 2 78806 95882
0 36596 5 1 1 36595
0 36597 7 1 2 69921 36596
0 36598 7 1 2 36594 36597
0 36599 5 1 1 36598
0 36600 7 1 2 67694 97370
0 36601 7 1 2 36599 36600
0 36602 7 1 2 104170 36601
0 36603 5 1 1 36602
0 36604 7 1 2 101354 81965
0 36605 7 1 2 75887 36604
0 36606 5 1 1 36605
0 36607 7 1 2 36603 36606
0 36608 5 1 1 36607
0 36609 7 1 2 73187 36608
0 36610 5 1 1 36609
0 36611 7 1 2 71677 90153
0 36612 5 1 1 36611
0 36613 7 1 2 36612 86634
0 36614 5 1 1 36613
0 36615 7 1 2 70214 36614
0 36616 5 1 1 36615
0 36617 7 2 2 68446 102311
0 36618 7 1 2 73188 104172
0 36619 5 1 1 36618
0 36620 7 1 2 36616 36619
0 36621 5 1 1 36620
0 36622 7 1 2 76329 36621
0 36623 5 1 1 36622
0 36624 7 1 2 97775 76786
0 36625 5 1 1 36624
0 36626 7 1 2 99589 36625
0 36627 5 1 1 36626
0 36628 7 1 2 70215 36627
0 36629 5 1 1 36628
0 36630 7 1 2 72710 95898
0 36631 7 1 2 36629 36630
0 36632 7 1 2 36623 36631
0 36633 5 1 1 36632
0 36634 7 2 2 66575 79965
0 36635 5 1 1 104174
0 36636 7 1 2 77940 104175
0 36637 5 1 1 36636
0 36638 7 1 2 36637 89973
0 36639 5 1 1 36638
0 36640 7 1 2 69545 36639
0 36641 7 1 2 36633 36640
0 36642 5 1 1 36641
0 36643 7 1 2 36610 36642
0 36644 7 1 2 36590 36643
0 36645 5 1 1 36644
0 36646 7 1 2 71111 36645
0 36647 5 1 1 36646
0 36648 7 1 2 81747 78924
0 36649 5 2 1 36648
0 36650 7 1 2 97347 104176
0 36651 5 1 1 36650
0 36652 7 1 2 65158 36651
0 36653 5 1 1 36652
0 36654 7 1 2 101764 99000
0 36655 5 1 1 36654
0 36656 7 1 2 73189 36655
0 36657 5 1 1 36656
0 36658 7 1 2 36653 36657
0 36659 5 1 1 36658
0 36660 7 1 2 67695 36659
0 36661 5 1 1 36660
0 36662 7 3 2 95358 92756
0 36663 5 1 1 104178
0 36664 7 1 2 70216 104179
0 36665 5 1 1 36664
0 36666 7 1 2 36661 36665
0 36667 5 1 1 36666
0 36668 7 1 2 71112 36667
0 36669 5 1 1 36668
0 36670 7 1 2 86308 92258
0 36671 5 1 1 36670
0 36672 7 1 2 36663 36671
0 36673 5 1 1 36672
0 36674 7 1 2 83189 36673
0 36675 5 1 1 36674
0 36676 7 1 2 36669 36675
0 36677 5 1 1 36676
0 36678 7 1 2 97408 36677
0 36679 5 1 1 36678
0 36680 7 1 2 74552 99231
0 36681 5 1 1 36680
0 36682 7 1 2 83849 75856
0 36683 7 1 2 84256 36682
0 36684 5 1 1 36683
0 36685 7 1 2 36681 36684
0 36686 5 1 1 36685
0 36687 7 1 2 64817 36686
0 36688 5 1 1 36687
0 36689 7 1 2 91949 99232
0 36690 5 1 1 36689
0 36691 7 1 2 36688 36690
0 36692 5 1 1 36691
0 36693 7 1 2 87648 36692
0 36694 5 1 1 36693
0 36695 7 2 2 64818 75851
0 36696 5 1 1 104181
0 36697 7 1 2 25597 36696
0 36698 5 1 1 36697
0 36699 7 1 2 83850 36698
0 36700 5 1 1 36699
0 36701 7 1 2 82027 92781
0 36702 5 1 1 36701
0 36703 7 1 2 36700 36702
0 36704 5 1 1 36703
0 36705 7 1 2 103752 36704
0 36706 5 1 1 36705
0 36707 7 1 2 36694 36706
0 36708 5 1 1 36707
0 36709 7 1 2 67696 36708
0 36710 5 1 1 36709
0 36711 7 1 2 84135 83396
0 36712 5 1 1 36711
0 36713 7 1 2 83550 83158
0 36714 7 1 2 3822 36713
0 36715 5 1 1 36714
0 36716 7 1 2 36712 36715
0 36717 5 1 1 36716
0 36718 7 1 2 68682 36717
0 36719 5 1 1 36718
0 36720 7 1 2 74553 78026
0 36721 7 1 2 86445 36720
0 36722 5 1 1 36721
0 36723 7 1 2 36719 36722
0 36724 5 1 1 36723
0 36725 7 1 2 68098 36724
0 36726 5 1 1 36725
0 36727 7 1 2 74554 97519
0 36728 5 1 1 36727
0 36729 7 1 2 36726 36728
0 36730 5 1 1 36729
0 36731 7 1 2 81976 36730
0 36732 5 1 1 36731
0 36733 7 1 2 36710 36732
0 36734 7 1 2 36679 36733
0 36735 7 1 2 36647 36734
0 36736 5 1 1 36735
0 36737 7 1 2 67360 36736
0 36738 5 1 1 36737
0 36739 7 2 2 96145 95490
0 36740 7 1 2 71438 104183
0 36741 5 1 1 36740
0 36742 7 1 2 97807 36741
0 36743 5 1 1 36742
0 36744 7 1 2 71678 36743
0 36745 5 1 1 36744
0 36746 7 1 2 75692 94726
0 36747 5 1 1 36746
0 36748 7 1 2 36745 36747
0 36749 5 1 1 36748
0 36750 7 1 2 70217 36749
0 36751 5 1 1 36750
0 36752 7 1 2 74967 104173
0 36753 5 1 1 36752
0 36754 7 1 2 36751 36753
0 36755 5 1 1 36754
0 36756 7 1 2 69922 36755
0 36757 5 1 1 36756
0 36758 7 3 2 70218 83153
0 36759 7 1 2 104185 95711
0 36760 5 1 1 36759
0 36761 7 1 2 36757 36760
0 36762 5 1 1 36761
0 36763 7 1 2 103667 36762
0 36764 5 1 1 36763
0 36765 7 1 2 36738 36764
0 36766 5 1 1 36765
0 36767 7 1 2 104151 36766
0 36768 5 1 1 36767
0 36769 7 1 2 69923 20677
0 36770 5 1 1 36769
0 36771 7 2 2 94198 36770
0 36772 7 1 2 70485 104188
0 36773 5 1 1 36772
0 36774 7 1 2 86322 89252
0 36775 5 1 1 36774
0 36776 7 1 2 36773 36775
0 36777 5 1 1 36776
0 36778 7 1 2 97280 36777
0 36779 5 1 1 36778
0 36780 7 1 2 83513 92667
0 36781 5 1 1 36780
0 36782 7 2 2 82934 81530
0 36783 5 1 1 104190
0 36784 7 1 2 36781 36783
0 36785 5 1 1 36784
0 36786 7 1 2 65456 36785
0 36787 5 1 1 36786
0 36788 7 1 2 65159 74890
0 36789 5 1 1 36788
0 36790 7 1 2 101401 36789
0 36791 5 1 1 36790
0 36792 7 1 2 81531 36791
0 36793 5 1 1 36792
0 36794 7 1 2 36787 36793
0 36795 7 1 2 36779 36794
0 36796 5 1 1 36795
0 36797 7 1 2 66346 36796
0 36798 5 1 1 36797
0 36799 7 1 2 81418 80906
0 36800 5 1 1 36799
0 36801 7 1 2 79910 89057
0 36802 5 1 1 36801
0 36803 7 1 2 103656 94697
0 36804 5 1 1 36803
0 36805 7 1 2 73975 36804
0 36806 5 1 1 36805
0 36807 7 1 2 92991 36806
0 36808 7 1 2 36802 36807
0 36809 5 1 1 36808
0 36810 7 1 2 67697 36809
0 36811 5 1 1 36810
0 36812 7 1 2 36800 36811
0 36813 5 1 1 36812
0 36814 7 1 2 64437 36813
0 36815 5 1 1 36814
0 36816 7 1 2 36798 36815
0 36817 5 1 1 36816
0 36818 7 1 2 73190 36817
0 36819 5 1 1 36818
0 36820 7 1 2 87455 95227
0 36821 5 1 1 36820
0 36822 7 2 2 80100 86478
0 36823 7 1 2 76599 104192
0 36824 5 1 1 36823
0 36825 7 1 2 36821 36824
0 36826 5 1 1 36825
0 36827 7 1 2 73762 36826
0 36828 5 1 1 36827
0 36829 7 2 2 76229 83374
0 36830 5 1 1 104194
0 36831 7 1 2 36828 36830
0 36832 5 1 1 36831
0 36833 7 1 2 67698 36832
0 36834 5 1 1 36833
0 36835 7 1 2 71844 94877
0 36836 5 1 1 36835
0 36837 7 1 2 75090 36836
0 36838 5 1 1 36837
0 36839 7 1 2 85017 36838
0 36840 5 1 1 36839
0 36841 7 1 2 80101 83940
0 36842 5 1 1 36841
0 36843 7 1 2 36840 36842
0 36844 5 1 1 36843
0 36845 7 1 2 77103 36844
0 36846 5 1 1 36845
0 36847 7 1 2 100645 101732
0 36848 5 1 1 36847
0 36849 7 1 2 73763 36848
0 36850 5 1 1 36849
0 36851 7 1 2 69924 83383
0 36852 5 1 1 36851
0 36853 7 1 2 71439 36852
0 36854 5 1 1 36853
0 36855 7 1 2 36850 36854
0 36856 5 1 1 36855
0 36857 7 1 2 85018 36856
0 36858 5 1 1 36857
0 36859 7 1 2 36846 36858
0 36860 7 1 2 36834 36859
0 36861 5 1 1 36860
0 36862 7 1 2 64438 36861
0 36863 5 1 1 36862
0 36864 7 1 2 36819 36863
0 36865 5 1 1 36864
0 36866 7 1 2 72428 36865
0 36867 5 1 1 36866
0 36868 7 4 2 99155 84459
0 36869 5 1 1 104196
0 36870 7 2 2 82247 95042
0 36871 7 1 2 104197 104200
0 36872 5 1 1 36871
0 36873 7 1 2 36867 36872
0 36874 5 1 1 36873
0 36875 7 1 2 66034 36874
0 36876 5 1 1 36875
0 36877 7 2 2 84407 99264
0 36878 7 1 2 104201 104202
0 36879 5 1 1 36878
0 36880 7 1 2 36876 36879
0 36881 5 1 1 36880
0 36882 7 1 2 103887 36881
0 36883 5 1 1 36882
0 36884 7 2 2 98113 103340
0 36885 7 1 2 75834 104204
0 36886 5 1 1 36885
0 36887 7 1 2 102550 99086
0 36888 7 1 2 84334 36887
0 36889 5 1 1 36888
0 36890 7 1 2 36886 36889
0 36891 5 1 1 36890
0 36892 7 1 2 77371 36891
0 36893 5 1 1 36892
0 36894 7 1 2 101182 18045
0 36895 5 4 1 36894
0 36896 7 2 2 100820 104206
0 36897 5 1 1 104210
0 36898 7 1 2 104152 104211
0 36899 5 1 1 36898
0 36900 7 1 2 36893 36899
0 36901 5 1 1 36900
0 36902 7 1 2 71679 36901
0 36903 5 1 1 36902
0 36904 7 1 2 91509 102589
0 36905 5 1 1 36904
0 36906 7 1 2 36897 36905
0 36907 5 1 1 36906
0 36908 7 1 2 70219 104153
0 36909 7 1 2 36907 36908
0 36910 5 1 1 36909
0 36911 7 1 2 36903 36910
0 36912 5 1 1 36911
0 36913 7 1 2 69925 36912
0 36914 5 1 1 36913
0 36915 7 1 2 96802 82152
0 36916 5 1 1 36915
0 36917 7 1 2 76051 81472
0 36918 7 1 2 75474 36917
0 36919 5 1 1 36918
0 36920 7 1 2 36916 36919
0 36921 5 1 1 36920
0 36922 7 1 2 71113 36921
0 36923 5 1 1 36922
0 36924 7 1 2 83139 92268
0 36925 7 1 2 81263 36924
0 36926 5 1 1 36925
0 36927 7 1 2 36923 36926
0 36928 5 1 1 36927
0 36929 7 1 2 103912 36928
0 36930 5 1 1 36929
0 36931 7 1 2 36914 36930
0 36932 5 1 1 36931
0 36933 7 1 2 85632 36932
0 36934 5 1 1 36933
0 36935 7 1 2 36883 36934
0 36936 7 1 2 36768 36935
0 36937 5 1 1 36936
0 36938 7 1 2 85530 36937
0 36939 5 1 1 36938
0 36940 7 1 2 86061 102160
0 36941 5 2 1 36940
0 36942 7 1 2 76488 87832
0 36943 5 1 1 36942
0 36944 7 1 2 104212 36943
0 36945 5 2 1 36944
0 36946 7 1 2 78140 104214
0 36947 5 1 1 36946
0 36948 7 1 2 76330 87288
0 36949 5 1 1 36948
0 36950 7 1 2 86951 36949
0 36951 5 1 1 36950
0 36952 7 1 2 76331 86812
0 36953 5 1 1 36952
0 36954 7 1 2 82320 36953
0 36955 5 1 1 36954
0 36956 7 1 2 36951 36955
0 36957 5 1 1 36956
0 36958 7 1 2 76600 36957
0 36959 5 1 1 36958
0 36960 7 1 2 88313 6265
0 36961 7 1 2 94698 36960
0 36962 5 1 1 36961
0 36963 7 1 2 73976 36962
0 36964 5 1 1 36963
0 36965 7 1 2 89058 95896
0 36966 5 1 1 36965
0 36967 7 1 2 648 36966
0 36968 7 1 2 36964 36967
0 36969 5 1 1 36968
0 36970 7 1 2 73191 36969
0 36971 5 1 1 36970
0 36972 7 1 2 36959 36971
0 36973 5 1 1 36972
0 36974 7 1 2 100500 36973
0 36975 5 1 1 36974
0 36976 7 1 2 36947 36975
0 36977 5 1 1 36976
0 36978 7 1 2 67209 36977
0 36979 5 1 1 36978
0 36980 7 2 2 95692 104186
0 36981 5 2 1 104216
0 36982 7 3 2 68099 94750
0 36983 5 2 1 104220
0 36984 7 1 2 71680 104184
0 36985 5 1 1 36984
0 36986 7 1 2 104223 36985
0 36987 5 1 1 36986
0 36988 7 1 2 70220 36987
0 36989 5 1 1 36988
0 36990 7 1 2 71681 94751
0 36991 5 1 1 36990
0 36992 7 1 2 36991 90008
0 36993 5 3 1 36992
0 36994 7 1 2 68100 104225
0 36995 5 1 1 36994
0 36996 7 1 2 36989 36995
0 36997 5 1 1 36996
0 36998 7 1 2 69926 36997
0 36999 5 1 1 36998
0 37000 7 1 2 104218 36999
0 37001 5 3 1 37000
0 37002 7 1 2 69927 104217
0 37003 5 1 1 37002
0 37004 7 1 2 66347 37003
0 37005 5 1 1 37004
0 37006 7 2 2 104228 37005
0 37007 7 1 2 103801 104231
0 37008 5 1 1 37007
0 37009 7 1 2 36979 37008
0 37010 5 1 1 37009
0 37011 7 1 2 67699 37010
0 37012 5 1 1 37011
0 37013 7 1 2 83247 80538
0 37014 5 1 1 37013
0 37015 7 1 2 87248 93920
0 37016 7 1 2 92974 37015
0 37017 5 1 1 37016
0 37018 7 1 2 71440 37017
0 37019 5 1 1 37018
0 37020 7 1 2 99583 99888
0 37021 7 1 2 37019 37020
0 37022 5 1 1 37021
0 37023 7 1 2 68101 37022
0 37024 5 1 1 37023
0 37025 7 1 2 37014 37024
0 37026 5 1 1 37025
0 37027 7 1 2 70486 37026
0 37028 5 1 1 37027
0 37029 7 1 2 76332 101696
0 37030 5 2 1 37029
0 37031 7 1 2 80165 104233
0 37032 5 1 1 37031
0 37033 7 1 2 83070 37032
0 37034 5 1 1 37033
0 37035 7 1 2 100861 37034
0 37036 7 1 2 37028 37035
0 37037 5 1 1 37036
0 37038 7 1 2 64439 37037
0 37039 5 1 1 37038
0 37040 7 1 2 77964 92204
0 37041 5 1 1 37040
0 37042 7 1 2 79253 37041
0 37043 5 1 1 37042
0 37044 7 1 2 64819 37043
0 37045 5 1 1 37044
0 37046 7 1 2 76418 98638
0 37047 5 1 1 37046
0 37048 7 1 2 37045 37047
0 37049 5 1 1 37048
0 37050 7 1 2 68102 37049
0 37051 5 1 1 37050
0 37052 7 1 2 81362 78837
0 37053 5 1 1 37052
0 37054 7 1 2 37051 37053
0 37055 5 1 1 37054
0 37056 7 1 2 82987 37055
0 37057 5 1 1 37056
0 37058 7 1 2 79070 81383
0 37059 5 1 1 37058
0 37060 7 1 2 84556 100638
0 37061 5 1 1 37060
0 37062 7 1 2 37059 37061
0 37063 5 1 1 37062
0 37064 7 1 2 73764 37063
0 37065 5 1 1 37064
0 37066 7 1 2 79578 83477
0 37067 5 1 1 37066
0 37068 7 1 2 66348 83159
0 37069 7 1 2 94727 37068
0 37070 5 1 1 37069
0 37071 7 1 2 37067 37070
0 37072 5 1 1 37071
0 37073 7 1 2 82118 37072
0 37074 5 1 1 37073
0 37075 7 1 2 37065 37074
0 37076 5 1 1 37075
0 37077 7 1 2 82012 37076
0 37078 5 1 1 37077
0 37079 7 1 2 37057 37078
0 37080 7 1 2 37039 37079
0 37081 5 1 1 37080
0 37082 7 1 2 66035 37081
0 37083 5 1 1 37082
0 37084 7 1 2 88352 93269
0 37085 5 1 1 37084
0 37086 7 1 2 80329 102332
0 37087 5 1 1 37086
0 37088 7 1 2 37085 37087
0 37089 5 1 1 37088
0 37090 7 1 2 76230 82604
0 37091 7 1 2 37089 37090
0 37092 5 1 1 37091
0 37093 7 1 2 37083 37092
0 37094 5 1 1 37093
0 37095 7 1 2 67210 101055
0 37096 7 1 2 37094 37095
0 37097 5 1 1 37096
0 37098 7 1 2 37012 37097
0 37099 5 1 1 37098
0 37100 7 1 2 67361 37099
0 37101 5 1 1 37100
0 37102 7 1 2 92630 103396
0 37103 5 1 1 37102
0 37104 7 1 2 66576 93169
0 37105 5 1 1 37104
0 37106 7 1 2 37103 37105
0 37107 5 1 1 37106
0 37108 7 1 2 78032 37107
0 37109 5 1 1 37108
0 37110 7 1 2 91464 37109
0 37111 5 1 1 37110
0 37112 7 1 2 73765 37111
0 37113 5 1 1 37112
0 37114 7 1 2 66577 10223
0 37115 5 1 1 37114
0 37116 7 1 2 70221 102977
0 37117 7 1 2 37115 37116
0 37118 5 1 1 37117
0 37119 7 1 2 33144 37118
0 37120 5 1 1 37119
0 37121 7 1 2 82248 37120
0 37122 5 1 1 37121
0 37123 7 1 2 103555 4367
0 37124 5 1 1 37123
0 37125 7 1 2 37122 37124
0 37126 5 1 1 37125
0 37127 7 1 2 69546 37126
0 37128 5 1 1 37127
0 37129 7 1 2 37113 37128
0 37130 5 1 1 37129
0 37131 7 1 2 70487 37130
0 37132 5 1 1 37131
0 37133 7 1 2 79828 103623
0 37134 5 1 1 37133
0 37135 7 1 2 77571 90933
0 37136 5 1 1 37135
0 37137 7 1 2 33942 37136
0 37138 5 1 1 37137
0 37139 7 1 2 93681 37138
0 37140 5 1 1 37139
0 37141 7 1 2 37134 37140
0 37142 5 1 1 37141
0 37143 7 1 2 82988 37142
0 37144 5 1 1 37143
0 37145 7 1 2 75981 102904
0 37146 5 1 1 37145
0 37147 7 1 2 103552 37146
0 37148 5 1 1 37147
0 37149 7 1 2 67700 92992
0 37150 5 2 1 37149
0 37151 7 1 2 86768 87815
0 37152 7 1 2 104235 37151
0 37153 7 1 2 37148 37152
0 37154 5 1 1 37153
0 37155 7 1 2 37144 37154
0 37156 5 1 1 37155
0 37157 7 1 2 69547 37156
0 37158 5 1 1 37157
0 37159 7 1 2 37132 37158
0 37160 5 1 1 37159
0 37161 7 1 2 71114 37160
0 37162 5 1 1 37161
0 37163 7 3 2 69548 81419
0 37164 5 1 1 104237
0 37165 7 1 2 104238 82864
0 37166 5 1 1 37165
0 37167 7 1 2 95213 104226
0 37168 5 1 1 37167
0 37169 7 1 2 37166 37168
0 37170 5 1 1 37169
0 37171 7 1 2 77542 37170
0 37172 5 1 1 37171
0 37173 7 1 2 37162 37172
0 37174 5 1 1 37173
0 37175 7 1 2 67211 99387
0 37176 7 1 2 37174 37175
0 37177 5 1 1 37176
0 37178 7 1 2 37101 37177
0 37179 5 1 1 37178
0 37180 7 1 2 75773 37179
0 37181 5 1 1 37180
0 37182 7 2 2 95204 97164
0 37183 7 1 2 103479 104240
0 37184 5 1 1 37183
0 37185 7 1 2 81748 97903
0 37186 5 1 1 37185
0 37187 7 1 2 72429 95201
0 37188 5 1 1 37187
0 37189 7 1 2 65160 98501
0 37190 7 1 2 37188 37189
0 37191 5 1 1 37190
0 37192 7 1 2 37186 37191
0 37193 5 1 1 37192
0 37194 7 1 2 85093 37193
0 37195 5 1 1 37194
0 37196 7 1 2 37184 37195
0 37197 5 1 1 37196
0 37198 7 1 2 69928 37197
0 37199 5 1 1 37198
0 37200 7 1 2 78807 74336
0 37201 7 1 2 104241 37200
0 37202 5 1 1 37201
0 37203 7 1 2 37199 37202
0 37204 5 1 1 37203
0 37205 7 1 2 71682 37204
0 37206 5 1 1 37205
0 37207 7 1 2 96815 99539
0 37208 7 1 2 103730 74344
0 37209 7 1 2 37207 37208
0 37210 5 1 1 37209
0 37211 7 1 2 37206 37210
0 37212 5 1 1 37211
0 37213 7 1 2 104154 37212
0 37214 5 1 1 37213
0 37215 7 3 2 77773 85428
0 37216 7 1 2 92384 104205
0 37217 7 1 2 104242 37216
0 37218 7 1 2 96578 37217
0 37219 5 1 1 37218
0 37220 7 1 2 37214 37219
0 37221 5 1 1 37220
0 37222 7 1 2 69214 37221
0 37223 5 1 1 37222
0 37224 7 1 2 103882 90262
0 37225 7 2 2 102536 37224
0 37226 7 1 2 81749 104245
0 37227 5 1 1 37226
0 37228 7 1 2 95509 75755
0 37229 7 1 2 82321 37228
0 37230 7 1 2 103896 37229
0 37231 5 1 1 37230
0 37232 7 1 2 37227 37231
0 37233 5 1 1 37232
0 37234 7 1 2 71683 37233
0 37235 5 1 1 37234
0 37236 7 1 2 96561 104246
0 37237 5 1 1 37236
0 37238 7 1 2 37235 37237
0 37239 5 1 1 37238
0 37240 7 1 2 93608 37239
0 37241 5 1 1 37240
0 37242 7 1 2 37223 37241
0 37243 5 1 1 37242
0 37244 7 1 2 68447 37243
0 37245 5 1 1 37244
0 37246 7 1 2 75930 91502
0 37247 5 2 1 37246
0 37248 7 1 2 85043 86872
0 37249 5 1 1 37248
0 37250 7 1 2 104247 37249
0 37251 5 1 1 37250
0 37252 7 1 2 66578 37251
0 37253 5 1 1 37252
0 37254 7 1 2 100826 97770
0 37255 5 1 1 37254
0 37256 7 1 2 81439 103188
0 37257 5 1 1 37256
0 37258 7 1 2 37255 37257
0 37259 5 1 1 37258
0 37260 7 1 2 66759 37259
0 37261 5 1 1 37260
0 37262 7 1 2 80082 81440
0 37263 7 1 2 83990 37262
0 37264 5 1 1 37263
0 37265 7 1 2 37261 37264
0 37266 7 1 2 37253 37265
0 37267 5 1 1 37266
0 37268 7 1 2 103914 37267
0 37269 5 1 1 37268
0 37270 7 1 2 102185 102392
0 37271 7 1 2 87456 37270
0 37272 7 1 2 90263 37271
0 37273 7 1 2 93010 37272
0 37274 5 1 1 37273
0 37275 7 1 2 37269 37274
0 37276 5 1 1 37275
0 37277 7 1 2 69215 37276
0 37278 5 1 1 37277
0 37279 7 2 2 64159 103888
0 37280 7 1 2 87457 104249
0 37281 7 1 2 90771 34085
0 37282 5 1 1 37281
0 37283 7 1 2 73766 98435
0 37284 5 1 1 37283
0 37285 7 1 2 97924 37284
0 37286 5 2 1 37285
0 37287 7 1 2 37282 104251
0 37288 7 1 2 37280 37287
0 37289 5 1 1 37288
0 37290 7 1 2 37278 37289
0 37291 5 1 1 37290
0 37292 7 1 2 83375 37291
0 37293 5 1 1 37292
0 37294 7 1 2 99639 93011
0 37295 5 1 1 37294
0 37296 7 2 2 93218 99021
0 37297 5 2 1 104253
0 37298 7 1 2 64160 104254
0 37299 5 1 1 37298
0 37300 7 1 2 37295 37299
0 37301 5 1 1 37300
0 37302 7 1 2 73767 37301
0 37303 5 1 1 37302
0 37304 7 1 2 92189 97697
0 37305 5 1 1 37304
0 37306 7 1 2 37303 37305
0 37307 5 1 1 37306
0 37308 7 1 2 103889 37307
0 37309 5 1 1 37308
0 37310 7 6 2 82451 104155
0 37311 7 1 2 101404 97127
0 37312 7 1 2 104257 37311
0 37313 5 1 1 37312
0 37314 7 1 2 37309 37313
0 37315 5 1 1 37314
0 37316 7 1 2 104193 37315
0 37317 5 1 1 37316
0 37318 7 1 2 37293 37317
0 37319 5 1 1 37318
0 37320 7 1 2 64820 37319
0 37321 5 1 1 37320
0 37322 7 2 2 67212 68103
0 37323 7 1 2 89756 104263
0 37324 7 1 2 100473 37323
0 37325 7 1 2 86946 104036
0 37326 7 1 2 37324 37325
0 37327 7 1 2 99601 37326
0 37328 5 1 1 37327
0 37329 7 1 2 37321 37328
0 37330 7 1 2 37245 37329
0 37331 5 1 1 37330
0 37332 7 1 2 77265 37331
0 37333 5 1 1 37332
0 37334 7 2 2 76489 97050
0 37335 5 5 1 104265
0 37336 7 2 2 68104 94284
0 37337 5 1 1 104272
0 37338 7 1 2 104266 104273
0 37339 5 1 1 37338
0 37340 7 1 2 73768 86110
0 37341 5 1 1 37340
0 37342 7 1 2 75091 101727
0 37343 5 1 1 37342
0 37344 7 1 2 74680 37343
0 37345 5 1 1 37344
0 37346 7 1 2 95901 37345
0 37347 7 1 2 37341 37346
0 37348 5 1 1 37347
0 37349 7 1 2 68105 37348
0 37350 5 1 1 37349
0 37351 7 1 2 103214 37350
0 37352 5 1 1 37351
0 37353 7 1 2 96755 37352
0 37354 5 1 1 37353
0 37355 7 1 2 37339 37354
0 37356 5 1 1 37355
0 37357 7 1 2 102500 37356
0 37358 5 1 1 37357
0 37359 7 4 2 74401 102164
0 37360 7 1 2 75018 104274
0 37361 5 1 1 37360
0 37362 7 1 2 75931 102246
0 37363 5 4 1 37362
0 37364 7 1 2 102168 104278
0 37365 5 2 1 37364
0 37366 7 1 2 74402 104282
0 37367 5 1 1 37366
0 37368 7 3 2 98114 95293
0 37369 7 1 2 82452 103310
0 37370 7 1 2 104284 37369
0 37371 5 1 1 37370
0 37372 7 1 2 37367 37371
0 37373 5 1 1 37372
0 37374 7 1 2 82274 37373
0 37375 5 1 1 37374
0 37376 7 1 2 37361 37375
0 37377 5 1 1 37376
0 37378 7 1 2 64821 37377
0 37379 5 1 1 37378
0 37380 7 1 2 104275 89967
0 37381 5 1 1 37380
0 37382 7 1 2 37379 37381
0 37383 5 1 1 37382
0 37384 7 1 2 73977 37383
0 37385 5 1 1 37384
0 37386 7 1 2 101997 77700
0 37387 5 1 1 37386
0 37388 7 1 2 102169 37387
0 37389 5 1 1 37388
0 37390 7 1 2 74403 37389
0 37391 5 1 1 37390
0 37392 7 3 2 82453 103240
0 37393 5 1 1 104287
0 37394 7 1 2 103644 104288
0 37395 5 1 1 37394
0 37396 7 1 2 37391 37395
0 37397 5 1 1 37396
0 37398 7 1 2 66349 37397
0 37399 5 1 1 37398
0 37400 7 1 2 87038 104276
0 37401 5 1 1 37400
0 37402 7 1 2 37399 37401
0 37403 5 1 1 37402
0 37404 7 1 2 64822 37403
0 37405 5 1 1 37404
0 37406 7 1 2 104277 93293
0 37407 5 1 1 37406
0 37408 7 1 2 37405 37407
0 37409 5 1 1 37408
0 37410 7 1 2 82322 37409
0 37411 5 1 1 37410
0 37412 7 1 2 37385 37411
0 37413 7 1 2 37358 37412
0 37414 5 1 1 37413
0 37415 7 1 2 77372 37414
0 37416 5 1 1 37415
0 37417 7 1 2 77572 81556
0 37418 7 1 2 88766 37417
0 37419 5 1 1 37418
0 37420 7 1 2 103558 37419
0 37421 5 1 1 37420
0 37422 7 1 2 73535 37421
0 37423 5 1 1 37422
0 37424 7 1 2 79829 85633
0 37425 5 1 1 37424
0 37426 7 2 2 76659 86062
0 37427 7 1 2 68448 104290
0 37428 5 1 1 37427
0 37429 7 1 2 37425 37428
0 37430 5 1 1 37429
0 37431 7 1 2 82249 37430
0 37432 5 1 1 37431
0 37433 7 1 2 37423 37432
0 37434 5 1 1 37433
0 37435 7 1 2 104007 37434
0 37436 5 1 1 37435
0 37437 7 1 2 37416 37436
0 37438 5 1 1 37437
0 37439 7 1 2 76906 37438
0 37440 5 1 1 37439
0 37441 7 1 2 78663 94330
0 37442 5 1 1 37441
0 37443 7 1 2 94161 37442
0 37444 5 1 1 37443
0 37445 7 1 2 104258 37444
0 37446 5 1 1 37445
0 37447 7 5 2 65832 104250
0 37448 7 1 2 82390 87649
0 37449 7 1 2 104292 37448
0 37450 5 1 1 37449
0 37451 7 1 2 37446 37450
0 37452 5 1 1 37451
0 37453 7 1 2 64823 37452
0 37454 5 1 1 37453
0 37455 7 1 2 99003 104259
0 37456 5 1 1 37455
0 37457 7 1 2 99935 104293
0 37458 5 1 1 37457
0 37459 7 1 2 37456 37458
0 37460 5 1 1 37459
0 37461 7 1 2 92771 37460
0 37462 5 1 1 37461
0 37463 7 1 2 37454 37462
0 37464 5 1 1 37463
0 37465 7 1 2 70222 37464
0 37466 5 1 1 37465
0 37467 7 2 2 103014 98062
0 37468 7 1 2 73536 104297
0 37469 5 1 1 37468
0 37470 7 1 2 85695 104294
0 37471 5 1 1 37470
0 37472 7 1 2 37469 37471
0 37473 5 1 1 37472
0 37474 7 1 2 73769 37473
0 37475 5 1 1 37474
0 37476 7 1 2 89790 104260
0 37477 5 1 1 37476
0 37478 7 1 2 37475 37477
0 37479 5 1 1 37478
0 37480 7 1 2 66579 37479
0 37481 5 1 1 37480
0 37482 7 1 2 73770 103048
0 37483 7 2 2 98154 37482
0 37484 7 1 2 89155 77774
0 37485 7 1 2 104299 37484
0 37486 5 1 1 37485
0 37487 7 1 2 37481 37486
0 37488 5 1 1 37487
0 37489 7 1 2 65161 37488
0 37490 5 1 1 37489
0 37491 7 1 2 87514 75835
0 37492 7 1 2 104300 37491
0 37493 5 1 1 37492
0 37494 7 1 2 37490 37493
0 37495 5 1 1 37494
0 37496 7 1 2 84408 37495
0 37497 5 1 1 37496
0 37498 7 1 2 37466 37497
0 37499 5 1 1 37498
0 37500 7 1 2 101942 37499
0 37501 5 1 1 37500
0 37502 7 1 2 64440 99907
0 37503 5 1 1 37502
0 37504 7 2 2 64824 37503
0 37505 5 1 1 104301
0 37506 7 1 2 26114 103415
0 37507 5 2 1 37506
0 37508 7 1 2 69929 104303
0 37509 5 1 1 37508
0 37510 7 1 2 69549 82717
0 37511 5 1 1 37510
0 37512 7 1 2 37509 37511
0 37513 7 1 2 37505 37512
0 37514 5 1 1 37513
0 37515 7 1 2 104261 37514
0 37516 5 1 1 37515
0 37517 7 1 2 103890 93080
0 37518 7 1 2 99896 37517
0 37519 5 1 1 37518
0 37520 7 1 2 37516 37519
0 37521 5 1 1 37520
0 37522 7 1 2 70488 37521
0 37523 5 1 1 37522
0 37524 7 1 2 69930 99892
0 37525 5 1 1 37524
0 37526 7 2 2 69550 79911
0 37527 5 2 1 104305
0 37528 7 1 2 104097 104307
0 37529 7 1 2 37525 37528
0 37530 5 1 1 37529
0 37531 7 1 2 104295 37530
0 37532 5 1 1 37531
0 37533 7 1 2 64825 94965
0 37534 5 1 1 37533
0 37535 7 2 2 99567 104156
0 37536 7 1 2 98642 94868
0 37537 7 1 2 104309 37536
0 37538 7 1 2 37534 37537
0 37539 5 1 1 37538
0 37540 7 1 2 37532 37539
0 37541 7 1 2 37523 37540
0 37542 5 1 1 37541
0 37543 7 1 2 71115 37542
0 37544 5 1 1 37543
0 37545 7 1 2 73537 79032
0 37546 5 1 1 37545
0 37547 7 1 2 83652 37546
0 37548 5 3 1 37547
0 37549 7 1 2 104296 104311
0 37550 5 1 1 37549
0 37551 7 1 2 100023 104298
0 37552 5 1 1 37551
0 37553 7 1 2 37550 37552
0 37554 5 1 1 37553
0 37555 7 1 2 68683 37554
0 37556 5 1 1 37555
0 37557 7 1 2 88857 103891
0 37558 7 1 2 93081 37557
0 37559 5 1 1 37558
0 37560 7 1 2 37556 37559
0 37561 5 1 1 37560
0 37562 7 1 2 71845 37561
0 37563 5 1 1 37562
0 37564 7 4 2 98326 92128
0 37565 7 1 2 103721 103015
0 37566 7 1 2 104314 37565
0 37567 5 1 1 37566
0 37568 7 1 2 82119 103892
0 37569 7 1 2 84429 37568
0 37570 5 1 1 37569
0 37571 7 1 2 37567 37570
0 37572 5 1 1 37571
0 37573 7 1 2 86651 37572
0 37574 5 1 1 37573
0 37575 7 1 2 37563 37574
0 37576 5 1 1 37575
0 37577 7 1 2 83190 37576
0 37578 5 1 1 37577
0 37579 7 1 2 77174 104262
0 37580 5 1 1 37579
0 37581 7 1 2 77469 95632
0 37582 7 2 2 74404 101573
0 37583 7 1 2 104318 95769
0 37584 7 1 2 37581 37583
0 37585 5 1 1 37584
0 37586 7 1 2 37580 37585
0 37587 5 1 1 37586
0 37588 7 1 2 64826 37587
0 37589 5 1 1 37588
0 37590 7 1 2 36136 15501
0 37591 5 1 1 37590
0 37592 7 1 2 95337 104310
0 37593 7 1 2 37591 37592
0 37594 5 1 1 37593
0 37595 7 1 2 37589 37594
0 37596 5 1 1 37595
0 37597 7 1 2 82989 37596
0 37598 5 1 1 37597
0 37599 7 1 2 37578 37598
0 37600 7 1 2 37544 37599
0 37601 5 1 1 37600
0 37602 7 1 2 72430 37601
0 37603 5 1 1 37602
0 37604 7 1 2 72166 100084
0 37605 7 1 2 102004 37604
0 37606 7 1 2 102085 37605
0 37607 5 1 1 37606
0 37608 7 1 2 37603 37607
0 37609 5 1 1 37608
0 37610 7 1 2 93012 37609
0 37611 5 1 1 37610
0 37612 7 1 2 37501 37611
0 37613 7 1 2 37440 37612
0 37614 7 1 2 37333 37613
0 37615 7 1 2 37181 37614
0 37616 7 1 2 36939 37615
0 37617 5 1 1 37616
0 37618 7 1 2 74038 37617
0 37619 5 1 1 37618
0 37620 7 1 2 36492 37619
0 37621 7 1 2 35827 37620
0 37622 7 1 2 33984 37621
0 37623 5 1 1 37622
0 37624 7 1 2 102267 37623
0 37625 5 1 1 37624
0 37626 7 1 2 68996 6110
0 37627 5 1 1 37626
0 37628 7 1 2 63909 16826
0 37629 5 1 1 37628
0 37630 7 8 2 37627 37629
0 37631 7 1 2 65162 13131
0 37632 5 1 1 37631
0 37633 7 1 2 13251 37632
0 37634 5 1 1 37633
0 37635 7 3 2 66036 84460
0 37636 7 1 2 85456 104328
0 37637 5 1 1 37636
0 37638 7 2 2 64161 66037
0 37639 5 1 1 104331
0 37640 7 1 2 92340 37639
0 37641 7 1 2 101513 37640
0 37642 5 1 1 37641
0 37643 7 1 2 37637 37642
0 37644 5 1 1 37643
0 37645 7 1 2 37634 37644
0 37646 5 1 1 37645
0 37647 7 2 2 70843 84461
0 37648 5 1 1 104333
0 37649 7 1 2 93750 104334
0 37650 5 1 1 37649
0 37651 7 1 2 65833 83706
0 37652 7 1 2 91743 37651
0 37653 5 1 1 37652
0 37654 7 1 2 37650 37653
0 37655 5 1 1 37654
0 37656 7 1 2 104332 37655
0 37657 5 1 1 37656
0 37658 7 1 2 37646 37657
0 37659 5 1 1 37658
0 37660 7 1 2 72711 37659
0 37661 5 1 1 37660
0 37662 7 3 2 96005 96032
0 37663 5 1 1 104335
0 37664 7 1 2 78576 101977
0 37665 7 1 2 104336 37664
0 37666 5 1 1 37665
0 37667 7 1 2 37661 37666
0 37668 5 1 1 37667
0 37669 7 1 2 66350 37668
0 37670 5 1 1 37669
0 37671 7 2 2 74681 94761
0 37672 5 1 1 104338
0 37673 7 1 2 73771 89376
0 37674 5 1 1 37673
0 37675 7 1 2 37672 37674
0 37676 5 2 1 37675
0 37677 7 1 2 81532 104340
0 37678 5 1 1 37677
0 37679 7 3 2 82120 98983
0 37680 7 1 2 103507 104342
0 37681 5 1 1 37680
0 37682 7 1 2 37678 37681
0 37683 5 1 1 37682
0 37684 7 1 2 101978 37683
0 37685 5 1 1 37684
0 37686 7 1 2 37670 37685
0 37687 5 1 1 37686
0 37688 7 1 2 73192 37687
0 37689 5 1 1 37688
0 37690 7 2 2 90107 93449
0 37691 5 1 1 104345
0 37692 7 1 2 65457 104346
0 37693 5 1 1 37692
0 37694 7 1 2 88691 81033
0 37695 5 1 1 37694
0 37696 7 1 2 37693 37695
0 37697 5 1 1 37696
0 37698 7 1 2 65834 37697
0 37699 5 1 1 37698
0 37700 7 1 2 89608 83294
0 37701 7 1 2 103875 37700
0 37702 5 1 1 37701
0 37703 7 1 2 37699 37702
0 37704 5 1 1 37703
0 37705 7 1 2 72712 37704
0 37706 5 1 1 37705
0 37707 7 1 2 81399 96105
0 37708 5 1 1 37707
0 37709 7 1 2 37706 37708
0 37710 5 1 1 37709
0 37711 7 1 2 64162 37710
0 37712 5 1 1 37711
0 37713 7 2 2 78577 93142
0 37714 7 1 2 86546 93120
0 37715 7 1 2 101318 37714
0 37716 7 1 2 104347 37715
0 37717 5 1 1 37716
0 37718 7 1 2 37712 37717
0 37719 5 1 1 37718
0 37720 7 1 2 76231 37719
0 37721 5 1 1 37720
0 37722 7 1 2 37689 37721
0 37723 5 1 1 37722
0 37724 7 1 2 78225 37723
0 37725 5 1 1 37724
0 37726 7 1 2 83582 97343
0 37727 5 1 1 37726
0 37728 7 1 2 66760 94163
0 37729 5 1 1 37728
0 37730 7 1 2 37727 37729
0 37731 5 1 1 37730
0 37732 7 1 2 92570 37731
0 37733 5 1 1 37732
0 37734 7 3 2 83816 98860
0 37735 7 1 2 74174 82683
0 37736 7 1 2 104349 37735
0 37737 5 1 1 37736
0 37738 7 1 2 37733 37737
0 37739 5 1 1 37738
0 37740 7 1 2 66038 37739
0 37741 5 1 1 37740
0 37742 7 1 2 71116 94382
0 37743 7 1 2 95303 37742
0 37744 5 1 1 37743
0 37745 7 1 2 37741 37744
0 37746 5 1 1 37745
0 37747 7 1 2 93049 99309
0 37748 7 1 2 37746 37747
0 37749 5 1 1 37748
0 37750 7 1 2 37725 37749
0 37751 5 1 1 37750
0 37752 7 1 2 67362 37751
0 37753 5 1 1 37752
0 37754 7 2 2 101995 81190
0 37755 7 1 2 87677 104352
0 37756 5 1 1 37755
0 37757 7 1 2 77875 80122
0 37758 5 2 1 37757
0 37759 7 1 2 34264 104354
0 37760 5 1 1 37759
0 37761 7 1 2 71441 37760
0 37762 5 1 1 37761
0 37763 7 1 2 70223 84388
0 37764 5 1 1 37763
0 37765 7 1 2 37762 37764
0 37766 5 1 1 37765
0 37767 7 1 2 64441 37766
0 37768 5 1 1 37767
0 37769 7 1 2 70224 74154
0 37770 5 1 1 37769
0 37771 7 1 2 75287 74156
0 37772 7 1 2 77589 37771
0 37773 5 1 1 37772
0 37774 7 1 2 37770 37773
0 37775 5 1 1 37774
0 37776 7 1 2 81237 37775
0 37777 5 1 1 37776
0 37778 7 1 2 37768 37777
0 37779 5 1 1 37778
0 37780 7 1 2 73538 37779
0 37781 5 1 1 37780
0 37782 7 1 2 101672 92429
0 37783 5 1 1 37782
0 37784 7 1 2 37781 37783
0 37785 5 1 1 37784
0 37786 7 1 2 85141 37785
0 37787 5 1 1 37786
0 37788 7 1 2 37756 37787
0 37789 5 1 1 37788
0 37790 7 1 2 64163 37789
0 37791 5 1 1 37790
0 37792 7 1 2 74356 101893
0 37793 7 1 2 104353 37792
0 37794 5 1 1 37793
0 37795 7 1 2 37791 37794
0 37796 5 1 1 37795
0 37797 7 1 2 72713 37796
0 37798 5 1 1 37797
0 37799 7 2 2 101555 78226
0 37800 7 1 2 104356 84266
0 37801 5 1 1 37800
0 37802 7 1 2 37798 37801
0 37803 5 1 1 37802
0 37804 7 1 2 73772 37803
0 37805 5 1 1 37804
0 37806 7 2 2 92806 91002
0 37807 7 1 2 92524 104358
0 37808 5 1 1 37807
0 37809 7 1 2 37805 37808
0 37810 5 1 1 37809
0 37811 7 1 2 80715 37810
0 37812 5 1 1 37811
0 37813 7 1 2 95548 95233
0 37814 5 1 1 37813
0 37815 7 1 2 15451 37814
0 37816 5 1 1 37815
0 37817 7 1 2 81007 83274
0 37818 5 1 1 37817
0 37819 7 2 2 81097 37818
0 37820 7 1 2 37816 104360
0 37821 5 1 1 37820
0 37822 7 2 2 86218 76707
0 37823 5 2 1 104362
0 37824 7 1 2 78227 104363
0 37825 5 1 1 37824
0 37826 7 1 2 95549 92487
0 37827 5 1 1 37826
0 37828 7 1 2 37825 37827
0 37829 5 1 1 37828
0 37830 7 1 2 87701 37829
0 37831 5 1 1 37830
0 37832 7 1 2 81034 96064
0 37833 5 1 1 37832
0 37834 7 1 2 37831 37833
0 37835 5 1 1 37834
0 37836 7 1 2 64827 37835
0 37837 5 1 1 37836
0 37838 7 1 2 87669 76787
0 37839 7 1 2 95850 37838
0 37840 5 1 1 37839
0 37841 7 1 2 37837 37840
0 37842 5 1 1 37841
0 37843 7 1 2 66351 37842
0 37844 5 1 1 37843
0 37845 7 1 2 37821 37844
0 37846 5 1 1 37845
0 37847 7 1 2 72714 37846
0 37848 5 1 1 37847
0 37849 7 1 2 93934 92009
0 37850 5 1 1 37849
0 37851 7 1 2 3745 37850
0 37852 5 1 1 37851
0 37853 7 1 2 95214 91003
0 37854 7 1 2 37852 37853
0 37855 5 1 1 37854
0 37856 7 1 2 37848 37855
0 37857 5 1 1 37856
0 37858 7 1 2 64164 37857
0 37859 5 1 1 37858
0 37860 7 1 2 99119 84984
0 37861 7 1 2 84469 37860
0 37862 5 1 1 37861
0 37863 7 1 2 70844 37862
0 37864 7 1 2 37859 37863
0 37865 7 1 2 37812 37864
0 37866 5 1 1 37865
0 37867 7 6 2 93609 85081
0 37868 5 2 1 104366
0 37869 7 1 2 72715 85389
0 37870 5 1 1 37869
0 37871 7 1 2 104372 37870
0 37872 5 1 1 37871
0 37873 7 1 2 83591 37872
0 37874 5 1 1 37873
0 37875 7 1 2 80023 93093
0 37876 5 1 1 37875
0 37877 7 1 2 86025 90098
0 37878 5 1 1 37877
0 37879 7 1 2 66580 101653
0 37880 5 1 1 37879
0 37881 7 1 2 37878 37880
0 37882 5 1 1 37881
0 37883 7 1 2 64442 86708
0 37884 7 1 2 37882 37883
0 37885 5 1 1 37884
0 37886 7 1 2 37876 37885
0 37887 5 1 1 37886
0 37888 7 1 2 69216 37887
0 37889 5 1 1 37888
0 37890 7 1 2 37874 37889
0 37891 5 1 1 37890
0 37892 7 1 2 73539 37891
0 37893 5 1 1 37892
0 37894 7 1 2 64443 89708
0 37895 5 1 1 37894
0 37896 7 1 2 93619 37895
0 37897 5 1 1 37896
0 37898 7 1 2 74192 95241
0 37899 5 1 1 37898
0 37900 7 1 2 37897 37899
0 37901 5 1 1 37900
0 37902 7 1 2 65458 37901
0 37903 5 1 1 37902
0 37904 7 1 2 76232 87846
0 37905 5 2 1 37904
0 37906 7 2 2 73193 87515
0 37907 7 1 2 65163 104376
0 37908 5 1 1 37907
0 37909 7 1 2 104374 37908
0 37910 5 1 1 37909
0 37911 7 1 2 74193 37910
0 37912 5 1 1 37911
0 37913 7 3 2 76490 78126
0 37914 5 1 1 104378
0 37915 7 3 2 69217 66352
0 37916 7 2 2 84462 104381
0 37917 5 1 1 104384
0 37918 7 1 2 37914 37917
0 37919 5 1 1 37918
0 37920 7 1 2 80419 37919
0 37921 5 1 1 37920
0 37922 7 2 2 70489 84035
0 37923 7 1 2 68449 100257
0 37924 7 1 2 104386 37923
0 37925 5 1 1 37924
0 37926 7 1 2 37921 37925
0 37927 7 1 2 37912 37926
0 37928 7 1 2 37903 37927
0 37929 5 1 1 37928
0 37930 7 1 2 67701 37929
0 37931 5 1 1 37930
0 37932 7 1 2 74856 92086
0 37933 5 1 1 37932
0 37934 7 1 2 82063 83275
0 37935 7 1 2 37933 37934
0 37936 5 1 1 37935
0 37937 7 1 2 94716 96528
0 37938 7 1 2 37936 37937
0 37939 5 1 1 37938
0 37940 7 3 2 69218 80024
0 37941 7 1 2 95476 104388
0 37942 5 1 1 37941
0 37943 7 1 2 66039 37942
0 37944 7 1 2 37939 37943
0 37945 7 1 2 37931 37944
0 37946 7 1 2 37893 37945
0 37947 5 1 1 37946
0 37948 7 3 2 73194 79855
0 37949 7 1 2 79040 94986
0 37950 5 1 1 37949
0 37951 7 1 2 104391 37950
0 37952 5 1 1 37951
0 37953 7 1 2 88692 79282
0 37954 5 1 1 37953
0 37955 7 1 2 37952 37954
0 37956 5 1 1 37955
0 37957 7 1 2 71442 37956
0 37958 5 1 1 37957
0 37959 7 1 2 82056 19103
0 37960 5 1 1 37959
0 37961 7 1 2 37958 37960
0 37962 5 1 1 37961
0 37963 7 1 2 67702 37962
0 37964 5 1 1 37963
0 37965 7 1 2 80631 101416
0 37966 5 1 1 37965
0 37967 7 2 2 71684 83397
0 37968 7 1 2 74905 104394
0 37969 5 1 1 37968
0 37970 7 1 2 37966 37969
0 37971 5 1 1 37970
0 37972 7 1 2 68684 37971
0 37973 5 2 1 37972
0 37974 7 1 2 69931 86111
0 37975 5 1 1 37974
0 37976 7 1 2 104396 37975
0 37977 5 1 1 37976
0 37978 7 1 2 81473 37977
0 37979 5 1 1 37978
0 37980 7 1 2 37964 37979
0 37981 5 1 1 37980
0 37982 7 1 2 64165 37981
0 37983 5 1 1 37982
0 37984 7 1 2 86035 83361
0 37985 5 1 1 37984
0 37986 7 1 2 69551 37985
0 37987 5 1 1 37986
0 37988 7 1 2 99315 14151
0 37989 7 1 2 37987 37988
0 37990 5 1 1 37989
0 37991 7 1 2 71117 37990
0 37992 7 1 2 37983 37991
0 37993 5 1 1 37992
0 37994 7 1 2 91004 37993
0 37995 7 1 2 37947 37994
0 37996 5 1 1 37995
0 37997 7 1 2 65164 75082
0 37998 5 1 1 37997
0 37999 7 1 2 82180 37998
0 38000 5 2 1 37999
0 38001 7 1 2 66040 104398
0 38002 5 1 1 38001
0 38003 7 1 2 38002 6214
0 38004 5 1 1 38003
0 38005 7 1 2 66581 38004
0 38006 5 1 1 38005
0 38007 7 1 2 66353 81115
0 38008 5 1 1 38007
0 38009 7 1 2 38006 38008
0 38010 5 1 1 38009
0 38011 7 1 2 64444 38010
0 38012 5 1 1 38011
0 38013 7 2 2 69552 78319
0 38014 7 1 2 104400 80323
0 38015 5 1 1 38014
0 38016 7 1 2 38012 38015
0 38017 5 1 1 38016
0 38018 7 1 2 99573 38017
0 38019 5 1 1 38018
0 38020 7 1 2 88678 101315
0 38021 5 1 1 38020
0 38022 7 1 2 101311 38021
0 38023 5 1 1 38022
0 38024 7 1 2 70225 38023
0 38025 5 1 1 38024
0 38026 7 3 2 76708 88879
0 38027 7 1 2 66582 104399
0 38028 5 1 1 38027
0 38029 7 1 2 66354 82121
0 38030 5 1 1 38029
0 38031 7 1 2 38028 38030
0 38032 5 1 1 38031
0 38033 7 1 2 104402 38032
0 38034 5 1 1 38033
0 38035 7 1 2 38025 38034
0 38036 5 1 1 38035
0 38037 7 1 2 64166 38036
0 38038 5 1 1 38037
0 38039 7 1 2 67703 38038
0 38040 7 1 2 38019 38039
0 38041 5 1 1 38040
0 38042 7 1 2 27733 95104
0 38043 5 1 1 38042
0 38044 7 1 2 88401 38043
0 38045 5 1 1 38044
0 38046 7 1 2 86330 38045
0 38047 5 1 1 38046
0 38048 7 1 2 81035 38047
0 38049 5 1 1 38048
0 38050 7 2 2 78664 86036
0 38051 5 1 1 104405
0 38052 7 2 2 81264 80123
0 38053 7 1 2 104406 104407
0 38054 5 1 1 38053
0 38055 7 1 2 38049 38054
0 38056 5 1 1 38055
0 38057 7 1 2 69219 38056
0 38058 5 1 1 38057
0 38059 7 1 2 101014 80907
0 38060 5 1 1 38059
0 38061 7 2 2 69220 81036
0 38062 7 1 2 75288 97932
0 38063 7 1 2 104409 38062
0 38064 5 1 1 38063
0 38065 7 1 2 38060 38064
0 38066 5 1 1 38065
0 38067 7 1 2 71443 38066
0 38068 5 1 1 38067
0 38069 7 1 2 72716 38068
0 38070 7 1 2 38058 38069
0 38071 5 1 1 38070
0 38072 7 1 2 73195 38071
0 38073 7 1 2 38041 38072
0 38074 5 1 1 38073
0 38075 7 1 2 81505 104367
0 38076 5 1 1 38075
0 38077 7 1 2 68450 93094
0 38078 7 1 2 93126 38077
0 38079 5 1 1 38078
0 38080 7 1 2 38076 38079
0 38081 5 1 1 38080
0 38082 7 1 2 66761 38081
0 38083 5 1 1 38082
0 38084 7 1 2 76688 93121
0 38085 7 1 2 103266 38084
0 38086 5 1 1 38085
0 38087 7 1 2 38083 38086
0 38088 5 1 1 38087
0 38089 7 1 2 65459 38088
0 38090 5 1 1 38089
0 38091 7 1 2 88478 94433
0 38092 5 1 1 38091
0 38093 7 1 2 99316 38092
0 38094 5 1 1 38093
0 38095 7 1 2 38090 38094
0 38096 5 1 1 38095
0 38097 7 1 2 81037 38096
0 38098 5 1 1 38097
0 38099 7 1 2 81506 84101
0 38100 5 1 1 38099
0 38101 7 1 2 74682 82208
0 38102 5 1 1 38101
0 38103 7 1 2 38100 38102
0 38104 5 1 1 38103
0 38105 7 1 2 81750 38104
0 38106 5 1 1 38105
0 38107 7 1 2 100752 81966
0 38108 7 1 2 101835 38107
0 38109 5 1 1 38108
0 38110 7 1 2 38106 38109
0 38111 5 1 1 38110
0 38112 7 1 2 101015 38111
0 38113 5 1 1 38112
0 38114 7 1 2 38098 38113
0 38115 7 1 2 38074 38114
0 38116 5 1 1 38115
0 38117 7 1 2 85142 38116
0 38118 5 1 1 38117
0 38119 7 1 2 65835 38118
0 38120 7 1 2 37996 38119
0 38121 5 1 1 38120
0 38122 7 1 2 72431 38121
0 38123 7 1 2 37866 38122
0 38124 5 1 1 38123
0 38125 7 1 2 37753 38124
0 38126 5 1 1 38125
0 38127 7 1 2 72264 38126
0 38128 5 1 1 38127
0 38129 7 3 2 86547 83044
0 38130 7 1 2 95934 104411
0 38131 5 1 1 38130
0 38132 7 1 2 23937 93944
0 38133 5 1 1 38132
0 38134 7 1 2 65460 38133
0 38135 5 1 1 38134
0 38136 7 1 2 65165 93690
0 38137 5 1 1 38136
0 38138 7 1 2 38135 38137
0 38139 5 1 1 38138
0 38140 7 1 2 78228 38139
0 38141 5 1 1 38140
0 38142 7 2 2 101846 96171
0 38143 7 1 2 77300 104414
0 38144 5 1 1 38143
0 38145 7 1 2 87702 91005
0 38146 5 1 1 38145
0 38147 7 1 2 83223 78349
0 38148 7 1 2 93147 38147
0 38149 5 1 1 38148
0 38150 7 1 2 38146 38149
0 38151 5 1 1 38150
0 38152 7 1 2 80420 38151
0 38153 5 1 1 38152
0 38154 7 1 2 38144 38153
0 38155 7 1 2 38141 38154
0 38156 5 1 1 38155
0 38157 7 1 2 73196 38156
0 38158 5 1 1 38157
0 38159 7 1 2 38131 38158
0 38160 5 1 1 38159
0 38161 7 1 2 101998 103746
0 38162 7 1 2 38160 38161
0 38163 5 1 1 38162
0 38164 7 1 2 38128 38163
0 38165 5 1 1 38164
0 38166 7 1 2 67123 38165
0 38167 5 1 1 38166
0 38168 7 3 2 89929 78350
0 38169 7 2 2 101883 104416
0 38170 7 2 2 69553 84339
0 38171 7 1 2 100538 104421
0 38172 5 1 1 38171
0 38173 7 1 2 88402 101000
0 38174 5 1 1 38173
0 38175 7 1 2 38172 38174
0 38176 5 1 1 38175
0 38177 7 1 2 104419 38176
0 38178 5 1 1 38177
0 38179 7 5 2 68872 92488
0 38180 7 1 2 70845 98115
0 38181 7 1 2 103034 38180
0 38182 7 1 2 104423 38181
0 38183 5 1 1 38182
0 38184 7 1 2 100768 92976
0 38185 5 1 1 38184
0 38186 7 2 2 73197 104424
0 38187 5 1 1 104428
0 38188 7 1 2 67363 104429
0 38189 5 1 1 38188
0 38190 7 1 2 38185 38189
0 38191 5 1 1 38190
0 38192 7 1 2 65836 85634
0 38193 7 1 2 38191 38192
0 38194 5 1 1 38193
0 38195 7 1 2 38183 38194
0 38196 5 1 1 38195
0 38197 7 1 2 69932 38196
0 38198 5 1 1 38197
0 38199 7 1 2 38178 38198
0 38200 5 1 1 38199
0 38201 7 1 2 71444 38200
0 38202 5 1 1 38201
0 38203 7 1 2 81284 77880
0 38204 5 1 1 38203
0 38205 7 1 2 82171 38204
0 38206 5 1 1 38205
0 38207 7 1 2 73198 95102
0 38208 5 1 1 38207
0 38209 7 1 2 38206 38208
0 38210 5 1 1 38209
0 38211 7 1 2 88369 38210
0 38212 5 1 1 38211
0 38213 7 1 2 86219 79199
0 38214 5 1 1 38213
0 38215 7 1 2 65166 94902
0 38216 5 1 1 38215
0 38217 7 1 2 38214 38216
0 38218 5 1 1 38217
0 38219 7 1 2 77952 38218
0 38220 5 1 1 38219
0 38221 7 1 2 88875 38220
0 38222 7 1 2 38212 38221
0 38223 5 1 1 38222
0 38224 7 1 2 97882 38223
0 38225 5 1 1 38224
0 38226 7 3 2 80716 81038
0 38227 7 3 2 83817 104430
0 38228 7 1 2 73540 103210
0 38229 7 1 2 104433 38228
0 38230 5 1 1 38229
0 38231 7 1 2 38225 38230
0 38232 5 1 1 38231
0 38233 7 1 2 85143 38232
0 38234 5 1 1 38233
0 38235 7 4 2 73199 89043
0 38236 5 1 1 104436
0 38237 7 1 2 88370 89226
0 38238 5 1 1 38237
0 38239 7 1 2 38238 104375
0 38240 7 1 2 38236 38239
0 38241 5 1 1 38240
0 38242 7 1 2 93074 91006
0 38243 7 1 2 38241 38242
0 38244 5 1 1 38243
0 38245 7 1 2 38234 38244
0 38246 5 1 1 38245
0 38247 7 1 2 67364 38246
0 38248 5 1 1 38247
0 38249 7 3 2 71118 89087
0 38250 7 1 2 74345 90009
0 38251 7 1 2 104440 38250
0 38252 7 1 2 72432 75756
0 38253 7 1 2 85635 38252
0 38254 7 1 2 86517 38253
0 38255 7 1 2 38251 38254
0 38256 5 1 1 38255
0 38257 7 1 2 38248 38256
0 38258 7 1 2 38202 38257
0 38259 5 1 1 38258
0 38260 7 1 2 67704 38259
0 38261 5 1 1 38260
0 38262 7 1 2 86328 80102
0 38263 5 1 1 38262
0 38264 7 1 2 99606 92010
0 38265 5 1 1 38264
0 38266 7 1 2 38263 38265
0 38267 5 1 1 38266
0 38268 7 1 2 38267 91051
0 38269 5 1 1 38268
0 38270 7 4 2 76233 91007
0 38271 7 1 2 73200 104443
0 38272 5 1 1 38271
0 38273 7 1 2 38269 38272
0 38274 5 1 1 38273
0 38275 7 1 2 81039 38274
0 38276 5 1 1 38275
0 38277 7 1 2 71119 89258
0 38278 7 1 2 101794 38277
0 38279 5 1 1 38278
0 38280 7 1 2 66041 74857
0 38281 7 1 2 95069 38280
0 38282 5 1 1 38281
0 38283 7 1 2 38279 38282
0 38284 5 1 1 38283
0 38285 7 1 2 78229 38284
0 38286 5 1 1 38285
0 38287 7 1 2 84409 91104
0 38288 7 1 2 96182 38287
0 38289 5 1 1 38288
0 38290 7 1 2 38286 38289
0 38291 5 1 1 38290
0 38292 7 1 2 75932 38291
0 38293 5 1 1 38292
0 38294 7 1 2 38276 38293
0 38295 5 1 1 38294
0 38296 7 1 2 67365 38295
0 38297 5 1 1 38296
0 38298 7 2 2 97954 78320
0 38299 7 1 2 74155 104447
0 38300 5 1 1 38299
0 38301 7 1 2 73201 99258
0 38302 5 1 1 38301
0 38303 7 1 2 38300 38302
0 38304 5 1 1 38303
0 38305 7 1 2 69554 38304
0 38306 5 1 1 38305
0 38307 7 1 2 104448 95456
0 38308 5 1 1 38307
0 38309 7 1 2 38306 38308
0 38310 5 1 1 38309
0 38311 7 1 2 94065 85104
0 38312 7 1 2 38310 38311
0 38313 5 1 1 38312
0 38314 7 4 2 90895 76394
0 38315 5 1 1 104449
0 38316 7 1 2 72433 101268
0 38317 7 1 2 104450 38316
0 38318 5 1 1 38317
0 38319 7 1 2 38313 38318
0 38320 5 1 1 38319
0 38321 7 1 2 80717 38320
0 38322 5 1 1 38321
0 38323 7 1 2 80632 91008
0 38324 7 3 2 72434 74793
0 38325 7 1 2 97648 104453
0 38326 7 1 2 38323 38325
0 38327 5 1 1 38326
0 38328 7 1 2 38322 38327
0 38329 7 1 2 38297 38328
0 38330 5 1 1 38329
0 38331 7 1 2 96082 38330
0 38332 5 1 1 38331
0 38333 7 1 2 38261 38332
0 38334 5 1 1 38333
0 38335 7 1 2 69221 38334
0 38336 5 1 1 38335
0 38337 7 2 2 88403 75083
0 38338 5 1 1 104456
0 38339 7 1 2 90719 75757
0 38340 7 2 2 104457 38339
0 38341 5 1 1 104458
0 38342 7 1 2 96756 104459
0 38343 5 1 1 38342
0 38344 7 1 2 18024 104267
0 38345 5 1 1 38344
0 38346 7 4 2 76358 78174
0 38347 5 1 1 104460
0 38348 7 1 2 86677 104461
0 38349 7 1 2 38345 38348
0 38350 5 1 1 38349
0 38351 7 1 2 38343 38350
0 38352 5 1 1 38351
0 38353 7 1 2 71120 38352
0 38354 5 1 1 38353
0 38355 7 2 2 88404 84490
0 38356 7 2 2 98781 104464
0 38357 7 1 2 100035 104466
0 38358 5 1 1 38357
0 38359 7 1 2 38354 38358
0 38360 5 1 1 38359
0 38361 7 1 2 69555 38360
0 38362 5 1 1 38361
0 38363 7 2 2 64445 80835
0 38364 7 1 2 68873 104468
0 38365 7 1 2 104467 38364
0 38366 5 1 1 38365
0 38367 7 1 2 38362 38366
0 38368 5 1 1 38367
0 38369 7 1 2 65837 38368
0 38370 5 1 1 38369
0 38371 7 2 2 97051 82568
0 38372 5 1 1 104470
0 38373 7 2 2 72717 78578
0 38374 7 1 2 97739 104472
0 38375 5 1 1 38374
0 38376 7 1 2 38372 38375
0 38377 5 1 1 38376
0 38378 7 1 2 64446 38377
0 38379 5 1 1 38378
0 38380 7 1 2 89913 97074
0 38381 5 1 1 38380
0 38382 7 1 2 38379 38381
0 38383 5 1 1 38382
0 38384 7 1 2 80718 38383
0 38385 5 1 1 38384
0 38386 7 1 2 83045 95313
0 38387 7 1 2 98221 38386
0 38388 5 1 1 38387
0 38389 7 1 2 38385 38388
0 38390 5 1 1 38389
0 38391 7 1 2 99742 90069
0 38392 7 1 2 38390 38391
0 38393 5 1 1 38392
0 38394 7 1 2 38370 38393
0 38395 5 1 1 38394
0 38396 7 1 2 69222 38395
0 38397 5 1 1 38396
0 38398 7 1 2 98217 87104
0 38399 7 1 2 86520 38398
0 38400 5 1 1 38399
0 38401 7 1 2 38341 38400
0 38402 5 1 1 38401
0 38403 7 1 2 100104 101094
0 38404 7 1 2 38402 38403
0 38405 5 1 1 38404
0 38406 7 1 2 38397 38405
0 38407 5 1 1 38406
0 38408 7 1 2 75416 38407
0 38409 5 1 1 38408
0 38410 7 1 2 77175 104252
0 38411 5 1 1 38410
0 38412 7 1 2 103596 38411
0 38413 5 1 1 38412
0 38414 7 1 2 69223 38413
0 38415 5 1 1 38414
0 38416 7 1 2 103601 38415
0 38417 5 1 1 38416
0 38418 7 1 2 86709 38417
0 38419 5 1 1 38418
0 38420 7 2 2 96757 81040
0 38421 5 1 1 104474
0 38422 7 1 2 102837 104475
0 38423 5 1 1 38422
0 38424 7 1 2 38419 38423
0 38425 5 1 1 38424
0 38426 7 1 2 38425 96142
0 38427 5 1 1 38426
0 38428 7 1 2 102319 98057
0 38429 7 1 2 90654 97296
0 38430 7 1 2 38428 38429
0 38431 5 1 1 38430
0 38432 7 1 2 38427 38431
0 38433 5 1 1 38432
0 38434 7 1 2 66355 38433
0 38435 5 1 1 38434
0 38436 7 1 2 85457 101173
0 38437 5 1 1 38436
0 38438 7 1 2 104115 38437
0 38439 5 1 1 38438
0 38440 7 1 2 92977 97202
0 38441 7 1 2 38439 38440
0 38442 5 1 1 38441
0 38443 7 1 2 38435 38442
0 38444 5 1 1 38443
0 38445 7 1 2 87361 38444
0 38446 5 1 1 38445
0 38447 7 1 2 68451 100705
0 38448 5 1 1 38447
0 38449 7 1 2 86151 38448
0 38450 5 1 1 38449
0 38451 7 1 2 101324 38450
0 38452 5 1 1 38451
0 38453 7 1 2 23200 104355
0 38454 5 1 1 38453
0 38455 7 1 2 69556 38454
0 38456 5 1 1 38455
0 38457 7 1 2 71685 104469
0 38458 5 1 1 38457
0 38459 7 1 2 38456 38458
0 38460 5 1 1 38459
0 38461 7 1 2 71445 38460
0 38462 5 1 1 38461
0 38463 7 1 2 75933 101539
0 38464 5 1 1 38463
0 38465 7 1 2 38462 38464
0 38466 5 1 1 38465
0 38467 7 1 2 73541 38466
0 38468 5 1 1 38467
0 38469 7 2 2 71121 80025
0 38470 7 1 2 78771 104476
0 38471 5 1 1 38470
0 38472 7 1 2 38468 38471
0 38473 5 1 1 38472
0 38474 7 1 2 88405 38473
0 38475 5 1 1 38474
0 38476 7 1 2 38452 38475
0 38477 5 1 1 38476
0 38478 7 1 2 85144 38477
0 38479 5 1 1 38478
0 38480 7 1 2 104444 82570
0 38481 5 1 1 38480
0 38482 7 1 2 38479 38481
0 38483 5 1 1 38482
0 38484 7 2 2 99449 92807
0 38485 7 1 2 38483 104478
0 38486 5 1 1 38485
0 38487 7 1 2 38446 38486
0 38488 7 1 2 38409 38487
0 38489 7 1 2 38336 38488
0 38490 5 1 1 38489
0 38491 7 1 2 67213 38490
0 38492 5 1 1 38491
0 38493 7 1 2 84057 95757
0 38494 7 2 2 67366 92352
0 38495 7 1 2 84030 104480
0 38496 7 1 2 38493 38495
0 38497 7 1 2 103802 38496
0 38498 5 1 1 38497
0 38499 7 1 2 38492 38498
0 38500 5 1 1 38499
0 38501 7 1 2 72167 38500
0 38502 5 1 1 38501
0 38503 7 1 2 73202 103181
0 38504 5 1 1 38503
0 38505 7 2 2 86972 38504
0 38506 5 1 1 104482
0 38507 7 1 2 99407 38506
0 38508 5 1 1 38507
0 38509 7 1 2 84844 83823
0 38510 5 2 1 38509
0 38511 7 1 2 104484 80486
0 38512 5 1 1 38511
0 38513 7 1 2 98436 93378
0 38514 7 1 2 38512 38513
0 38515 5 1 1 38514
0 38516 7 1 2 97904 95168
0 38517 5 2 1 38516
0 38518 7 1 2 100378 104454
0 38519 5 1 1 38518
0 38520 7 1 2 104486 38519
0 38521 5 1 1 38520
0 38522 7 1 2 69224 38521
0 38523 5 1 1 38522
0 38524 7 1 2 99461 88460
0 38525 5 1 1 38524
0 38526 7 1 2 38523 38525
0 38527 5 1 1 38526
0 38528 7 1 2 80719 38527
0 38529 5 1 1 38528
0 38530 7 1 2 38515 38529
0 38531 7 1 2 38508 38530
0 38532 5 1 1 38531
0 38533 7 1 2 78508 38532
0 38534 5 1 1 38533
0 38535 7 1 2 80720 88461
0 38536 5 1 1 38535
0 38537 7 1 2 104483 38536
0 38538 5 1 1 38537
0 38539 7 1 2 102320 85392
0 38540 7 1 2 38538 38539
0 38541 5 1 1 38540
0 38542 7 1 2 38534 38541
0 38543 5 1 1 38542
0 38544 7 1 2 102682 38543
0 38545 5 1 1 38544
0 38546 7 1 2 81369 86973
0 38547 5 2 1 38546
0 38548 7 1 2 98502 77373
0 38549 5 1 1 38548
0 38550 7 2 2 98611 74068
0 38551 5 2 1 104490
0 38552 7 1 2 38549 104492
0 38553 5 1 1 38552
0 38554 7 1 2 64167 38553
0 38555 5 1 1 38554
0 38556 7 1 2 19240 38555
0 38557 5 1 1 38556
0 38558 7 1 2 104488 38557
0 38559 5 1 1 38558
0 38560 7 1 2 77374 98384
0 38561 5 1 1 38560
0 38562 7 1 2 98374 98523
0 38563 5 1 1 38562
0 38564 7 1 2 38561 38563
0 38565 5 1 1 38564
0 38566 7 1 2 64168 38565
0 38567 5 1 1 38566
0 38568 7 1 2 98375 98732
0 38569 5 1 1 38568
0 38570 7 1 2 38567 38569
0 38571 5 1 1 38570
0 38572 7 1 2 81894 38571
0 38573 5 1 1 38572
0 38574 7 1 2 80633 103501
0 38575 5 1 1 38574
0 38576 7 1 2 38573 38575
0 38577 5 1 1 38576
0 38578 7 1 2 82708 38577
0 38579 5 1 1 38578
0 38580 7 1 2 38559 38579
0 38581 5 1 1 38580
0 38582 7 1 2 72718 38581
0 38583 5 1 1 38582
0 38584 7 2 2 81751 73978
0 38585 5 3 1 104494
0 38586 7 2 2 82709 104496
0 38587 5 1 1 104499
0 38588 7 1 2 97569 104500
0 38589 7 1 2 92894 38588
0 38590 5 1 1 38589
0 38591 7 1 2 38583 38590
0 38592 5 1 1 38591
0 38593 7 1 2 102625 38592
0 38594 5 1 1 38593
0 38595 7 1 2 38545 38594
0 38596 5 1 1 38595
0 38597 7 1 2 70226 38596
0 38598 5 1 1 38597
0 38599 7 3 2 73203 86983
0 38600 7 1 2 102853 104501
0 38601 5 1 1 38600
0 38602 7 2 2 66762 102665
0 38603 7 1 2 83487 104504
0 38604 5 1 1 38603
0 38605 7 1 2 38601 38604
0 38606 5 1 1 38605
0 38607 7 1 2 72435 38606
0 38608 5 1 1 38607
0 38609 7 2 2 81895 85531
0 38610 7 7 2 72168 103294
0 38611 7 1 2 81363 104508
0 38612 7 1 2 104506 38611
0 38613 5 1 1 38612
0 38614 7 1 2 38608 38613
0 38615 5 1 1 38614
0 38616 7 1 2 68685 38615
0 38617 5 1 1 38616
0 38618 7 3 2 73204 83154
0 38619 5 1 1 104515
0 38620 7 2 2 89727 104516
0 38621 7 1 2 100907 103295
0 38622 7 1 2 104518 38621
0 38623 5 1 1 38622
0 38624 7 1 2 38617 38623
0 38625 5 1 1 38624
0 38626 7 1 2 78509 38625
0 38627 5 1 1 38626
0 38628 7 4 2 82454 98222
0 38629 5 1 1 104520
0 38630 7 1 2 102683 104521
0 38631 5 1 1 38630
0 38632 7 1 2 98748 103354
0 38633 5 1 1 38632
0 38634 7 1 2 38631 38633
0 38635 5 1 1 38634
0 38636 7 1 2 86063 38635
0 38637 5 1 1 38636
0 38638 7 3 2 65838 67124
0 38639 7 2 2 101556 104524
0 38640 7 1 2 72265 100983
0 38641 7 1 2 104527 38640
0 38642 5 1 1 38641
0 38643 7 1 2 38637 38642
0 38644 5 1 1 38643
0 38645 7 1 2 72719 38644
0 38646 5 1 1 38645
0 38647 7 3 2 81896 81041
0 38648 5 1 1 104529
0 38649 7 1 2 78542 103355
0 38650 7 1 2 104530 38649
0 38651 5 1 1 38650
0 38652 7 1 2 38646 38651
0 38653 5 1 1 38652
0 38654 7 1 2 81364 38653
0 38655 5 1 1 38654
0 38656 7 1 2 38627 38655
0 38657 7 1 2 38598 38656
0 38658 5 1 1 38657
0 38659 7 1 2 85145 38658
0 38660 5 1 1 38659
0 38661 7 1 2 86868 102733
0 38662 5 1 1 38661
0 38663 7 1 2 100118 102770
0 38664 5 1 1 38663
0 38665 7 1 2 38662 38664
0 38666 5 1 1 38665
0 38667 7 1 2 66042 38666
0 38668 5 1 1 38667
0 38669 7 5 2 69557 72169
0 38670 7 2 2 71122 67214
0 38671 7 5 2 104532 104537
0 38672 7 1 2 98503 86781
0 38673 7 1 2 104539 38672
0 38674 5 1 1 38673
0 38675 7 1 2 38668 38674
0 38676 5 1 1 38675
0 38677 7 1 2 64169 38676
0 38678 5 1 1 38677
0 38679 7 1 2 98504 99809
0 38680 5 1 1 38679
0 38681 7 1 2 104493 38680
0 38682 5 1 1 38681
0 38683 7 1 2 68686 38682
0 38684 5 1 1 38683
0 38685 7 1 2 29061 38684
0 38686 5 1 1 38685
0 38687 7 1 2 67215 38686
0 38688 5 1 1 38687
0 38689 7 4 2 69558 67367
0 38690 7 1 2 72266 95338
0 38691 7 1 2 104544 38690
0 38692 7 1 2 88384 38691
0 38693 5 1 1 38692
0 38694 7 1 2 38688 38693
0 38695 5 1 1 38694
0 38696 7 1 2 102791 38695
0 38697 5 1 1 38696
0 38698 7 1 2 38678 38697
0 38699 5 1 1 38698
0 38700 7 1 2 68452 38699
0 38701 5 1 1 38700
0 38702 7 1 2 100107 34804
0 38703 5 1 1 38702
0 38704 7 1 2 98505 38703
0 38705 5 1 1 38704
0 38706 7 1 2 99462 81110
0 38707 5 1 1 38706
0 38708 7 1 2 101031 38707
0 38709 7 1 2 38705 38708
0 38710 5 1 1 38709
0 38711 7 1 2 102684 38710
0 38712 5 1 1 38711
0 38713 7 1 2 103049 97475
0 38714 7 1 2 101979 38713
0 38715 5 1 1 38714
0 38716 7 1 2 38712 38715
0 38717 5 1 1 38716
0 38718 7 1 2 86678 38717
0 38719 5 1 1 38718
0 38720 7 1 2 38701 38719
0 38721 5 1 1 38720
0 38722 7 1 2 74555 38721
0 38723 5 1 1 38722
0 38724 7 2 2 77176 102229
0 38725 7 1 2 78020 102827
0 38726 7 1 2 104548 38725
0 38727 5 1 1 38726
0 38728 7 1 2 38723 38727
0 38729 5 1 1 38728
0 38730 7 1 2 82028 38729
0 38731 5 1 1 38730
0 38732 7 1 2 94862 104509
0 38733 5 1 1 38732
0 38734 7 1 2 102742 38733
0 38735 5 1 1 38734
0 38736 7 1 2 65461 38735
0 38737 5 1 1 38736
0 38738 7 1 2 80421 102734
0 38739 5 2 1 38738
0 38740 7 1 2 98176 102707
0 38741 5 1 1 38740
0 38742 7 1 2 104550 38741
0 38743 7 1 2 38737 38742
0 38744 5 1 1 38743
0 38745 7 1 2 68106 38744
0 38746 5 1 1 38745
0 38747 7 1 2 87215 102810
0 38748 5 1 1 38747
0 38749 7 1 2 82416 102856
0 38750 7 1 2 102368 38749
0 38751 5 1 1 38750
0 38752 7 1 2 38748 38751
0 38753 7 1 2 38746 38752
0 38754 5 1 1 38753
0 38755 7 1 2 64170 38754
0 38756 5 1 1 38755
0 38757 7 1 2 98506 102799
0 38758 7 1 2 102425 38757
0 38759 5 1 1 38758
0 38760 7 1 2 38756 38759
0 38761 5 1 1 38760
0 38762 7 1 2 81042 38761
0 38763 5 1 1 38762
0 38764 7 1 2 67705 38763
0 38765 7 1 2 38731 38764
0 38766 5 1 1 38765
0 38767 7 1 2 82581 104107
0 38768 5 1 1 38767
0 38769 7 1 2 102424 89851
0 38770 7 1 2 97498 38769
0 38771 5 1 1 38770
0 38772 7 1 2 77177 38771
0 38773 5 1 1 38772
0 38774 7 1 2 38768 38773
0 38775 5 1 1 38774
0 38776 7 1 2 102763 38775
0 38777 5 1 1 38776
0 38778 7 1 2 65462 27761
0 38779 5 1 1 38778
0 38780 7 1 2 33586 96595
0 38781 5 1 1 38780
0 38782 7 1 2 64447 38781
0 38783 5 1 1 38782
0 38784 7 1 2 38779 38783
0 38785 5 1 1 38784
0 38786 7 1 2 98992 38785
0 38787 5 1 1 38786
0 38788 7 1 2 77992 98459
0 38789 7 1 2 102426 38788
0 38790 5 1 1 38789
0 38791 7 1 2 38787 38790
0 38792 5 1 1 38791
0 38793 7 1 2 102626 38792
0 38794 5 1 1 38793
0 38795 7 1 2 64171 38794
0 38796 7 1 2 38777 38795
0 38797 5 1 1 38796
0 38798 7 1 2 85696 103599
0 38799 5 1 1 38798
0 38800 7 2 2 71846 98177
0 38801 7 1 2 82417 104552
0 38802 5 1 1 38801
0 38803 7 1 2 81752 102818
0 38804 5 1 1 38803
0 38805 7 1 2 38802 38804
0 38806 5 1 1 38805
0 38807 7 1 2 101385 38806
0 38808 5 1 1 38807
0 38809 7 1 2 38799 38808
0 38810 5 1 1 38809
0 38811 7 1 2 102685 38810
0 38812 5 1 1 38811
0 38813 7 1 2 85697 102857
0 38814 7 1 2 96106 38813
0 38815 5 1 1 38814
0 38816 7 1 2 38812 38815
0 38817 5 1 1 38816
0 38818 7 1 2 68107 38817
0 38819 5 1 1 38818
0 38820 7 1 2 98437 102370
0 38821 5 1 1 38820
0 38822 7 1 2 97905 97512
0 38823 5 1 1 38822
0 38824 7 1 2 38821 38823
0 38825 5 1 1 38824
0 38826 7 1 2 65463 38825
0 38827 5 1 1 38826
0 38828 7 1 2 98438 85636
0 38829 7 1 2 87643 38828
0 38830 5 1 1 38829
0 38831 7 1 2 38827 38830
0 38832 5 1 1 38831
0 38833 7 1 2 75417 38832
0 38834 5 1 1 38833
0 38835 7 1 2 95047 102453
0 38836 5 1 1 38835
0 38837 7 2 2 72436 100379
0 38838 5 1 1 104554
0 38839 7 1 2 88430 104555
0 38840 5 1 1 38839
0 38841 7 1 2 38836 38840
0 38842 5 1 1 38841
0 38843 7 1 2 65464 38842
0 38844 5 1 1 38843
0 38845 7 2 2 94863 84036
0 38846 5 1 1 104556
0 38847 7 1 2 103561 104557
0 38848 5 1 1 38847
0 38849 7 1 2 97906 82122
0 38850 5 1 1 38849
0 38851 7 1 2 70846 104455
0 38852 5 1 1 38851
0 38853 7 1 2 38850 38852
0 38854 5 1 1 38853
0 38855 7 1 2 80634 38854
0 38856 5 1 1 38855
0 38857 7 1 2 38848 38856
0 38858 7 1 2 38844 38857
0 38859 7 1 2 38834 38858
0 38860 5 1 1 38859
0 38861 7 1 2 104540 38860
0 38862 5 1 1 38861
0 38863 7 2 2 77375 102764
0 38864 5 1 1 104558
0 38865 7 1 2 74794 104559
0 38866 5 1 1 38865
0 38867 7 1 2 98385 104541
0 38868 7 1 2 81512 38867
0 38869 5 1 1 38868
0 38870 7 1 2 38866 38869
0 38871 5 1 1 38870
0 38872 7 1 2 81897 38871
0 38873 5 1 1 38872
0 38874 7 1 2 69225 38873
0 38875 7 1 2 38862 38874
0 38876 7 1 2 38819 38875
0 38877 5 1 1 38876
0 38878 7 1 2 38797 38877
0 38879 5 1 1 38878
0 38880 7 1 2 72720 38879
0 38881 5 1 1 38880
0 38882 7 1 2 78230 38881
0 38883 7 1 2 38766 38882
0 38884 5 1 1 38883
0 38885 7 1 2 38660 38884
0 38886 5 1 1 38885
0 38887 7 1 2 76333 38886
0 38888 5 1 1 38887
0 38889 7 4 2 77693 85812
0 38890 7 2 2 85146 104560
0 38891 5 1 1 104564
0 38892 7 1 2 38891 96067
0 38893 5 1 1 38892
0 38894 7 1 2 77376 38893
0 38895 5 1 1 38894
0 38896 7 1 2 78047 78231
0 38897 7 1 2 94361 38896
0 38898 5 1 1 38897
0 38899 7 1 2 38895 38898
0 38900 5 1 1 38899
0 38901 7 1 2 102735 38900
0 38902 5 1 1 38901
0 38903 7 1 2 98961 103825
0 38904 5 1 1 38903
0 38905 7 2 2 86390 85105
0 38906 7 1 2 90227 104566
0 38907 5 1 1 38906
0 38908 7 1 2 38904 38907
0 38909 5 2 1 38908
0 38910 7 1 2 81898 104568
0 38911 5 1 1 38910
0 38912 7 1 2 85698 78232
0 38913 5 2 1 38912
0 38914 7 1 2 85147 20736
0 38915 7 1 2 97945 38914
0 38916 5 1 1 38915
0 38917 7 1 2 104570 38916
0 38918 5 1 1 38917
0 38919 7 1 2 77178 38918
0 38920 5 1 1 38919
0 38921 7 1 2 38911 38920
0 38922 5 1 1 38921
0 38923 7 1 2 97907 38922
0 38924 5 1 1 38923
0 38925 7 6 2 68453 81043
0 38926 7 1 2 82029 104572
0 38927 5 1 1 38926
0 38928 7 1 2 77179 91088
0 38929 5 1 1 38928
0 38930 7 1 2 38927 38929
0 38931 5 1 1 38930
0 38932 7 1 2 72437 38931
0 38933 5 1 1 38932
0 38934 7 1 2 89914 98590
0 38935 5 2 1 38934
0 38936 7 1 2 38933 104578
0 38937 5 1 1 38936
0 38938 7 1 2 80635 38937
0 38939 5 1 1 38938
0 38940 7 2 2 87053 98591
0 38941 7 1 2 78579 104580
0 38942 5 1 1 38941
0 38943 7 1 2 98288 87684
0 38944 5 1 1 38943
0 38945 7 1 2 38942 38944
0 38946 5 1 1 38945
0 38947 7 1 2 80721 38946
0 38948 5 1 1 38947
0 38949 7 1 2 98274 104561
0 38950 5 1 1 38949
0 38951 7 1 2 76162 102129
0 38952 7 1 2 104403 38951
0 38953 5 1 1 38952
0 38954 7 1 2 38950 38953
0 38955 7 1 2 38948 38954
0 38956 7 1 2 38939 38955
0 38957 5 1 1 38956
0 38958 7 1 2 85148 38957
0 38959 5 1 1 38958
0 38960 7 2 2 68108 76622
0 38961 7 1 2 103278 78233
0 38962 7 1 2 104582 38961
0 38963 5 1 1 38962
0 38964 7 2 2 99714 79109
0 38965 7 1 2 79733 79520
0 38966 7 1 2 104584 38965
0 38967 5 1 1 38966
0 38968 7 1 2 38963 38967
0 38969 5 1 1 38968
0 38970 7 1 2 81899 38969
0 38971 5 1 1 38970
0 38972 7 1 2 85699 98259
0 38973 5 1 1 38972
0 38974 7 2 2 88420 78048
0 38975 5 1 1 104586
0 38976 7 1 2 98178 104587
0 38977 5 1 1 38976
0 38978 7 1 2 38973 38977
0 38979 5 1 1 38978
0 38980 7 1 2 78234 38979
0 38981 5 1 1 38980
0 38982 7 1 2 38971 38981
0 38983 7 1 2 38959 38982
0 38984 5 1 1 38983
0 38985 7 1 2 70847 38984
0 38986 5 1 1 38985
0 38987 7 1 2 38924 38986
0 38988 5 1 1 38987
0 38989 7 1 2 102686 38988
0 38990 5 1 1 38989
0 38991 7 1 2 38902 38990
0 38992 5 1 1 38991
0 38993 7 1 2 69226 38992
0 38994 5 1 1 38993
0 38995 7 1 2 87249 97601
0 38996 5 3 1 38995
0 38997 7 1 2 101779 104588
0 38998 5 1 1 38997
0 38999 7 1 2 102758 91009
0 39000 7 1 2 38998 38999
0 39001 5 1 1 39000
0 39002 7 3 2 65839 92129
0 39003 7 1 2 68874 100154
0 39004 7 2 2 104591 39003
0 39005 7 1 2 98376 104594
0 39006 7 1 2 101766 39005
0 39007 5 1 1 39006
0 39008 7 1 2 39001 39007
0 39009 5 1 1 39008
0 39010 7 1 2 64172 39009
0 39011 5 1 1 39010
0 39012 7 2 2 102800 91010
0 39013 7 1 2 94190 94880
0 39014 5 1 1 39013
0 39015 7 1 2 97908 39014
0 39016 5 1 1 39015
0 39017 7 1 2 84340 99029
0 39018 7 1 2 87616 39017
0 39019 5 1 1 39018
0 39020 7 1 2 39016 39019
0 39021 5 1 1 39020
0 39022 7 1 2 104596 39021
0 39023 5 1 1 39022
0 39024 7 1 2 39011 39023
0 39025 5 1 1 39024
0 39026 7 1 2 68109 39025
0 39027 5 1 1 39026
0 39028 7 2 2 99408 102687
0 39029 7 1 2 74556 104598
0 39030 5 1 1 39029
0 39031 7 1 2 68687 83029
0 39032 7 1 2 102780 39031
0 39033 5 1 1 39032
0 39034 7 1 2 39030 39033
0 39035 5 1 1 39034
0 39036 7 1 2 74795 95854
0 39037 7 1 2 39035 39036
0 39038 5 1 1 39037
0 39039 7 1 2 39027 39038
0 39040 5 1 1 39039
0 39041 7 1 2 77470 39040
0 39042 5 1 1 39041
0 39043 7 2 2 74683 77266
0 39044 7 1 2 85637 95054
0 39045 5 1 1 39044
0 39046 7 1 2 104600 39045
0 39047 5 1 1 39046
0 39048 7 1 2 85746 96071
0 39049 5 1 1 39048
0 39050 7 1 2 39047 39049
0 39051 5 1 1 39050
0 39052 7 1 2 73205 39051
0 39053 5 1 1 39052
0 39054 7 1 2 86686 77377
0 39055 5 1 1 39054
0 39056 7 1 2 39053 39055
0 39057 5 1 1 39056
0 39058 7 1 2 102653 39057
0 39059 5 1 1 39058
0 39060 7 4 2 70848 104542
0 39061 5 1 1 104602
0 39062 7 1 2 85700 104603
0 39063 5 1 1 39062
0 39064 7 1 2 39059 39063
0 39065 5 1 1 39064
0 39066 7 1 2 78235 39065
0 39067 5 1 1 39066
0 39068 7 4 2 67125 103065
0 39069 7 2 2 90070 96107
0 39070 7 1 2 104606 104610
0 39071 5 1 1 39070
0 39072 7 1 2 102609 104569
0 39073 5 1 1 39072
0 39074 7 1 2 39071 39073
0 39075 5 1 1 39074
0 39076 7 1 2 81900 39075
0 39077 5 1 1 39076
0 39078 7 2 2 73773 95888
0 39079 7 1 2 104604 104612
0 39080 5 1 1 39079
0 39081 7 1 2 87281 104040
0 39082 7 1 2 92036 39081
0 39083 5 1 1 39082
0 39084 7 1 2 39080 39083
0 39085 5 1 1 39084
0 39086 7 1 2 73542 39085
0 39087 5 1 1 39086
0 39088 7 2 2 66043 102627
0 39089 7 1 2 95525 104614
0 39090 5 1 1 39089
0 39091 7 1 2 39061 39090
0 39092 5 1 1 39091
0 39093 7 1 2 104562 39092
0 39094 5 1 1 39093
0 39095 7 5 2 71123 72170
0 39096 7 2 2 102353 104616
0 39097 7 1 2 102134 96725
0 39098 7 1 2 104621 39097
0 39099 5 1 1 39098
0 39100 7 1 2 39094 39099
0 39101 7 1 2 39087 39100
0 39102 5 1 1 39101
0 39103 7 1 2 85149 39102
0 39104 5 1 1 39103
0 39105 7 1 2 39077 39104
0 39106 7 1 2 39067 39105
0 39107 5 1 1 39106
0 39108 7 1 2 67368 39107
0 39109 5 1 1 39108
0 39110 7 1 2 97883 104565
0 39111 5 1 1 39110
0 39112 7 1 2 77471 38975
0 39113 5 1 1 39112
0 39114 7 1 2 70849 96065
0 39115 7 1 2 39113 39114
0 39116 5 1 1 39115
0 39117 7 1 2 39111 39116
0 39118 5 1 1 39117
0 39119 7 1 2 103356 39118
0 39120 5 1 1 39119
0 39121 7 1 2 39109 39120
0 39122 5 1 1 39121
0 39123 7 1 2 64173 39122
0 39124 5 1 1 39123
0 39125 7 1 2 78236 104599
0 39126 5 1 1 39125
0 39127 7 3 2 100155 97476
0 39128 7 1 2 74405 85106
0 39129 7 1 2 96803 39128
0 39130 7 1 2 104623 39129
0 39131 5 1 1 39130
0 39132 7 1 2 39126 39131
0 39133 5 1 1 39132
0 39134 7 1 2 104583 39133
0 39135 5 1 1 39134
0 39136 7 1 2 96960 103050
0 39137 7 1 2 97864 39136
0 39138 7 4 2 73206 74102
0 39139 7 1 2 104417 104626
0 39140 7 1 2 39137 39139
0 39141 5 1 1 39140
0 39142 7 1 2 39135 39141
0 39143 5 1 1 39142
0 39144 7 1 2 73774 39143
0 39145 5 1 1 39144
0 39146 7 1 2 93709 102708
0 39147 7 2 2 72438 79734
0 39148 7 1 2 92497 104630
0 39149 7 1 2 39146 39148
0 39150 5 1 1 39149
0 39151 7 1 2 39145 39150
0 39152 5 1 1 39151
0 39153 7 1 2 84845 39152
0 39154 5 1 1 39153
0 39155 7 1 2 39124 39154
0 39156 7 1 2 39042 39155
0 39157 7 1 2 38994 39156
0 39158 5 1 1 39157
0 39159 7 1 2 90812 39158
0 39160 5 1 1 39159
0 39161 7 1 2 64828 80422
0 39162 5 3 1 39161
0 39163 7 1 2 86230 104632
0 39164 5 1 1 39163
0 39165 7 1 2 77613 39164
0 39166 5 1 1 39165
0 39167 7 1 2 77675 83583
0 39168 5 1 1 39167
0 39169 7 1 2 39166 39168
0 39170 5 1 1 39169
0 39171 7 1 2 82200 39170
0 39172 5 1 1 39171
0 39173 7 1 2 100474 104343
0 39174 5 1 1 39173
0 39175 7 1 2 39172 39174
0 39176 5 1 1 39175
0 39177 7 1 2 70227 39176
0 39178 5 1 1 39177
0 39179 7 1 2 67706 93509
0 39180 7 1 2 103504 39179
0 39181 5 1 1 39180
0 39182 7 1 2 39178 39181
0 39183 5 1 1 39182
0 39184 7 1 2 78237 39183
0 39185 5 1 1 39184
0 39186 7 1 2 80083 95270
0 39187 7 1 2 94398 39186
0 39188 7 1 2 91973 39187
0 39189 5 1 1 39188
0 39190 7 1 2 39185 39189
0 39191 5 1 1 39190
0 39192 7 1 2 100112 39191
0 39193 5 1 1 39192
0 39194 7 1 2 29051 104268
0 39195 5 4 1 39194
0 39196 7 1 2 104420 104635
0 39197 5 1 1 39196
0 39198 7 1 2 78175 99273
0 39199 7 1 2 90509 39198
0 39200 7 1 2 101365 39199
0 39201 5 1 1 39200
0 39202 7 1 2 39197 39201
0 39203 5 1 1 39202
0 39204 7 1 2 84743 39203
0 39205 5 1 1 39204
0 39206 7 1 2 72721 95431
0 39207 5 1 1 39206
0 39208 7 5 2 67707 78580
0 39209 7 1 2 92165 104639
0 39210 5 1 1 39209
0 39211 7 1 2 39207 39210
0 39212 5 1 1 39211
0 39213 7 1 2 66763 98032
0 39214 7 1 2 39212 39213
0 39215 5 1 1 39214
0 39216 7 1 2 82030 82172
0 39217 5 1 1 39216
0 39218 7 1 2 101669 39217
0 39219 5 1 1 39218
0 39220 7 1 2 66356 97052
0 39221 7 1 2 39219 39220
0 39222 5 1 1 39221
0 39223 7 1 2 39215 39222
0 39224 5 1 1 39223
0 39225 7 1 2 91011 39224
0 39226 5 1 1 39225
0 39227 7 1 2 39205 39226
0 39228 5 1 1 39227
0 39229 7 1 2 65465 39228
0 39230 5 1 1 39229
0 39231 7 1 2 39193 39230
0 39232 5 1 1 39231
0 39233 7 1 2 102654 39232
0 39234 5 1 1 39233
0 39235 7 2 2 70228 100380
0 39236 7 1 2 102688 97203
0 39237 7 1 2 91012 39236
0 39238 7 1 2 104644 39237
0 39239 7 1 2 87362 92201
0 39240 7 1 2 39238 39239
0 39241 5 1 1 39240
0 39242 7 1 2 39234 39241
0 39243 5 1 1 39242
0 39244 7 1 2 64174 39243
0 39245 5 1 1 39244
0 39246 7 1 2 94489 96677
0 39247 5 1 1 39246
0 39248 7 1 2 39247 84011
0 39249 5 1 1 39248
0 39250 7 1 2 80636 81376
0 39251 5 1 1 39250
0 39252 7 1 2 71686 104613
0 39253 5 1 1 39252
0 39254 7 1 2 39251 39253
0 39255 5 1 1 39254
0 39256 7 1 2 84102 39255
0 39257 5 1 1 39256
0 39258 7 1 2 39249 39257
0 39259 5 1 1 39258
0 39260 7 1 2 70229 39259
0 39261 5 1 1 39260
0 39262 7 1 2 90842 104337
0 39263 5 1 1 39262
0 39264 7 1 2 81377 84012
0 39265 5 1 1 39264
0 39266 7 1 2 101422 92668
0 39267 5 1 1 39266
0 39268 7 1 2 39265 39267
0 39269 5 1 1 39268
0 39270 7 1 2 80637 39269
0 39271 5 1 1 39270
0 39272 7 1 2 39263 39271
0 39273 7 1 2 39261 39272
0 39274 5 1 1 39273
0 39275 7 1 2 98439 39274
0 39276 5 1 1 39275
0 39277 7 1 2 80855 84103
0 39278 7 1 2 102470 39277
0 39279 7 1 2 87363 39278
0 39280 5 1 1 39279
0 39281 7 1 2 39276 39280
0 39282 5 1 1 39281
0 39283 7 1 2 104597 39282
0 39284 5 1 1 39283
0 39285 7 1 2 39245 39284
0 39286 5 1 1 39285
0 39287 7 1 2 77472 39286
0 39288 5 1 1 39287
0 39289 7 1 2 21946 104373
0 39290 5 2 1 39289
0 39291 7 1 2 71124 94362
0 39292 5 1 1 39291
0 39293 7 1 2 97504 39292
0 39294 5 1 1 39293
0 39295 7 1 2 89776 39294
0 39296 5 1 1 39295
0 39297 7 1 2 98303 101703
0 39298 5 1 1 39297
0 39299 7 1 2 94313 100801
0 39300 5 1 1 39299
0 39301 7 1 2 39298 39300
0 39302 5 1 1 39301
0 39303 7 1 2 68110 39302
0 39304 5 1 1 39303
0 39305 7 1 2 81044 104563
0 39306 5 1 1 39305
0 39307 7 1 2 39304 39306
0 39308 5 1 1 39307
0 39309 7 1 2 85150 39308
0 39310 5 1 1 39309
0 39311 7 1 2 39296 39310
0 39312 5 1 1 39311
0 39313 7 1 2 102736 39312
0 39314 5 1 1 39313
0 39315 7 2 2 66764 77311
0 39316 7 1 2 77976 104648
0 39317 5 1 1 39316
0 39318 7 1 2 99805 39317
0 39319 5 1 1 39318
0 39320 7 1 2 68454 39319
0 39321 5 1 1 39320
0 39322 7 1 2 82854 93779
0 39323 5 1 1 39322
0 39324 7 1 2 66044 39323
0 39325 5 1 1 39324
0 39326 7 2 2 39321 39325
0 39327 5 1 1 104650
0 39328 7 1 2 68111 39327
0 39329 5 1 1 39328
0 39330 7 1 2 99843 82686
0 39331 5 1 1 39330
0 39332 7 1 2 68455 39331
0 39333 5 1 1 39332
0 39334 7 1 2 81119 39333
0 39335 5 2 1 39334
0 39336 7 1 2 68112 104652
0 39337 5 1 1 39336
0 39338 7 1 2 99845 39337
0 39339 5 1 1 39338
0 39340 7 1 2 81901 39339
0 39341 5 1 1 39340
0 39342 7 1 2 77876 87998
0 39343 5 1 1 39342
0 39344 7 1 2 81008 39343
0 39345 5 1 1 39344
0 39346 7 1 2 85701 39345
0 39347 5 1 1 39346
0 39348 7 1 2 88414 92871
0 39349 5 1 1 39348
0 39350 7 1 2 97505 39349
0 39351 5 1 1 39350
0 39352 7 1 2 73207 39351
0 39353 5 1 1 39352
0 39354 7 1 2 39347 39353
0 39355 7 1 2 39341 39354
0 39356 7 1 2 39329 39355
0 39357 5 1 1 39356
0 39358 7 1 2 78238 39357
0 39359 5 1 1 39358
0 39360 7 1 2 88406 83376
0 39361 5 1 1 39360
0 39362 7 1 2 104425 97946
0 39363 7 1 2 39361 39362
0 39364 5 1 1 39363
0 39365 7 1 2 39359 39364
0 39366 5 1 1 39365
0 39367 7 1 2 102759 39366
0 39368 5 1 1 39367
0 39369 7 1 2 39314 39368
0 39370 5 1 1 39369
0 39371 7 1 2 104646 39370
0 39372 5 1 1 39371
0 39373 7 1 2 81618 101932
0 39374 5 1 1 39373
0 39375 7 1 2 69933 103880
0 39376 7 1 2 39374 39375
0 39377 5 1 1 39376
0 39378 7 1 2 21573 39377
0 39379 5 1 1 39378
0 39380 7 1 2 104462 39379
0 39381 5 1 1 39380
0 39382 7 1 2 103348 104640
0 39383 7 1 2 104585 39382
0 39384 5 1 1 39383
0 39385 7 1 2 39381 39384
0 39386 5 1 1 39385
0 39387 7 1 2 64175 39386
0 39388 5 1 1 39387
0 39389 7 1 2 78786 95012
0 39390 5 1 1 39389
0 39391 7 1 2 72439 74194
0 39392 7 1 2 91503 39391
0 39393 7 1 2 90071 39392
0 39394 7 1 2 39390 39393
0 39395 5 1 1 39394
0 39396 7 1 2 39388 39395
0 39397 5 1 1 39396
0 39398 7 1 2 66045 39397
0 39399 5 1 1 39398
0 39400 7 1 2 93046 101602
0 39401 7 1 2 89597 39400
0 39402 7 1 2 104636 39401
0 39403 5 1 1 39402
0 39404 7 1 2 39399 39403
0 39405 5 1 1 39404
0 39406 7 1 2 102655 39405
0 39407 5 1 1 39406
0 39408 7 2 2 93710 97197
0 39409 7 1 2 98668 104654
0 39410 7 1 2 81088 39409
0 39411 5 1 1 39410
0 39412 7 1 2 64176 76689
0 39413 7 1 2 80124 98552
0 39414 7 1 2 39412 39413
0 39415 7 1 2 91013 39414
0 39416 5 1 1 39415
0 39417 7 1 2 39411 39416
0 39418 5 1 1 39417
0 39419 7 4 2 71446 87803
0 39420 7 1 2 102709 104656
0 39421 7 1 2 39418 39420
0 39422 5 1 1 39421
0 39423 7 1 2 39407 39422
0 39424 5 1 1 39423
0 39425 7 1 2 84846 39424
0 39426 5 1 1 39425
0 39427 7 1 2 39372 39426
0 39428 7 1 2 39288 39427
0 39429 7 1 2 39160 39428
0 39430 7 1 2 38888 39429
0 39431 7 1 2 38502 39430
0 39432 7 1 2 102803 99120
0 39433 7 2 2 78913 39432
0 39434 7 1 2 95592 104660
0 39435 5 1 1 39434
0 39436 7 1 2 92757 78239
0 39437 5 1 1 39436
0 39438 7 2 2 91072 81400
0 39439 7 1 2 68875 87927
0 39440 7 1 2 104662 39439
0 39441 5 1 1 39440
0 39442 7 1 2 39437 39441
0 39443 5 1 1 39442
0 39444 7 1 2 64829 39443
0 39445 5 1 1 39444
0 39446 7 5 2 78176 84373
0 39447 7 1 2 76119 104664
0 39448 5 1 1 39447
0 39449 7 1 2 39445 39448
0 39450 5 1 1 39449
0 39451 7 1 2 73775 99640
0 39452 7 1 2 39450 39451
0 39453 5 1 1 39452
0 39454 7 1 2 39435 39453
0 39455 5 1 1 39454
0 39456 7 1 2 102628 39455
0 39457 5 1 1 39456
0 39458 7 2 2 104026 77775
0 39459 7 1 2 100578 92600
0 39460 7 1 2 103291 39459
0 39461 7 1 2 104669 39460
0 39462 5 1 1 39461
0 39463 7 1 2 39457 39462
0 39464 5 1 1 39463
0 39465 7 1 2 65167 39464
0 39466 5 1 1 39465
0 39467 7 1 2 77806 82777
0 39468 7 1 2 101585 39467
0 39469 7 2 2 76163 92353
0 39470 7 1 2 104624 104671
0 39471 7 1 2 39468 39470
0 39472 5 1 1 39471
0 39473 7 1 2 39466 39472
0 39474 5 1 1 39473
0 39475 7 1 2 66583 39474
0 39476 5 1 1 39475
0 39477 7 2 2 98139 102629
0 39478 7 3 2 78177 85019
0 39479 7 1 2 86294 104675
0 39480 7 1 2 104673 39479
0 39481 7 1 2 100908 39480
0 39482 5 1 1 39481
0 39483 7 1 2 39476 39482
0 39484 5 1 1 39483
0 39485 7 1 2 84847 39484
0 39486 5 1 1 39485
0 39487 7 1 2 83905 102630
0 39488 7 1 2 80218 39487
0 39489 7 1 2 104637 39488
0 39490 5 1 1 39489
0 39491 7 1 2 103056 97850
0 39492 7 1 2 102869 39491
0 39493 5 1 1 39492
0 39494 7 1 2 39490 39493
0 39495 5 1 1 39494
0 39496 7 1 2 74684 39495
0 39497 5 1 1 39496
0 39498 7 1 2 73208 103684
0 39499 5 1 1 39498
0 39500 7 1 2 104487 39499
0 39501 5 1 1 39500
0 39502 7 1 2 64177 39501
0 39503 5 1 1 39502
0 39504 7 1 2 78744 98652
0 39505 5 1 1 39504
0 39506 7 1 2 39503 39505
0 39507 5 1 1 39506
0 39508 7 1 2 66765 39507
0 39509 5 1 1 39508
0 39510 7 1 2 76788 97698
0 39511 5 1 1 39510
0 39512 7 1 2 39509 39511
0 39513 5 1 1 39512
0 39514 7 1 2 71447 39513
0 39515 5 1 1 39514
0 39516 7 1 2 74858 78905
0 39517 7 1 2 97699 39516
0 39518 5 1 1 39517
0 39519 7 1 2 39515 39518
0 39520 5 1 1 39519
0 39521 7 1 2 65466 39520
0 39522 5 1 1 39521
0 39523 7 1 2 97909 80210
0 39524 7 1 2 84122 39523
0 39525 7 1 2 78914 39524
0 39526 5 1 1 39525
0 39527 7 1 2 39522 39526
0 39528 5 1 1 39527
0 39529 7 1 2 72722 39528
0 39530 5 1 1 39529
0 39531 7 1 2 96961 74881
0 39532 5 1 1 39531
0 39533 7 3 2 72440 80722
0 39534 7 1 2 69227 104678
0 39535 5 1 1 39534
0 39536 7 1 2 39532 39535
0 39537 5 1 1 39536
0 39538 7 1 2 73209 39537
0 39539 5 1 1 39538
0 39540 7 5 2 73543 96918
0 39541 7 1 2 86769 104681
0 39542 5 1 1 39541
0 39543 7 1 2 39539 39542
0 39544 5 1 1 39543
0 39545 7 1 2 76234 39544
0 39546 5 1 1 39545
0 39547 7 2 2 66766 76601
0 39548 5 1 1 104686
0 39549 7 2 2 77676 104687
0 39550 7 1 2 101982 104688
0 39551 5 1 1 39550
0 39552 7 1 2 39546 39551
0 39553 5 1 1 39552
0 39554 7 1 2 82551 39553
0 39555 5 1 1 39554
0 39556 7 1 2 39530 39555
0 39557 5 1 1 39556
0 39558 7 1 2 102631 39557
0 39559 5 1 1 39558
0 39560 7 2 2 72723 74859
0 39561 7 1 2 100639 104690
0 39562 5 1 1 39561
0 39563 7 1 2 88407 92719
0 39564 5 1 1 39563
0 39565 7 1 2 39562 39564
0 39566 5 1 1 39565
0 39567 7 1 2 82455 102719
0 39568 7 1 2 39566 39567
0 39569 5 1 1 39568
0 39570 7 1 2 39559 39569
0 39571 5 1 1 39570
0 39572 7 1 2 75289 39571
0 39573 5 1 1 39572
0 39574 7 1 2 39497 39573
0 39575 5 1 1 39574
0 39576 7 1 2 78240 39575
0 39577 5 1 1 39576
0 39578 7 1 2 39486 39577
0 39579 5 1 1 39578
0 39580 7 1 2 77267 39579
0 39581 5 1 1 39580
0 39582 7 2 2 98179 100947
0 39583 7 1 2 102204 104692
0 39584 5 1 1 39583
0 39585 7 1 2 98188 104426
0 39586 5 1 1 39585
0 39587 7 1 2 39584 39586
0 39588 5 1 1 39587
0 39589 7 1 2 85532 39588
0 39590 5 1 1 39589
0 39591 7 1 2 92367 95593
0 39592 7 1 2 104693 39591
0 39593 5 1 1 39592
0 39594 7 1 2 39590 39593
0 39595 5 1 1 39594
0 39596 7 1 2 65467 39595
0 39597 5 1 1 39596
0 39598 7 2 2 100909 81045
0 39599 7 1 2 99030 85151
0 39600 7 1 2 104694 39599
0 39601 5 1 1 39600
0 39602 7 1 2 39597 39601
0 39603 5 1 1 39602
0 39604 7 1 2 73776 39603
0 39605 5 1 1 39604
0 39606 7 1 2 99559 92571
0 39607 5 1 1 39606
0 39608 7 1 2 99602 91740
0 39609 5 1 1 39608
0 39610 7 1 2 39607 39609
0 39611 5 1 1 39610
0 39612 7 1 2 72441 104427
0 39613 7 1 2 39611 39612
0 39614 5 1 1 39613
0 39615 7 1 2 39605 39614
0 39616 5 1 1 39615
0 39617 7 1 2 72267 39616
0 39618 5 1 1 39617
0 39619 7 1 2 100425 80320
0 39620 7 1 2 100948 39619
0 39621 7 1 2 101359 104348
0 39622 7 1 2 39620 39621
0 39623 5 1 1 39622
0 39624 7 1 2 39618 39623
0 39625 5 1 1 39624
0 39626 7 1 2 67126 39625
0 39627 5 1 1 39626
0 39628 7 2 2 77523 90233
0 39629 7 1 2 78581 104696
0 39630 5 1 1 39629
0 39631 7 1 2 68688 82605
0 39632 5 1 1 39631
0 39633 7 1 2 86144 39632
0 39634 5 1 1 39633
0 39635 7 1 2 70490 39634
0 39636 5 1 1 39635
0 39637 7 1 2 80543 82123
0 39638 5 2 1 39637
0 39639 7 1 2 39636 104698
0 39640 5 1 1 39639
0 39641 7 1 2 81046 39640
0 39642 5 1 1 39641
0 39643 7 1 2 39630 39642
0 39644 5 1 1 39643
0 39645 7 1 2 93711 74250
0 39646 7 1 2 102415 39645
0 39647 7 1 2 39644 39646
0 39648 5 1 1 39647
0 39649 7 1 2 39627 39648
0 39650 5 1 1 39649
0 39651 7 1 2 73210 39650
0 39652 5 1 1 39651
0 39653 7 2 2 102231 102858
0 39654 5 1 1 104700
0 39655 7 1 2 102419 94501
0 39656 5 1 1 39655
0 39657 7 1 2 39654 39656
0 39658 5 1 1 39657
0 39659 7 5 2 73544 81047
0 39660 7 1 2 75148 93712
0 39661 7 1 2 78351 39660
0 39662 7 1 2 104702 39661
0 39663 7 1 2 39658 39662
0 39664 5 1 1 39663
0 39665 7 1 2 72724 39664
0 39666 7 1 2 39652 39665
0 39667 5 1 1 39666
0 39668 7 2 2 77378 102859
0 39669 5 1 1 104707
0 39670 7 1 2 86906 104708
0 39671 5 1 1 39670
0 39672 7 1 2 102720 80914
0 39673 5 1 1 39672
0 39674 7 1 2 39671 39673
0 39675 5 1 1 39674
0 39676 7 1 2 73545 39675
0 39677 5 1 1 39676
0 39678 7 1 2 86026 77180
0 39679 7 1 2 102371 102721
0 39680 7 1 2 39678 39679
0 39681 5 1 1 39680
0 39682 7 1 2 39677 39681
0 39683 5 1 1 39682
0 39684 7 1 2 85533 39683
0 39685 5 1 1 39684
0 39686 7 2 2 72442 95339
0 39687 7 4 2 67216 73777
0 39688 7 1 2 104533 104711
0 39689 7 1 2 104709 39688
0 39690 5 1 1 39689
0 39691 7 1 2 38864 39690
0 39692 5 1 1 39691
0 39693 7 1 2 69228 39692
0 39694 5 1 1 39693
0 39695 7 2 2 98236 102632
0 39696 7 1 2 93511 104715
0 39697 5 1 1 39696
0 39698 7 1 2 39694 39697
0 39699 5 1 1 39698
0 39700 7 1 2 66767 39699
0 39701 5 1 1 39700
0 39702 7 1 2 78301 102771
0 39703 5 1 1 39702
0 39704 7 1 2 39701 39703
0 39705 5 1 1 39704
0 39706 7 1 2 68456 39705
0 39707 5 1 1 39706
0 39708 7 1 2 73778 99633
0 39709 7 1 2 89757 39708
0 39710 7 1 2 98733 39709
0 39711 5 1 1 39710
0 39712 7 1 2 39707 39711
0 39713 5 1 1 39712
0 39714 7 1 2 65468 39713
0 39715 5 1 1 39714
0 39716 7 1 2 82935 102737
0 39717 5 1 1 39716
0 39718 7 1 2 67369 101445
0 39719 7 1 2 102727 39718
0 39720 5 1 1 39719
0 39721 7 1 2 39717 39720
0 39722 5 1 1 39721
0 39723 7 1 2 70491 39722
0 39724 5 1 1 39723
0 39725 7 1 2 72171 94864
0 39726 7 2 2 99702 39725
0 39727 5 1 1 104717
0 39728 7 1 2 68457 104718
0 39729 5 1 1 39728
0 39730 7 1 2 39724 39729
0 39731 5 1 1 39730
0 39732 7 1 2 101319 39731
0 39733 5 1 1 39732
0 39734 7 1 2 39715 39733
0 39735 5 1 1 39734
0 39736 7 1 2 73211 39735
0 39737 5 1 1 39736
0 39738 7 1 2 39685 39737
0 39739 5 1 1 39738
0 39740 7 1 2 85152 39739
0 39741 5 1 1 39740
0 39742 7 2 2 82606 104712
0 39743 7 1 2 74251 92494
0 39744 7 1 2 93601 39743
0 39745 7 1 2 104719 39744
0 39746 5 1 1 39745
0 39747 7 1 2 76858 104319
0 39748 7 1 2 87110 39747
0 39749 5 1 1 39748
0 39750 7 1 2 39746 39749
0 39751 5 1 1 39750
0 39752 7 1 2 65469 39751
0 39753 5 1 1 39752
0 39754 7 1 2 102372 102633
0 39755 7 1 2 84430 91014
0 39756 7 1 2 39754 39755
0 39757 5 1 1 39756
0 39758 7 1 2 93768 102393
0 39759 7 3 2 79354 39758
0 39760 7 1 2 68689 104721
0 39761 7 1 2 83464 39760
0 39762 5 1 1 39761
0 39763 7 1 2 39757 39762
0 39764 7 1 2 39753 39763
0 39765 5 1 1 39764
0 39766 7 1 2 68113 39765
0 39767 5 1 1 39766
0 39768 7 1 2 98801 83404
0 39769 7 1 2 83461 39768
0 39770 5 1 1 39769
0 39771 7 2 2 102689 103201
0 39772 7 1 2 95637 85153
0 39773 7 1 2 104724 39772
0 39774 7 1 2 39770 39773
0 39775 5 1 1 39774
0 39776 7 1 2 39767 39775
0 39777 5 1 1 39776
0 39778 7 1 2 72443 39777
0 39779 5 1 1 39778
0 39780 7 1 2 85458 78241
0 39781 7 1 2 86984 39780
0 39782 5 1 1 39781
0 39783 7 1 2 85534 85612
0 39784 7 1 2 91105 39783
0 39785 5 1 1 39784
0 39786 7 1 2 39782 39785
0 39787 5 1 1 39786
0 39788 7 1 2 73779 39787
0 39789 5 1 1 39788
0 39790 7 2 2 79982 96172
0 39791 7 3 2 75758 104726
0 39792 7 1 2 97841 104728
0 39793 5 1 1 39792
0 39794 7 1 2 39789 39793
0 39795 5 1 1 39794
0 39796 7 1 2 68114 39795
0 39797 5 1 1 39796
0 39798 7 3 2 81238 90072
0 39799 5 2 1 104731
0 39800 7 1 2 85535 80638
0 39801 7 1 2 104732 39800
0 39802 5 1 1 39801
0 39803 7 1 2 39797 39802
0 39804 5 1 1 39803
0 39805 7 1 2 102772 39804
0 39806 5 1 1 39805
0 39807 7 1 2 39779 39806
0 39808 5 1 1 39807
0 39809 7 1 2 71125 39808
0 39810 5 1 1 39809
0 39811 7 1 2 103059 104725
0 39812 5 1 1 39811
0 39813 7 1 2 78582 104505
0 39814 5 1 1 39813
0 39815 7 1 2 39812 39814
0 39816 5 1 1 39815
0 39817 7 1 2 70492 39816
0 39818 5 1 1 39817
0 39819 7 2 2 102467 94869
0 39820 7 1 2 89396 104736
0 39821 5 1 1 39820
0 39822 7 1 2 86231 102666
0 39823 5 1 1 39822
0 39824 7 1 2 103016 89397
0 39825 5 1 1 39824
0 39826 7 1 2 39823 39825
0 39827 5 1 1 39826
0 39828 7 1 2 87567 39827
0 39829 5 1 1 39828
0 39830 7 1 2 39821 39829
0 39831 5 1 1 39830
0 39832 7 1 2 73546 39831
0 39833 5 1 1 39832
0 39834 7 1 2 39818 39833
0 39835 5 1 1 39834
0 39836 7 1 2 85154 39835
0 39837 5 1 1 39836
0 39838 7 1 2 67217 87655
0 39839 7 1 2 104670 39838
0 39840 5 1 1 39839
0 39841 7 1 2 39837 39840
0 39842 5 1 1 39841
0 39843 7 1 2 67370 39842
0 39844 5 1 1 39843
0 39845 7 1 2 85442 90010
0 39846 7 1 2 78242 39845
0 39847 5 1 1 39846
0 39848 7 1 2 65470 97671
0 39849 7 1 2 104415 39848
0 39850 5 1 1 39849
0 39851 7 1 2 39847 39850
0 39852 5 1 1 39851
0 39853 7 1 2 103357 39852
0 39854 5 1 1 39853
0 39855 7 1 2 39844 39854
0 39856 5 1 1 39855
0 39857 7 1 2 77379 39856
0 39858 5 1 1 39857
0 39859 7 1 2 39810 39858
0 39860 5 1 1 39859
0 39861 7 1 2 66584 39860
0 39862 5 1 1 39861
0 39863 7 1 2 70850 87568
0 39864 7 1 2 104510 39863
0 39865 5 1 1 39864
0 39866 7 1 2 93143 102860
0 39867 5 1 1 39866
0 39868 7 1 2 39727 39867
0 39869 7 1 2 104551 39868
0 39870 7 1 2 39865 39869
0 39871 5 1 1 39870
0 39872 7 1 2 73547 39871
0 39873 5 1 1 39872
0 39874 7 1 2 73212 102765
0 39875 5 1 1 39874
0 39876 7 1 2 73780 104701
0 39877 5 1 1 39876
0 39878 7 1 2 39875 39877
0 39879 7 1 2 39873 39878
0 39880 5 1 1 39879
0 39881 7 3 2 78178 96519
0 39882 7 1 2 98343 104738
0 39883 7 1 2 39880 39882
0 39884 5 1 1 39883
0 39885 7 1 2 67708 39884
0 39886 7 1 2 39862 39885
0 39887 7 1 2 39741 39886
0 39888 5 1 1 39887
0 39889 7 1 2 65168 39888
0 39890 7 1 2 39667 39889
0 39891 5 1 1 39890
0 39892 7 1 2 77285 90073
0 39893 7 1 2 94483 39892
0 39894 5 1 1 39893
0 39895 7 1 2 6304 39894
0 39896 5 1 1 39895
0 39897 7 1 2 101005 39896
0 39898 5 1 1 39897
0 39899 7 1 2 87458 78243
0 39900 5 1 1 39899
0 39901 7 1 2 88730 85155
0 39902 5 1 1 39901
0 39903 7 1 2 39900 39902
0 39904 5 1 1 39903
0 39905 7 1 2 73781 39904
0 39906 5 1 1 39905
0 39907 7 1 2 68115 94271
0 39908 5 1 1 39907
0 39909 7 1 2 78244 39908
0 39910 5 1 1 39909
0 39911 7 1 2 39906 39910
0 39912 5 1 1 39911
0 39913 7 1 2 101320 39912
0 39914 5 1 1 39913
0 39915 7 1 2 39898 39914
0 39916 5 1 1 39915
0 39917 7 1 2 73548 39916
0 39918 5 1 1 39917
0 39919 7 1 2 84911 85156
0 39920 5 1 1 39919
0 39921 7 1 2 91029 39920
0 39922 5 1 1 39921
0 39923 7 1 2 66585 39922
0 39924 5 1 1 39923
0 39925 7 2 2 80723 78245
0 39926 5 4 1 104741
0 39927 7 1 2 39924 104743
0 39928 5 1 1 39927
0 39929 7 1 2 73213 39928
0 39930 5 1 1 39929
0 39931 7 1 2 86770 95935
0 39932 5 1 1 39931
0 39933 7 1 2 39930 39932
0 39934 5 1 1 39933
0 39935 7 1 2 74195 39934
0 39936 5 1 1 39935
0 39937 7 1 2 74130 79056
0 39938 7 1 2 78179 39937
0 39939 7 1 2 85376 39938
0 39940 5 1 1 39939
0 39941 7 1 2 39936 39940
0 39942 5 1 1 39941
0 39943 7 1 2 66046 39942
0 39944 5 1 1 39943
0 39945 7 1 2 39918 39944
0 39946 5 1 1 39945
0 39947 7 1 2 72444 39946
0 39948 5 1 1 39947
0 39949 7 1 2 102236 104357
0 39950 5 1 1 39949
0 39951 7 1 2 39948 39950
0 39952 5 1 1 39951
0 39953 7 1 2 102656 39952
0 39954 5 1 1 39953
0 39955 7 2 2 64448 87125
0 39956 7 1 2 104747 104553
0 39957 5 1 1 39956
0 39958 7 1 2 79983 76623
0 39959 7 1 2 103834 39958
0 39960 5 1 1 39959
0 39961 7 1 2 39957 39960
0 39962 5 1 1 39961
0 39963 7 1 2 91052 39962
0 39964 5 1 1 39963
0 39965 7 1 2 67371 87656
0 39966 7 1 2 96060 39965
0 39967 5 1 1 39966
0 39968 7 1 2 39964 39967
0 39969 5 1 1 39968
0 39970 7 1 2 73214 39969
0 39971 5 1 1 39970
0 39972 7 1 2 77881 38051
0 39973 5 1 1 39972
0 39974 7 1 2 98275 91015
0 39975 7 1 2 39973 39974
0 39976 5 1 1 39975
0 39977 7 1 2 39971 39976
0 39978 5 1 1 39977
0 39979 7 1 2 69229 39978
0 39980 5 1 1 39979
0 39981 7 1 2 77181 93769
0 39982 7 1 2 95443 39981
0 39983 7 1 2 102518 39982
0 39984 5 1 1 39983
0 39985 7 1 2 39980 39984
0 39986 5 1 1 39985
0 39987 7 1 2 102610 39986
0 39988 5 1 1 39987
0 39989 7 1 2 39954 39988
0 39990 5 1 1 39989
0 39991 7 1 2 67709 39990
0 39992 5 1 1 39991
0 39993 7 1 2 103753 91053
0 39994 5 1 1 39993
0 39995 7 1 2 39994 104571
0 39996 5 1 1 39995
0 39997 7 1 2 81048 39996
0 39998 5 1 1 39997
0 39999 7 2 2 77524 79110
0 40000 7 1 2 87159 104749
0 40001 7 1 2 95836 40000
0 40002 5 1 1 40001
0 40003 7 1 2 39998 40002
0 40004 5 1 1 40003
0 40005 7 1 2 102843 40004
0 40006 5 1 1 40005
0 40007 7 1 2 88693 78380
0 40008 5 1 1 40007
0 40009 7 1 2 80423 80993
0 40010 5 1 1 40009
0 40011 7 1 2 40008 40010
0 40012 5 1 1 40011
0 40013 7 1 2 104722 40012
0 40014 5 1 1 40013
0 40015 7 1 2 40006 40014
0 40016 5 1 1 40015
0 40017 7 1 2 97165 40016
0 40018 5 1 1 40017
0 40019 7 1 2 88679 81212
0 40020 5 2 1 40019
0 40021 7 1 2 83676 104751
0 40022 5 1 1 40021
0 40023 7 1 2 40022 104723
0 40024 5 1 1 40023
0 40025 7 3 2 98829 75759
0 40026 7 2 2 104534 104753
0 40027 7 1 2 71847 103017
0 40028 7 1 2 102338 40027
0 40029 7 1 2 104756 40028
0 40030 5 1 1 40029
0 40031 7 1 2 40024 40030
0 40032 5 1 1 40031
0 40033 7 1 2 98407 40032
0 40034 5 1 1 40033
0 40035 7 1 2 64449 85382
0 40036 7 1 2 97987 96175
0 40037 7 1 2 40035 40036
0 40038 5 1 1 40037
0 40039 7 1 2 68876 84136
0 40040 7 1 2 87582 40039
0 40041 5 1 1 40040
0 40042 7 1 2 91030 40041
0 40043 5 1 1 40042
0 40044 7 7 2 73215 81049
0 40045 5 1 1 104758
0 40046 7 1 2 72725 104759
0 40047 7 1 2 40043 40046
0 40048 5 1 1 40047
0 40049 7 1 2 40038 40048
0 40050 5 1 1 40049
0 40051 7 1 2 103358 40050
0 40052 5 1 1 40051
0 40053 7 1 2 77877 102822
0 40054 7 1 2 99066 40053
0 40055 7 1 2 104757 40054
0 40056 5 1 1 40055
0 40057 7 1 2 40052 40056
0 40058 5 1 1 40057
0 40059 7 1 2 73549 40058
0 40060 5 1 1 40059
0 40061 7 3 2 81753 104760
0 40062 5 1 1 104765
0 40063 7 4 2 99634 91242
0 40064 7 1 2 78246 104768
0 40065 7 1 2 104766 40064
0 40066 5 1 1 40065
0 40067 7 1 2 40060 40066
0 40068 5 1 1 40067
0 40069 7 1 2 85536 40068
0 40070 5 1 1 40069
0 40071 7 1 2 40034 40070
0 40072 7 1 2 40018 40071
0 40073 7 1 2 39992 40072
0 40074 7 1 2 39891 40073
0 40075 5 1 1 40074
0 40076 7 1 2 76602 40075
0 40077 5 1 1 40076
0 40078 7 1 2 39581 40077
0 40079 7 1 2 89665 36635
0 40080 5 1 1 40079
0 40081 7 1 2 65169 40080
0 40082 5 1 1 40081
0 40083 7 1 2 40082 656
0 40084 5 1 1 40083
0 40085 7 1 2 96083 40084
0 40086 5 1 1 40085
0 40087 7 2 2 67710 93219
0 40088 5 1 1 104772
0 40089 7 1 2 78745 104773
0 40090 5 1 1 40089
0 40091 7 1 2 40086 40090
0 40092 5 1 1 40091
0 40093 7 1 2 81050 40092
0 40094 5 1 1 40093
0 40095 7 2 2 67711 97884
0 40096 7 1 2 100248 104774
0 40097 5 1 1 40096
0 40098 7 1 2 40094 40097
0 40099 5 1 1 40098
0 40100 7 1 2 69230 40099
0 40101 5 1 1 40100
0 40102 7 1 2 100249 101046
0 40103 5 1 1 40102
0 40104 7 2 2 85537 78510
0 40105 5 1 1 104776
0 40106 7 1 2 74196 93542
0 40107 5 1 1 40106
0 40108 7 1 2 40105 40107
0 40109 5 2 1 40108
0 40110 7 1 2 104778 92173
0 40111 5 1 1 40110
0 40112 7 1 2 83272 83749
0 40113 5 1 1 40112
0 40114 7 1 2 92886 40113
0 40115 5 1 1 40114
0 40116 7 1 2 64178 40115
0 40117 5 1 1 40116
0 40118 7 1 2 40117 10339
0 40119 5 1 1 40118
0 40120 7 1 2 70851 40119
0 40121 5 1 1 40120
0 40122 7 1 2 66357 104777
0 40123 5 1 1 40122
0 40124 7 1 2 40121 40123
0 40125 5 1 1 40124
0 40126 7 1 2 80940 40125
0 40127 5 1 1 40126
0 40128 7 1 2 40111 40127
0 40129 5 1 1 40128
0 40130 7 1 2 68116 40129
0 40131 5 1 1 40130
0 40132 7 1 2 40103 40131
0 40133 7 1 2 40101 40132
0 40134 5 1 1 40133
0 40135 7 1 2 67372 40134
0 40136 5 1 1 40135
0 40137 7 2 2 71448 95614
0 40138 7 2 2 74069 104780
0 40139 7 1 2 80941 97085
0 40140 7 1 2 104782 40139
0 40141 5 1 1 40140
0 40142 7 1 2 40136 40141
0 40143 5 1 1 40142
0 40144 7 1 2 103062 40143
0 40145 5 1 1 40144
0 40146 7 2 2 99265 91243
0 40147 7 1 2 97999 104784
0 40148 5 1 1 40147
0 40149 7 2 2 67373 84184
0 40150 7 1 2 99307 84272
0 40151 7 1 2 104786 40150
0 40152 5 1 1 40151
0 40153 7 1 2 40148 40152
0 40154 5 1 1 40153
0 40155 7 1 2 69231 40154
0 40156 5 1 1 40155
0 40157 7 2 2 74406 97477
0 40158 7 1 2 78459 83863
0 40159 5 1 1 40158
0 40160 7 1 2 67712 95457
0 40161 5 1 1 40160
0 40162 7 1 2 92887 40161
0 40163 7 1 2 40159 40162
0 40164 5 1 1 40163
0 40165 7 1 2 104788 40164
0 40166 5 1 1 40165
0 40167 7 1 2 40156 40166
0 40168 5 1 1 40167
0 40169 7 1 2 80942 40168
0 40170 5 1 1 40169
0 40171 7 1 2 19821 92812
0 40172 5 1 1 40171
0 40173 7 2 2 78447 40172
0 40174 7 1 2 64450 104790
0 40175 5 1 1 40174
0 40176 7 1 2 78127 83750
0 40177 5 1 1 40176
0 40178 7 1 2 40175 40177
0 40179 5 1 1 40178
0 40180 7 1 2 92174 40179
0 40181 5 1 1 40180
0 40182 7 1 2 79562 93488
0 40183 7 1 2 84410 40182
0 40184 7 1 2 104641 40183
0 40185 5 1 1 40184
0 40186 7 1 2 40181 40185
0 40187 5 1 1 40186
0 40188 7 1 2 72445 104525
0 40189 7 1 2 40187 40188
0 40190 5 1 1 40189
0 40191 7 1 2 40170 40190
0 40192 5 1 1 40191
0 40193 7 1 2 68117 40192
0 40194 5 1 1 40193
0 40195 7 3 2 71126 83991
0 40196 5 2 1 104792
0 40197 7 1 2 78448 104795
0 40198 5 5 1 40197
0 40199 7 1 2 92790 37648
0 40200 5 1 1 40199
0 40201 7 2 2 14791 40200
0 40202 7 1 2 64179 104802
0 40203 5 1 1 40202
0 40204 7 1 2 76334 6252
0 40205 5 1 1 40204
0 40206 7 1 2 102218 40205
0 40207 5 1 1 40206
0 40208 7 1 2 40203 40207
0 40209 5 1 1 40208
0 40210 7 1 2 73216 40209
0 40211 5 1 1 40210
0 40212 7 1 2 102219 89486
0 40213 5 1 1 40212
0 40214 7 1 2 40211 40213
0 40215 5 1 1 40214
0 40216 7 1 2 104797 40215
0 40217 5 1 1 40216
0 40218 7 1 2 85459 104793
0 40219 7 1 2 90884 40218
0 40220 5 1 1 40219
0 40221 7 1 2 93443 102051
0 40222 7 1 2 87204 40221
0 40223 5 1 1 40222
0 40224 7 1 2 40220 40223
0 40225 5 1 1 40224
0 40226 7 1 2 73550 40225
0 40227 5 1 1 40226
0 40228 7 2 2 77070 83992
0 40229 5 2 1 104804
0 40230 7 1 2 98815 104806
0 40231 5 2 1 40230
0 40232 7 1 2 64180 104808
0 40233 5 1 1 40232
0 40234 7 1 2 83993 103837
0 40235 5 1 1 40234
0 40236 7 1 2 40233 40235
0 40237 5 2 1 40236
0 40238 7 1 2 83285 104810
0 40239 5 1 1 40238
0 40240 7 1 2 68690 74175
0 40241 7 1 2 93559 93122
0 40242 7 1 2 40240 40241
0 40243 7 1 2 79966 40242
0 40244 5 1 1 40243
0 40245 7 1 2 40239 40244
0 40246 7 1 2 40227 40245
0 40247 5 1 1 40246
0 40248 7 1 2 64451 40247
0 40249 5 1 1 40248
0 40250 7 1 2 69559 100253
0 40251 7 1 2 104811 40250
0 40252 5 1 1 40251
0 40253 7 1 2 40249 40252
0 40254 7 1 2 40217 40253
0 40255 5 1 1 40254
0 40256 7 1 2 72446 40255
0 40257 5 1 1 40256
0 40258 7 1 2 81051 97702
0 40259 7 1 2 100254 40258
0 40260 5 1 1 40259
0 40261 7 1 2 40257 40260
0 40262 5 1 1 40261
0 40263 7 1 2 67127 40262
0 40264 5 1 1 40263
0 40265 7 1 2 40194 40264
0 40266 5 1 1 40265
0 40267 7 1 2 72268 40266
0 40268 5 1 1 40267
0 40269 7 1 2 40145 40268
0 40270 5 1 1 40269
0 40271 7 1 2 85157 40270
0 40272 5 1 1 40271
0 40273 7 1 2 93620 99319
0 40274 7 1 2 85158 104642
0 40275 7 1 2 40273 40274
0 40276 5 1 1 40275
0 40277 7 2 2 65170 87884
0 40278 5 1 1 104812
0 40279 7 1 2 100910 104813
0 40280 7 1 2 89747 40279
0 40281 5 1 1 40280
0 40282 7 1 2 40276 40281
0 40283 5 1 1 40282
0 40284 7 1 2 102784 40283
0 40285 5 1 1 40284
0 40286 7 1 2 71449 67218
0 40287 7 1 2 102747 40286
0 40288 7 1 2 104042 40287
0 40289 7 1 2 91016 93273
0 40290 7 1 2 40288 40289
0 40291 5 1 1 40290
0 40292 7 1 2 40285 40291
0 40293 5 1 1 40292
0 40294 7 1 2 77268 40293
0 40295 5 1 1 40294
0 40296 7 1 2 76235 81116
0 40297 5 1 1 40296
0 40298 7 1 2 71127 77055
0 40299 5 1 1 40298
0 40300 7 1 2 82793 40299
0 40301 7 1 2 100833 40300
0 40302 5 1 1 40301
0 40303 7 1 2 40297 40302
0 40304 5 1 1 40303
0 40305 7 1 2 85443 40304
0 40306 5 1 1 40305
0 40307 7 1 2 80257 78060
0 40308 5 1 1 40307
0 40309 7 1 2 2975 40308
0 40310 5 1 1 40309
0 40311 7 1 2 65840 40310
0 40312 5 1 1 40311
0 40313 7 1 2 95135 77071
0 40314 5 1 1 40313
0 40315 7 1 2 73551 40314
0 40316 7 1 2 40312 40315
0 40317 5 1 1 40316
0 40318 7 1 2 96125 92331
0 40319 5 1 1 40318
0 40320 7 1 2 65171 40319
0 40321 5 1 1 40320
0 40322 7 1 2 76603 97885
0 40323 5 1 1 40322
0 40324 7 2 2 64452 94839
0 40325 7 1 2 77590 104814
0 40326 5 1 1 40325
0 40327 7 1 2 68458 40326
0 40328 7 1 2 40323 40327
0 40329 7 1 2 40321 40328
0 40330 5 1 1 40329
0 40331 7 1 2 64181 40330
0 40332 7 1 2 40317 40331
0 40333 5 1 1 40332
0 40334 7 1 2 40306 40333
0 40335 5 1 1 40334
0 40336 7 1 2 102634 40335
0 40337 5 1 1 40336
0 40338 7 1 2 83017 80281
0 40339 5 1 1 40338
0 40340 7 1 2 66586 76628
0 40341 5 1 1 40340
0 40342 7 1 2 40339 40341
0 40343 5 1 1 40342
0 40344 7 1 2 102844 40343
0 40345 5 1 1 40344
0 40346 7 1 2 40337 40345
0 40347 5 1 1 40346
0 40348 7 1 2 72447 40347
0 40349 5 1 1 40348
0 40350 7 1 2 100122 81507
0 40351 5 1 1 40350
0 40352 7 2 2 70852 68459
0 40353 7 2 2 74685 78291
0 40354 5 1 1 104818
0 40355 7 1 2 76491 40354
0 40356 5 1 1 40355
0 40357 7 1 2 101016 40356
0 40358 5 1 1 40357
0 40359 7 1 2 93621 81052
0 40360 5 1 1 40359
0 40361 7 1 2 40358 40360
0 40362 5 1 1 40361
0 40363 7 1 2 104816 40362
0 40364 5 1 1 40363
0 40365 7 1 2 40351 40364
0 40366 5 1 1 40365
0 40367 7 1 2 102773 40366
0 40368 5 1 1 40367
0 40369 7 1 2 40349 40368
0 40370 5 1 1 40369
0 40371 7 1 2 72726 40370
0 40372 5 1 1 40371
0 40373 7 4 2 64182 67219
0 40374 7 1 2 80253 104820
0 40375 5 1 1 40374
0 40376 7 1 2 76492 100139
0 40377 7 1 2 100763 40376
0 40378 5 1 1 40377
0 40379 7 1 2 40375 40378
0 40380 5 1 1 40379
0 40381 7 1 2 68460 40380
0 40382 5 1 1 40381
0 40383 7 3 2 100165 76941
0 40384 7 1 2 75418 99673
0 40385 7 1 2 104824 40384
0 40386 5 1 1 40385
0 40387 7 1 2 40382 40386
0 40388 5 1 1 40387
0 40389 7 1 2 67374 40388
0 40390 5 1 1 40389
0 40391 7 1 2 100426 81508
0 40392 7 1 2 103267 40391
0 40393 5 1 1 40392
0 40394 7 1 2 40390 40393
0 40395 5 1 1 40394
0 40396 7 1 2 69560 40395
0 40397 5 1 1 40396
0 40398 7 2 2 67375 84527
0 40399 7 1 2 96241 104827
0 40400 5 1 1 40399
0 40401 7 1 2 95136 104682
0 40402 5 1 1 40401
0 40403 7 1 2 40400 40402
0 40404 5 1 1 40403
0 40405 7 1 2 71128 40404
0 40406 5 1 1 40405
0 40407 7 1 2 64183 102804
0 40408 7 1 2 101741 40407
0 40409 5 1 1 40408
0 40410 7 1 2 40406 40409
0 40411 5 1 1 40410
0 40412 7 1 2 67220 40411
0 40413 5 1 1 40412
0 40414 7 1 2 40397 40413
0 40415 5 1 1 40414
0 40416 7 1 2 70853 40415
0 40417 5 1 1 40416
0 40418 7 1 2 100427 93757
0 40419 7 1 2 104783 40418
0 40420 5 1 1 40419
0 40421 7 1 2 40417 40420
0 40422 5 1 1 40421
0 40423 7 1 2 84619 40422
0 40424 5 1 1 40423
0 40425 7 1 2 40372 40424
0 40426 5 1 1 40425
0 40427 7 1 2 68118 40426
0 40428 5 1 1 40427
0 40429 7 1 2 67376 104543
0 40430 5 2 1 40429
0 40431 7 1 2 101281 102861
0 40432 5 1 1 40431
0 40433 7 1 2 104829 40432
0 40434 5 1 1 40433
0 40435 7 1 2 85538 40434
0 40436 5 1 1 40435
0 40437 7 2 2 69232 100134
0 40438 7 2 2 102690 104831
0 40439 5 1 1 104833
0 40440 7 1 2 102673 40439
0 40441 5 1 1 40440
0 40442 7 1 2 72448 80282
0 40443 7 1 2 40441 40442
0 40444 5 1 1 40443
0 40445 7 1 2 40436 40444
0 40446 5 1 1 40445
0 40447 7 1 2 72727 40446
0 40448 5 1 1 40447
0 40449 7 2 2 101138 103268
0 40450 5 1 1 104835
0 40451 7 1 2 102611 104836
0 40452 5 1 1 40451
0 40453 7 1 2 40448 40452
0 40454 5 1 1 40453
0 40455 7 1 2 73217 40454
0 40456 5 1 1 40455
0 40457 7 2 2 65841 100428
0 40458 5 3 1 104837
0 40459 7 3 2 70854 100085
0 40460 5 2 1 104842
0 40461 7 1 2 68691 104843
0 40462 5 1 1 40461
0 40463 7 1 2 104839 40462
0 40464 5 1 1 40463
0 40465 7 2 2 67713 104617
0 40466 7 1 2 104781 104847
0 40467 7 1 2 40464 40466
0 40468 5 1 1 40467
0 40469 7 1 2 40456 40468
0 40470 5 1 1 40469
0 40471 7 1 2 81310 40470
0 40472 5 1 1 40471
0 40473 7 1 2 40428 40472
0 40474 5 1 1 40473
0 40475 7 1 2 78247 40474
0 40476 5 1 1 40475
0 40477 7 1 2 40295 40476
0 40478 7 1 2 40272 40477
0 40479 5 1 1 40478
0 40480 7 1 2 81902 40479
0 40481 5 1 1 40480
0 40482 7 1 2 76164 104665
0 40483 5 1 1 40482
0 40484 7 1 2 83751 91079
0 40485 5 1 1 40484
0 40486 7 1 2 40483 40485
0 40487 5 1 1 40486
0 40488 7 1 2 66768 40487
0 40489 5 1 1 40488
0 40490 7 1 2 78180 96875
0 40491 5 1 1 40490
0 40492 7 1 2 40489 40491
0 40493 5 1 1 40492
0 40494 7 1 2 65471 40493
0 40495 5 1 1 40494
0 40496 7 1 2 80424 87384
0 40497 5 1 1 40496
0 40498 7 1 2 96596 40497
0 40499 5 1 1 40498
0 40500 7 1 2 104666 40499
0 40501 5 1 1 40500
0 40502 7 1 2 40495 40501
0 40503 5 1 1 40502
0 40504 7 1 2 73552 40503
0 40505 5 1 1 40504
0 40506 7 1 2 98977 96159
0 40507 5 1 1 40506
0 40508 7 1 2 40505 40507
0 40509 5 1 1 40508
0 40510 7 1 2 64453 40509
0 40511 5 1 1 40510
0 40512 7 1 2 100465 86647
0 40513 5 1 1 40512
0 40514 7 1 2 87126 82250
0 40515 7 1 2 78248 40514
0 40516 7 1 2 40513 40515
0 40517 5 1 1 40516
0 40518 7 1 2 67377 40517
0 40519 7 1 2 40511 40518
0 40520 5 1 1 40519
0 40521 7 2 2 80125 85159
0 40522 7 1 2 68119 104849
0 40523 5 1 1 40522
0 40524 7 1 2 77473 90655
0 40525 5 1 1 40524
0 40526 7 1 2 40523 40525
0 40527 5 1 1 40526
0 40528 7 1 2 78583 40527
0 40529 5 1 1 40528
0 40530 7 1 2 87999 76789
0 40531 7 1 2 90074 40530
0 40532 5 1 1 40531
0 40533 7 1 2 40529 40532
0 40534 5 1 1 40533
0 40535 7 1 2 66769 40534
0 40536 5 1 1 40535
0 40537 7 1 2 64454 18627
0 40538 5 1 1 40537
0 40539 7 1 2 91017 40538
0 40540 7 1 2 101683 40539
0 40541 5 1 1 40540
0 40542 7 1 2 40536 40541
0 40543 5 1 1 40542
0 40544 7 1 2 71687 40543
0 40545 5 1 1 40544
0 40546 7 1 2 83509 74882
0 40547 5 1 1 40546
0 40548 7 1 2 89777 40547
0 40549 5 1 1 40548
0 40550 7 1 2 88462 90075
0 40551 7 1 2 88784 40550
0 40552 5 1 1 40551
0 40553 7 1 2 40549 40552
0 40554 5 1 1 40553
0 40555 7 1 2 77474 40554
0 40556 5 1 1 40555
0 40557 7 2 2 71129 82357
0 40558 5 1 1 104851
0 40559 7 1 2 70230 80051
0 40560 5 1 1 40559
0 40561 7 1 2 40558 40560
0 40562 5 1 1 40561
0 40563 7 1 2 89778 40562
0 40564 5 1 1 40563
0 40565 7 1 2 40556 40564
0 40566 7 1 2 40545 40565
0 40567 5 1 1 40566
0 40568 7 1 2 65472 40567
0 40569 5 1 1 40568
0 40570 7 1 2 68877 93450
0 40571 7 1 2 101849 40570
0 40572 5 1 1 40571
0 40573 7 1 2 95870 7756
0 40574 5 1 1 40573
0 40575 7 1 2 90004 40574
0 40576 5 1 1 40575
0 40577 7 1 2 7814 40576
0 40578 5 1 1 40577
0 40579 7 1 2 66047 82650
0 40580 7 1 2 40578 40579
0 40581 5 1 1 40580
0 40582 7 1 2 40572 40581
0 40583 5 1 1 40582
0 40584 7 1 2 68120 40583
0 40585 5 1 1 40584
0 40586 7 1 2 103413 91106
0 40587 5 1 1 40586
0 40588 7 1 2 78249 97662
0 40589 5 1 1 40588
0 40590 7 1 2 40587 40589
0 40591 5 1 1 40590
0 40592 7 1 2 85768 40591
0 40593 5 1 1 40592
0 40594 7 1 2 40585 40593
0 40595 7 1 2 40569 40594
0 40596 5 1 1 40595
0 40597 7 1 2 67714 40596
0 40598 5 1 1 40597
0 40599 7 2 2 77475 91018
0 40600 7 2 2 87061 104853
0 40601 5 1 1 104855
0 40602 7 1 2 66048 2556
0 40603 5 2 1 40602
0 40604 7 1 2 91107 104857
0 40605 5 1 1 40604
0 40606 7 1 2 71130 80639
0 40607 7 1 2 98669 91882
0 40608 7 1 2 79682 40607
0 40609 7 1 2 40606 40608
0 40610 5 1 1 40609
0 40611 7 1 2 40605 40610
0 40612 7 1 2 40601 40611
0 40613 5 1 1 40612
0 40614 7 1 2 68461 40613
0 40615 5 1 1 40614
0 40616 7 1 2 81903 75760
0 40617 7 1 2 104441 40616
0 40618 5 1 1 40617
0 40619 7 1 2 40615 40618
0 40620 5 1 1 40619
0 40621 7 1 2 85020 40620
0 40622 5 1 1 40621
0 40623 7 1 2 97967 40622
0 40624 7 1 2 40598 40623
0 40625 5 1 1 40624
0 40626 7 1 2 40520 40625
0 40627 5 1 1 40626
0 40628 7 1 2 82873 76690
0 40629 7 1 2 90076 40628
0 40630 5 1 1 40629
0 40631 7 1 2 95871 40630
0 40632 5 1 1 40631
0 40633 7 1 2 73218 40632
0 40634 5 1 1 40633
0 40635 7 1 2 104418 83227
0 40636 5 1 1 40635
0 40637 7 1 2 40634 40636
0 40638 5 1 1 40637
0 40639 7 1 2 66049 40638
0 40640 5 1 1 40639
0 40641 7 1 2 87987 90077
0 40642 7 1 2 97791 40641
0 40643 5 1 1 40642
0 40644 7 1 2 40640 40643
0 40645 5 1 1 40644
0 40646 7 1 2 96758 40645
0 40647 5 1 1 40646
0 40648 7 1 2 71688 86352
0 40649 7 1 2 104567 40648
0 40650 5 1 1 40649
0 40651 7 1 2 38315 40650
0 40652 5 1 1 40651
0 40653 7 1 2 97177 40652
0 40654 5 1 1 40653
0 40655 7 1 2 40647 40654
0 40656 5 1 1 40655
0 40657 7 1 2 84848 40656
0 40658 5 1 1 40657
0 40659 7 1 2 75419 97527
0 40660 5 1 1 40659
0 40661 7 1 2 26534 40660
0 40662 5 1 1 40661
0 40663 7 1 2 65473 40662
0 40664 5 1 1 40663
0 40665 7 1 2 40664 96856
0 40666 5 1 1 40665
0 40667 7 1 2 78250 40666
0 40668 5 1 1 40667
0 40669 7 1 2 94533 84557
0 40670 5 1 1 40669
0 40671 7 1 2 90222 40670
0 40672 5 1 1 40671
0 40673 7 1 2 81754 40672
0 40674 5 1 1 40673
0 40675 7 2 2 82627 81213
0 40676 5 1 1 104859
0 40677 7 1 2 97797 40676
0 40678 7 1 2 40674 40677
0 40679 5 1 1 40678
0 40680 7 1 2 85160 40679
0 40681 5 1 1 40680
0 40682 7 1 2 40668 40681
0 40683 5 1 1 40682
0 40684 7 1 2 98408 40683
0 40685 5 1 1 40684
0 40686 7 1 2 40658 40685
0 40687 7 1 2 40627 40686
0 40688 5 1 1 40687
0 40689 7 1 2 85807 79120
0 40690 5 1 1 40689
0 40691 7 1 2 73219 11412
0 40692 5 1 1 40691
0 40693 7 1 2 40692 3824
0 40694 5 1 1 40693
0 40695 7 1 2 78251 40694
0 40696 5 1 1 40695
0 40697 7 1 2 40690 40696
0 40698 5 1 1 40697
0 40699 7 1 2 66050 40698
0 40700 5 1 1 40699
0 40701 7 1 2 77269 88422
0 40702 5 1 1 40701
0 40703 7 1 2 66051 94884
0 40704 5 1 1 40703
0 40705 7 1 2 40702 40704
0 40706 5 1 1 40705
0 40707 7 1 2 78252 40706
0 40708 5 1 1 40707
0 40709 7 1 2 80724 104761
0 40710 5 1 1 40709
0 40711 7 1 2 84849 77270
0 40712 7 1 2 92647 40711
0 40713 5 1 1 40712
0 40714 7 1 2 40710 40713
0 40715 5 1 1 40714
0 40716 7 1 2 73782 40715
0 40717 5 1 1 40716
0 40718 7 3 2 65172 83906
0 40719 7 1 2 80321 104861
0 40720 5 1 1 40719
0 40721 7 1 2 40045 40720
0 40722 5 1 1 40721
0 40723 7 1 2 81755 40722
0 40724 5 1 1 40723
0 40725 7 1 2 40717 40724
0 40726 5 1 1 40725
0 40727 7 1 2 85161 40726
0 40728 5 1 1 40727
0 40729 7 1 2 40708 40728
0 40730 5 1 1 40729
0 40731 7 1 2 73553 40730
0 40732 5 1 1 40731
0 40733 7 1 2 89212 84771
0 40734 5 1 1 40733
0 40735 7 1 2 74796 40734
0 40736 5 1 1 40735
0 40737 7 1 2 65474 96891
0 40738 7 1 2 17758 40737
0 40739 5 1 1 40738
0 40740 7 1 2 40736 40739
0 40741 5 1 1 40740
0 40742 7 1 2 104739 40741
0 40743 5 1 1 40742
0 40744 7 1 2 40732 40743
0 40745 7 1 2 40700 40744
0 40746 5 1 1 40745
0 40747 7 1 2 72728 40746
0 40748 5 1 1 40747
0 40749 7 1 2 99810 92259
0 40750 7 1 2 79121 40749
0 40751 5 3 1 40750
0 40752 7 1 2 40748 104864
0 40753 5 1 1 40752
0 40754 7 1 2 72449 40753
0 40755 5 1 1 40754
0 40756 7 1 2 70855 40755
0 40757 5 1 1 40756
0 40758 7 1 2 102635 40757
0 40759 7 1 2 40688 40758
0 40760 5 1 1 40759
0 40761 7 2 2 97938 85162
0 40762 7 1 2 78511 104867
0 40763 5 1 1 40762
0 40764 7 1 2 78485 94364
0 40765 5 1 1 40764
0 40766 7 1 2 87062 97687
0 40767 5 1 1 40766
0 40768 7 1 2 40765 40767
0 40769 5 1 1 40768
0 40770 7 1 2 78253 40769
0 40771 5 1 1 40770
0 40772 7 1 2 40763 40771
0 40773 5 1 1 40772
0 40774 7 1 2 68121 40773
0 40775 5 1 1 40774
0 40776 7 2 2 86391 94920
0 40777 7 1 2 97933 104869
0 40778 5 1 1 40777
0 40779 7 1 2 77476 97502
0 40780 5 1 1 40779
0 40781 7 1 2 81904 97663
0 40782 5 1 1 40781
0 40783 7 1 2 40782 98367
0 40784 7 1 2 40780 40783
0 40785 5 1 1 40784
0 40786 7 1 2 78254 40785
0 40787 5 1 1 40786
0 40788 7 1 2 40778 40787
0 40789 5 1 1 40788
0 40790 7 1 2 87804 40789
0 40791 5 1 1 40790
0 40792 7 1 2 40775 40791
0 40793 5 1 1 40792
0 40794 7 1 2 102760 40793
0 40795 5 1 1 40794
0 40796 7 1 2 64184 40795
0 40797 7 1 2 40760 40796
0 40798 5 1 1 40797
0 40799 7 2 2 68122 89044
0 40800 5 2 1 104871
0 40801 7 1 2 73220 83570
0 40802 5 1 1 40801
0 40803 7 1 2 104873 40802
0 40804 7 1 2 97523 40803
0 40805 5 1 1 40804
0 40806 7 1 2 71131 40805
0 40807 5 1 1 40806
0 40808 7 2 2 94045 86245
0 40809 7 1 2 69561 104875
0 40810 5 1 1 40809
0 40811 7 1 2 40810 87172
0 40812 5 1 1 40811
0 40813 7 1 2 75420 40812
0 40814 5 1 1 40813
0 40815 7 1 2 87670 95151
0 40816 5 1 1 40815
0 40817 7 1 2 40816 97525
0 40818 7 1 2 40814 40817
0 40819 7 1 2 40807 40818
0 40820 5 1 1 40819
0 40821 7 1 2 78255 40820
0 40822 5 1 1 40821
0 40823 7 1 2 81053 97943
0 40824 5 1 1 40823
0 40825 7 1 2 90218 97531
0 40826 5 1 1 40825
0 40827 7 1 2 40824 40826
0 40828 5 1 1 40827
0 40829 7 1 2 85163 40828
0 40830 5 1 1 40829
0 40831 7 1 2 40822 40830
0 40832 5 1 1 40831
0 40833 7 1 2 67715 40832
0 40834 5 1 1 40833
0 40835 7 1 2 97939 104870
0 40836 5 1 1 40835
0 40837 7 1 2 68462 104856
0 40838 5 1 1 40837
0 40839 7 1 2 40836 40838
0 40840 5 1 1 40839
0 40841 7 1 2 85021 40840
0 40842 5 1 1 40841
0 40843 7 1 2 40834 40842
0 40844 5 1 1 40843
0 40845 7 1 2 97910 40844
0 40846 5 1 1 40845
0 40847 7 1 2 77004 91019
0 40848 7 1 2 102819 40847
0 40849 5 1 1 40848
0 40850 7 2 2 97106 96399
0 40851 7 1 2 83907 79111
0 40852 7 1 2 104877 40851
0 40853 5 1 1 40852
0 40854 7 1 2 40849 40853
0 40855 5 1 1 40854
0 40856 7 1 2 67716 40855
0 40857 5 1 1 40856
0 40858 7 7 2 68692 85022
0 40859 7 1 2 89088 104878
0 40860 7 1 2 104879 40859
0 40861 5 1 1 40860
0 40862 7 1 2 40857 40861
0 40863 5 1 1 40862
0 40864 7 1 2 71132 40863
0 40865 5 1 1 40864
0 40866 7 2 2 89089 79521
0 40867 7 1 2 100971 90991
0 40868 7 1 2 104886 40867
0 40869 5 1 1 40868
0 40870 7 1 2 40865 40869
0 40871 5 1 1 40870
0 40872 7 1 2 84850 40871
0 40873 5 1 1 40872
0 40874 7 1 2 73221 103637
0 40875 5 1 1 40874
0 40876 7 1 2 104874 40875
0 40877 5 1 1 40876
0 40878 7 1 2 78256 40877
0 40879 5 1 1 40878
0 40880 7 1 2 88818 104729
0 40881 5 1 1 40880
0 40882 7 1 2 40879 40881
0 40883 5 1 1 40882
0 40884 7 1 2 98409 40883
0 40885 5 1 1 40884
0 40886 7 1 2 87805 97510
0 40887 5 1 1 40886
0 40888 7 1 2 90934 95152
0 40889 5 1 1 40888
0 40890 7 1 2 40887 40889
0 40891 5 1 1 40890
0 40892 7 1 2 69562 40891
0 40893 5 1 1 40892
0 40894 7 4 2 67717 79735
0 40895 7 1 2 83398 76709
0 40896 7 1 2 104888 40895
0 40897 5 1 1 40896
0 40898 7 1 2 40893 40897
0 40899 5 1 1 40898
0 40900 7 1 2 78257 40899
0 40901 5 1 1 40900
0 40902 7 1 2 67718 104876
0 40903 5 1 1 40902
0 40904 7 1 2 40903 98949
0 40905 5 1 1 40904
0 40906 7 1 2 104451 40905
0 40907 5 1 1 40906
0 40908 7 2 2 67719 74797
0 40909 7 1 2 97562 79122
0 40910 7 1 2 104892 40909
0 40911 5 1 1 40910
0 40912 7 1 2 40907 40911
0 40913 5 1 1 40912
0 40914 7 1 2 75421 40913
0 40915 5 1 1 40914
0 40916 7 1 2 83908 78258
0 40917 5 1 1 40916
0 40918 7 1 2 104734 40917
0 40919 5 1 1 40918
0 40920 7 1 2 80234 40919
0 40921 5 1 1 40920
0 40922 7 2 2 68123 77125
0 40923 7 1 2 91108 104894
0 40924 5 1 1 40923
0 40925 7 1 2 40921 40924
0 40926 5 1 1 40925
0 40927 7 1 2 80640 40926
0 40928 5 1 1 40927
0 40929 7 1 2 75031 103826
0 40930 5 1 1 40929
0 40931 7 1 2 40928 40930
0 40932 5 1 1 40931
0 40933 7 1 2 81905 78460
0 40934 7 1 2 40932 40933
0 40935 5 1 1 40934
0 40936 7 1 2 97324 91704
0 40937 7 1 2 104750 40936
0 40938 7 1 2 104895 40937
0 40939 5 1 1 40938
0 40940 7 1 2 72450 40939
0 40941 7 1 2 40935 40940
0 40942 7 1 2 40915 40941
0 40943 7 1 2 40901 40942
0 40944 5 1 1 40943
0 40945 7 1 2 85780 96179
0 40946 5 1 1 40945
0 40947 7 1 2 66052 104868
0 40948 5 1 1 40947
0 40949 7 1 2 40946 40948
0 40950 5 1 1 40949
0 40951 7 1 2 68124 40950
0 40952 5 1 1 40951
0 40953 7 1 2 68463 95856
0 40954 5 1 1 40953
0 40955 7 1 2 77005 40954
0 40956 5 1 1 40955
0 40957 7 1 2 84257 40956
0 40958 5 1 1 40957
0 40959 7 1 2 95942 90203
0 40960 5 1 1 40959
0 40961 7 1 2 81906 104463
0 40962 5 1 1 40961
0 40963 7 1 2 40960 40962
0 40964 5 1 1 40963
0 40965 7 1 2 40958 40964
0 40966 5 1 1 40965
0 40967 7 1 2 40952 40966
0 40968 5 1 1 40967
0 40969 7 1 2 64455 40968
0 40970 5 1 1 40969
0 40971 7 1 2 86967 104740
0 40972 5 1 1 40971
0 40973 7 1 2 89915 104730
0 40974 5 1 1 40973
0 40975 7 1 2 40972 40974
0 40976 5 1 1 40975
0 40977 7 1 2 74686 40976
0 40978 5 1 1 40977
0 40979 7 1 2 73783 89916
0 40980 7 1 2 85655 40979
0 40981 7 1 2 91020 40980
0 40982 5 1 1 40981
0 40983 7 1 2 40978 40982
0 40984 7 1 2 40970 40983
0 40985 5 1 1 40984
0 40986 7 1 2 72729 40985
0 40987 5 1 1 40986
0 40988 7 1 2 67378 104865
0 40989 7 1 2 40987 40988
0 40990 5 1 1 40989
0 40991 7 1 2 40944 40990
0 40992 5 1 1 40991
0 40993 7 1 2 40885 40992
0 40994 5 1 1 40993
0 40995 7 1 2 70856 40994
0 40996 5 1 1 40995
0 40997 7 1 2 40873 40996
0 40998 7 1 2 40846 40997
0 40999 5 1 1 40998
0 41000 7 1 2 102691 40999
0 41001 5 1 1 41000
0 41002 7 2 2 97955 83729
0 41003 5 1 1 104896
0 41004 7 1 2 98237 81401
0 41005 5 1 1 41004
0 41006 7 1 2 41003 41005
0 41007 5 1 1 41006
0 41008 7 1 2 69563 41007
0 41009 5 1 1 41008
0 41010 7 2 2 67379 95294
0 41011 7 1 2 78381 104898
0 41012 5 1 1 41011
0 41013 7 1 2 41009 41012
0 41014 5 1 1 41013
0 41015 7 1 2 74687 41014
0 41016 5 1 1 41015
0 41017 7 1 2 98223 104643
0 41018 5 1 1 41017
0 41019 7 1 2 41016 41018
0 41020 5 1 1 41019
0 41021 7 1 2 73222 41020
0 41022 5 1 1 41021
0 41023 7 2 2 75422 78512
0 41024 7 1 2 98033 104900
0 41025 5 1 1 41024
0 41026 7 1 2 41022 41025
0 41027 5 1 1 41026
0 41028 7 1 2 85164 41027
0 41029 5 1 1 41028
0 41030 7 1 2 95801 103827
0 41031 7 1 2 104126 41030
0 41032 5 1 1 41031
0 41033 7 1 2 41029 41032
0 41034 5 1 1 41033
0 41035 7 1 2 70857 41034
0 41036 5 1 1 41035
0 41037 7 1 2 68125 96155
0 41038 5 1 1 41037
0 41039 7 1 2 104735 41038
0 41040 5 1 1 41039
0 41041 7 1 2 78486 104030
0 41042 7 1 2 41040 41041
0 41043 5 1 1 41042
0 41044 7 1 2 41036 41043
0 41045 5 1 1 41044
0 41046 7 1 2 102692 41045
0 41047 5 1 1 41046
0 41048 7 1 2 103828 104601
0 41049 5 1 1 41048
0 41050 7 1 2 38187 41049
0 41051 5 1 1 41050
0 41052 7 1 2 102738 104473
0 41053 7 1 2 41051 41052
0 41054 5 1 1 41053
0 41055 7 1 2 41047 41054
0 41056 5 1 1 41055
0 41057 7 1 2 80725 41056
0 41058 5 1 1 41057
0 41059 7 1 2 81907 104653
0 41060 5 1 1 41059
0 41061 7 1 2 104651 41060
0 41062 5 1 1 41061
0 41063 7 1 2 73223 41062
0 41064 5 1 1 41063
0 41065 7 1 2 101566 89045
0 41066 5 1 1 41065
0 41067 7 1 2 41064 41066
0 41068 5 1 1 41067
0 41069 7 1 2 78259 41068
0 41070 5 1 1 41069
0 41071 7 1 2 101704 92648
0 41072 5 1 1 41071
0 41073 7 1 2 40062 41072
0 41074 5 1 1 41073
0 41075 7 1 2 73554 41074
0 41076 5 1 1 41075
0 41077 7 1 2 77380 85808
0 41078 5 1 1 41077
0 41079 7 1 2 41076 41078
0 41080 5 1 1 41079
0 41081 7 1 2 85165 41080
0 41082 5 1 1 41081
0 41083 7 1 2 41070 41082
0 41084 5 1 1 41083
0 41085 7 1 2 72730 41084
0 41086 5 1 1 41085
0 41087 7 1 2 104866 41086
0 41088 5 1 1 41087
0 41089 7 1 2 102739 41088
0 41090 5 1 1 41089
0 41091 7 1 2 69233 41090
0 41092 7 1 2 41058 41091
0 41093 7 1 2 41001 41092
0 41094 5 1 1 41093
0 41095 7 1 2 97409 41094
0 41096 7 1 2 40798 41095
0 41097 5 1 1 41096
0 41098 7 1 2 40481 41097
0 41099 7 1 2 40078 41098
0 41100 7 1 2 39431 41099
0 41101 7 1 2 84528 83994
0 41102 7 1 2 102740 41101
0 41103 5 1 1 41102
0 41104 7 1 2 98377 103926
0 41105 5 1 1 41104
0 41106 7 1 2 68464 104844
0 41107 5 1 1 41106
0 41108 7 1 2 41105 41107
0 41109 5 1 1 41108
0 41110 7 1 2 90863 102792
0 41111 7 1 2 41109 41110
0 41112 5 1 1 41111
0 41113 7 1 2 41103 41112
0 41114 5 1 1 41113
0 41115 7 1 2 71848 41114
0 41116 5 1 1 41115
0 41117 7 1 2 69564 95297
0 41118 5 3 1 41117
0 41119 7 1 2 66770 104902
0 41120 5 1 1 41119
0 41121 7 1 2 16210 41120
0 41122 5 1 1 41121
0 41123 7 1 2 98189 102667
0 41124 7 1 2 41122 41123
0 41125 5 1 1 41124
0 41126 7 1 2 41116 41125
0 41127 5 1 1 41126
0 41128 7 1 2 71133 41127
0 41129 5 1 1 41128
0 41130 7 1 2 80994 102378
0 41131 5 1 1 41130
0 41132 7 5 2 68693 90234
0 41133 5 2 1 104905
0 41134 7 1 2 102375 104910
0 41135 5 1 1 41134
0 41136 7 1 2 67720 76626
0 41137 7 1 2 41135 41136
0 41138 5 1 1 41137
0 41139 7 1 2 41131 41138
0 41140 5 1 1 41139
0 41141 7 1 2 102725 41140
0 41142 5 1 1 41141
0 41143 7 1 2 41129 41142
0 41144 5 1 1 41143
0 41145 7 1 2 76493 41144
0 41146 5 1 1 41145
0 41147 7 1 2 98253 36869
0 41148 5 1 1 41147
0 41149 7 1 2 104344 41148
0 41150 5 1 1 41149
0 41151 7 1 2 82173 103717
0 41152 7 1 2 102385 41151
0 41153 5 1 1 41152
0 41154 7 1 2 41150 41153
0 41155 5 1 1 41154
0 41156 7 1 2 64185 41155
0 41157 5 1 1 41156
0 41158 7 2 2 72731 84364
0 41159 5 2 1 104912
0 41160 7 1 2 99189 82124
0 41161 7 1 2 104913 41160
0 41162 5 1 1 41161
0 41163 7 1 2 41157 41162
0 41164 5 1 1 41163
0 41165 7 1 2 102657 41164
0 41166 5 1 1 41165
0 41167 7 1 2 67721 104203
0 41168 5 1 1 41167
0 41169 7 1 2 103848 41168
0 41170 5 2 1 41169
0 41171 7 1 2 77731 104737
0 41172 5 1 1 41171
0 41173 7 1 2 71849 102668
0 41174 7 1 2 86663 41173
0 41175 5 1 1 41174
0 41176 7 1 2 41172 41175
0 41177 5 1 1 41176
0 41178 7 1 2 104916 41177
0 41179 5 1 1 41178
0 41180 7 1 2 80425 102636
0 41181 7 1 2 101980 41180
0 41182 7 1 2 104638 41181
0 41183 5 1 1 41182
0 41184 7 2 2 76494 101193
0 41185 5 3 1 104918
0 41186 7 2 2 100579 102130
0 41187 5 1 1 104923
0 41188 7 1 2 104920 41187
0 41189 5 2 1 41188
0 41190 7 1 2 95638 104622
0 41191 7 1 2 104925 41190
0 41192 5 1 1 41191
0 41193 7 1 2 41183 41192
0 41194 5 1 1 41193
0 41195 7 1 2 75423 41194
0 41196 5 1 1 41195
0 41197 7 1 2 41179 41196
0 41198 7 1 2 41166 41197
0 41199 7 1 2 41146 41198
0 41200 5 1 1 41199
0 41201 7 1 2 78260 41200
0 41202 5 1 1 41201
0 41203 7 1 2 80968 102479
0 41204 5 1 1 41203
0 41205 7 1 2 84163 88780
0 41206 5 1 1 41205
0 41207 7 1 2 41204 41206
0 41208 5 2 1 41207
0 41209 7 1 2 103614 104927
0 41210 5 1 1 41209
0 41211 7 1 2 99523 84529
0 41212 7 1 2 86117 41211
0 41213 5 1 1 41212
0 41214 7 1 2 41210 41213
0 41215 5 1 1 41214
0 41216 7 1 2 83752 41215
0 41217 5 1 1 41216
0 41218 7 1 2 98399 104928
0 41219 5 1 1 41218
0 41220 7 1 2 99524 83730
0 41221 7 1 2 92178 41220
0 41222 5 1 1 41221
0 41223 7 1 2 41219 41222
0 41224 5 1 1 41223
0 41225 7 1 2 74197 41224
0 41226 5 1 1 41225
0 41227 7 2 2 78128 96759
0 41228 5 1 1 104929
0 41229 7 1 2 99719 81150
0 41230 7 1 2 104930 41229
0 41231 5 1 1 41230
0 41232 7 1 2 41226 41231
0 41233 7 1 2 41217 41232
0 41234 5 1 1 41233
0 41235 7 1 2 67221 41234
0 41236 5 1 1 41235
0 41237 7 2 2 95615 101547
0 41238 7 1 2 70231 102165
0 41239 7 1 2 104931 41238
0 41240 5 1 1 41239
0 41241 7 1 2 41236 41240
0 41242 5 1 1 41241
0 41243 7 1 2 70858 41242
0 41244 5 1 1 41243
0 41245 7 2 2 67222 97053
0 41246 7 1 2 92842 104933
0 41247 7 1 2 104932 41246
0 41248 5 1 1 41247
0 41249 7 1 2 41244 41248
0 41250 5 1 1 41249
0 41251 7 1 2 72172 41250
0 41252 5 1 1 41251
0 41253 7 1 2 101742 102710
0 41254 7 1 2 104481 41253
0 41255 5 1 1 41254
0 41256 7 1 2 67128 83995
0 41257 7 1 2 103311 41256
0 41258 7 1 2 104491 41257
0 41259 5 1 1 41258
0 41260 7 1 2 41255 41259
0 41261 5 1 1 41260
0 41262 7 1 2 64186 41261
0 41263 5 1 1 41262
0 41264 7 1 2 104840 104845
0 41265 5 1 1 41264
0 41266 7 1 2 78394 41265
0 41267 5 1 1 41266
0 41268 7 1 2 102247 74346
0 41269 5 1 1 41268
0 41270 7 1 2 41267 41269
0 41271 5 1 1 41270
0 41272 7 1 2 77182 41271
0 41273 5 1 1 41272
0 41274 7 1 2 99156 100580
0 41275 7 1 2 96121 41274
0 41276 5 1 1 41275
0 41277 7 1 2 41273 41276
0 41278 5 1 1 41277
0 41279 7 1 2 68465 102793
0 41280 7 1 2 41278 41279
0 41281 5 1 1 41280
0 41282 7 1 2 41263 41281
0 41283 5 1 1 41282
0 41284 7 1 2 71850 41283
0 41285 5 1 1 41284
0 41286 7 1 2 99031 75062
0 41287 7 1 2 104834 41286
0 41288 7 1 2 78513 41287
0 41289 5 1 1 41288
0 41290 7 1 2 41285 41289
0 41291 5 1 1 41290
0 41292 7 1 2 75424 41291
0 41293 5 1 1 41292
0 41294 7 1 2 100489 101273
0 41295 5 1 1 41294
0 41296 7 1 2 84085 74860
0 41297 7 1 2 98249 41296
0 41298 5 1 1 41297
0 41299 7 1 2 41295 41298
0 41300 5 1 1 41299
0 41301 7 1 2 64187 41300
0 41302 5 1 1 41301
0 41303 7 1 2 71450 103835
0 41304 7 1 2 104819 41303
0 41305 5 1 1 41304
0 41306 7 1 2 41302 41305
0 41307 5 1 1 41306
0 41308 7 1 2 102394 91244
0 41309 7 1 2 41307 41308
0 41310 5 1 1 41309
0 41311 7 1 2 41293 41310
0 41312 7 1 2 41252 41311
0 41313 5 1 1 41312
0 41314 7 1 2 85166 41313
0 41315 5 1 1 41314
0 41316 7 1 2 41202 41315
0 41317 5 1 1 41316
0 41318 7 1 2 70493 41317
0 41319 5 1 1 41318
0 41320 7 1 2 31425 75702
0 41321 5 5 1 41320
0 41322 7 1 2 104897 104935
0 41323 5 1 1 41322
0 41324 7 1 2 68466 88329
0 41325 5 1 1 41324
0 41326 7 1 2 92961 41325
0 41327 5 1 1 41326
0 41328 7 1 2 98400 41327
0 41329 5 1 1 41328
0 41330 7 1 2 41323 41329
0 41331 5 1 1 41330
0 41332 7 1 2 64456 41331
0 41333 5 1 1 41332
0 41334 7 1 2 87235 101174
0 41335 5 1 1 41334
0 41336 7 1 2 102146 83753
0 41337 5 1 1 41336
0 41338 7 1 2 41335 41337
0 41339 5 1 1 41338
0 41340 7 1 2 98612 41339
0 41341 5 1 1 41340
0 41342 7 1 2 41333 41341
0 41343 5 1 1 41342
0 41344 7 1 2 66771 41343
0 41345 5 1 1 41344
0 41346 7 1 2 103844 80109
0 41347 5 1 1 41346
0 41348 7 1 2 41345 41347
0 41349 5 1 1 41348
0 41350 7 1 2 69234 41349
0 41351 5 1 1 41350
0 41352 7 1 2 99688 75032
0 41353 7 1 2 93531 41352
0 41354 5 1 1 41353
0 41355 7 1 2 41351 41354
0 41356 5 1 1 41355
0 41357 7 1 2 70859 41356
0 41358 5 1 1 41357
0 41359 7 2 2 91431 84521
0 41360 7 1 2 103615 92354
0 41361 7 1 2 104940 41360
0 41362 5 1 1 41361
0 41363 7 1 2 41358 41362
0 41364 5 1 1 41363
0 41365 7 1 2 85167 41364
0 41366 5 1 1 41365
0 41367 7 2 2 85082 92385
0 41368 5 1 1 104942
0 41369 7 1 2 86959 104943
0 41370 5 1 1 41369
0 41371 7 1 2 104645 95299
0 41372 5 1 1 41371
0 41373 7 1 2 41370 41372
0 41374 5 1 1 41373
0 41375 7 4 2 95283 98613
0 41376 7 1 2 78261 104944
0 41377 7 1 2 41374 41376
0 41378 5 1 1 41377
0 41379 7 1 2 41366 41378
0 41380 5 1 1 41379
0 41381 7 1 2 67223 41380
0 41382 5 1 1 41381
0 41383 7 1 2 87250 95868
0 41384 5 1 1 41383
0 41385 7 1 2 68467 91060
0 41386 5 1 1 41385
0 41387 7 1 2 41384 41386
0 41388 5 1 1 41387
0 41389 7 1 2 100572 101194
0 41390 7 1 2 41388 41389
0 41391 5 1 1 41390
0 41392 7 1 2 41382 41391
0 41393 5 1 1 41392
0 41394 7 1 2 72173 41393
0 41395 5 1 1 41394
0 41396 7 1 2 82137 86239
0 41397 5 1 1 41396
0 41398 7 1 2 6981 41397
0 41399 5 1 1 41398
0 41400 7 1 2 78262 41399
0 41401 5 1 1 41400
0 41402 7 1 2 78896 84674
0 41403 5 1 1 41402
0 41404 7 1 2 79283 81402
0 41405 5 1 1 41404
0 41406 7 1 2 41403 41405
0 41407 5 1 1 41406
0 41408 7 1 2 84711 90078
0 41409 7 1 2 41407 41408
0 41410 5 1 1 41409
0 41411 7 1 2 41401 41410
0 41412 5 1 1 41411
0 41413 7 1 2 73784 41412
0 41414 5 1 1 41413
0 41415 7 1 2 64830 7342
0 41416 5 2 1 41415
0 41417 7 1 2 68468 104948
0 41418 5 1 1 41417
0 41419 7 1 2 41418 80818
0 41420 5 1 1 41419
0 41421 7 1 2 66358 41420
0 41422 5 3 1 41421
0 41423 7 1 2 92962 104950
0 41424 5 1 1 41423
0 41425 7 1 2 81533 41424
0 41426 5 1 1 41425
0 41427 7 1 2 103839 104951
0 41428 5 1 1 41427
0 41429 7 1 2 81474 41428
0 41430 5 1 1 41429
0 41431 7 1 2 41426 41430
0 41432 5 1 1 41431
0 41433 7 1 2 85168 41432
0 41434 5 1 1 41433
0 41435 7 1 2 41414 41434
0 41436 5 1 1 41435
0 41437 7 1 2 71134 41436
0 41438 5 1 1 41437
0 41439 7 1 2 87563 78897
0 41440 5 1 1 41439
0 41441 7 1 2 69934 96854
0 41442 5 1 1 41441
0 41443 7 1 2 41440 41442
0 41444 5 1 1 41443
0 41445 7 1 2 71451 41444
0 41446 5 1 1 41445
0 41447 7 1 2 104952 41446
0 41448 5 1 1 41447
0 41449 7 1 2 90079 92939
0 41450 7 1 2 41448 41449
0 41451 5 1 1 41450
0 41452 7 1 2 41438 41451
0 41453 5 1 1 41452
0 41454 7 1 2 72451 41453
0 41455 5 1 1 41454
0 41456 7 1 2 94644 87111
0 41457 5 1 1 41456
0 41458 7 1 2 80426 85169
0 41459 7 1 2 104936 41458
0 41460 5 1 1 41459
0 41461 7 1 2 41457 41460
0 41462 5 1 1 41461
0 41463 7 1 2 103845 41462
0 41464 5 1 1 41463
0 41465 7 1 2 41455 41464
0 41466 5 1 1 41465
0 41467 7 1 2 102612 41466
0 41468 5 1 1 41467
0 41469 7 1 2 26055 101642
0 41470 5 1 1 41469
0 41471 7 1 2 71452 41470
0 41472 5 1 1 41471
0 41473 7 1 2 82607 83328
0 41474 5 2 1 41473
0 41475 7 1 2 41472 104953
0 41476 5 1 1 41475
0 41477 7 1 2 104769 104611
0 41478 7 1 2 41476 41477
0 41479 5 1 1 41478
0 41480 7 1 2 69235 41479
0 41481 7 1 2 41468 41480
0 41482 5 1 1 41481
0 41483 7 1 2 78514 104937
0 41484 5 1 1 41483
0 41485 7 1 2 73555 77114
0 41486 7 1 2 99140 41485
0 41487 5 1 1 41486
0 41488 7 1 2 41484 41487
0 41489 5 1 1 41488
0 41490 7 1 2 96176 41489
0 41491 5 1 1 41490
0 41492 7 1 2 103652 37691
0 41493 5 1 1 41492
0 41494 7 1 2 71453 41493
0 41495 5 1 1 41494
0 41496 7 1 2 68469 99830
0 41497 5 1 1 41496
0 41498 7 1 2 76495 101713
0 41499 5 1 1 41498
0 41500 7 1 2 41497 41499
0 41501 5 1 1 41500
0 41502 7 1 2 82990 41501
0 41503 5 1 1 41502
0 41504 7 1 2 41495 41503
0 41505 5 1 1 41504
0 41506 7 1 2 67722 41505
0 41507 5 1 1 41506
0 41508 7 1 2 90759 104903
0 41509 5 1 1 41508
0 41510 7 1 2 95314 91093
0 41511 5 1 1 41510
0 41512 7 1 2 41509 41511
0 41513 5 1 1 41512
0 41514 7 1 2 68470 41513
0 41515 5 1 1 41514
0 41516 7 1 2 66772 81475
0 41517 7 1 2 92739 41516
0 41518 5 1 1 41517
0 41519 7 1 2 41515 41518
0 41520 5 1 1 41519
0 41521 7 1 2 71135 41520
0 41522 5 1 1 41521
0 41523 7 1 2 92772 75693
0 41524 7 1 2 103701 41523
0 41525 5 1 1 41524
0 41526 7 1 2 41522 41525
0 41527 7 1 2 41507 41526
0 41528 5 1 1 41527
0 41529 7 1 2 78263 41528
0 41530 5 1 1 41529
0 41531 7 1 2 41491 41530
0 41532 5 1 1 41531
0 41533 7 1 2 72452 41532
0 41534 5 1 1 41533
0 41535 7 1 2 103467 96184
0 41536 5 1 1 41535
0 41537 7 1 2 84164 79123
0 41538 5 1 1 41537
0 41539 7 1 2 41536 41538
0 41540 5 1 1 41539
0 41541 7 1 2 78584 41540
0 41542 5 1 1 41541
0 41543 7 1 2 95789 104445
0 41544 5 1 1 41543
0 41545 7 1 2 41542 41544
0 41546 5 1 1 41545
0 41547 7 1 2 97752 41546
0 41548 5 1 1 41547
0 41549 7 1 2 41534 41548
0 41550 5 1 1 41549
0 41551 7 1 2 102658 41550
0 41552 5 1 1 41551
0 41553 7 1 2 95352 95315
0 41554 7 1 2 78264 104511
0 41555 7 1 2 41553 41554
0 41556 7 1 2 87617 41555
0 41557 5 1 1 41556
0 41558 7 1 2 64188 41557
0 41559 7 1 2 41552 41558
0 41560 5 1 1 41559
0 41561 7 1 2 65475 41560
0 41562 7 1 2 41482 41561
0 41563 5 1 1 41562
0 41564 7 1 2 76236 93781
0 41565 5 1 1 41564
0 41566 7 1 2 41565 94180
0 41567 5 1 1 41566
0 41568 7 1 2 68471 41567
0 41569 5 1 1 41568
0 41570 7 1 2 92740 95107
0 41571 5 1 1 41570
0 41572 7 1 2 41569 41571
0 41573 5 1 1 41572
0 41574 7 1 2 98460 102637
0 41575 7 1 2 41573 41574
0 41576 5 1 1 41575
0 41577 7 1 2 83458 97604
0 41578 5 1 1 41577
0 41579 7 1 2 100821 102774
0 41580 7 1 2 41578 41579
0 41581 5 1 1 41580
0 41582 7 1 2 41576 41581
0 41583 5 1 1 41582
0 41584 7 1 2 104667 41583
0 41585 5 1 1 41584
0 41586 7 1 2 87251 80974
0 41587 5 2 1 41586
0 41588 7 1 2 92176 104955
0 41589 5 1 1 41588
0 41590 7 1 2 80641 41589
0 41591 5 1 1 41590
0 41592 7 1 2 81756 104938
0 41593 5 1 1 41592
0 41594 7 1 2 1356 41593
0 41595 7 1 2 41591 41594
0 41596 5 1 1 41595
0 41597 7 1 2 78515 41596
0 41598 5 1 1 41597
0 41599 7 3 2 82608 97771
0 41600 5 1 1 104957
0 41601 7 1 2 80235 98986
0 41602 5 1 1 41601
0 41603 7 1 2 41600 41602
0 41604 5 1 1 41603
0 41605 7 1 2 69935 81092
0 41606 7 1 2 41604 41605
0 41607 5 1 1 41606
0 41608 7 1 2 41598 41607
0 41609 5 1 1 41608
0 41610 7 1 2 102775 41609
0 41611 5 1 1 41610
0 41612 7 2 2 77056 79208
0 41613 5 1 1 104960
0 41614 7 1 2 75703 41613
0 41615 5 1 1 41614
0 41616 7 2 2 98763 102693
0 41617 7 1 2 41615 104962
0 41618 5 1 1 41617
0 41619 7 2 2 64831 92584
0 41620 7 1 2 103312 97478
0 41621 7 1 2 104964 41620
0 41622 5 1 1 41621
0 41623 7 1 2 41618 41622
0 41624 5 1 1 41623
0 41625 7 1 2 81054 41624
0 41626 5 1 1 41625
0 41627 7 1 2 92549 104512
0 41628 7 1 2 104939 41627
0 41629 5 1 1 41628
0 41630 7 1 2 41626 41629
0 41631 5 1 1 41630
0 41632 7 1 2 88371 41631
0 41633 5 1 1 41632
0 41634 7 1 2 99032 87885
0 41635 7 1 2 102638 41634
0 41636 7 1 2 74861 91135
0 41637 7 1 2 95243 41636
0 41638 7 1 2 41635 41637
0 41639 5 1 1 41638
0 41640 7 1 2 41633 41639
0 41641 7 1 2 41611 41640
0 41642 5 1 1 41641
0 41643 7 1 2 85170 41642
0 41644 5 1 1 41643
0 41645 7 1 2 41585 41644
0 41646 5 1 1 41645
0 41647 7 1 2 85539 41646
0 41648 5 1 1 41647
0 41649 7 1 2 76604 78453
0 41650 5 1 1 41649
0 41651 7 2 2 71454 83739
0 41652 5 1 1 104966
0 41653 7 1 2 71689 41652
0 41654 7 1 2 41650 41653
0 41655 5 1 1 41654
0 41656 7 1 2 66359 104794
0 41657 5 1 1 41656
0 41658 7 1 2 41655 41657
0 41659 5 1 1 41658
0 41660 7 1 2 70232 41659
0 41661 5 1 1 41660
0 41662 7 2 2 71136 80084
0 41663 7 1 2 83996 104968
0 41664 5 1 1 41663
0 41665 7 1 2 41661 41664
0 41666 5 1 1 41665
0 41667 7 1 2 69565 41666
0 41668 5 1 1 41667
0 41669 7 1 2 76496 83754
0 41670 5 1 1 41669
0 41671 7 1 2 34688 41670
0 41672 5 1 1 41671
0 41673 7 1 2 90244 41672
0 41674 5 1 1 41673
0 41675 7 1 2 41668 41674
0 41676 5 1 1 41675
0 41677 7 1 2 64189 41676
0 41678 5 1 1 41677
0 41679 7 1 2 99986 96837
0 41680 5 1 1 41679
0 41681 7 1 2 41678 41680
0 41682 5 1 1 41681
0 41683 7 1 2 98190 104595
0 41684 7 1 2 41682 41683
0 41685 5 1 1 41684
0 41686 7 1 2 41648 41685
0 41687 7 1 2 41563 41686
0 41688 7 1 2 41395 41687
0 41689 7 1 2 41319 41688
0 41690 5 1 1 41689
0 41691 7 1 2 68126 41690
0 41692 5 1 1 41691
0 41693 7 1 2 75475 85171
0 41694 5 1 1 41693
0 41695 7 1 2 91031 41694
0 41696 5 3 1 41695
0 41697 7 1 2 84675 104970
0 41698 5 1 1 41697
0 41699 7 1 2 92631 91021
0 41700 5 1 1 41699
0 41701 7 1 2 41698 41700
0 41702 5 1 1 41701
0 41703 7 1 2 68472 41702
0 41704 5 1 1 41703
0 41705 7 1 2 93634 92985
0 41706 5 1 1 41705
0 41707 7 1 2 81403 78265
0 41708 5 1 1 41707
0 41709 7 1 2 41706 41708
0 41710 5 1 1 41709
0 41711 7 1 2 70233 41710
0 41712 5 1 1 41711
0 41713 7 1 2 41704 41712
0 41714 5 1 1 41713
0 41715 7 1 2 76497 41714
0 41716 5 1 1 41715
0 41717 7 4 2 67723 76395
0 41718 7 1 2 90896 96242
0 41719 7 1 2 104973 41718
0 41720 5 1 1 41719
0 41721 7 1 2 41716 41720
0 41722 5 1 1 41721
0 41723 7 1 2 68127 41722
0 41724 5 1 1 41723
0 41725 7 1 2 74798 81612
0 41726 7 1 2 92998 41725
0 41727 5 1 1 41726
0 41728 7 1 2 41724 41727
0 41729 5 1 1 41728
0 41730 7 1 2 81908 41729
0 41731 5 1 1 41730
0 41732 7 1 2 95773 84676
0 41733 5 1 1 41732
0 41734 7 1 2 67724 94367
0 41735 5 1 1 41734
0 41736 7 1 2 41733 41735
0 41737 5 1 1 41736
0 41738 7 1 2 85172 41737
0 41739 5 1 1 41738
0 41740 7 1 2 67725 91022
0 41741 7 1 2 101807 41740
0 41742 5 1 1 41741
0 41743 7 1 2 41739 41742
0 41744 5 1 1 41743
0 41745 7 1 2 70234 41744
0 41746 5 1 1 41745
0 41747 7 1 2 86926 101805
0 41748 5 1 1 41747
0 41749 7 1 2 78266 41748
0 41750 5 1 1 41749
0 41751 7 1 2 91883 79112
0 41752 7 1 2 97326 41751
0 41753 5 1 1 41752
0 41754 7 1 2 41750 41753
0 41755 5 1 1 41754
0 41756 7 1 2 67726 41755
0 41757 5 1 1 41756
0 41758 7 1 2 41746 41757
0 41759 5 1 1 41758
0 41760 7 1 2 68128 41759
0 41761 5 1 1 41760
0 41762 7 1 2 104397 89855
0 41763 5 1 1 41762
0 41764 7 1 2 41763 95571
0 41765 5 1 1 41764
0 41766 7 1 2 41761 41765
0 41767 5 1 1 41766
0 41768 7 1 2 76498 41767
0 41769 5 1 1 41768
0 41770 7 1 2 41731 41769
0 41771 5 1 1 41770
0 41772 7 1 2 102801 41771
0 41773 5 1 1 41772
0 41774 7 1 2 95779 88296
0 41775 5 1 1 41774
0 41776 7 1 2 95983 41775
0 41777 5 1 1 41776
0 41778 7 1 2 81183 102999
0 41779 5 1 1 41778
0 41780 7 1 2 84912 41779
0 41781 5 1 1 41780
0 41782 7 1 2 66360 88853
0 41783 5 1 1 41782
0 41784 7 1 2 81757 79305
0 41785 5 1 1 41784
0 41786 7 1 2 81909 77631
0 41787 5 1 1 41786
0 41788 7 2 2 65173 41787
0 41789 7 1 2 41785 104977
0 41790 5 1 1 41789
0 41791 7 1 2 41783 41790
0 41792 7 1 2 41781 41791
0 41793 5 1 1 41792
0 41794 7 1 2 85173 41793
0 41795 5 1 1 41794
0 41796 7 1 2 41777 41795
0 41797 5 1 1 41796
0 41798 7 1 2 73224 41797
0 41799 5 1 1 41798
0 41800 7 1 2 86451 5570
0 41801 7 1 2 84925 41800
0 41802 5 1 1 41801
0 41803 7 1 2 74688 90080
0 41804 7 1 2 41802 41803
0 41805 5 1 1 41804
0 41806 7 1 2 86466 90081
0 41807 5 1 1 41806
0 41808 7 1 2 96157 41807
0 41809 7 1 2 41805 41808
0 41810 5 1 1 41809
0 41811 7 1 2 64832 41810
0 41812 5 1 1 41811
0 41813 7 1 2 84576 95785
0 41814 7 1 2 90665 41813
0 41815 5 1 1 41814
0 41816 7 1 2 41812 41815
0 41817 7 1 2 41799 41816
0 41818 5 1 1 41817
0 41819 7 1 2 75019 41818
0 41820 5 1 1 41819
0 41821 7 1 2 76605 104341
0 41822 5 1 1 41821
0 41823 7 1 2 95786 103408
0 41824 5 1 1 41823
0 41825 7 1 2 86255 83071
0 41826 5 1 1 41825
0 41827 7 1 2 41824 41826
0 41828 7 1 2 41822 41827
0 41829 5 1 1 41828
0 41830 7 1 2 78267 41829
0 41831 5 1 1 41830
0 41832 7 1 2 41820 41831
0 41833 5 1 1 41832
0 41834 7 1 2 64457 41833
0 41835 5 1 1 41834
0 41836 7 1 2 90219 96177
0 41837 5 1 1 41836
0 41838 7 1 2 90120 78268
0 41839 5 1 1 41838
0 41840 7 1 2 41837 41839
0 41841 5 1 1 41840
0 41842 7 1 2 65476 41841
0 41843 5 1 1 41842
0 41844 7 1 2 94033 95444
0 41845 5 1 1 41844
0 41846 7 1 2 41843 41845
0 41847 5 1 1 41846
0 41848 7 1 2 81300 41847
0 41849 5 1 1 41848
0 41850 7 1 2 67727 41849
0 41851 7 1 2 41835 41850
0 41852 5 1 1 41851
0 41853 7 2 2 81758 78321
0 41854 5 1 1 104979
0 41855 7 1 2 68129 41854
0 41856 5 1 1 41855
0 41857 7 1 2 104053 41856
0 41858 5 1 1 41857
0 41859 7 1 2 5584 41858
0 41860 5 1 1 41859
0 41861 7 1 2 69566 41860
0 41862 5 1 1 41861
0 41863 7 1 2 82874 74862
0 41864 5 2 1 41863
0 41865 7 1 2 79931 104981
0 41866 5 2 1 41865
0 41867 7 1 2 64833 104983
0 41868 5 1 1 41867
0 41869 7 1 2 41868 12387
0 41870 5 1 1 41869
0 41871 7 1 2 66773 41870
0 41872 5 1 1 41871
0 41873 7 1 2 103734 95583
0 41874 5 1 1 41873
0 41875 7 1 2 41872 41874
0 41876 5 1 1 41875
0 41877 7 1 2 65477 41876
0 41878 5 1 1 41877
0 41879 7 1 2 64458 86620
0 41880 5 1 1 41879
0 41881 7 1 2 103419 6992
0 41882 5 1 1 41881
0 41883 7 1 2 70494 41882
0 41884 5 1 1 41883
0 41885 7 1 2 41880 41884
0 41886 7 1 2 41878 41885
0 41887 5 1 1 41886
0 41888 7 1 2 68130 41887
0 41889 5 1 1 41888
0 41890 7 1 2 41862 41889
0 41891 5 1 1 41890
0 41892 7 1 2 66361 41891
0 41893 5 1 1 41892
0 41894 7 1 2 80427 104860
0 41895 5 1 1 41894
0 41896 7 1 2 69567 103454
0 41897 5 1 1 41896
0 41898 7 1 2 41895 41897
0 41899 5 1 1 41898
0 41900 7 1 2 71455 41899
0 41901 5 1 1 41900
0 41902 7 2 2 66774 78778
0 41903 7 1 2 80026 104985
0 41904 5 1 1 41903
0 41905 7 1 2 41901 41904
0 41906 5 1 1 41905
0 41907 7 1 2 65478 41906
0 41908 5 1 1 41907
0 41909 7 1 2 84772 102920
0 41910 5 1 1 41909
0 41911 7 1 2 41910 79258
0 41912 5 1 1 41911
0 41913 7 1 2 41908 41912
0 41914 5 1 1 41913
0 41915 7 1 2 65174 41914
0 41916 5 1 1 41915
0 41917 7 1 2 75786 86140
0 41918 5 1 1 41917
0 41919 7 1 2 104954 41918
0 41920 5 1 1 41919
0 41921 7 1 2 65479 41920
0 41922 5 1 1 41921
0 41923 7 1 2 93941 95187
0 41924 5 1 1 41923
0 41925 7 1 2 41922 41924
0 41926 5 1 1 41925
0 41927 7 1 2 81214 41926
0 41928 5 1 1 41927
0 41929 7 2 2 69568 96006
0 41930 7 1 2 86220 79234
0 41931 7 1 2 104987 41930
0 41932 5 1 1 41931
0 41933 7 1 2 41928 41932
0 41934 7 1 2 41916 41933
0 41935 7 1 2 41893 41934
0 41936 5 1 1 41935
0 41937 7 1 2 85174 41936
0 41938 5 1 1 41937
0 41939 7 1 2 100534 104187
0 41940 5 1 1 41939
0 41941 7 1 2 73556 97802
0 41942 5 1 1 41941
0 41943 7 1 2 81251 41942
0 41944 5 1 1 41943
0 41945 7 1 2 64834 41944
0 41946 5 1 1 41945
0 41947 7 1 2 41940 41946
0 41948 5 1 1 41947
0 41949 7 1 2 89748 41948
0 41950 5 1 1 41949
0 41951 7 1 2 96592 89613
0 41952 5 1 1 41951
0 41953 7 1 2 94728 79124
0 41954 5 1 1 41953
0 41955 7 1 2 41952 41954
0 41956 5 1 1 41955
0 41957 7 1 2 75063 41956
0 41958 5 1 1 41957
0 41959 7 1 2 79033 79113
0 41960 7 1 2 101843 41959
0 41961 5 1 1 41960
0 41962 7 1 2 41958 41961
0 41963 5 1 1 41962
0 41964 7 1 2 75425 41963
0 41965 5 1 1 41964
0 41966 7 1 2 72732 41965
0 41967 7 1 2 41950 41966
0 41968 7 1 2 41938 41967
0 41969 5 1 1 41968
0 41970 7 1 2 64190 41969
0 41971 7 1 2 41852 41970
0 41972 5 1 1 41971
0 41973 7 1 2 89174 90082
0 41974 5 1 1 41973
0 41975 7 1 2 78280 41974
0 41976 5 1 1 41975
0 41977 7 1 2 74198 96019
0 41978 7 1 2 81301 41977
0 41979 7 1 2 41976 41978
0 41980 5 1 1 41979
0 41981 7 1 2 41972 41980
0 41982 5 1 1 41981
0 41983 7 1 2 102639 41982
0 41984 5 1 1 41983
0 41985 7 1 2 41773 41984
0 41986 5 1 1 41985
0 41987 7 1 2 66053 41986
0 41988 5 1 1 41987
0 41989 7 1 2 84104 104971
0 41990 5 1 1 41989
0 41991 7 1 2 736 41990
0 41992 5 1 1 41991
0 41993 7 1 2 64459 41992
0 41994 5 1 1 41993
0 41995 7 1 2 81476 95984
0 41996 5 1 1 41995
0 41997 7 1 2 41994 41996
0 41998 5 1 1 41997
0 41999 7 1 2 69236 41998
0 42000 5 1 1 41999
0 42001 7 1 2 69569 104368
0 42002 7 1 2 104972 42001
0 42003 5 1 1 42002
0 42004 7 1 2 42000 42003
0 42005 5 1 1 42004
0 42006 7 1 2 71137 42005
0 42007 5 1 1 42006
0 42008 7 1 2 104974 74362
0 42009 7 1 2 79438 42008
0 42010 5 1 1 42009
0 42011 7 1 2 42007 42010
0 42012 5 1 1 42011
0 42013 7 1 2 68131 42012
0 42014 5 1 1 42013
0 42015 7 1 2 69570 100835
0 42016 7 1 2 104359 42015
0 42017 5 1 1 42016
0 42018 7 1 2 42014 42017
0 42019 5 1 1 42018
0 42020 7 1 2 81910 42019
0 42021 5 1 1 42020
0 42022 7 1 2 98971 104369
0 42023 5 1 1 42022
0 42024 7 1 2 99560 85023
0 42025 5 2 1 42024
0 42026 7 1 2 42023 104989
0 42027 5 1 1 42026
0 42028 7 1 2 75426 42027
0 42029 5 1 1 42028
0 42030 7 1 2 84258 104370
0 42031 5 1 1 42030
0 42032 7 1 2 104990 42031
0 42033 5 1 1 42032
0 42034 7 1 2 68694 42033
0 42035 5 1 1 42034
0 42036 7 1 2 42029 42035
0 42037 5 1 1 42036
0 42038 7 1 2 77183 42037
0 42039 5 1 1 42038
0 42040 7 1 2 94717 82201
0 42041 7 1 2 79750 42040
0 42042 5 1 1 42041
0 42043 7 1 2 42039 42042
0 42044 5 1 1 42043
0 42045 7 1 2 104854 42044
0 42046 5 1 1 42045
0 42047 7 1 2 92808 78061
0 42048 7 1 2 97825 42047
0 42049 5 1 1 42048
0 42050 7 1 2 96881 42049
0 42051 5 1 1 42050
0 42052 7 1 2 100937 85175
0 42053 7 1 2 42051 42052
0 42054 5 1 1 42053
0 42055 7 1 2 42046 42054
0 42056 7 1 2 42021 42055
0 42057 5 1 1 42056
0 42058 7 1 2 102694 42057
0 42059 5 1 1 42058
0 42060 7 1 2 103236 91245
0 42061 7 1 2 85176 42060
0 42062 7 1 2 92959 42061
0 42063 5 1 1 42062
0 42064 7 1 2 76499 74357
0 42065 7 1 2 102695 42064
0 42066 7 1 2 104975 42065
0 42067 5 1 1 42066
0 42068 7 1 2 42063 42067
0 42069 5 1 1 42068
0 42070 7 1 2 64460 42069
0 42071 5 1 1 42070
0 42072 7 1 2 67728 93344
0 42073 7 2 2 67224 75824
0 42074 7 1 2 103381 104991
0 42075 7 1 2 42072 42074
0 42076 5 1 1 42075
0 42077 7 1 2 42071 42076
0 42078 5 1 1 42077
0 42079 7 1 2 68132 42078
0 42080 5 1 1 42079
0 42081 7 1 2 74358 85083
0 42082 7 1 2 102135 42081
0 42083 7 1 2 87084 75836
0 42084 7 1 2 42082 42083
0 42085 5 1 1 42084
0 42086 7 1 2 42080 42085
0 42087 5 1 1 42086
0 42088 7 1 2 84913 42087
0 42089 5 1 1 42088
0 42090 7 2 2 75934 82275
0 42091 5 2 1 104993
0 42092 7 1 2 78959 84259
0 42093 5 1 1 42092
0 42094 7 1 2 81759 42093
0 42095 5 1 1 42094
0 42096 7 1 2 75982 42095
0 42097 5 1 1 42096
0 42098 7 1 2 64835 42097
0 42099 5 1 1 42098
0 42100 7 1 2 104995 42099
0 42101 5 1 1 42100
0 42102 7 4 2 75761 102640
0 42103 7 1 2 78413 104997
0 42104 7 1 2 84535 42103
0 42105 7 1 2 42101 42104
0 42106 5 1 1 42105
0 42107 7 1 2 42089 42106
0 42108 7 1 2 42059 42107
0 42109 5 1 1 42108
0 42110 7 1 2 68473 42109
0 42111 5 1 1 42110
0 42112 7 1 2 79538 101847
0 42113 7 1 2 103333 104607
0 42114 7 1 2 42112 42113
0 42115 5 1 1 42114
0 42116 7 1 2 74557 74359
0 42117 7 1 2 104264 42116
0 42118 7 1 2 75837 42117
0 42119 5 1 1 42118
0 42120 7 1 2 42115 42119
0 42121 5 1 1 42120
0 42122 7 1 2 69571 42121
0 42123 5 1 1 42122
0 42124 7 1 2 73225 79591
0 42125 5 1 1 42124
0 42126 7 1 2 42125 79867
0 42127 5 1 1 42126
0 42128 7 1 2 72269 93047
0 42129 7 1 2 79010 42128
0 42130 7 1 2 98170 42129
0 42131 7 1 2 42127 42130
0 42132 5 1 1 42131
0 42133 7 1 2 42123 42132
0 42134 5 1 1 42133
0 42135 7 1 2 81760 42134
0 42136 5 1 1 42135
0 42137 7 1 2 64191 102641
0 42138 7 1 2 104446 42137
0 42139 7 1 2 94968 42138
0 42140 5 1 1 42139
0 42141 7 3 2 67006 102696
0 42142 7 1 2 84491 93713
0 42143 7 1 2 105001 42142
0 42144 7 1 2 91143 42143
0 42145 7 1 2 89179 42144
0 42146 5 1 1 42145
0 42147 7 1 2 42140 42146
0 42148 7 1 2 42136 42147
0 42149 5 1 1 42148
0 42150 7 1 2 78414 42149
0 42151 5 1 1 42150
0 42152 7 1 2 68133 100595
0 42153 5 1 1 42152
0 42154 7 1 2 65480 93954
0 42155 5 1 1 42154
0 42156 7 1 2 70235 18262
0 42157 7 1 2 42155 42156
0 42158 5 1 1 42157
0 42159 7 1 2 42153 42158
0 42160 5 1 1 42159
0 42161 7 1 2 104379 42160
0 42162 5 1 1 42161
0 42163 7 1 2 80040 83522
0 42164 5 1 1 42163
0 42165 7 1 2 66362 42164
0 42166 5 1 1 42165
0 42167 7 1 2 73557 99493
0 42168 5 1 1 42167
0 42169 7 1 2 42166 42168
0 42170 5 1 1 42169
0 42171 7 1 2 73226 42170
0 42172 5 1 1 42171
0 42173 7 1 2 99512 86246
0 42174 5 1 1 42173
0 42175 7 1 2 100716 42174
0 42176 7 1 2 42172 42175
0 42177 5 1 1 42176
0 42178 7 1 2 69237 42177
0 42179 5 1 1 42178
0 42180 7 1 2 42162 42179
0 42181 5 1 1 42180
0 42182 7 1 2 78269 42181
0 42183 5 1 1 42182
0 42184 7 1 2 91061 104380
0 42185 7 1 2 89180 42184
0 42186 5 1 1 42185
0 42187 7 1 2 42183 42186
0 42188 5 1 1 42187
0 42189 7 1 2 102697 42188
0 42190 5 1 1 42189
0 42191 7 1 2 103229 103455
0 42192 7 1 2 104998 84536
0 42193 7 1 2 42191 42192
0 42194 5 1 1 42193
0 42195 7 1 2 42190 42194
0 42196 5 1 1 42195
0 42197 7 1 2 71138 42196
0 42198 5 1 1 42197
0 42199 7 1 2 96237 102642
0 42200 7 1 2 101464 42199
0 42201 5 1 1 42200
0 42202 7 1 2 99694 80466
0 42203 7 1 2 96726 102698
0 42204 7 1 2 42202 42203
0 42205 7 1 2 97315 42204
0 42206 5 1 1 42205
0 42207 7 1 2 42201 42206
0 42208 5 1 1 42207
0 42209 7 1 2 89749 42208
0 42210 5 1 1 42209
0 42211 7 1 2 42198 42210
0 42212 5 1 1 42211
0 42213 7 1 2 67729 42212
0 42214 5 1 1 42213
0 42215 7 1 2 42151 42214
0 42216 7 1 2 42111 42215
0 42217 7 1 2 41988 42216
0 42218 5 1 1 42217
0 42219 7 1 2 98507 42218
0 42220 5 1 1 42219
0 42221 7 1 2 41692 42220
0 42222 7 1 2 41100 42221
0 42223 7 1 2 38167 42222
0 42224 5 1 1 42223
0 42225 7 1 2 104320 42224
0 42226 5 1 1 42225
0 42227 7 1 2 37625 42226
0 42228 7 1 2 32991 42227
0 42229 7 1 2 30055 42228
0 42230 7 1 2 25995 42229
0 42231 5 1 1 42230
0 42232 7 1 2 99358 42231
0 42233 5 1 1 42232
0 42234 7 2 2 75935 97740
0 42235 5 2 1 105004
0 42236 7 1 2 101099 105006
0 42237 5 6 1 42236
0 42238 7 1 2 64461 105008
0 42239 5 1 1 42238
0 42240 7 1 2 99174 80995
0 42241 5 1 1 42240
0 42242 7 1 2 42239 42241
0 42243 5 1 1 42242
0 42244 7 1 2 69936 42243
0 42245 5 1 1 42244
0 42246 7 1 2 102040 104477
0 42247 5 1 1 42246
0 42248 7 1 2 42245 42247
0 42249 5 1 1 42248
0 42250 7 1 2 82323 42249
0 42251 5 1 1 42250
0 42252 7 1 2 96649 96258
0 42253 5 1 1 42252
0 42254 7 3 2 71139 80726
0 42255 7 1 2 103166 105014
0 42256 5 1 1 42255
0 42257 7 1 2 42253 42256
0 42258 5 1 1 42257
0 42259 7 1 2 69572 42258
0 42260 5 1 1 42259
0 42261 7 3 2 64462 81138
0 42262 7 2 2 97563 105017
0 42263 5 1 1 105020
0 42264 7 1 2 71456 105021
0 42265 5 1 1 42264
0 42266 7 1 2 42260 42265
0 42267 5 1 1 42266
0 42268 7 1 2 98116 42267
0 42269 5 1 1 42268
0 42270 7 1 2 42251 42269
0 42271 5 1 1 42270
0 42272 7 1 2 79147 42271
0 42273 5 1 1 42272
0 42274 7 1 2 65175 102238
0 42275 5 1 1 42274
0 42276 7 1 2 96653 98276
0 42277 5 1 1 42276
0 42278 7 1 2 42275 42277
0 42279 5 1 1 42278
0 42280 7 1 2 76606 42279
0 42281 5 1 1 42280
0 42282 7 1 2 98238 101518
0 42283 5 1 1 42282
0 42284 7 1 2 104579 42283
0 42285 5 1 1 42284
0 42286 7 1 2 80727 42285
0 42287 5 1 1 42286
0 42288 7 1 2 82324 99259
0 42289 5 1 1 42288
0 42290 7 1 2 65176 98277
0 42291 5 1 1 42290
0 42292 7 1 2 42289 42291
0 42293 5 1 1 42292
0 42294 7 1 2 73227 42293
0 42295 5 1 1 42294
0 42296 7 1 2 42287 42295
0 42297 7 1 2 42281 42296
0 42298 5 1 1 42297
0 42299 7 1 2 78878 42298
0 42300 5 1 1 42299
0 42301 7 1 2 67730 42300
0 42302 7 1 2 42273 42301
0 42303 5 1 1 42302
0 42304 7 1 2 80126 99175
0 42305 5 1 1 42304
0 42306 7 2 2 84965 99157
0 42307 7 1 2 73228 105022
0 42308 5 1 1 42307
0 42309 7 1 2 42305 42308
0 42310 5 1 1 42309
0 42311 7 1 2 65481 42310
0 42312 5 1 1 42311
0 42313 7 1 2 99176 94471
0 42314 5 1 1 42313
0 42315 7 1 2 105007 42314
0 42316 5 1 1 42315
0 42317 7 1 2 65177 42316
0 42318 5 1 1 42317
0 42319 7 1 2 42312 42318
0 42320 5 1 1 42319
0 42321 7 1 2 69937 42320
0 42322 5 1 1 42321
0 42323 7 1 2 97556 103508
0 42324 7 1 2 97235 42323
0 42325 5 1 1 42324
0 42326 7 1 2 42322 42325
0 42327 5 1 1 42326
0 42328 7 1 2 94913 42327
0 42329 5 1 1 42328
0 42330 7 1 2 97128 98902
0 42331 7 1 2 100007 42330
0 42332 7 1 2 104024 42331
0 42333 5 1 1 42332
0 42334 7 1 2 72733 42333
0 42335 7 1 2 42329 42334
0 42336 5 1 1 42335
0 42337 7 1 2 69238 42336
0 42338 7 1 2 42303 42337
0 42339 5 1 1 42338
0 42340 7 1 2 85476 42339
0 42341 5 1 1 42340
0 42342 7 2 2 68134 103905
0 42343 7 1 2 80728 79457
0 42344 5 1 1 42343
0 42345 7 4 2 71955 82325
0 42346 7 1 2 90720 87963
0 42347 7 1 2 105026 42346
0 42348 5 1 1 42347
0 42349 7 1 2 42344 42348
0 42350 5 1 1 42349
0 42351 7 1 2 67731 42350
0 42352 5 1 1 42351
0 42353 7 1 2 72734 104087
0 42354 7 1 2 105027 42353
0 42355 5 1 1 42354
0 42356 7 1 2 42352 42355
0 42357 5 1 1 42356
0 42358 7 1 2 71457 42357
0 42359 5 1 1 42358
0 42360 7 1 2 86323 92632
0 42361 7 1 2 103806 42360
0 42362 5 1 1 42361
0 42363 7 1 2 42359 42362
0 42364 5 1 1 42363
0 42365 7 1 2 105024 42364
0 42366 5 1 1 42365
0 42367 7 1 2 82501 42366
0 42368 5 1 1 42367
0 42369 7 1 2 68997 42368
0 42370 7 1 2 42341 42369
0 42371 5 1 1 42370
0 42372 7 2 2 74316 92411
0 42373 7 1 2 102244 74039
0 42374 7 1 2 105030 42373
0 42375 7 1 2 103742 42374
0 42376 5 1 1 42375
0 42377 7 1 2 42371 42376
0 42378 5 1 1 42377
0 42379 7 1 2 66587 42378
0 42380 5 1 1 42379
0 42381 7 1 2 69573 101943
0 42382 5 1 1 42381
0 42383 7 1 2 81534 102482
0 42384 5 1 1 42383
0 42385 7 1 2 42382 42384
0 42386 5 2 1 42385
0 42387 7 1 2 64836 105032
0 42388 5 1 1 42387
0 42389 7 2 2 92927 97465
0 42390 5 1 1 105034
0 42391 7 1 2 69574 105035
0 42392 5 1 1 42391
0 42393 7 1 2 42388 42392
0 42394 5 1 1 42393
0 42395 7 1 2 82991 42394
0 42396 5 1 1 42395
0 42397 7 3 2 72453 76960
0 42398 5 1 1 105036
0 42399 7 1 2 84744 104657
0 42400 7 1 2 105037 42399
0 42401 5 1 1 42400
0 42402 7 1 2 42396 42401
0 42403 5 1 1 42402
0 42404 7 1 2 79148 42403
0 42405 5 1 1 42404
0 42406 7 1 2 93467 99274
0 42407 5 1 1 42406
0 42408 7 1 2 101933 42407
0 42409 5 1 1 42408
0 42410 7 1 2 79665 83584
0 42411 7 1 2 42409 42410
0 42412 5 1 1 42411
0 42413 7 1 2 42405 42412
0 42414 5 1 1 42413
0 42415 7 1 2 66054 42414
0 42416 5 1 1 42415
0 42417 7 3 2 72735 79175
0 42418 5 1 1 105039
0 42419 7 1 2 90702 105040
0 42420 5 1 1 42419
0 42421 7 1 2 93013 104949
0 42422 5 1 1 42421
0 42423 7 1 2 101412 42422
0 42424 7 1 2 42420 42423
0 42425 5 1 1 42424
0 42426 7 1 2 90897 97220
0 42427 7 1 2 42425 42426
0 42428 5 1 1 42427
0 42429 7 1 2 42416 42428
0 42430 5 1 1 42429
0 42431 7 1 2 70860 42430
0 42432 5 1 1 42431
0 42433 7 2 2 74968 83997
0 42434 5 3 1 105042
0 42435 7 1 2 90772 105044
0 42436 5 2 1 42435
0 42437 7 1 2 69575 105047
0 42438 5 1 1 42437
0 42439 7 2 2 68695 81477
0 42440 5 1 1 105049
0 42441 7 1 2 78449 42440
0 42442 5 1 1 42441
0 42443 7 1 2 79176 42442
0 42444 5 1 1 42443
0 42445 7 1 2 42438 42444
0 42446 5 2 1 42445
0 42447 7 2 2 67380 92423
0 42448 7 1 2 94971 105053
0 42449 7 1 2 105051 42448
0 42450 5 1 1 42449
0 42451 7 1 2 42432 42450
0 42452 5 1 1 42451
0 42453 7 1 2 70236 42452
0 42454 5 1 1 42453
0 42455 7 1 2 101944 104906
0 42456 5 2 1 42455
0 42457 7 1 2 103562 93028
0 42458 5 1 1 42457
0 42459 7 1 2 105055 42458
0 42460 5 1 1 42459
0 42461 7 1 2 70861 42460
0 42462 5 1 1 42461
0 42463 7 2 2 93220 84295
0 42464 5 2 1 105057
0 42465 7 1 2 100789 105058
0 42466 5 1 1 42465
0 42467 7 1 2 42462 42466
0 42468 5 1 1 42467
0 42469 7 1 2 69938 42468
0 42470 5 1 1 42469
0 42471 7 3 2 87806 103563
0 42472 7 1 2 95510 80027
0 42473 7 1 2 105061 42472
0 42474 5 1 1 42473
0 42475 7 1 2 42470 42474
0 42476 5 1 1 42475
0 42477 7 1 2 78879 42476
0 42478 5 1 1 42477
0 42479 7 1 2 42454 42478
0 42480 5 1 1 42479
0 42481 7 1 2 69239 42480
0 42482 5 1 1 42481
0 42483 7 1 2 74558 105052
0 42484 5 1 1 42483
0 42485 7 1 2 7745 42484
0 42486 5 1 1 42485
0 42487 7 1 2 99463 94972
0 42488 7 1 2 42486 42487
0 42489 5 1 1 42488
0 42490 7 1 2 42482 42489
0 42491 5 1 1 42490
0 42492 7 1 2 70495 42491
0 42493 5 1 1 42492
0 42494 7 1 2 68696 102953
0 42495 7 1 2 86495 42494
0 42496 5 1 1 42495
0 42497 7 1 2 81911 79666
0 42498 5 1 1 42497
0 42499 7 1 2 42496 42498
0 42500 5 1 1 42499
0 42501 7 1 2 70237 42500
0 42502 5 1 1 42501
0 42503 7 1 2 76237 102308
0 42504 5 1 1 42503
0 42505 7 1 2 78880 42504
0 42506 5 1 1 42505
0 42507 7 1 2 42502 42506
0 42508 5 1 1 42507
0 42509 7 1 2 69576 42508
0 42510 5 1 1 42509
0 42511 7 1 2 76500 82308
0 42512 7 1 2 85373 42511
0 42513 5 1 1 42512
0 42514 7 1 2 42510 42513
0 42515 5 1 1 42514
0 42516 7 1 2 72736 42515
0 42517 5 1 1 42516
0 42518 7 1 2 101861 104066
0 42519 5 1 1 42518
0 42520 7 1 2 87964 79683
0 42521 7 1 2 103164 42520
0 42522 5 1 1 42521
0 42523 7 1 2 42519 42522
0 42524 5 1 1 42523
0 42525 7 2 2 67732 42524
0 42526 7 1 2 92928 105064
0 42527 5 1 1 42526
0 42528 7 1 2 42517 42527
0 42529 5 1 1 42528
0 42530 7 1 2 98440 42529
0 42531 5 1 1 42530
0 42532 7 5 2 72737 81912
0 42533 7 4 2 88380 105066
0 42534 7 1 2 99297 100016
0 42535 7 1 2 102969 42534
0 42536 7 1 2 105071 42535
0 42537 5 1 1 42536
0 42538 7 2 2 68697 95416
0 42539 7 2 2 90650 86611
0 42540 7 1 2 80467 105077
0 42541 7 1 2 105075 42540
0 42542 5 1 1 42541
0 42543 7 1 2 64837 105065
0 42544 5 1 1 42543
0 42545 7 1 2 42542 42544
0 42546 5 1 1 42545
0 42547 7 1 2 98508 76335
0 42548 7 1 2 42546 42547
0 42549 5 1 1 42548
0 42550 7 1 2 42537 42549
0 42551 7 1 2 42531 42550
0 42552 5 1 1 42551
0 42553 7 1 2 68135 42552
0 42554 5 1 1 42553
0 42555 7 1 2 97410 78881
0 42556 5 1 1 42555
0 42557 7 1 2 81268 83861
0 42558 5 10 1 42557
0 42559 7 2 2 91198 105079
0 42560 7 1 2 70641 96173
0 42561 7 1 2 105089 42560
0 42562 5 1 1 42561
0 42563 7 1 2 42556 42562
0 42564 5 1 1 42563
0 42565 7 1 2 70496 42564
0 42566 5 1 1 42565
0 42567 7 1 2 91805 85191
0 42568 7 1 2 105090 42567
0 42569 5 1 1 42568
0 42570 7 1 2 42566 42569
0 42571 5 1 1 42570
0 42572 7 1 2 87807 42571
0 42573 5 1 1 42572
0 42574 7 1 2 70497 80268
0 42575 7 1 2 83585 42574
0 42576 5 1 1 42575
0 42577 7 1 2 81913 93226
0 42578 5 1 1 42577
0 42579 7 1 2 42576 42578
0 42580 5 1 1 42579
0 42581 7 1 2 95420 42580
0 42582 5 1 1 42581
0 42583 7 1 2 42573 42582
0 42584 5 1 1 42583
0 42585 7 1 2 70238 42584
0 42586 5 1 1 42585
0 42587 7 2 2 81761 91450
0 42588 5 1 1 105091
0 42589 7 1 2 104658 105092
0 42590 5 2 1 42589
0 42591 7 1 2 76607 102309
0 42592 5 1 1 42591
0 42593 7 1 2 89234 42592
0 42594 5 1 1 42593
0 42595 7 1 2 95021 42594
0 42596 5 1 1 42595
0 42597 7 1 2 69577 42596
0 42598 5 1 1 42597
0 42599 7 1 2 105093 42598
0 42600 5 1 1 42599
0 42601 7 1 2 78882 42600
0 42602 5 1 1 42601
0 42603 7 1 2 42586 42602
0 42604 5 1 1 42603
0 42605 7 1 2 98441 42604
0 42606 5 1 1 42605
0 42607 7 1 2 91831 80203
0 42608 7 1 2 80269 42607
0 42609 7 1 2 97229 105078
0 42610 7 1 2 42608 42609
0 42611 5 1 1 42610
0 42612 7 1 2 42606 42611
0 42613 7 1 2 42554 42612
0 42614 5 1 1 42613
0 42615 7 1 2 69240 42614
0 42616 5 1 1 42615
0 42617 7 3 2 97720 78996
0 42618 7 1 2 80028 105095
0 42619 5 1 1 42618
0 42620 7 1 2 78181 76978
0 42621 7 1 2 103510 42620
0 42622 5 1 1 42621
0 42623 7 1 2 42619 42622
0 42624 5 1 1 42623
0 42625 7 1 2 72738 42624
0 42626 5 1 1 42625
0 42627 7 3 2 67733 76809
0 42628 7 1 2 79413 79114
0 42629 7 1 2 105098 42628
0 42630 5 1 1 42629
0 42631 7 1 2 42626 42630
0 42632 5 1 1 42631
0 42633 7 1 2 80642 42632
0 42634 5 1 1 42633
0 42635 7 1 2 83804 84677
0 42636 7 1 2 95437 42635
0 42637 5 1 1 42636
0 42638 7 1 2 42634 42637
0 42639 5 1 1 42638
0 42640 7 1 2 71458 42639
0 42641 5 1 1 42640
0 42642 7 1 2 64463 82745
0 42643 5 2 1 42642
0 42644 7 1 2 95183 95421
0 42645 7 1 2 105101 42644
0 42646 5 1 1 42645
0 42647 7 1 2 42641 42646
0 42648 5 1 1 42647
0 42649 7 1 2 70239 42648
0 42650 5 1 1 42649
0 42651 7 3 2 68136 98912
0 42652 7 1 2 78322 79531
0 42653 7 1 2 105103 42652
0 42654 5 1 1 42653
0 42655 7 1 2 42650 42654
0 42656 5 1 1 42655
0 42657 7 1 2 102301 42656
0 42658 5 1 1 42657
0 42659 7 1 2 42616 42658
0 42660 5 1 1 42659
0 42661 7 1 2 71140 42660
0 42662 5 1 1 42661
0 42663 7 1 2 85024 79669
0 42664 5 1 1 42663
0 42665 7 1 2 74906 104889
0 42666 7 1 2 79526 42665
0 42667 5 1 1 42666
0 42668 7 1 2 42664 42667
0 42669 5 1 1 42668
0 42670 7 1 2 71459 42669
0 42671 5 1 1 42670
0 42672 7 1 2 87928 90992
0 42673 7 1 2 79686 42672
0 42674 5 1 1 42673
0 42675 7 1 2 42671 42674
0 42676 5 1 1 42675
0 42677 7 1 2 99275 42676
0 42678 5 1 1 42677
0 42679 7 1 2 82404 97166
0 42680 5 1 1 42679
0 42681 7 1 2 83909 101155
0 42682 5 1 1 42681
0 42683 7 1 2 42680 42682
0 42684 5 1 1 42683
0 42685 7 3 2 64838 71956
0 42686 7 1 2 79687 105106
0 42687 7 1 2 42684 42686
0 42688 5 1 1 42687
0 42689 7 1 2 42678 42688
0 42690 5 1 1 42689
0 42691 7 1 2 69578 42690
0 42692 5 1 1 42691
0 42693 7 2 2 90876 98224
0 42694 5 1 1 105109
0 42695 7 2 2 86091 85107
0 42696 7 1 2 84185 105111
0 42697 7 1 2 105110 42696
0 42698 5 1 1 42697
0 42699 7 1 2 42692 42698
0 42700 5 1 1 42699
0 42701 7 1 2 69241 102354
0 42702 7 1 2 42700 42701
0 42703 5 1 1 42702
0 42704 7 1 2 42662 42703
0 42705 7 1 2 42493 42704
0 42706 5 1 1 42705
0 42707 7 1 2 68998 42706
0 42708 5 1 1 42707
0 42709 7 1 2 42380 42708
0 42710 5 1 1 42709
0 42711 7 1 2 73857 42710
0 42712 5 1 1 42711
0 42713 7 1 2 39548 92652
0 42714 5 1 1 42713
0 42715 7 1 2 95022 42714
0 42716 5 1 1 42715
0 42717 7 1 2 69579 42716
0 42718 5 1 1 42717
0 42719 7 1 2 71851 80270
0 42720 7 1 2 97659 42719
0 42721 5 1 1 42720
0 42722 7 1 2 93229 42721
0 42723 5 1 1 42722
0 42724 7 1 2 72739 42723
0 42725 5 1 1 42724
0 42726 7 1 2 103167 98913
0 42727 5 1 1 42726
0 42728 7 1 2 42725 42727
0 42729 5 1 1 42728
0 42730 7 1 2 68137 42729
0 42731 5 1 1 42730
0 42732 7 1 2 105094 42731
0 42733 7 1 2 42718 42732
0 42734 5 1 1 42733
0 42735 7 1 2 71141 42734
0 42736 5 1 1 42735
0 42737 7 1 2 75427 103689
0 42738 7 1 2 90760 42737
0 42739 5 1 1 42738
0 42740 7 1 2 42736 42739
0 42741 5 1 1 42740
0 42742 7 1 2 72454 42741
0 42743 5 1 1 42742
0 42744 7 1 2 97301 92505
0 42745 5 1 1 42744
0 42746 7 1 2 78415 42745
0 42747 5 1 1 42746
0 42748 7 2 2 80367 92190
0 42749 5 1 1 105113
0 42750 7 1 2 71690 105114
0 42751 5 1 1 42750
0 42752 7 1 2 42747 42751
0 42753 5 1 1 42752
0 42754 7 1 2 69580 42753
0 42755 5 1 1 42754
0 42756 7 1 2 77088 93164
0 42757 5 1 1 42756
0 42758 7 1 2 101398 42757
0 42759 5 1 1 42758
0 42760 7 1 2 92503 42759
0 42761 5 1 1 42760
0 42762 7 1 2 42755 42761
0 42763 5 1 1 42762
0 42764 7 1 2 72455 42763
0 42765 5 1 1 42764
0 42766 7 1 2 80368 100417
0 42767 7 1 2 93496 42766
0 42768 5 1 1 42767
0 42769 7 1 2 42765 42768
0 42770 5 1 1 42769
0 42771 7 1 2 70240 42770
0 42772 5 1 1 42771
0 42773 7 2 2 75983 78416
0 42774 7 1 2 80500 105115
0 42775 5 1 1 42774
0 42776 7 1 2 77715 101394
0 42777 5 1 1 42776
0 42778 7 1 2 42775 42777
0 42779 5 1 1 42778
0 42780 7 1 2 98614 42779
0 42781 5 1 1 42780
0 42782 7 1 2 97682 91047
0 42783 5 1 1 42782
0 42784 7 1 2 99146 42783
0 42785 5 1 1 42784
0 42786 7 1 2 80369 42785
0 42787 5 1 1 42786
0 42788 7 2 2 71142 93014
0 42789 5 1 1 105117
0 42790 7 1 2 70241 105118
0 42791 5 1 1 42790
0 42792 7 2 2 72740 89452
0 42793 5 1 1 105119
0 42794 7 1 2 90773 42793
0 42795 5 1 1 42794
0 42796 7 1 2 78062 42795
0 42797 5 1 1 42796
0 42798 7 1 2 42791 42797
0 42799 7 1 2 42787 42798
0 42800 5 1 1 42799
0 42801 7 1 2 72456 42800
0 42802 5 1 1 42801
0 42803 7 1 2 105056 42802
0 42804 5 1 1 42803
0 42805 7 1 2 69939 42804
0 42806 5 1 1 42805
0 42807 7 1 2 42781 42806
0 42808 7 1 2 42772 42807
0 42809 5 1 1 42808
0 42810 7 1 2 70498 42809
0 42811 5 1 1 42810
0 42812 7 1 2 42743 42811
0 42813 5 1 1 42812
0 42814 7 1 2 69242 42813
0 42815 5 1 1 42814
0 42816 7 1 2 85477 42815
0 42817 5 1 1 42816
0 42818 7 1 2 75630 101067
0 42819 5 1 1 42818
0 42820 7 1 2 103664 42819
0 42821 5 1 1 42820
0 42822 7 1 2 74559 42821
0 42823 5 1 1 42822
0 42824 7 1 2 67734 90502
0 42825 5 1 1 42824
0 42826 7 1 2 42823 42825
0 42827 5 1 1 42826
0 42828 7 1 2 80643 42827
0 42829 5 1 1 42828
0 42830 7 1 2 100560 105104
0 42831 5 1 1 42830
0 42832 7 1 2 42829 42831
0 42833 5 1 1 42832
0 42834 7 1 2 71460 42833
0 42835 5 1 1 42834
0 42836 7 1 2 101159 81333
0 42837 5 1 1 42836
0 42838 7 1 2 67735 42837
0 42839 5 1 1 42838
0 42840 7 1 2 91617 83998
0 42841 5 1 1 42840
0 42842 7 1 2 42839 42841
0 42843 5 1 1 42842
0 42844 7 1 2 102439 42843
0 42845 5 1 1 42844
0 42846 7 1 2 42835 42845
0 42847 5 1 1 42846
0 42848 7 1 2 67381 42847
0 42849 5 1 1 42848
0 42850 7 1 2 82502 42849
0 42851 5 1 1 42850
0 42852 7 1 2 90345 42851
0 42853 7 1 2 42817 42852
0 42854 5 1 1 42853
0 42855 7 2 2 93015 84411
0 42856 5 1 1 105121
0 42857 7 1 2 92773 104659
0 42858 5 1 1 42857
0 42859 7 1 2 42856 42858
0 42860 5 1 1 42859
0 42861 7 1 2 69581 42860
0 42862 5 1 1 42861
0 42863 7 2 2 85084 78382
0 42864 5 1 1 105123
0 42865 7 1 2 78746 105124
0 42866 5 1 1 42865
0 42867 7 1 2 42862 42866
0 42868 5 2 1 42867
0 42869 7 1 2 84851 105125
0 42870 5 1 1 42869
0 42871 7 3 2 101519 81055
0 42872 7 1 2 103328 105127
0 42873 5 1 1 42872
0 42874 7 1 2 42870 42873
0 42875 5 1 1 42874
0 42876 7 1 2 68698 42875
0 42877 5 1 1 42876
0 42878 7 1 2 101086 105128
0 42879 5 1 1 42878
0 42880 7 1 2 42877 42879
0 42881 5 1 1 42880
0 42882 7 1 2 72457 42881
0 42883 5 1 1 42882
0 42884 7 3 2 86064 84678
0 42885 7 1 2 66055 99168
0 42886 7 1 2 105130 42885
0 42887 5 1 1 42886
0 42888 7 1 2 42883 42887
0 42889 5 1 1 42888
0 42890 7 1 2 70862 42889
0 42891 5 1 1 42890
0 42892 7 1 2 74969 103906
0 42893 7 2 2 105131 42892
0 42894 7 1 2 92341 105133
0 42895 5 1 1 42894
0 42896 7 1 2 42891 42895
0 42897 5 1 1 42896
0 42898 7 1 2 69243 42897
0 42899 5 1 1 42898
0 42900 7 1 2 103740 105134
0 42901 5 1 1 42900
0 42902 7 1 2 42899 42901
0 42903 5 1 1 42902
0 42904 7 1 2 94083 105112
0 42905 7 1 2 42903 42904
0 42906 5 1 1 42905
0 42907 7 1 2 42854 42906
0 42908 5 1 1 42907
0 42909 7 1 2 63910 42908
0 42910 5 1 1 42909
0 42911 7 1 2 100008 89265
0 42912 7 1 2 90346 42911
0 42913 5 1 1 42912
0 42914 7 1 2 67382 42913
0 42915 5 1 1 42914
0 42916 7 6 2 78182 89582
0 42917 5 1 1 105135
0 42918 7 2 2 68878 88985
0 42919 5 1 1 105141
0 42920 7 1 2 42917 42919
0 42921 5 1 1 42920
0 42922 7 1 2 80370 89745
0 42923 5 1 1 42922
0 42924 7 1 2 32293 42923
0 42925 5 1 1 42924
0 42926 7 1 2 68138 42925
0 42927 5 1 1 42926
0 42928 7 1 2 76501 95032
0 42929 5 1 1 42928
0 42930 7 1 2 42927 42929
0 42931 5 1 1 42930
0 42932 7 1 2 42921 42931
0 42933 5 1 1 42932
0 42934 7 5 2 68879 88077
0 42935 7 1 2 68139 82326
0 42936 5 1 1 42935
0 42937 7 1 2 15430 42936
0 42938 5 1 1 42937
0 42939 7 1 2 105080 42938
0 42940 5 1 1 42939
0 42941 7 1 2 80729 88000
0 42942 7 1 2 101167 42941
0 42943 5 1 1 42942
0 42944 7 1 2 42940 42943
0 42945 5 1 1 42944
0 42946 7 1 2 105143 42945
0 42947 5 1 1 42946
0 42948 7 1 2 42933 42947
0 42949 5 1 1 42948
0 42950 7 1 2 67736 42949
0 42951 5 1 1 42950
0 42952 7 1 2 83505 83974
0 42953 5 2 1 42952
0 42954 7 1 2 65178 100753
0 42955 5 1 1 42954
0 42956 7 1 2 105148 42955
0 42957 5 1 1 42956
0 42958 7 4 2 94234 91171
0 42959 7 1 2 97721 81967
0 42960 7 1 2 92315 42959
0 42961 7 1 2 105150 42960
0 42962 7 1 2 42957 42961
0 42963 5 1 1 42962
0 42964 7 1 2 72458 42963
0 42965 7 1 2 42951 42964
0 42966 5 1 1 42965
0 42967 7 1 2 42915 42966
0 42968 5 1 1 42967
0 42969 7 1 2 71143 42968
0 42970 5 1 1 42969
0 42971 7 1 2 82327 105033
0 42972 5 1 1 42971
0 42973 7 1 2 84165 104138
0 42974 7 1 2 97344 42973
0 42975 5 1 1 42974
0 42976 7 1 2 42972 42975
0 42977 5 1 1 42976
0 42978 7 1 2 94639 42977
0 42979 5 1 1 42978
0 42980 7 1 2 80166 98764
0 42981 7 2 2 96654 42980
0 42982 7 3 2 89546 96251
0 42983 7 4 2 77908 105156
0 42984 7 1 2 105154 105159
0 42985 5 1 1 42984
0 42986 7 1 2 42979 42985
0 42987 5 1 1 42986
0 42988 7 1 2 68880 42987
0 42989 5 1 1 42988
0 42990 7 1 2 64464 105155
0 42991 7 1 2 105136 42990
0 42992 5 1 1 42991
0 42993 7 1 2 66056 42992
0 42994 7 1 2 42989 42993
0 42995 5 1 1 42994
0 42996 7 1 2 69244 42995
0 42997 7 1 2 42970 42996
0 42998 5 1 1 42997
0 42999 7 1 2 85478 42998
0 43000 5 1 1 42999
0 43001 7 4 2 94074 90317
0 43002 5 1 1 105163
0 43003 7 1 2 101862 105164
0 43004 5 1 1 43003
0 43005 7 1 2 64465 91929
0 43006 7 1 2 105028 43005
0 43007 5 1 1 43006
0 43008 7 1 2 43004 43007
0 43009 5 1 1 43008
0 43010 7 1 2 67737 43009
0 43011 5 1 1 43010
0 43012 7 1 2 81478 91930
0 43013 7 1 2 105029 43012
0 43014 5 1 1 43013
0 43015 7 1 2 43011 43014
0 43016 5 1 1 43015
0 43017 7 1 2 68881 43016
0 43018 5 1 1 43017
0 43019 7 1 2 64839 98914
0 43020 7 1 2 105137 43019
0 43021 5 1 1 43020
0 43022 7 1 2 43018 43021
0 43023 5 1 1 43022
0 43024 7 1 2 71461 43023
0 43025 5 1 1 43024
0 43026 7 2 2 67738 90336
0 43027 7 1 2 78323 98887
0 43028 7 1 2 105167 43027
0 43029 5 1 1 43028
0 43030 7 1 2 43025 43029
0 43031 5 1 1 43030
0 43032 7 1 2 105025 43031
0 43033 5 1 1 43032
0 43034 7 1 2 82503 43033
0 43035 5 1 1 43034
0 43036 7 1 2 63911 43035
0 43037 7 1 2 43000 43036
0 43038 5 1 1 43037
0 43039 7 1 2 84323 84463
0 43040 7 1 2 105031 43039
0 43041 7 1 2 103743 43040
0 43042 7 1 2 90337 43041
0 43043 5 1 1 43042
0 43044 7 1 2 43038 43043
0 43045 5 1 1 43044
0 43046 7 1 2 66588 43045
0 43047 5 1 1 43046
0 43048 7 1 2 42910 43047
0 43049 7 1 2 42712 43048
0 43050 5 1 1 43049
0 43051 7 1 2 73558 43050
0 43052 5 1 1 43051
0 43053 7 1 2 70242 104227
0 43054 5 1 1 43053
0 43055 7 1 2 12053 43054
0 43056 5 2 1 43055
0 43057 7 1 2 90044 105169
0 43058 5 1 1 43057
0 43059 7 1 2 70499 80453
0 43060 5 1 1 43059
0 43061 7 1 2 87703 101367
0 43062 7 1 2 43060 43061
0 43063 5 1 1 43062
0 43064 7 1 2 77543 43063
0 43065 5 1 1 43064
0 43066 7 1 2 43058 43065
0 43067 5 1 1 43066
0 43068 7 1 2 103668 43067
0 43069 5 1 1 43068
0 43070 7 1 2 78598 76419
0 43071 5 1 1 43070
0 43072 7 1 2 90021 43071
0 43073 5 1 1 43072
0 43074 7 1 2 75428 43073
0 43075 5 1 1 43074
0 43076 7 2 2 65482 95048
0 43077 5 1 1 105171
0 43078 7 1 2 81285 100887
0 43079 7 2 2 105172 43078
0 43080 5 1 1 105173
0 43081 7 1 2 43075 43080
0 43082 5 1 1 43081
0 43083 7 1 2 68140 43082
0 43084 5 1 1 43083
0 43085 7 1 2 75694 94939
0 43086 5 1 1 43085
0 43087 7 1 2 43084 43086
0 43088 5 1 1 43087
0 43089 7 1 2 72741 43088
0 43090 5 1 1 43089
0 43091 7 1 2 87816 105045
0 43092 5 2 1 43091
0 43093 7 1 2 66057 105175
0 43094 5 1 1 43093
0 43095 7 2 2 75429 75695
0 43096 5 1 1 105177
0 43097 7 1 2 97297 105178
0 43098 5 1 1 43097
0 43099 7 1 2 70500 43098
0 43100 7 1 2 43094 43099
0 43101 5 1 1 43100
0 43102 7 1 2 92741 92758
0 43103 5 1 1 43102
0 43104 7 1 2 65483 43103
0 43105 5 1 1 43104
0 43106 7 1 2 71852 43105
0 43107 7 1 2 43101 43106
0 43108 5 1 1 43107
0 43109 7 1 2 43090 43108
0 43110 5 1 1 43109
0 43111 7 1 2 69940 43110
0 43112 5 1 1 43111
0 43113 7 1 2 83975 104798
0 43114 5 1 1 43113
0 43115 7 1 2 100897 96529
0 43116 5 1 1 43115
0 43117 7 1 2 43114 43116
0 43118 5 1 1 43117
0 43119 7 1 2 71853 43118
0 43120 5 1 1 43119
0 43121 7 1 2 71144 95049
0 43122 5 1 1 43121
0 43123 7 1 2 77115 75696
0 43124 5 1 1 43123
0 43125 7 1 2 43122 43124
0 43126 5 1 1 43125
0 43127 7 1 2 65484 43126
0 43128 5 1 1 43127
0 43129 7 2 2 70501 94472
0 43130 5 1 1 105179
0 43131 7 1 2 68474 105180
0 43132 5 1 1 43131
0 43133 7 1 2 43128 43132
0 43134 5 1 1 43133
0 43135 7 1 2 72742 43134
0 43136 5 1 1 43135
0 43137 7 1 2 43120 43136
0 43138 5 1 1 43137
0 43139 7 1 2 68141 43138
0 43140 5 1 1 43139
0 43141 7 1 2 87182 105116
0 43142 5 1 1 43141
0 43143 7 1 2 71854 90763
0 43144 5 1 1 43143
0 43145 7 1 2 105046 43144
0 43146 5 1 1 43145
0 43147 7 1 2 64840 43146
0 43148 5 1 1 43147
0 43149 7 1 2 88712 78422
0 43150 5 1 1 43149
0 43151 7 1 2 79736 14465
0 43152 7 1 2 43150 43151
0 43153 5 1 1 43152
0 43154 7 1 2 70502 43153
0 43155 7 1 2 43148 43154
0 43156 5 1 1 43155
0 43157 7 2 2 80371 74970
0 43158 5 1 1 105181
0 43159 7 1 2 27168 43158
0 43160 5 1 1 43159
0 43161 7 1 2 72743 43160
0 43162 5 1 1 43161
0 43163 7 1 2 65485 42749
0 43164 7 1 2 43162 43163
0 43165 5 1 1 43164
0 43166 7 1 2 68475 43165
0 43167 7 1 2 43156 43166
0 43168 5 1 1 43167
0 43169 7 1 2 43142 43168
0 43170 5 1 1 43169
0 43171 7 1 2 75430 43170
0 43172 5 1 1 43171
0 43173 7 1 2 77116 90764
0 43174 5 1 1 43173
0 43175 7 3 2 71145 81420
0 43176 5 1 1 105183
0 43177 7 1 2 81286 105184
0 43178 5 1 1 43177
0 43179 7 1 2 43174 43178
0 43180 5 1 1 43179
0 43181 7 1 2 84852 43180
0 43182 5 1 1 43181
0 43183 7 1 2 72744 105174
0 43184 5 1 1 43183
0 43185 7 1 2 103577 43184
0 43186 5 1 1 43185
0 43187 7 1 2 71146 43186
0 43188 5 1 1 43187
0 43189 7 1 2 43182 43188
0 43190 7 1 2 43172 43189
0 43191 7 1 2 43140 43190
0 43192 7 1 2 43112 43191
0 43193 5 1 1 43192
0 43194 7 1 2 69582 43193
0 43195 5 1 1 43194
0 43196 7 1 2 94987 43077
0 43197 5 1 1 43196
0 43198 7 1 2 90942 43197
0 43199 5 1 1 43198
0 43200 7 1 2 84798 86755
0 43201 5 1 1 43200
0 43202 7 1 2 90943 43201
0 43203 5 1 1 43202
0 43204 7 1 2 988 43203
0 43205 5 1 1 43204
0 43206 7 1 2 75431 43205
0 43207 5 1 1 43206
0 43208 7 1 2 65486 1882
0 43209 5 1 1 43208
0 43210 7 1 2 70503 84718
0 43211 5 1 1 43210
0 43212 7 1 2 81311 43211
0 43213 7 1 2 43209 43212
0 43214 5 1 1 43213
0 43215 7 1 2 43207 43214
0 43216 7 1 2 43199 43215
0 43217 5 1 1 43216
0 43218 7 1 2 72745 43217
0 43219 5 1 1 43218
0 43220 7 1 2 74689 105048
0 43221 5 1 1 43220
0 43222 7 1 2 64466 105176
0 43223 5 1 1 43222
0 43224 7 1 2 64467 43096
0 43225 5 1 1 43224
0 43226 7 1 2 97298 43225
0 43227 5 1 1 43226
0 43228 7 1 2 43223 43227
0 43229 7 1 2 43221 43228
0 43230 5 1 1 43229
0 43231 7 1 2 70504 43230
0 43232 5 1 1 43231
0 43233 7 1 2 68699 82031
0 43234 5 1 1 43233
0 43235 7 1 2 7721 43234
0 43236 5 1 1 43235
0 43237 7 1 2 68476 43236
0 43238 5 1 1 43237
0 43239 7 1 2 90939 43238
0 43240 5 1 1 43239
0 43241 7 1 2 86274 96530
0 43242 7 1 2 43240 43241
0 43243 5 1 1 43242
0 43244 7 1 2 43232 43243
0 43245 5 1 1 43244
0 43246 7 1 2 71855 43245
0 43247 5 1 1 43246
0 43248 7 1 2 43219 43247
0 43249 5 1 1 43248
0 43250 7 1 2 71147 43249
0 43251 5 1 1 43250
0 43252 7 2 2 74971 87127
0 43253 5 1 1 105186
0 43254 7 3 2 64468 95271
0 43255 5 1 1 105188
0 43256 7 1 2 105187 105189
0 43257 5 1 1 43256
0 43258 7 1 2 103692 2947
0 43259 5 1 1 43258
0 43260 7 1 2 78705 43259
0 43261 5 1 1 43260
0 43262 7 1 2 82391 98953
0 43263 5 1 1 43262
0 43264 7 1 2 77614 90453
0 43265 5 1 1 43264
0 43266 7 1 2 43263 43265
0 43267 7 1 2 43261 43266
0 43268 5 1 1 43267
0 43269 7 1 2 71462 43268
0 43270 5 1 1 43269
0 43271 7 1 2 66058 87833
0 43272 5 1 1 43271
0 43273 7 1 2 81334 43272
0 43274 5 1 1 43273
0 43275 7 1 2 84186 43274
0 43276 5 1 1 43275
0 43277 7 1 2 43270 43276
0 43278 5 1 1 43277
0 43279 7 1 2 84853 43278
0 43280 5 1 1 43279
0 43281 7 1 2 43257 43280
0 43282 7 1 2 43251 43281
0 43283 5 1 1 43282
0 43284 7 1 2 69941 43283
0 43285 5 1 1 43284
0 43286 7 1 2 101064 103859
0 43287 5 1 1 43286
0 43288 7 1 2 78467 43287
0 43289 5 1 1 43288
0 43290 7 1 2 75984 43289
0 43291 5 1 1 43290
0 43292 7 1 2 90765 94962
0 43293 5 1 1 43292
0 43294 7 1 2 43291 43293
0 43295 5 1 1 43294
0 43296 7 1 2 69942 43295
0 43297 5 1 1 43296
0 43298 7 5 2 71148 74972
0 43299 7 1 2 81479 105191
0 43300 5 1 1 43299
0 43301 7 1 2 84414 81167
0 43302 5 1 1 43301
0 43303 7 1 2 69583 43302
0 43304 5 1 1 43303
0 43305 7 1 2 68477 96028
0 43306 5 1 1 43305
0 43307 7 1 2 79254 43306
0 43308 5 1 1 43307
0 43309 7 1 2 98941 43308
0 43310 5 1 1 43309
0 43311 7 1 2 43304 43310
0 43312 5 1 1 43311
0 43313 7 1 2 67739 43312
0 43314 5 1 1 43313
0 43315 7 1 2 43300 43314
0 43316 7 1 2 43297 43315
0 43317 5 1 1 43316
0 43318 7 1 2 80730 43317
0 43319 5 1 1 43318
0 43320 7 1 2 95085 81535
0 43321 5 1 1 43320
0 43322 7 1 2 76420 97281
0 43323 7 1 2 88787 43322
0 43324 5 1 1 43323
0 43325 7 1 2 43321 43324
0 43326 5 1 1 43325
0 43327 7 1 2 98942 43326
0 43328 5 1 1 43327
0 43329 7 1 2 80904 76942
0 43330 7 1 2 97783 43329
0 43331 7 1 2 89374 43330
0 43332 5 1 1 43331
0 43333 7 1 2 43328 43332
0 43334 7 1 2 43319 43333
0 43335 7 1 2 43285 43334
0 43336 7 1 2 43195 43335
0 43337 5 1 1 43336
0 43338 7 1 2 67383 43337
0 43339 5 1 1 43338
0 43340 7 1 2 43069 43339
0 43341 5 2 1 43340
0 43342 7 1 2 78883 105196
0 43343 5 1 1 43342
0 43344 7 3 2 83329 97282
0 43345 5 1 1 105198
0 43346 7 2 2 4037 43345
0 43347 5 1 1 105201
0 43348 7 1 2 64469 105202
0 43349 5 1 1 43348
0 43350 7 1 2 69584 40278
0 43351 5 1 1 43350
0 43352 7 1 2 67384 43351
0 43353 7 1 2 43349 43352
0 43354 5 1 1 43353
0 43355 7 1 2 91432 97075
0 43356 5 1 1 43355
0 43357 7 1 2 43354 43356
0 43358 5 1 1 43357
0 43359 7 1 2 105192 43358
0 43360 5 1 1 43359
0 43361 7 1 2 76961 99987
0 43362 7 1 2 101077 43361
0 43363 5 1 1 43362
0 43364 7 1 2 43360 43363
0 43365 5 1 1 43364
0 43366 7 1 2 86065 43365
0 43367 5 1 1 43366
0 43368 7 4 2 67385 84679
0 43369 7 2 2 76421 94473
0 43370 7 1 2 101667 105207
0 43371 7 1 2 105203 43370
0 43372 5 1 1 43371
0 43373 7 1 2 43367 43372
0 43374 5 1 1 43373
0 43375 7 1 2 68478 43374
0 43376 5 1 1 43375
0 43377 7 1 2 81985 99950
0 43378 7 1 2 87071 43377
0 43379 7 1 2 105204 43378
0 43380 5 1 1 43379
0 43381 7 1 2 43376 43380
0 43382 5 2 1 43381
0 43383 7 1 2 79149 105209
0 43384 5 1 1 43383
0 43385 7 1 2 43343 43384
0 43386 5 1 1 43385
0 43387 7 1 2 85540 43386
0 43388 5 1 1 43387
0 43389 7 1 2 86679 92669
0 43390 5 2 1 43389
0 43391 7 1 2 67740 95225
0 43392 5 1 1 43391
0 43393 7 1 2 105211 43392
0 43394 5 1 1 43393
0 43395 7 1 2 64470 43394
0 43396 5 1 1 43395
0 43397 7 1 2 83057 100754
0 43398 5 1 1 43397
0 43399 7 1 2 100071 43398
0 43400 5 1 1 43399
0 43401 7 1 2 75432 43400
0 43402 5 1 1 43401
0 43403 7 1 2 84792 91744
0 43404 5 1 1 43403
0 43405 7 1 2 80041 43404
0 43406 7 1 2 43402 43405
0 43407 5 1 1 43406
0 43408 7 1 2 93095 43407
0 43409 5 1 1 43408
0 43410 7 1 2 43396 43409
0 43411 5 1 1 43410
0 43412 7 1 2 73229 43411
0 43413 5 1 1 43412
0 43414 7 1 2 81145 88649
0 43415 5 1 1 43414
0 43416 7 1 2 78956 82138
0 43417 5 1 1 43416
0 43418 7 1 2 43415 43417
0 43419 5 1 1 43418
0 43420 7 1 2 64471 43419
0 43421 5 1 1 43420
0 43422 7 1 2 79967 84680
0 43423 5 1 1 43422
0 43424 7 1 2 64472 105041
0 43425 5 1 1 43424
0 43426 7 1 2 43423 43425
0 43427 5 1 1 43426
0 43428 7 1 2 80731 43427
0 43429 5 1 1 43428
0 43430 7 1 2 43421 43429
0 43431 7 1 2 43413 43430
0 43432 5 1 1 43431
0 43433 7 1 2 66059 43432
0 43434 5 1 1 43433
0 43435 7 1 2 87886 90940
0 43436 7 1 2 105015 43435
0 43437 5 1 1 43436
0 43438 7 1 2 81158 92289
0 43439 5 1 1 43438
0 43440 7 1 2 67386 43439
0 43441 7 1 2 43437 43440
0 43442 7 1 2 43434 43441
0 43443 5 1 1 43442
0 43444 7 1 2 86985 83837
0 43445 5 1 1 43444
0 43446 7 1 2 90019 101888
0 43447 5 1 1 43446
0 43448 7 1 2 69943 43447
0 43449 5 1 1 43448
0 43450 7 1 2 71463 101587
0 43451 5 1 1 43450
0 43452 7 1 2 43449 43451
0 43453 5 1 1 43452
0 43454 7 1 2 73230 43453
0 43455 5 1 1 43454
0 43456 7 1 2 99623 94385
0 43457 5 1 1 43456
0 43458 7 1 2 64841 81441
0 43459 7 1 2 43457 43458
0 43460 5 1 1 43459
0 43461 7 1 2 43455 43460
0 43462 5 1 1 43461
0 43463 7 1 2 65179 43462
0 43464 5 1 1 43463
0 43465 7 1 2 85996 33600
0 43466 5 1 1 43465
0 43467 7 1 2 69585 43466
0 43468 5 1 1 43467
0 43469 7 1 2 75433 76032
0 43470 5 1 1 43469
0 43471 7 1 2 103481 43470
0 43472 5 1 1 43471
0 43473 7 1 2 84793 43472
0 43474 5 1 1 43473
0 43475 7 1 2 43468 43474
0 43476 5 1 1 43475
0 43477 7 1 2 64842 43476
0 43478 5 1 1 43477
0 43479 7 1 2 80732 90045
0 43480 5 1 1 43479
0 43481 7 1 2 86680 101126
0 43482 5 1 1 43481
0 43483 7 1 2 43480 43482
0 43484 5 1 1 43483
0 43485 7 1 2 64473 43484
0 43486 5 1 1 43485
0 43487 7 1 2 67741 43486
0 43488 7 1 2 43478 43487
0 43489 7 1 2 43464 43488
0 43490 5 1 1 43489
0 43491 7 1 2 64843 81625
0 43492 5 1 1 43491
0 43493 7 1 2 519 43492
0 43494 5 1 1 43493
0 43495 7 1 2 68142 43494
0 43496 5 1 1 43495
0 43497 7 2 2 76660 81239
0 43498 5 1 1 105213
0 43499 7 1 2 43496 43498
0 43500 5 1 1 43499
0 43501 7 1 2 81914 43500
0 43502 5 1 1 43501
0 43503 7 1 2 74690 90877
0 43504 5 1 1 43503
0 43505 7 1 2 69586 43504
0 43506 5 1 1 43505
0 43507 7 1 2 99879 43506
0 43508 5 2 1 43507
0 43509 7 1 2 95025 105215
0 43510 5 1 1 43509
0 43511 7 1 2 81762 81552
0 43512 5 1 1 43511
0 43513 7 1 2 99952 81252
0 43514 5 1 1 43513
0 43515 7 1 2 86681 43514
0 43516 5 1 1 43515
0 43517 7 1 2 43512 43516
0 43518 5 1 1 43517
0 43519 7 1 2 75434 43518
0 43520 5 1 1 43519
0 43521 7 1 2 43510 43520
0 43522 7 1 2 43502 43521
0 43523 5 1 1 43522
0 43524 7 1 2 68479 43523
0 43525 5 1 1 43524
0 43526 7 1 2 74827 91479
0 43527 5 1 1 43526
0 43528 7 1 2 102156 43527
0 43529 5 1 1 43528
0 43530 7 1 2 81763 43529
0 43531 5 1 1 43530
0 43532 7 2 2 80372 79259
0 43533 5 1 1 105217
0 43534 7 1 2 80900 105218
0 43535 5 1 1 43534
0 43536 7 1 2 72746 43535
0 43537 7 1 2 43531 43536
0 43538 7 1 2 43525 43537
0 43539 5 1 1 43538
0 43540 7 1 2 43490 43539
0 43541 5 1 1 43540
0 43542 7 1 2 43445 43541
0 43543 5 1 1 43542
0 43544 7 1 2 71149 43543
0 43545 5 1 1 43544
0 43546 7 1 2 80544 78033
0 43547 5 1 1 43546
0 43548 7 1 2 105212 43547
0 43549 5 1 1 43548
0 43550 7 1 2 66060 43549
0 43551 5 1 1 43550
0 43552 7 3 2 81915 83649
0 43553 5 1 1 105219
0 43554 7 1 2 97283 105220
0 43555 5 1 1 43554
0 43556 7 1 2 43551 43555
0 43557 5 1 1 43556
0 43558 7 1 2 71464 43557
0 43559 5 1 1 43558
0 43560 7 1 2 78437 102979
0 43561 5 1 1 43560
0 43562 7 1 2 43559 43561
0 43563 5 1 1 43562
0 43564 7 1 2 68143 43563
0 43565 5 1 1 43564
0 43566 7 1 2 94940 89440
0 43567 5 1 1 43566
0 43568 7 1 2 43567 43253
0 43569 5 1 1 43568
0 43570 7 1 2 69944 43569
0 43571 5 1 1 43570
0 43572 7 2 2 76422 88645
0 43573 5 1 1 105222
0 43574 7 1 2 70505 90766
0 43575 5 1 1 43574
0 43576 7 1 2 43573 43575
0 43577 7 1 2 43571 43576
0 43578 5 1 1 43577
0 43579 7 1 2 91745 43578
0 43580 5 1 1 43579
0 43581 7 1 2 76423 87821
0 43582 5 1 1 43581
0 43583 7 1 2 67742 79999
0 43584 5 1 1 43583
0 43585 7 1 2 43582 43584
0 43586 5 1 1 43585
0 43587 7 1 2 69945 43586
0 43588 5 1 1 43587
0 43589 7 1 2 85068 43588
0 43590 7 1 2 43580 43589
0 43591 5 1 1 43590
0 43592 7 1 2 66775 43591
0 43593 5 1 1 43592
0 43594 7 1 2 43565 43593
0 43595 5 1 1 43594
0 43596 7 1 2 69587 43595
0 43597 5 1 1 43596
0 43598 7 1 2 90774 16131
0 43599 5 1 1 43598
0 43600 7 1 2 79034 43599
0 43601 5 1 1 43600
0 43602 7 1 2 88680 104018
0 43603 5 1 1 43602
0 43604 7 1 2 43601 43603
0 43605 5 1 1 43604
0 43606 7 1 2 68480 43605
0 43607 5 1 1 43606
0 43608 7 1 2 70506 83983
0 43609 5 1 1 43608
0 43610 7 1 2 86896 84009
0 43611 7 1 2 43609 43610
0 43612 5 1 1 43611
0 43613 7 1 2 43607 43612
0 43614 5 1 1 43613
0 43615 7 1 2 69588 43614
0 43616 5 1 1 43615
0 43617 7 3 2 69946 87128
0 43618 7 1 2 84712 84296
0 43619 7 1 2 105224 43618
0 43620 5 1 1 43619
0 43621 7 1 2 43616 43620
0 43622 5 1 1 43621
0 43623 7 1 2 75435 43622
0 43624 5 1 1 43623
0 43625 7 1 2 99874 83399
0 43626 5 1 1 43625
0 43627 7 1 2 43533 43626
0 43628 5 1 1 43627
0 43629 7 1 2 70507 43628
0 43630 5 1 1 43629
0 43631 7 1 2 86682 81240
0 43632 5 1 1 43631
0 43633 7 1 2 76424 95875
0 43634 5 1 1 43633
0 43635 7 1 2 43632 43634
0 43636 7 1 2 43630 43635
0 43637 5 1 1 43636
0 43638 7 1 2 103699 43637
0 43639 5 1 1 43638
0 43640 7 1 2 72459 43639
0 43641 7 1 2 43624 43640
0 43642 7 1 2 43597 43641
0 43643 7 1 2 43545 43642
0 43644 5 1 1 43643
0 43645 7 2 2 43443 43644
0 43646 7 1 2 78884 105227
0 43647 5 1 1 43646
0 43648 7 2 2 64844 101945
0 43649 5 1 1 105229
0 43650 7 1 2 43649 42390
0 43651 5 3 1 43650
0 43652 7 3 2 65180 80373
0 43653 5 3 1 105234
0 43654 7 1 2 97605 105237
0 43655 5 1 1 43654
0 43656 7 1 2 105231 43655
0 43657 5 1 1 43656
0 43658 7 1 2 93816 99624
0 43659 5 1 1 43658
0 43660 7 1 2 95407 105062
0 43661 7 1 2 43659 43660
0 43662 5 1 1 43661
0 43663 7 1 2 43657 43662
0 43664 5 1 1 43663
0 43665 7 1 2 66061 43664
0 43666 5 1 1 43665
0 43667 7 2 2 93803 103564
0 43668 7 1 2 105122 105240
0 43669 5 1 1 43668
0 43670 7 1 2 43666 43669
0 43671 5 1 1 43670
0 43672 7 1 2 68481 43671
0 43673 5 1 1 43672
0 43674 7 1 2 77977 101678
0 43675 7 1 2 105232 43674
0 43676 5 1 1 43675
0 43677 7 1 2 69589 43676
0 43678 7 1 2 43673 43677
0 43679 5 1 1 43678
0 43680 7 1 2 90703 92670
0 43681 5 1 1 43680
0 43682 7 1 2 37663 43681
0 43683 5 1 1 43682
0 43684 7 1 2 70243 43683
0 43685 5 1 1 43684
0 43686 7 1 2 96558 105238
0 43687 5 1 1 43686
0 43688 7 1 2 82139 43687
0 43689 5 1 1 43688
0 43690 7 1 2 43685 43689
0 43691 5 1 1 43690
0 43692 7 1 2 68482 43691
0 43693 5 1 1 43692
0 43694 7 2 2 64845 74907
0 43695 7 1 2 71691 96033
0 43696 7 1 2 105242 43695
0 43697 5 1 1 43696
0 43698 7 1 2 43693 43697
0 43699 5 1 1 43698
0 43700 7 1 2 105009 43699
0 43701 5 1 1 43700
0 43702 7 1 2 88708 87834
0 43703 5 1 1 43702
0 43704 7 1 2 71692 93275
0 43705 5 1 1 43704
0 43706 7 1 2 43703 43705
0 43707 5 1 1 43706
0 43708 7 1 2 65487 43707
0 43709 5 1 1 43708
0 43710 7 1 2 86221 77716
0 43711 5 1 1 43710
0 43712 7 1 2 102362 43711
0 43713 5 1 1 43712
0 43714 7 1 2 83534 43713
0 43715 5 1 1 43714
0 43716 7 1 2 43709 43715
0 43717 5 1 1 43716
0 43718 7 1 2 80836 97054
0 43719 7 1 2 43717 43718
0 43720 5 1 1 43719
0 43721 7 1 2 64474 43720
0 43722 7 1 2 43701 43721
0 43723 5 1 1 43722
0 43724 7 1 2 79150 43723
0 43725 7 1 2 43679 43724
0 43726 5 1 1 43725
0 43727 7 1 2 43647 43726
0 43728 5 1 1 43727
0 43729 7 1 2 82456 43728
0 43730 5 1 1 43729
0 43731 7 1 2 96962 74560
0 43732 7 1 2 74070 43731
0 43733 7 1 2 80152 43732
0 43734 5 1 1 43733
0 43735 7 1 2 75936 91433
0 43736 5 1 1 43735
0 43737 7 1 2 68144 103168
0 43738 5 1 1 43737
0 43739 7 1 2 43736 43738
0 43740 5 1 1 43739
0 43741 7 1 2 66062 99754
0 43742 7 1 2 43740 43741
0 43743 5 1 1 43742
0 43744 7 1 2 43734 43743
0 43745 5 1 1 43744
0 43746 7 1 2 69590 43745
0 43747 5 1 1 43746
0 43748 7 1 2 64846 105010
0 43749 5 1 1 43748
0 43750 7 1 2 80837 102041
0 43751 5 1 1 43750
0 43752 7 1 2 43749 43751
0 43753 5 1 1 43752
0 43754 7 1 2 77993 92824
0 43755 7 1 2 43753 43754
0 43756 5 1 1 43755
0 43757 7 1 2 43747 43756
0 43758 5 1 1 43757
0 43759 7 1 2 104079 43758
0 43760 5 1 1 43759
0 43761 7 5 2 67387 80211
0 43762 5 1 1 105244
0 43763 7 2 2 93057 105245
0 43764 7 1 2 80183 105249
0 43765 5 1 1 43764
0 43766 7 3 2 96919 84341
0 43767 7 1 2 75985 86705
0 43768 5 1 1 43767
0 43769 7 1 2 68145 89816
0 43770 5 1 1 43769
0 43771 7 1 2 43768 43770
0 43772 5 1 1 43771
0 43773 7 1 2 105251 43772
0 43774 5 1 1 43773
0 43775 7 1 2 43765 43774
0 43776 5 2 1 43775
0 43777 7 1 2 71150 105254
0 43778 5 1 1 43777
0 43779 7 1 2 92774 91048
0 43780 5 1 1 43779
0 43781 7 1 2 66363 105214
0 43782 5 1 1 43781
0 43783 7 1 2 43780 43782
0 43784 5 1 1 43783
0 43785 7 1 2 105252 43784
0 43786 5 1 1 43785
0 43787 7 1 2 43778 43786
0 43788 5 1 1 43787
0 43789 7 1 2 78885 43788
0 43790 5 1 1 43789
0 43791 7 1 2 43760 43790
0 43792 5 1 1 43791
0 43793 7 1 2 68483 43792
0 43794 5 1 1 43793
0 43795 7 1 2 72460 99568
0 43796 7 1 2 99970 43795
0 43797 7 1 2 87551 43796
0 43798 5 1 1 43797
0 43799 7 1 2 74071 105246
0 43800 7 1 2 99875 43799
0 43801 5 1 1 43800
0 43802 7 1 2 43798 43801
0 43803 5 1 1 43802
0 43804 7 1 2 69947 43803
0 43805 5 1 1 43804
0 43806 7 1 2 99320 105193
0 43807 7 1 2 105247 43806
0 43808 5 1 1 43807
0 43809 7 1 2 43805 43808
0 43810 5 1 1 43809
0 43811 7 1 2 97293 43810
0 43812 5 1 1 43811
0 43813 7 1 2 43794 43812
0 43814 5 1 1 43813
0 43815 7 1 2 67743 43814
0 43816 5 1 1 43815
0 43817 7 3 2 69948 93758
0 43818 5 1 1 105256
0 43819 7 2 2 79596 77909
0 43820 7 1 2 105005 105259
0 43821 5 1 1 43820
0 43822 7 1 2 103812 94345
0 43823 7 1 2 105011 43822
0 43824 5 1 1 43823
0 43825 7 1 2 43821 43824
0 43826 5 1 1 43825
0 43827 7 1 2 105257 43826
0 43828 5 1 1 43827
0 43829 7 1 2 74561 105260
0 43830 5 1 1 43829
0 43831 7 2 2 70508 86507
0 43832 7 2 2 71957 105261
0 43833 7 1 2 95873 105263
0 43834 5 1 1 43833
0 43835 7 1 2 43830 43834
0 43836 5 1 1 43835
0 43837 7 1 2 74799 99249
0 43838 7 1 2 43836 43837
0 43839 5 1 1 43838
0 43840 7 1 2 43828 43839
0 43841 5 1 1 43840
0 43842 7 1 2 101056 43841
0 43843 5 1 1 43842
0 43844 7 1 2 43816 43843
0 43845 5 1 1 43844
0 43846 7 1 2 82992 43845
0 43847 5 1 1 43846
0 43848 7 1 2 90046 80822
0 43849 5 1 1 43848
0 43850 7 1 2 80153 80454
0 43851 5 1 1 43850
0 43852 7 1 2 43849 43851
0 43853 5 2 1 43852
0 43854 7 1 2 78886 105265
0 43855 5 1 1 43854
0 43856 7 1 2 76826 75592
0 43857 7 1 2 86843 86100
0 43858 7 1 2 43856 43857
0 43859 5 1 1 43858
0 43860 7 1 2 43855 43859
0 43861 5 1 1 43860
0 43862 7 6 2 67744 97911
0 43863 7 2 2 101006 105267
0 43864 7 1 2 43861 105273
0 43865 5 1 1 43864
0 43866 7 1 2 43847 43865
0 43867 7 1 2 43730 43866
0 43868 7 1 2 43388 43867
0 43869 5 1 1 43868
0 43870 7 1 2 68999 43869
0 43871 5 1 1 43870
0 43872 7 2 2 93264 98964
0 43873 7 2 2 89633 93070
0 43874 7 1 2 65606 105277
0 43875 7 1 2 105275 43874
0 43876 5 1 1 43875
0 43877 7 2 2 71151 103546
0 43878 7 1 2 90952 102954
0 43879 7 1 2 105279 43878
0 43880 5 1 1 43879
0 43881 7 1 2 43876 43880
0 43882 5 1 1 43881
0 43883 7 1 2 68882 43882
0 43884 5 1 1 43883
0 43885 7 1 2 84611 99244
0 43886 7 1 2 105276 43885
0 43887 5 1 1 43886
0 43888 7 1 2 43884 43887
0 43889 5 1 1 43888
0 43890 7 1 2 64192 43889
0 43891 5 1 1 43890
0 43892 7 1 2 70863 105012
0 43893 5 1 1 43892
0 43894 7 1 2 98943 103473
0 43895 5 1 1 43894
0 43896 7 1 2 43893 43895
0 43897 5 2 1 43896
0 43898 7 2 2 68883 93733
0 43899 7 1 2 87868 91705
0 43900 7 1 2 105283 43899
0 43901 7 1 2 105281 43900
0 43902 5 1 1 43901
0 43903 7 1 2 43891 43902
0 43904 5 1 1 43903
0 43905 7 1 2 64475 43904
0 43906 5 1 1 43905
0 43907 7 2 2 99298 85025
0 43908 7 1 2 104136 105285
0 43909 5 1 1 43908
0 43910 7 2 2 84297 99266
0 43911 7 1 2 101957 105287
0 43912 5 1 1 43911
0 43913 7 1 2 66063 102344
0 43914 5 1 1 43913
0 43915 7 1 2 71152 104255
0 43916 5 1 1 43915
0 43917 7 1 2 69949 43916
0 43918 7 1 2 43914 43917
0 43919 5 1 1 43918
0 43920 7 1 2 43912 43919
0 43921 5 1 1 43920
0 43922 7 1 2 69245 43921
0 43923 5 1 1 43922
0 43924 7 1 2 43909 43923
0 43925 5 1 1 43924
0 43926 7 1 2 79151 89124
0 43927 7 1 2 43925 43926
0 43928 5 1 1 43927
0 43929 7 1 2 43906 43928
0 43930 5 1 1 43929
0 43931 7 1 2 81764 43930
0 43932 5 1 1 43931
0 43933 7 1 2 89270 101951
0 43934 5 2 1 43933
0 43935 7 2 2 67388 82457
0 43936 7 1 2 101863 79390
0 43937 7 1 2 105291 43936
0 43938 7 1 2 105289 43937
0 43939 5 1 1 43938
0 43940 7 1 2 43932 43939
0 43941 5 1 1 43940
0 43942 7 1 2 65181 43941
0 43943 5 1 1 43942
0 43944 7 1 2 97803 104917
0 43945 5 2 1 43944
0 43946 7 1 2 103864 90945
0 43947 5 1 1 43946
0 43948 7 1 2 105293 43947
0 43949 5 1 1 43948
0 43950 7 2 2 70864 97330
0 43951 7 1 2 66883 79381
0 43952 7 1 2 105295 43951
0 43953 7 1 2 43949 43952
0 43954 5 1 1 43953
0 43955 7 1 2 43943 43954
0 43956 5 1 1 43955
0 43957 7 1 2 73979 43956
0 43958 5 1 1 43957
0 43959 7 1 2 43871 43958
0 43960 5 1 1 43959
0 43961 7 1 2 73858 43960
0 43962 5 1 1 43961
0 43963 7 1 2 82458 105228
0 43964 5 1 1 43963
0 43965 7 1 2 85541 105197
0 43966 5 1 1 43965
0 43967 7 1 2 105266 105274
0 43968 5 1 1 43967
0 43969 7 1 2 68484 105255
0 43970 5 1 1 43969
0 43971 7 1 2 99881 105250
0 43972 5 1 1 43971
0 43973 7 1 2 43970 43972
0 43974 5 1 1 43973
0 43975 7 1 2 71153 43974
0 43976 5 1 1 43975
0 43977 7 1 2 81312 80000
0 43978 5 1 1 43977
0 43979 7 1 2 81335 43978
0 43980 5 1 1 43979
0 43981 7 1 2 105258 43980
0 43982 5 1 1 43981
0 43983 7 1 2 69591 81165
0 43984 5 1 1 43983
0 43985 7 1 2 43982 43984
0 43986 5 1 1 43985
0 43987 7 1 2 105253 43986
0 43988 5 1 1 43987
0 43989 7 1 2 43976 43988
0 43990 5 1 1 43989
0 43991 7 1 2 67745 43990
0 43992 5 1 1 43991
0 43993 7 2 2 73231 102905
0 43994 5 1 1 105297
0 43995 7 1 2 99569 77072
0 43996 7 1 2 101908 43995
0 43997 7 1 2 105298 43996
0 43998 5 1 1 43997
0 43999 7 1 2 43992 43998
0 44000 5 1 1 43999
0 44001 7 1 2 82993 44000
0 44002 5 1 1 44001
0 44003 7 1 2 43968 44002
0 44004 7 1 2 43966 44003
0 44005 7 1 2 43964 44004
0 44006 5 1 1 44005
0 44007 7 1 2 90347 44006
0 44008 5 1 1 44007
0 44009 7 1 2 105013 43347
0 44010 5 1 1 44009
0 44011 7 1 2 69950 80127
0 44012 7 1 2 105288 44011
0 44013 5 1 1 44012
0 44014 7 1 2 44010 44013
0 44015 5 1 1 44014
0 44016 7 1 2 64476 44015
0 44017 5 1 1 44016
0 44018 7 1 2 65182 105233
0 44019 5 1 1 44018
0 44020 7 1 2 100605 105063
0 44021 5 1 1 44020
0 44022 7 1 2 44019 44021
0 44023 5 1 1 44022
0 44024 7 1 2 80996 44023
0 44025 5 1 1 44024
0 44026 7 1 2 44017 44025
0 44027 5 1 1 44026
0 44028 7 1 2 82459 44027
0 44029 5 1 1 44028
0 44030 7 1 2 78129 99087
0 44031 7 1 2 104941 44030
0 44032 5 1 1 44031
0 44033 7 1 2 44029 44032
0 44034 5 1 1 44033
0 44035 7 1 2 86066 44034
0 44036 5 1 1 44035
0 44037 7 1 2 72461 105129
0 44038 5 1 1 44037
0 44039 7 1 2 44038 42694
0 44040 5 1 1 44039
0 44041 7 1 2 67746 44040
0 44042 5 1 1 44041
0 44043 7 1 2 87890 99250
0 44044 5 1 1 44043
0 44045 7 1 2 44042 44044
0 44046 5 2 1 44045
0 44047 7 1 2 97602 105299
0 44048 5 1 1 44047
0 44049 7 1 2 105241 105126
0 44050 5 1 1 44049
0 44051 7 1 2 44048 44050
0 44052 5 1 1 44051
0 44053 7 1 2 82460 44052
0 44054 5 1 1 44053
0 44055 7 1 2 44036 44054
0 44056 5 1 1 44055
0 44057 7 1 2 68485 44056
0 44058 5 1 1 44057
0 44059 7 3 2 69246 84342
0 44060 7 1 2 101679 105301
0 44061 7 1 2 105300 44060
0 44062 5 1 1 44061
0 44063 7 1 2 85542 105210
0 44064 5 1 1 44063
0 44065 7 1 2 44062 44064
0 44066 7 1 2 44058 44065
0 44067 5 1 1 44066
0 44068 7 1 2 105144 44067
0 44069 5 1 1 44068
0 44070 7 1 2 44008 44069
0 44071 5 1 1 44070
0 44072 7 1 2 63912 44071
0 44073 5 1 1 44072
0 44074 7 1 2 93804 105290
0 44075 5 1 1 44074
0 44076 7 1 2 99104 81536
0 44077 5 1 1 44076
0 44078 7 1 2 44075 44077
0 44079 5 1 1 44078
0 44080 7 1 2 67389 44079
0 44081 5 1 1 44080
0 44082 7 1 2 105294 44081
0 44083 5 1 1 44082
0 44084 7 1 2 93113 44083
0 44085 5 1 1 44084
0 44086 7 4 2 64193 84464
0 44087 7 2 2 75519 105304
0 44088 7 1 2 95316 98117
0 44089 7 1 2 93425 44088
0 44090 7 1 2 105308 44089
0 44091 5 1 1 44090
0 44092 7 1 2 44085 44091
0 44093 5 1 1 44092
0 44094 7 1 2 90348 44093
0 44095 5 1 1 44094
0 44096 7 2 2 74973 74072
0 44097 5 1 1 105310
0 44098 7 1 2 103978 44097
0 44099 5 3 1 44098
0 44100 7 1 2 69247 105312
0 44101 5 1 1 44100
0 44102 7 1 2 85460 105194
0 44103 5 1 1 44102
0 44104 7 1 2 44101 44103
0 44105 5 1 1 44104
0 44106 7 1 2 105205 44105
0 44107 5 1 1 44106
0 44108 7 3 2 82461 97055
0 44109 7 2 2 68146 81093
0 44110 5 1 1 105318
0 44111 7 1 2 105315 105319
0 44112 5 1 1 44111
0 44113 7 1 2 44107 44112
0 44114 5 1 1 44113
0 44115 7 1 2 69951 44114
0 44116 5 1 1 44115
0 44117 7 1 2 95639 74337
0 44118 7 1 2 102044 44117
0 44119 5 1 1 44118
0 44120 7 1 2 44116 44119
0 44121 5 1 1 44120
0 44122 7 1 2 94466 98873
0 44123 7 1 2 44121 44122
0 44124 5 1 1 44123
0 44125 7 1 2 44095 44124
0 44126 5 1 1 44125
0 44127 7 1 2 73980 44126
0 44128 5 1 1 44127
0 44129 7 1 2 67129 44128
0 44130 7 1 2 44073 44129
0 44131 7 1 2 43962 44130
0 44132 7 1 2 43052 44131
0 44133 5 1 1 44132
0 44134 7 2 2 78183 96385
0 44135 5 1 1 105320
0 44136 7 2 2 73859 77035
0 44137 5 1 1 105322
0 44138 7 1 2 68884 105323
0 44139 5 1 1 44138
0 44140 7 2 2 44135 44139
0 44141 5 4 1 105324
0 44142 7 1 2 88381 101208
0 44143 5 1 1 44142
0 44144 7 2 2 80733 82875
0 44145 5 1 1 105330
0 44146 7 1 2 68486 44145
0 44147 7 1 2 44143 44146
0 44148 5 1 1 44147
0 44149 7 1 2 66589 96650
0 44150 5 1 1 44149
0 44151 7 1 2 73559 101503
0 44152 7 1 2 44150 44151
0 44153 5 1 1 44152
0 44154 7 1 2 44148 44153
0 44155 5 1 1 44154
0 44156 7 1 2 69952 44155
0 44157 5 1 1 44156
0 44158 7 1 2 104171 44157
0 44159 5 1 1 44158
0 44160 7 1 2 72747 44159
0 44161 5 1 1 44160
0 44162 7 1 2 69592 92007
0 44163 5 1 1 44162
0 44164 7 1 2 85702 44163
0 44165 5 1 1 44164
0 44166 7 3 2 81765 74691
0 44167 7 1 2 81176 105332
0 44168 5 1 1 44167
0 44169 7 1 2 67747 44168
0 44170 7 1 2 44165 44169
0 44171 5 1 1 44170
0 44172 7 1 2 44161 44171
0 44173 5 1 1 44172
0 44174 7 1 2 64477 83330
0 44175 7 1 2 87364 44174
0 44176 5 1 1 44175
0 44177 7 1 2 44173 44176
0 44178 5 1 1 44177
0 44179 7 1 2 105326 44178
0 44180 5 1 1 44179
0 44181 7 1 2 64847 104304
0 44182 5 1 1 44181
0 44183 7 1 2 86256 86652
0 44184 5 1 1 44183
0 44185 7 1 2 44182 44184
0 44186 5 1 1 44185
0 44187 7 1 2 67748 44186
0 44188 5 1 1 44187
0 44189 7 1 2 104014 104166
0 44190 5 1 1 44189
0 44191 7 1 2 44188 44190
0 44192 5 1 1 44191
0 44193 7 1 2 70509 44192
0 44194 5 1 1 44193
0 44195 7 1 2 83006 92633
0 44196 7 1 2 100024 44195
0 44197 5 1 1 44196
0 44198 7 1 2 44194 44197
0 44199 5 1 1 44198
0 44200 7 1 2 88078 44199
0 44201 5 1 1 44200
0 44202 7 1 2 85703 101854
0 44203 5 1 1 44202
0 44204 7 2 2 67749 85704
0 44205 5 1 1 105335
0 44206 7 1 2 87650 92671
0 44207 5 1 1 44206
0 44208 7 1 2 44205 44207
0 44209 7 1 2 44203 44208
0 44210 5 1 1 44209
0 44211 7 1 2 88986 44210
0 44212 5 1 1 44211
0 44213 7 1 2 44201 44212
0 44214 5 1 1 44213
0 44215 7 1 2 64478 44214
0 44216 5 1 1 44215
0 44217 7 3 2 87651 90935
0 44218 5 1 1 105337
0 44219 7 1 2 67750 89046
0 44220 5 1 1 44219
0 44221 7 1 2 44218 44220
0 44222 5 2 1 44221
0 44223 7 1 2 64848 105340
0 44224 5 1 1 44223
0 44225 7 1 2 73560 88773
0 44226 5 1 1 44225
0 44227 7 1 2 71693 100795
0 44228 7 1 2 44226 44227
0 44229 5 1 1 44228
0 44230 7 1 2 100845 44229
0 44231 5 1 1 44230
0 44232 7 1 2 92672 44231
0 44233 5 1 1 44232
0 44234 7 1 2 44224 44233
0 44235 5 1 1 44234
0 44236 7 1 2 88987 44235
0 44237 5 1 1 44236
0 44238 7 1 2 44216 44237
0 44239 5 1 1 44238
0 44240 7 1 2 87410 44239
0 44241 5 1 1 44240
0 44242 7 1 2 44180 44241
0 44243 5 1 1 44242
0 44244 7 1 2 71465 44243
0 44245 5 1 1 44244
0 44246 7 3 2 66884 98080
0 44247 7 3 2 71694 96443
0 44248 5 1 1 105345
0 44249 7 1 2 101504 44248
0 44250 5 2 1 44249
0 44251 7 2 2 98564 105348
0 44252 5 1 1 105350
0 44253 7 1 2 64849 87657
0 44254 5 2 1 44253
0 44255 7 1 2 28401 81537
0 44256 7 1 2 105352 44255
0 44257 5 1 1 44256
0 44258 7 1 2 44252 44257
0 44259 5 1 1 44258
0 44260 7 1 2 105342 44259
0 44261 5 1 1 44260
0 44262 7 1 2 44245 44261
0 44263 5 1 1 44262
0 44264 7 1 2 68147 44263
0 44265 5 1 1 44264
0 44266 7 1 2 76336 105351
0 44267 5 1 1 44266
0 44268 7 1 2 105081 105336
0 44269 5 1 1 44268
0 44270 7 1 2 44267 44269
0 44271 5 1 1 44270
0 44272 7 1 2 98081 44271
0 44273 5 1 1 44272
0 44274 7 1 2 76661 81480
0 44275 5 1 1 44274
0 44276 7 1 2 69593 78960
0 44277 5 2 1 44276
0 44278 7 1 2 92995 105354
0 44279 5 1 1 44278
0 44280 7 1 2 44275 44279
0 44281 5 1 1 44280
0 44282 7 1 2 86067 44281
0 44283 5 1 1 44282
0 44284 7 1 2 69953 104119
0 44285 5 1 1 44284
0 44286 7 1 2 44283 44285
0 44287 5 1 1 44286
0 44288 7 1 2 68487 44287
0 44289 5 1 1 44288
0 44290 7 1 2 81557 80908
0 44291 5 1 1 44290
0 44292 7 1 2 82140 85797
0 44293 5 1 1 44292
0 44294 7 1 2 44291 44293
0 44295 5 1 1 44294
0 44296 7 1 2 69594 44295
0 44297 5 1 1 44296
0 44298 7 1 2 44289 44297
0 44299 5 1 1 44298
0 44300 7 1 2 94084 79391
0 44301 5 1 1 44300
0 44302 7 1 2 98078 44301
0 44303 5 3 1 44302
0 44304 7 1 2 73232 105356
0 44305 7 1 2 44299 44304
0 44306 5 1 1 44305
0 44307 7 1 2 44273 44306
0 44308 5 1 1 44307
0 44309 7 1 2 66885 44308
0 44310 5 1 1 44309
0 44311 7 1 2 44265 44310
0 44312 5 1 1 44311
0 44313 7 1 2 71154 44312
0 44314 5 1 1 44313
0 44315 7 1 2 81995 74974
0 44316 5 2 1 44315
0 44317 7 1 2 66064 81241
0 44318 5 1 1 44317
0 44319 7 1 2 105359 44318
0 44320 5 2 1 44319
0 44321 7 1 2 68488 105361
0 44322 5 1 1 44321
0 44323 7 1 2 90220 80975
0 44324 5 1 1 44323
0 44325 7 1 2 44322 44324
0 44326 5 1 1 44325
0 44327 7 1 2 69954 44326
0 44328 5 1 1 44327
0 44329 7 1 2 87056 92088
0 44330 5 2 1 44329
0 44331 7 2 2 69595 105363
0 44332 5 1 1 105365
0 44333 7 1 2 82174 105366
0 44334 5 1 1 44333
0 44335 7 1 2 44328 44334
0 44336 5 1 1 44335
0 44337 7 1 2 67751 44336
0 44338 5 1 1 44337
0 44339 7 1 2 74975 1510
0 44340 7 1 2 81481 44339
0 44341 7 1 2 91746 44340
0 44342 5 1 1 44341
0 44343 7 1 2 44338 44342
0 44344 5 1 1 44343
0 44345 7 1 2 86068 44344
0 44346 5 1 1 44345
0 44347 7 1 2 83440 105043
0 44348 5 2 1 44347
0 44349 7 1 2 83400 92191
0 44350 5 1 1 44349
0 44351 7 1 2 105367 44350
0 44352 5 1 1 44351
0 44353 7 1 2 75436 44352
0 44354 5 1 1 44353
0 44355 7 1 2 99919 93470
0 44356 5 3 1 44355
0 44357 7 1 2 66065 105369
0 44358 5 1 1 44357
0 44359 7 1 2 82081 82202
0 44360 5 1 1 44359
0 44361 7 1 2 44358 44360
0 44362 5 1 1 44361
0 44363 7 1 2 66776 44362
0 44364 5 1 1 44363
0 44365 7 1 2 44354 44364
0 44366 5 1 1 44365
0 44367 7 1 2 65488 44366
0 44368 5 1 1 44367
0 44369 7 1 2 97340 81558
0 44370 5 1 1 44369
0 44371 7 1 2 71695 82671
0 44372 5 1 1 44371
0 44373 7 1 2 44370 44372
0 44374 5 1 1 44373
0 44375 7 1 2 81442 44374
0 44376 5 1 1 44375
0 44377 7 1 2 78450 44376
0 44378 5 1 1 44377
0 44379 7 1 2 71466 44378
0 44380 5 1 1 44379
0 44381 7 1 2 93203 44380
0 44382 5 1 1 44381
0 44383 7 1 2 73561 44382
0 44384 5 1 1 44383
0 44385 7 1 2 44368 44384
0 44386 5 1 1 44385
0 44387 7 1 2 76962 44386
0 44388 5 1 1 44387
0 44389 7 1 2 44346 44388
0 44390 5 1 1 44389
0 44391 7 2 2 66886 105357
0 44392 7 1 2 44390 105372
0 44393 5 1 1 44392
0 44394 7 1 2 44314 44393
0 44395 5 1 1 44394
0 44396 7 1 2 67390 44395
0 44397 5 1 1 44396
0 44398 7 1 2 77544 80943
0 44399 5 1 1 44398
0 44400 7 1 2 104213 44399
0 44401 5 1 1 44400
0 44402 7 1 2 105343 44401
0 44403 5 1 1 44402
0 44404 7 1 2 75582 90704
0 44405 7 2 2 90953 92316
0 44406 7 1 2 94674 91681
0 44407 7 1 2 105374 44406
0 44408 7 1 2 44404 44407
0 44409 5 1 1 44408
0 44410 7 1 2 44403 44409
0 44411 5 1 1 44410
0 44412 7 1 2 103669 44411
0 44413 5 1 1 44412
0 44414 7 1 2 44397 44413
0 44415 5 1 1 44414
0 44416 7 1 2 70865 44415
0 44417 5 1 1 44416
0 44418 7 3 2 69000 89583
0 44419 5 1 1 105376
0 44420 7 1 2 63808 105377
0 44421 5 1 1 44420
0 44422 7 1 2 63913 99322
0 44423 5 2 1 44422
0 44424 7 1 2 7108 105379
0 44425 7 1 2 44421 44424
0 44426 5 1 1 44425
0 44427 7 1 2 78487 104545
0 44428 7 1 2 44426 44427
0 44429 7 1 2 104215 44428
0 44430 5 1 1 44429
0 44431 7 1 2 77832 84465
0 44432 7 1 2 99323 44431
0 44433 5 1 1 44432
0 44434 7 1 2 84577 89634
0 44435 7 1 2 94339 44434
0 44436 5 1 1 44435
0 44437 7 1 2 91154 78334
0 44438 7 1 2 89584 44437
0 44439 5 1 1 44438
0 44440 7 1 2 44436 44439
0 44441 7 1 2 44433 44440
0 44442 5 1 1 44441
0 44443 7 2 2 85613 98360
0 44444 7 1 2 66066 77049
0 44445 7 1 2 105381 44444
0 44446 7 1 2 44442 44445
0 44447 5 1 1 44446
0 44448 7 1 2 44430 44447
0 44449 5 1 1 44448
0 44450 7 1 2 84228 44449
0 44451 5 1 1 44450
0 44452 7 1 2 44417 44451
0 44453 5 1 1 44452
0 44454 7 1 2 64194 44453
0 44455 5 1 1 44454
0 44456 7 1 2 87411 88988
0 44457 5 1 1 44456
0 44458 7 1 2 105325 44457
0 44459 5 1 1 44458
0 44460 7 1 2 100025 44459
0 44461 5 1 1 44460
0 44462 7 1 2 94548 73924
0 44463 7 1 2 87412 44462
0 44464 7 1 2 91415 44463
0 44465 5 1 1 44464
0 44466 7 1 2 44461 44465
0 44467 5 1 1 44466
0 44468 7 1 2 72748 44467
0 44469 5 1 1 44468
0 44470 7 1 2 87413 94347
0 44471 7 2 2 94138 96511
0 44472 7 1 2 84095 105383
0 44473 7 1 2 44470 44472
0 44474 5 1 1 44473
0 44475 7 1 2 44469 44474
0 44476 5 1 1 44475
0 44477 7 1 2 71856 44476
0 44478 5 1 1 44477
0 44479 7 1 2 83653 24653
0 44480 5 3 1 44479
0 44481 7 1 2 105076 105385
0 44482 7 1 2 98082 44481
0 44483 5 1 1 44482
0 44484 7 1 2 44478 44483
0 44485 5 1 1 44484
0 44486 7 1 2 70510 44485
0 44487 5 1 1 44486
0 44488 7 2 2 87105 104312
0 44489 7 1 2 83999 105388
0 44490 7 1 2 98083 44489
0 44491 5 1 1 44490
0 44492 7 1 2 44487 44491
0 44493 5 1 1 44492
0 44494 7 1 2 67391 44493
0 44495 5 1 1 44494
0 44496 7 1 2 96727 99276
0 44497 7 1 2 104083 44496
0 44498 7 1 2 92835 96351
0 44499 7 1 2 44497 44498
0 44500 5 1 1 44499
0 44501 7 1 2 44495 44500
0 44502 5 1 1 44501
0 44503 7 1 2 69248 44502
0 44504 5 1 1 44503
0 44505 7 1 2 70511 104546
0 44506 7 1 2 101878 44505
0 44507 7 2 2 80468 91172
0 44508 7 3 2 87414 92449
0 44509 7 1 2 98954 105392
0 44510 7 1 2 105390 44509
0 44511 7 1 2 44506 44510
0 44512 5 1 1 44511
0 44513 7 1 2 44504 44512
0 44514 5 1 1 44513
0 44515 7 1 2 70244 44514
0 44516 5 1 1 44515
0 44517 7 1 2 85705 105321
0 44518 5 1 1 44517
0 44519 7 1 2 8045 44137
0 44520 5 1 1 44519
0 44521 7 1 2 85706 44520
0 44522 5 1 1 44521
0 44523 7 2 2 100026 94603
0 44524 7 1 2 69001 87183
0 44525 7 1 2 105395 44524
0 44526 5 1 1 44525
0 44527 7 1 2 44522 44526
0 44528 5 1 1 44527
0 44529 7 1 2 68885 44528
0 44530 5 1 1 44529
0 44531 7 1 2 44518 44530
0 44532 5 1 1 44531
0 44533 7 1 2 74199 98765
0 44534 7 1 2 44532 44533
0 44535 5 1 1 44534
0 44536 7 1 2 44516 44535
0 44537 5 1 1 44536
0 44538 7 1 2 105313 44537
0 44539 5 1 1 44538
0 44540 7 1 2 101235 93016
0 44541 5 1 1 44540
0 44542 7 1 2 82392 93153
0 44543 5 1 1 44542
0 44544 7 1 2 44541 44543
0 44545 5 1 1 44544
0 44546 7 1 2 70866 44545
0 44547 5 1 1 44546
0 44548 7 1 2 2038 105059
0 44549 5 1 1 44548
0 44550 7 1 2 78053 44549
0 44551 5 1 1 44550
0 44552 7 1 2 44547 44551
0 44553 5 1 1 44552
0 44554 7 1 2 72462 44553
0 44555 5 1 1 44554
0 44556 7 1 2 78423 82090
0 44557 5 1 1 44556
0 44558 7 1 2 87552 44557
0 44559 5 1 1 44558
0 44560 7 1 2 66590 18238
0 44561 5 1 1 44560
0 44562 7 1 2 81990 81647
0 44563 7 1 2 44561 44562
0 44564 5 1 1 44563
0 44565 7 1 2 44559 44564
0 44566 5 1 1 44565
0 44567 7 1 2 97912 44566
0 44568 5 1 1 44567
0 44569 7 1 2 44555 44568
0 44570 5 1 1 44569
0 44571 7 1 2 69596 44570
0 44572 5 1 1 44571
0 44573 7 1 2 66067 104207
0 44574 5 1 1 44573
0 44575 7 1 2 98239 93154
0 44576 5 1 1 44575
0 44577 7 1 2 44574 44576
0 44578 5 1 1 44577
0 44579 7 1 2 70867 44578
0 44580 5 1 1 44579
0 44581 7 1 2 98180 105311
0 44582 5 1 1 44581
0 44583 7 1 2 44580 44582
0 44584 5 1 1 44583
0 44585 7 1 2 83635 44584
0 44586 5 1 1 44585
0 44587 7 1 2 82158 98157
0 44588 7 1 2 95517 44587
0 44589 5 1 1 44588
0 44590 7 1 2 44586 44589
0 44591 7 1 2 44572 44590
0 44592 5 1 1 44591
0 44593 7 1 2 71857 44592
0 44594 5 1 1 44593
0 44595 7 1 2 66068 93155
0 44596 5 1 1 44595
0 44597 7 1 2 6092 44596
0 44598 5 1 1 44597
0 44599 7 1 2 68489 44598
0 44600 5 1 1 44599
0 44601 7 1 2 66777 105120
0 44602 5 1 1 44601
0 44603 7 1 2 90775 44602
0 44604 5 1 1 44603
0 44605 7 1 2 81509 44604
0 44606 5 1 1 44605
0 44607 7 1 2 44600 44606
0 44608 5 1 1 44607
0 44609 7 1 2 69597 44608
0 44610 5 1 1 44609
0 44611 7 2 2 79250 84298
0 44612 5 1 1 105397
0 44613 7 1 2 91810 105398
0 44614 5 1 1 44613
0 44615 7 1 2 64479 93156
0 44616 5 1 1 44615
0 44617 7 1 2 65183 92192
0 44618 5 1 1 44617
0 44619 7 1 2 44616 44618
0 44620 5 1 1 44619
0 44621 7 1 2 68490 44620
0 44622 5 1 1 44621
0 44623 7 2 2 74743 81968
0 44624 5 1 1 105399
0 44625 7 1 2 87337 105400
0 44626 5 1 1 44625
0 44627 7 1 2 44622 44626
0 44628 5 1 1 44627
0 44629 7 1 2 71155 44628
0 44630 5 1 1 44629
0 44631 7 1 2 44614 44630
0 44632 7 1 2 44610 44631
0 44633 5 1 1 44632
0 44634 7 1 2 67392 44633
0 44635 5 1 1 44634
0 44636 7 1 2 102158 103670
0 44637 5 1 1 44636
0 44638 7 1 2 44635 44637
0 44639 5 1 1 44638
0 44640 7 1 2 65842 44639
0 44641 5 1 1 44640
0 44642 7 1 2 72749 80560
0 44643 5 1 1 44642
0 44644 7 1 2 13950 44643
0 44645 5 1 1 44644
0 44646 7 1 2 70245 44645
0 44647 5 1 1 44646
0 44648 7 1 2 71696 99141
0 44649 5 1 1 44648
0 44650 7 1 2 44647 44649
0 44651 5 1 1 44650
0 44652 7 1 2 82609 44651
0 44653 5 1 1 44652
0 44654 7 1 2 77184 103624
0 44655 5 1 1 44654
0 44656 7 1 2 44653 44655
0 44657 5 1 1 44656
0 44658 7 1 2 98442 44657
0 44659 5 1 1 44658
0 44660 7 1 2 44641 44659
0 44661 5 1 1 44660
0 44662 7 1 2 68700 44661
0 44663 5 1 1 44662
0 44664 7 1 2 44594 44663
0 44665 5 1 1 44664
0 44666 7 1 2 70512 44665
0 44667 5 1 1 44666
0 44668 7 1 2 82552 105182
0 44669 5 1 1 44668
0 44670 7 1 2 70868 87901
0 44671 5 1 1 44670
0 44672 7 1 2 44669 44671
0 44673 5 1 1 44672
0 44674 7 1 2 66069 44673
0 44675 5 1 1 44674
0 44676 7 1 2 71156 93157
0 44677 5 2 1 44676
0 44678 7 1 2 66591 91470
0 44679 5 1 1 44678
0 44680 7 1 2 105401 44679
0 44681 5 1 1 44680
0 44682 7 1 2 80374 44681
0 44683 5 1 1 44682
0 44684 7 1 2 71697 86897
0 44685 7 1 2 76945 44684
0 44686 5 1 1 44685
0 44687 7 1 2 44683 44686
0 44688 5 1 1 44687
0 44689 7 1 2 65843 44688
0 44690 5 1 1 44689
0 44691 7 1 2 44675 44690
0 44692 5 1 1 44691
0 44693 7 1 2 68491 44692
0 44694 5 1 1 44693
0 44695 7 2 2 85707 93468
0 44696 7 1 2 74073 105403
0 44697 5 1 1 44696
0 44698 7 1 2 44694 44697
0 44699 5 1 1 44698
0 44700 7 1 2 67393 44699
0 44701 5 1 1 44700
0 44702 7 1 2 85069 105402
0 44703 5 2 1 44702
0 44704 7 1 2 98443 73925
0 44705 7 1 2 105405 44704
0 44706 5 1 1 44705
0 44707 7 1 2 44701 44706
0 44708 5 1 1 44707
0 44709 7 1 2 64480 44708
0 44710 5 1 1 44709
0 44711 7 1 2 98481 95714
0 44712 5 1 1 44711
0 44713 7 2 2 72750 98509
0 44714 7 1 2 82358 79737
0 44715 5 1 1 44714
0 44716 7 1 2 80734 80797
0 44717 5 1 1 44716
0 44718 7 1 2 44715 44717
0 44719 5 1 1 44718
0 44720 7 1 2 105407 44719
0 44721 5 1 1 44720
0 44722 7 1 2 71157 44721
0 44723 7 1 2 44712 44722
0 44724 5 1 1 44723
0 44725 7 1 2 80204 97204
0 44726 5 1 1 44725
0 44727 7 1 2 38838 44726
0 44728 5 1 1 44727
0 44729 7 1 2 93158 44728
0 44730 5 1 1 44729
0 44731 7 2 2 65489 93221
0 44732 7 1 2 87338 99078
0 44733 7 1 2 105409 44732
0 44734 5 1 1 44733
0 44735 7 1 2 44730 44734
0 44736 5 1 1 44735
0 44737 7 1 2 68492 44736
0 44738 5 1 1 44737
0 44739 7 1 2 97913 105404
0 44740 5 1 1 44739
0 44741 7 1 2 66070 44740
0 44742 7 1 2 44738 44741
0 44743 5 1 1 44742
0 44744 7 1 2 44724 44743
0 44745 5 1 1 44744
0 44746 7 1 2 74809 104699
0 44747 5 1 1 44746
0 44748 7 1 2 105408 44747
0 44749 5 1 1 44748
0 44750 7 1 2 80531 103264
0 44751 5 1 1 44750
0 44752 7 1 2 44749 44751
0 44753 5 1 1 44752
0 44754 7 1 2 71158 44753
0 44755 5 1 1 44754
0 44756 7 1 2 82203 103815
0 44757 7 1 2 103102 44756
0 44758 5 1 1 44757
0 44759 7 1 2 44755 44758
0 44760 5 1 1 44759
0 44761 7 1 2 75437 44760
0 44762 5 1 1 44761
0 44763 7 1 2 66778 95405
0 44764 5 1 1 44763
0 44765 7 1 2 105368 44764
0 44766 5 1 1 44765
0 44767 7 1 2 97914 83113
0 44768 7 1 2 44766 44767
0 44769 5 1 1 44768
0 44770 7 1 2 44762 44769
0 44771 7 1 2 44745 44770
0 44772 5 1 1 44771
0 44773 7 1 2 69598 44772
0 44774 5 1 1 44773
0 44775 7 1 2 98444 93017
0 44776 5 1 1 44775
0 44777 7 1 2 104256 44776
0 44778 5 1 1 44777
0 44779 7 1 2 84113 100777
0 44780 5 1 1 44779
0 44781 7 1 2 97653 96456
0 44782 5 1 1 44781
0 44783 7 1 2 44780 44782
0 44784 5 1 1 44783
0 44785 7 1 2 44778 44784
0 44786 5 1 1 44785
0 44787 7 1 2 83535 92412
0 44788 7 1 2 101078 44787
0 44789 5 1 1 44788
0 44790 7 1 2 102461 30622
0 44791 5 1 1 44790
0 44792 7 1 2 81648 96531
0 44793 7 1 2 44791 44792
0 44794 5 1 1 44793
0 44795 7 1 2 44789 44794
0 44796 5 1 1 44795
0 44797 7 1 2 68701 97557
0 44798 7 1 2 44796 44797
0 44799 5 1 1 44798
0 44800 7 1 2 44786 44799
0 44801 7 1 2 44774 44800
0 44802 7 1 2 44710 44801
0 44803 7 1 2 44667 44802
0 44804 5 1 1 44803
0 44805 7 1 2 69955 44804
0 44806 5 1 1 44805
0 44807 7 2 2 68148 78383
0 44808 5 1 1 105411
0 44809 7 1 2 44332 44808
0 44810 5 1 1 44809
0 44811 7 1 2 87652 44810
0 44812 5 1 1 44811
0 44813 7 1 2 87704 74976
0 44814 5 1 1 44813
0 44815 7 1 2 78973 44814
0 44816 5 2 1 44815
0 44817 7 1 2 81766 105413
0 44818 5 1 1 44817
0 44819 7 1 2 75084 92649
0 44820 5 1 1 44819
0 44821 7 1 2 22716 44820
0 44822 7 1 2 44818 44821
0 44823 5 1 1 44822
0 44824 7 1 2 71159 44823
0 44825 5 1 1 44824
0 44826 7 1 2 44812 44825
0 44827 5 1 1 44826
0 44828 7 1 2 65844 44827
0 44829 5 1 1 44828
0 44830 7 1 2 73981 89970
0 44831 5 1 1 44830
0 44832 7 1 2 82309 75986
0 44833 5 1 1 44832
0 44834 7 1 2 99902 44833
0 44835 5 1 1 44834
0 44836 7 1 2 44831 44835
0 44837 5 1 1 44836
0 44838 7 1 2 98711 44837
0 44839 5 1 1 44838
0 44840 7 1 2 44829 44839
0 44841 5 1 1 44840
0 44842 7 1 2 64850 44841
0 44843 5 1 1 44842
0 44844 7 1 2 75020 89047
0 44845 5 1 1 44844
0 44846 7 1 2 66364 84243
0 44847 5 1 1 44846
0 44848 7 1 2 44845 44847
0 44849 5 1 1 44848
0 44850 7 1 2 98712 44849
0 44851 5 1 1 44850
0 44852 7 1 2 67752 44851
0 44853 7 1 2 44843 44852
0 44854 5 1 1 44853
0 44855 7 1 2 77807 105221
0 44856 5 1 1 44855
0 44857 7 1 2 71160 104060
0 44858 5 1 1 44857
0 44859 7 1 2 44856 44858
0 44860 5 1 1 44859
0 44861 7 1 2 75476 44860
0 44862 5 1 1 44861
0 44863 7 1 2 101260 44862
0 44864 5 1 1 44863
0 44865 7 1 2 93058 44864
0 44866 5 1 1 44865
0 44867 7 1 2 75092 101733
0 44868 5 1 1 44867
0 44869 7 1 2 93406 44868
0 44870 5 1 1 44869
0 44871 7 1 2 44866 44870
0 44872 5 1 1 44871
0 44873 7 1 2 68149 44872
0 44874 5 1 1 44873
0 44875 7 1 2 101506 98524
0 44876 5 1 1 44875
0 44877 7 2 2 66592 74338
0 44878 7 1 2 92430 105415
0 44879 5 1 1 44878
0 44880 7 1 2 44876 44879
0 44881 5 1 1 44880
0 44882 7 1 2 73562 44881
0 44883 5 1 1 44882
0 44884 7 1 2 93241 97649
0 44885 7 1 2 87653 44884
0 44886 5 1 1 44885
0 44887 7 1 2 72751 44886
0 44888 7 1 2 44883 44887
0 44889 7 1 2 44874 44888
0 44890 5 1 1 44889
0 44891 7 1 2 67394 44890
0 44892 7 1 2 44854 44891
0 44893 5 1 1 44892
0 44894 7 2 2 72752 84854
0 44895 5 1 1 105417
0 44896 7 1 2 81662 105418
0 44897 5 1 1 44896
0 44898 7 1 2 103559 44897
0 44899 5 1 1 44898
0 44900 7 1 2 73563 44899
0 44901 5 1 1 44900
0 44902 7 1 2 73233 105338
0 44903 5 1 1 44902
0 44904 7 1 2 44901 44903
0 44905 5 1 1 44904
0 44906 7 1 2 71161 44905
0 44907 5 1 1 44906
0 44908 7 2 2 100793 86069
0 44909 7 1 2 93018 105419
0 44910 5 1 1 44909
0 44911 7 1 2 44907 44910
0 44912 5 1 1 44911
0 44913 7 1 2 70869 44912
0 44914 5 1 1 44913
0 44915 7 1 2 77808 74074
0 44916 7 1 2 95387 44915
0 44917 7 1 2 95359 44916
0 44918 5 1 1 44917
0 44919 7 1 2 44914 44918
0 44920 5 1 1 44919
0 44921 7 1 2 69599 44920
0 44922 5 1 1 44921
0 44923 7 1 2 64851 95518
0 44924 7 1 2 104180 44923
0 44925 5 1 1 44924
0 44926 7 1 2 44922 44925
0 44927 5 1 1 44926
0 44928 7 1 2 72463 44927
0 44929 5 1 1 44928
0 44930 7 1 2 100313 99207
0 44931 5 1 1 44930
0 44932 7 1 2 65184 102525
0 44933 5 1 1 44932
0 44934 7 1 2 44931 44933
0 44935 5 1 1 44934
0 44936 7 1 2 64852 44935
0 44937 5 1 1 44936
0 44938 7 2 2 73564 89441
0 44939 7 1 2 71698 98474
0 44940 7 1 2 105421 44939
0 44941 5 1 1 44940
0 44942 7 1 2 44937 44941
0 44943 5 1 1 44942
0 44944 7 1 2 70870 44943
0 44945 5 1 1 44944
0 44946 7 1 2 83191 105054
0 44947 7 1 2 105422 44946
0 44948 5 1 1 44947
0 44949 7 1 2 44945 44948
0 44950 5 1 1 44949
0 44951 7 1 2 71162 44950
0 44952 5 1 1 44951
0 44953 7 1 2 100314 80029
0 44954 5 1 1 44953
0 44955 7 1 2 65185 79260
0 44956 5 1 1 44955
0 44957 7 1 2 44954 44956
0 44958 5 1 1 44957
0 44959 7 1 2 96760 77073
0 44960 7 1 2 44958 44959
0 44961 5 1 1 44960
0 44962 7 1 2 44952 44961
0 44963 5 1 1 44962
0 44964 7 1 2 80735 44963
0 44965 5 1 1 44964
0 44966 7 1 2 44929 44965
0 44967 7 1 2 44893 44966
0 44968 7 1 2 44806 44967
0 44969 5 1 1 44968
0 44970 7 1 2 105373 44969
0 44971 5 1 1 44970
0 44972 7 3 2 67753 93059
0 44973 7 1 2 98240 94632
0 44974 5 1 1 44973
0 44975 7 2 2 67395 90373
0 44976 7 1 2 79738 87929
0 44977 7 1 2 94149 44976
0 44978 7 1 2 105426 44977
0 44979 5 1 1 44978
0 44980 7 1 2 44974 44979
0 44981 5 1 1 44980
0 44982 7 1 2 105423 44981
0 44983 5 1 1 44982
0 44984 7 1 2 98241 91199
0 44985 7 1 2 85044 44984
0 44986 7 1 2 91410 93479
0 44987 7 1 2 44985 44986
0 44988 5 1 1 44987
0 44989 7 1 2 44983 44988
0 44990 5 1 1 44989
0 44991 7 1 2 74562 44990
0 44992 5 1 1 44991
0 44993 7 1 2 65186 84389
0 44994 5 1 1 44993
0 44995 7 1 2 105360 44994
0 44996 5 1 1 44995
0 44997 7 1 2 105268 44996
0 44998 5 1 1 44997
0 44999 7 2 2 81056 93159
0 45000 5 1 1 105428
0 45001 7 1 2 98510 105429
0 45002 5 1 1 45001
0 45003 7 1 2 97886 104208
0 45004 5 1 1 45003
0 45005 7 1 2 95376 98965
0 45006 5 1 1 45005
0 45007 7 1 2 45004 45006
0 45008 7 1 2 45002 45007
0 45009 7 1 2 44998 45008
0 45010 5 1 1 45009
0 45011 7 1 2 88989 45010
0 45012 5 1 1 45011
0 45013 7 1 2 44992 45012
0 45014 5 1 1 45013
0 45015 7 1 2 87415 45014
0 45016 5 1 1 45015
0 45017 7 1 2 99876 98615
0 45018 5 1 1 45017
0 45019 7 1 2 97129 105355
0 45020 5 1 1 45019
0 45021 7 1 2 45018 45020
0 45022 5 1 1 45021
0 45023 7 1 2 71163 45022
0 45024 5 1 1 45023
0 45025 7 1 2 67396 105362
0 45026 5 1 1 45025
0 45027 7 1 2 45024 45026
0 45028 5 1 1 45027
0 45029 7 1 2 67754 45028
0 45030 5 1 1 45029
0 45031 7 1 2 82573 44110
0 45032 5 1 1 45031
0 45033 7 1 2 96761 45032
0 45034 5 1 1 45033
0 45035 7 1 2 65845 45034
0 45036 7 1 2 45030 45035
0 45037 5 1 1 45036
0 45038 7 1 2 10425 45000
0 45039 5 1 1 45038
0 45040 7 1 2 72464 45039
0 45041 5 1 1 45040
0 45042 7 1 2 77381 104209
0 45043 5 1 1 45042
0 45044 7 1 2 70871 45043
0 45045 7 1 2 45041 45044
0 45046 5 1 1 45045
0 45047 7 1 2 105327 45046
0 45048 7 1 2 45037 45047
0 45049 5 1 1 45048
0 45050 7 1 2 45016 45049
0 45051 5 1 1 45050
0 45052 7 1 2 69956 95780
0 45053 7 1 2 45051 45052
0 45054 5 1 1 45053
0 45055 7 1 2 44971 45054
0 45056 5 1 1 45055
0 45057 7 1 2 69249 45056
0 45058 5 1 1 45057
0 45059 7 1 2 81482 105282
0 45060 5 1 1 45059
0 45061 7 2 2 95340 97056
0 45062 7 1 2 79261 105430
0 45063 5 1 1 45062
0 45064 7 1 2 45060 45063
0 45065 5 1 1 45064
0 45066 7 1 2 69250 45065
0 45067 5 1 1 45066
0 45068 7 1 2 100493 105286
0 45069 5 1 1 45068
0 45070 7 1 2 45067 45069
0 45071 5 1 1 45070
0 45072 7 1 2 79901 94274
0 45073 5 2 1 45072
0 45074 7 1 2 105328 105432
0 45075 5 1 1 45074
0 45076 7 1 2 84745 105396
0 45077 5 1 1 45076
0 45078 7 1 2 73982 88990
0 45079 5 1 1 45078
0 45080 7 1 2 45077 45079
0 45081 5 1 1 45080
0 45082 7 1 2 65490 45081
0 45083 5 1 1 45082
0 45084 7 1 2 69957 87143
0 45085 5 1 1 45084
0 45086 7 1 2 88991 45085
0 45087 5 1 1 45086
0 45088 7 2 2 80298 88043
0 45089 7 1 2 102940 94336
0 45090 7 1 2 105434 45089
0 45091 5 1 1 45090
0 45092 7 1 2 45087 45091
0 45093 7 1 2 45083 45092
0 45094 5 1 1 45093
0 45095 7 1 2 87416 45094
0 45096 5 1 1 45095
0 45097 7 1 2 45075 45096
0 45098 5 1 1 45097
0 45099 7 1 2 45071 45098
0 45100 5 1 1 45099
0 45101 7 1 2 72174 45100
0 45102 7 1 2 45058 45101
0 45103 7 1 2 44539 45102
0 45104 7 1 2 44455 45103
0 45105 5 1 1 45104
0 45106 7 1 2 44133 45105
0 45107 5 1 1 45106
0 45108 7 1 2 67755 91687
0 45109 5 2 1 45108
0 45110 7 1 2 80469 93635
0 45111 7 1 2 88079 45110
0 45112 5 1 1 45111
0 45113 7 1 2 105436 45112
0 45114 5 1 1 45113
0 45115 7 1 2 69958 45114
0 45116 5 1 1 45115
0 45117 7 2 2 87345 102942
0 45118 5 1 1 105438
0 45119 7 1 2 84585 94372
0 45120 7 1 2 45118 45119
0 45121 5 1 1 45120
0 45122 7 1 2 45116 45121
0 45123 5 1 1 45122
0 45124 7 1 2 68886 45123
0 45125 5 1 1 45124
0 45126 7 1 2 70513 105439
0 45127 5 1 1 45126
0 45128 7 1 2 67756 16036
0 45129 7 1 2 105138 45128
0 45130 7 1 2 45127 45129
0 45131 5 1 1 45130
0 45132 7 1 2 45125 45131
0 45133 5 1 1 45132
0 45134 7 1 2 70246 45133
0 45135 5 1 1 45134
0 45136 7 1 2 91832 102980
0 45137 7 1 2 105168 45136
0 45138 5 1 1 45137
0 45139 7 1 2 45135 45138
0 45140 5 1 1 45139
0 45141 7 1 2 68493 45140
0 45142 5 1 1 45141
0 45143 7 1 2 79694 91660
0 45144 7 2 2 84681 45143
0 45145 7 2 2 94671 90374
0 45146 7 1 2 105440 105442
0 45147 5 1 1 45146
0 45148 7 1 2 45147 105437
0 45149 5 1 1 45148
0 45150 7 1 2 70247 45149
0 45151 5 1 1 45150
0 45152 7 1 2 65689 78706
0 45153 7 1 2 84586 45152
0 45154 7 1 2 91724 45153
0 45155 5 1 1 45154
0 45156 7 1 2 45151 45155
0 45157 5 1 1 45156
0 45158 7 1 2 68887 45157
0 45159 5 1 1 45158
0 45160 7 1 2 67757 101777
0 45161 7 1 2 105139 45160
0 45162 5 1 1 45161
0 45163 7 1 2 45159 45162
0 45164 5 1 1 45163
0 45165 7 1 2 69959 45164
0 45166 5 1 1 45165
0 45167 7 1 2 84587 92205
0 45168 7 1 2 92517 45167
0 45169 5 1 1 45168
0 45170 7 1 2 45166 45169
0 45171 5 1 1 45170
0 45172 7 1 2 82994 45171
0 45173 5 1 1 45172
0 45174 7 1 2 1320 83523
0 45175 5 1 1 45174
0 45176 7 1 2 84588 45175
0 45177 7 1 2 90338 45176
0 45178 5 1 1 45177
0 45179 7 1 2 45173 45178
0 45180 7 1 2 45142 45179
0 45181 5 1 1 45180
0 45182 7 1 2 88229 45181
0 45183 5 1 1 45182
0 45184 7 1 2 88992 105386
0 45185 5 1 1 45184
0 45186 7 1 2 73926 79284
0 45187 5 2 1 45186
0 45188 7 1 2 69600 92989
0 45189 5 2 1 45188
0 45190 7 1 2 105444 105446
0 45191 5 3 1 45190
0 45192 7 2 2 70727 71858
0 45193 7 1 2 91938 105451
0 45194 7 1 2 105448 45193
0 45195 5 1 1 45194
0 45196 7 1 2 45185 45195
0 45197 5 1 1 45196
0 45198 7 1 2 68888 45197
0 45199 5 1 1 45198
0 45200 7 1 2 105140 105387
0 45201 5 1 1 45200
0 45202 7 1 2 45199 45201
0 45203 5 1 1 45202
0 45204 7 1 2 70514 45203
0 45205 5 1 1 45204
0 45206 7 1 2 90339 105389
0 45207 5 1 1 45206
0 45208 7 1 2 45205 45207
0 45209 5 1 1 45208
0 45210 7 1 2 80856 45209
0 45211 5 1 1 45210
0 45212 7 1 2 104306 90349
0 45213 5 1 1 45212
0 45214 7 1 2 45211 45213
0 45215 5 1 1 45214
0 45216 7 1 2 67758 45215
0 45217 5 1 1 45216
0 45218 7 1 2 98830 100931
0 45219 7 1 2 104691 95656
0 45220 7 1 2 105391 45219
0 45221 7 1 2 45218 45220
0 45222 5 1 1 45221
0 45223 7 1 2 45217 45222
0 45224 5 1 1 45223
0 45225 7 1 2 88582 45224
0 45226 5 1 1 45225
0 45227 7 1 2 84855 79209
0 45228 5 1 1 45227
0 45229 7 1 2 43553 45228
0 45230 5 2 1 45229
0 45231 7 1 2 80857 105453
0 45232 5 1 1 45231
0 45233 7 1 2 104308 45232
0 45234 5 1 1 45233
0 45235 7 1 2 81342 45234
0 45236 5 1 1 45235
0 45237 7 1 2 69960 86751
0 45238 5 1 1 45237
0 45239 7 1 2 104089 45238
0 45240 5 1 1 45239
0 45241 7 1 2 75438 45240
0 45242 5 1 1 45241
0 45243 7 1 2 80299 103195
0 45244 5 1 1 45243
0 45245 7 1 2 76662 87630
0 45246 5 1 1 45245
0 45247 7 1 2 64481 45246
0 45248 5 1 1 45247
0 45249 7 1 2 65491 45248
0 45250 5 1 1 45249
0 45251 7 1 2 45244 45250
0 45252 7 1 2 45242 45251
0 45253 5 1 1 45252
0 45254 7 1 2 80190 45253
0 45255 5 1 1 45254
0 45256 7 1 2 45236 45255
0 45257 5 1 1 45256
0 45258 7 1 2 66887 45257
0 45259 5 1 1 45258
0 45260 7 2 2 81139 87654
0 45261 7 1 2 94976 97251
0 45262 7 1 2 105455 45261
0 45263 5 1 1 45262
0 45264 7 1 2 45259 45263
0 45265 5 1 1 45264
0 45266 7 1 2 67759 45265
0 45267 5 1 1 45266
0 45268 7 2 2 89172 97245
0 45269 7 1 2 90721 89125
0 45270 7 1 2 95552 45269
0 45271 7 1 2 105457 45270
0 45272 5 1 1 45271
0 45273 7 1 2 45267 45272
0 45274 5 1 1 45273
0 45275 7 1 2 73860 45274
0 45276 5 1 1 45275
0 45277 7 1 2 45226 45276
0 45278 7 1 2 45183 45277
0 45279 5 1 1 45278
0 45280 7 1 2 99388 45279
0 45281 5 1 1 45280
0 45282 7 2 2 72753 77994
0 45283 5 1 1 105459
0 45284 7 3 2 88583 90350
0 45285 5 2 1 105461
0 45286 7 3 2 91451 88030
0 45287 7 1 2 66779 87749
0 45288 7 2 2 92130 89518
0 45289 7 1 2 45287 105469
0 45290 7 1 2 105466 45289
0 45291 5 1 1 45290
0 45292 7 1 2 105464 45291
0 45293 5 1 1 45292
0 45294 7 1 2 105460 45293
0 45295 5 1 1 45294
0 45296 7 1 2 92634 104526
0 45297 7 1 2 91695 45296
0 45298 7 2 2 76963 86404
0 45299 7 1 2 94413 105471
0 45300 7 1 2 45297 45299
0 45301 5 1 1 45300
0 45302 7 1 2 45295 45301
0 45303 5 1 1 45302
0 45304 7 1 2 67397 45303
0 45305 5 1 1 45304
0 45306 7 2 2 97057 96300
0 45307 7 1 2 89126 105473
0 45308 7 1 2 90351 45307
0 45309 5 1 1 45308
0 45310 7 1 2 45305 45309
0 45311 5 1 1 45310
0 45312 7 1 2 65492 45311
0 45313 5 1 1 45312
0 45314 7 2 2 75679 99208
0 45315 5 1 1 105475
0 45316 7 2 2 96762 96131
0 45317 7 1 2 64482 103365
0 45318 7 1 2 105477 45317
0 45319 5 1 1 45318
0 45320 7 1 2 45315 45319
0 45321 5 1 1 45320
0 45322 7 1 2 70872 45321
0 45323 5 1 1 45322
0 45324 7 1 2 70642 103757
0 45325 7 2 2 98882 45324
0 45326 7 1 2 91452 89127
0 45327 7 1 2 105479 45326
0 45328 5 1 1 45327
0 45329 7 1 2 45323 45328
0 45330 5 1 1 45329
0 45331 7 1 2 65493 45330
0 45332 5 1 1 45331
0 45333 7 1 2 94865 105476
0 45334 5 1 1 45333
0 45335 7 1 2 45332 45334
0 45336 5 1 1 45335
0 45337 7 1 2 68889 45336
0 45338 5 1 1 45337
0 45339 7 1 2 80736 96549
0 45340 7 1 2 95673 45339
0 45341 7 1 2 99209 45340
0 45342 5 1 1 45341
0 45343 7 1 2 45338 45342
0 45344 5 1 1 45343
0 45345 7 1 2 73861 45344
0 45346 5 1 1 45345
0 45347 7 1 2 94866 99210
0 45348 7 1 2 105462 45347
0 45349 5 1 1 45348
0 45350 7 1 2 45346 45349
0 45351 7 1 2 45313 45350
0 45352 5 1 1 45351
0 45353 7 1 2 69251 45352
0 45354 5 1 1 45353
0 45355 7 5 2 67130 73862
0 45356 7 1 2 100232 86405
0 45357 7 1 2 105481 45356
0 45358 5 1 1 45357
0 45359 7 1 2 92131 93846
0 45360 7 1 2 91173 45359
0 45361 7 1 2 92457 45360
0 45362 5 1 1 45361
0 45363 7 1 2 45358 45362
0 45364 5 1 1 45363
0 45365 7 2 2 79035 88001
0 45366 7 1 2 96550 98766
0 45367 7 1 2 105486 45366
0 45368 7 1 2 45364 45367
0 45369 5 1 1 45368
0 45370 7 1 2 45354 45369
0 45371 5 1 1 45370
0 45372 7 1 2 73983 45371
0 45373 5 1 1 45372
0 45374 7 1 2 35024 97549
0 45375 5 3 1 45374
0 45376 7 1 2 74563 105488
0 45377 5 1 1 45376
0 45378 7 1 2 69961 98933
0 45379 5 1 1 45378
0 45380 7 1 2 75439 100755
0 45381 5 1 1 45380
0 45382 7 1 2 103714 45381
0 45383 7 1 2 45379 45382
0 45384 7 1 2 45377 45383
0 45385 5 2 1 45384
0 45386 7 1 2 80191 105491
0 45387 5 1 1 45386
0 45388 7 2 2 81767 78707
0 45389 5 1 1 105493
0 45390 7 2 2 93909 45389
0 45391 5 1 1 105495
0 45392 7 1 2 69962 105496
0 45393 5 1 1 45392
0 45394 7 1 2 70248 77955
0 45395 7 1 2 105353 45394
0 45396 7 1 2 45393 45395
0 45397 5 1 1 45396
0 45398 7 2 2 68494 99497
0 45399 5 1 1 105497
0 45400 7 1 2 89856 45399
0 45401 7 1 2 45397 45400
0 45402 5 2 1 45401
0 45403 7 1 2 81343 105499
0 45404 5 1 1 45403
0 45405 7 1 2 45387 45404
0 45406 5 1 1 45405
0 45407 7 1 2 102052 45406
0 45408 5 1 1 45407
0 45409 7 1 2 64483 79912
0 45410 7 2 2 101057 45409
0 45411 7 1 2 81344 105501
0 45412 5 1 1 45411
0 45413 7 1 2 45408 45412
0 45414 5 1 1 45413
0 45415 7 1 2 66888 45414
0 45416 5 1 1 45415
0 45417 7 1 2 100911 87428
0 45418 7 1 2 96221 45417
0 45419 7 1 2 105132 45418
0 45420 5 1 1 45419
0 45421 7 1 2 45416 45420
0 45422 5 1 1 45421
0 45423 7 1 2 73863 45422
0 45424 5 1 1 45423
0 45425 7 1 2 79644 101864
0 45426 5 1 1 45425
0 45427 7 1 2 70249 45391
0 45428 5 1 1 45427
0 45429 7 1 2 64853 101637
0 45430 7 1 2 45428 45429
0 45431 5 1 1 45430
0 45432 7 1 2 79794 43818
0 45433 7 1 2 45431 45432
0 45434 5 1 1 45433
0 45435 7 1 2 45426 45434
0 45436 5 1 1 45435
0 45437 7 1 2 96328 45436
0 45438 5 1 1 45437
0 45439 7 2 2 80737 90289
0 45440 7 1 2 74040 92286
0 45441 7 1 2 105503 45440
0 45442 5 1 1 45441
0 45443 7 1 2 45438 45442
0 45444 5 1 1 45443
0 45445 7 1 2 67131 45444
0 45446 5 1 1 45445
0 45447 7 1 2 69067 94399
0 45448 7 1 2 100802 94598
0 45449 7 1 2 89809 45448
0 45450 7 1 2 45447 45449
0 45451 5 1 1 45450
0 45452 7 1 2 45446 45451
0 45453 5 1 1 45452
0 45454 7 2 2 72754 82504
0 45455 5 1 1 105505
0 45456 7 1 2 74430 16639
0 45457 7 2 2 45455 45456
0 45458 7 1 2 84653 105507
0 45459 7 1 2 45453 45458
0 45460 5 1 1 45459
0 45461 7 1 2 88584 105500
0 45462 5 1 1 45461
0 45463 7 1 2 88230 105492
0 45464 5 1 1 45463
0 45465 7 1 2 45462 45464
0 45466 5 1 1 45465
0 45467 7 1 2 102053 45466
0 45468 5 1 1 45467
0 45469 7 1 2 88585 105502
0 45470 5 1 1 45469
0 45471 7 1 2 45468 45470
0 45472 5 1 1 45471
0 45473 7 1 2 90352 45472
0 45474 5 1 1 45473
0 45475 7 2 2 88031 92317
0 45476 7 1 2 85543 81140
0 45477 7 1 2 105509 45476
0 45478 7 1 2 105441 45477
0 45479 7 1 2 98539 45478
0 45480 5 1 1 45479
0 45481 7 1 2 45474 45480
0 45482 7 1 2 45460 45481
0 45483 7 1 2 45424 45482
0 45484 5 1 1 45483
0 45485 7 1 2 67398 45484
0 45486 5 1 1 45485
0 45487 7 1 2 70728 97915
0 45488 7 1 2 89930 86406
0 45489 7 1 2 94235 90525
0 45490 7 1 2 45488 45489
0 45491 7 1 2 45487 45490
0 45492 5 1 1 45491
0 45493 7 1 2 87106 102459
0 45494 7 1 2 90340 45493
0 45495 5 1 1 45494
0 45496 7 1 2 45492 45495
0 45497 5 1 1 45496
0 45498 7 1 2 70515 45497
0 45499 5 1 1 45498
0 45500 7 1 2 82995 89090
0 45501 7 1 2 94242 45500
0 45502 7 1 2 94997 45501
0 45503 7 1 2 102295 45502
0 45504 5 1 1 45503
0 45505 7 1 2 45499 45504
0 45506 5 1 1 45505
0 45507 7 1 2 69252 45506
0 45508 5 1 1 45507
0 45509 7 2 2 69601 87184
0 45510 5 1 1 105511
0 45511 7 1 2 70873 102412
0 45512 7 1 2 93549 45511
0 45513 7 1 2 105512 45512
0 45514 5 1 1 45513
0 45515 7 1 2 45508 45514
0 45516 5 1 1 45515
0 45517 7 1 2 88586 45516
0 45518 5 1 1 45517
0 45519 7 2 2 69602 99409
0 45520 7 1 2 94085 94826
0 45521 7 1 2 96132 45520
0 45522 7 1 2 105513 45521
0 45523 5 1 1 45522
0 45524 7 1 2 45518 45523
0 45525 5 1 1 45524
0 45526 7 1 2 67760 45525
0 45527 5 1 1 45526
0 45528 7 1 2 83625 76890
0 45529 7 1 2 105478 45528
0 45530 5 1 1 45529
0 45531 7 2 2 99190 84635
0 45532 7 1 2 75807 86612
0 45533 7 1 2 105515 45532
0 45534 5 1 1 45533
0 45535 7 1 2 45530 45534
0 45536 5 1 1 45535
0 45537 7 1 2 68890 45536
0 45538 5 1 1 45537
0 45539 7 1 2 80300 97143
0 45540 7 1 2 105516 45539
0 45541 5 1 1 45540
0 45542 7 1 2 45538 45541
0 45543 5 1 1 45542
0 45544 7 1 2 70874 45543
0 45545 5 1 1 45544
0 45546 7 1 2 89091 76005
0 45547 7 1 2 105480 45546
0 45548 5 1 1 45547
0 45549 7 1 2 45545 45548
0 45550 5 1 1 45549
0 45551 7 1 2 69253 45550
0 45552 5 1 1 45551
0 45553 7 1 2 93598 103758
0 45554 7 3 2 69603 76891
0 45555 7 2 2 84324 86407
0 45556 7 1 2 105517 105520
0 45557 7 1 2 45553 45556
0 45558 5 1 1 45557
0 45559 7 1 2 45552 45558
0 45560 5 1 1 45559
0 45561 7 1 2 73864 45560
0 45562 5 1 1 45561
0 45563 7 1 2 99450 97180
0 45564 7 2 2 83295 86408
0 45565 7 1 2 99124 105522
0 45566 7 1 2 45563 45565
0 45567 7 1 2 94537 45566
0 45568 5 1 1 45567
0 45569 7 1 2 45562 45568
0 45570 7 1 2 45527 45569
0 45571 5 1 1 45570
0 45572 7 1 2 100027 45571
0 45573 5 1 1 45572
0 45574 7 1 2 45486 45573
0 45575 7 1 2 45373 45574
0 45576 7 1 2 45281 45575
0 45577 5 1 1 45576
0 45578 7 1 2 84398 45577
0 45579 5 1 1 45578
0 45580 7 1 2 91985 105449
0 45581 5 1 1 45580
0 45582 7 2 2 86613 89547
0 45583 7 4 2 63979 64854
0 45584 7 1 2 92373 105526
0 45585 7 1 2 105524 45584
0 45586 5 1 1 45585
0 45587 7 1 2 45581 45586
0 45588 5 1 1 45587
0 45589 7 1 2 65187 45588
0 45590 5 1 1 45589
0 45591 7 3 2 70516 88993
0 45592 7 1 2 101816 105530
0 45593 5 1 1 45592
0 45594 7 1 2 45590 45593
0 45595 5 1 1 45594
0 45596 7 1 2 71164 45595
0 45597 5 1 1 45596
0 45598 7 2 2 94150 91670
0 45599 7 1 2 93536 94998
0 45600 7 1 2 105533 45599
0 45601 5 1 1 45600
0 45602 7 1 2 86614 105527
0 45603 7 1 2 81510 45602
0 45604 7 1 2 92287 45603
0 45605 5 1 1 45604
0 45606 7 1 2 45601 45605
0 45607 5 1 1 45606
0 45608 7 1 2 69604 45607
0 45609 5 1 1 45608
0 45610 7 1 2 45597 45609
0 45611 5 1 1 45610
0 45612 7 1 2 87417 45611
0 45613 5 1 1 45612
0 45614 7 1 2 64855 97664
0 45615 5 1 1 45614
0 45616 7 1 2 64484 76624
0 45617 5 1 1 45616
0 45618 7 1 2 45615 45617
0 45619 5 1 1 45618
0 45620 7 1 2 70517 45619
0 45621 7 1 2 105329 45620
0 45622 5 1 1 45621
0 45623 7 1 2 45613 45622
0 45624 5 1 1 45623
0 45625 7 1 2 72175 45624
0 45626 5 1 1 45625
0 45627 7 1 2 103813 91638
0 45628 7 1 2 100901 45627
0 45629 7 1 2 96329 45628
0 45630 5 1 1 45629
0 45631 7 1 2 45626 45630
0 45632 5 1 1 45631
0 45633 7 1 2 67761 45632
0 45634 5 1 1 45633
0 45635 7 2 2 72176 76964
0 45636 7 3 2 74564 79815
0 45637 5 1 1 105537
0 45638 7 1 2 72755 105538
0 45639 7 1 2 105535 45638
0 45640 7 1 2 105344 45639
0 45641 5 1 1 45640
0 45642 7 1 2 45634 45641
0 45643 5 1 1 45642
0 45644 7 1 2 82996 45643
0 45645 5 1 1 45644
0 45646 7 1 2 75440 103103
0 45647 5 1 1 45646
0 45648 7 1 2 87354 45647
0 45649 5 1 1 45648
0 45650 7 1 2 80030 45649
0 45651 5 1 1 45650
0 45652 7 1 2 82797 100899
0 45653 5 1 1 45652
0 45654 7 1 2 80375 45653
0 45655 5 1 1 45654
0 45656 7 2 2 87252 88336
0 45657 5 1 1 105540
0 45658 7 1 2 80249 101388
0 45659 5 1 1 45658
0 45660 7 1 2 45657 45659
0 45661 5 3 1 45660
0 45662 7 1 2 81768 105542
0 45663 5 1 1 45662
0 45664 7 1 2 27963 45663
0 45665 7 1 2 45655 45664
0 45666 5 1 1 45665
0 45667 7 1 2 71165 45666
0 45668 5 1 1 45667
0 45669 7 1 2 45651 45668
0 45670 5 2 1 45669
0 45671 7 1 2 81345 105545
0 45672 5 1 1 45671
0 45673 7 1 2 91991 105016
0 45674 5 1 1 45673
0 45675 7 1 2 85598 96462
0 45676 7 1 2 97551 45675
0 45677 5 1 1 45676
0 45678 7 1 2 101381 45677
0 45679 5 1 1 45678
0 45680 7 1 2 45674 45679
0 45681 5 2 1 45680
0 45682 7 1 2 80192 105547
0 45683 5 1 1 45682
0 45684 7 1 2 45672 45683
0 45685 5 1 1 45684
0 45686 7 1 2 66889 45685
0 45687 5 1 1 45686
0 45688 7 1 2 80376 83566
0 45689 5 1 1 45688
0 45690 7 1 2 104589 45689
0 45691 5 1 1 45690
0 45692 7 1 2 79285 45691
0 45693 5 1 1 45692
0 45694 7 1 2 69605 89039
0 45695 5 1 1 45694
0 45696 7 1 2 104302 45695
0 45697 5 1 1 45696
0 45698 7 1 2 45693 45697
0 45699 5 1 1 45698
0 45700 7 2 2 91639 45699
0 45701 7 1 2 87429 105549
0 45702 5 1 1 45701
0 45703 7 1 2 45687 45702
0 45704 5 1 1 45703
0 45705 7 1 2 73865 45704
0 45706 5 1 1 45705
0 45707 7 1 2 88587 105546
0 45708 5 1 1 45707
0 45709 7 1 2 88231 105548
0 45710 5 1 1 45709
0 45711 7 1 2 45708 45710
0 45712 5 1 1 45711
0 45713 7 1 2 90353 45712
0 45714 5 1 1 45713
0 45715 7 4 2 91645 97160
0 45716 7 1 2 105550 105551
0 45717 5 1 1 45716
0 45718 7 1 2 99193 102906
0 45719 5 1 1 45718
0 45720 7 1 2 77382 104150
0 45721 5 1 1 45720
0 45722 7 3 2 64856 68702
0 45723 5 2 1 105555
0 45724 7 1 2 66780 105558
0 45725 5 1 1 45724
0 45726 7 1 2 45721 45725
0 45727 7 2 2 45719 45726
0 45728 7 1 2 79667 105482
0 45729 7 1 2 105560 45728
0 45730 5 1 1 45729
0 45731 7 1 2 81009 105447
0 45732 5 1 1 45731
0 45733 7 2 2 82269 45732
0 45734 7 1 2 86548 105562
0 45735 5 1 1 45734
0 45736 7 1 2 95514 104907
0 45737 7 1 2 100028 45736
0 45738 5 1 1 45737
0 45739 7 1 2 45735 45738
0 45740 5 1 1 45739
0 45741 7 1 2 91393 105510
0 45742 7 1 2 45740 45741
0 45743 5 1 1 45742
0 45744 7 1 2 45730 45743
0 45745 5 1 1 45744
0 45746 7 1 2 69002 45745
0 45747 5 1 1 45746
0 45748 7 1 2 88232 90354
0 45749 7 1 2 105561 45748
0 45750 5 1 1 45749
0 45751 7 1 2 45747 45750
0 45752 5 1 1 45751
0 45753 7 1 2 70518 45752
0 45754 5 1 1 45753
0 45755 7 1 2 45717 45754
0 45756 7 1 2 45714 45755
0 45757 7 1 2 45706 45756
0 45758 5 1 1 45757
0 45759 7 1 2 67762 45758
0 45760 5 1 1 45759
0 45761 7 2 2 96199 75536
0 45762 5 1 1 105564
0 45763 7 1 2 90341 105565
0 45764 5 1 1 45763
0 45765 7 1 2 80644 99288
0 45766 7 1 2 96833 45765
0 45767 5 1 1 45766
0 45768 7 1 2 45764 45767
0 45769 5 1 1 45768
0 45770 7 1 2 71166 45769
0 45771 5 1 1 45770
0 45772 7 1 2 69003 90342
0 45773 5 1 1 45772
0 45774 7 1 2 105380 45773
0 45775 5 1 1 45774
0 45776 7 1 2 69963 101230
0 45777 5 2 1 45776
0 45778 7 1 2 85638 78054
0 45779 5 1 1 45778
0 45780 7 1 2 105566 45779
0 45781 5 1 1 45780
0 45782 7 1 2 72177 45781
0 45783 7 1 2 45775 45782
0 45784 5 1 1 45783
0 45785 7 1 2 45771 45784
0 45786 5 1 1 45785
0 45787 7 1 2 66890 45786
0 45788 5 1 1 45787
0 45789 7 1 2 77732 91200
0 45790 7 1 2 94474 91661
0 45791 7 1 2 45789 45790
0 45792 7 1 2 102171 105375
0 45793 7 1 2 45791 45792
0 45794 5 1 1 45793
0 45795 7 1 2 45788 45794
0 45796 5 1 1 45795
0 45797 7 1 2 81483 45796
0 45798 5 1 1 45797
0 45799 7 1 2 105494 105483
0 45800 5 1 1 45799
0 45801 7 1 2 100803 76123
0 45802 7 1 2 90251 45801
0 45803 5 1 1 45802
0 45804 7 1 2 45800 45803
0 45805 5 1 1 45804
0 45806 7 1 2 69964 45805
0 45807 5 1 1 45806
0 45808 7 1 2 97776 94092
0 45809 7 1 2 96195 45808
0 45810 5 1 1 45809
0 45811 7 1 2 45807 45810
0 45812 5 1 1 45811
0 45813 7 1 2 70250 45812
0 45814 5 1 1 45813
0 45815 7 1 2 105498 105484
0 45816 5 1 1 45815
0 45817 7 1 2 45814 45816
0 45818 5 1 1 45817
0 45819 7 1 2 69004 45818
0 45820 5 1 1 45819
0 45821 7 1 2 79036 95973
0 45822 7 1 2 90252 45821
0 45823 7 1 2 80944 45822
0 45824 5 1 1 45823
0 45825 7 1 2 45820 45824
0 45826 5 1 1 45825
0 45827 7 1 2 94914 45826
0 45828 5 1 1 45827
0 45829 7 1 2 81146 92132
0 45830 7 2 2 76663 45829
0 45831 7 1 2 105552 105568
0 45832 5 1 1 45831
0 45833 7 1 2 105465 45832
0 45834 5 1 1 45833
0 45835 7 1 2 68495 45834
0 45836 5 1 1 45835
0 45837 7 2 2 71958 89354
0 45838 7 1 2 81141 105570
0 45839 7 1 2 105553 45838
0 45840 5 1 1 45839
0 45841 7 1 2 45836 45840
0 45842 5 1 1 45841
0 45843 7 1 2 69606 45842
0 45844 5 1 1 45843
0 45845 7 1 2 89953 105463
0 45846 5 1 1 45845
0 45847 7 1 2 104164 97704
0 45848 5 1 1 45847
0 45849 7 1 2 97258 105569
0 45850 5 1 1 45849
0 45851 7 1 2 45848 45850
0 45852 5 1 1 45851
0 45853 7 1 2 68496 45852
0 45854 5 1 1 45853
0 45855 7 1 2 90722 97646
0 45856 7 1 2 105571 45855
0 45857 5 1 1 45856
0 45858 7 1 2 45854 45857
0 45859 5 1 1 45858
0 45860 7 1 2 73866 45859
0 45861 5 1 1 45860
0 45862 7 1 2 45846 45861
0 45863 7 1 2 45844 45862
0 45864 5 1 1 45863
0 45865 7 1 2 86070 45864
0 45866 5 1 1 45865
0 45867 7 1 2 45828 45866
0 45868 5 1 1 45867
0 45869 7 1 2 83755 45868
0 45870 5 1 1 45869
0 45871 7 1 2 45798 45870
0 45872 7 1 2 45760 45871
0 45873 7 1 2 45645 45872
0 45874 5 1 1 45873
0 45875 7 1 2 67399 45874
0 45876 5 1 1 45875
0 45877 7 1 2 82505 45876
0 45878 5 1 1 45877
0 45879 7 1 2 68497 75680
0 45880 5 1 1 45879
0 45881 7 1 2 80377 97152
0 45882 7 1 2 104313 45881
0 45883 5 1 1 45882
0 45884 7 1 2 45880 45883
0 45885 5 1 1 45884
0 45886 7 1 2 70251 45885
0 45887 5 1 1 45886
0 45888 7 1 2 68498 80501
0 45889 5 1 1 45888
0 45890 7 1 2 64857 45889
0 45891 5 1 1 45890
0 45892 7 1 2 75681 45891
0 45893 5 1 1 45892
0 45894 7 1 2 45887 45893
0 45895 5 1 1 45894
0 45896 7 1 2 68891 45895
0 45897 5 1 1 45896
0 45898 7 1 2 71859 97573
0 45899 5 1 1 45898
0 45900 7 1 2 75156 90981
0 45901 5 1 1 45900
0 45902 7 1 2 45899 45901
0 45903 5 1 1 45902
0 45904 7 1 2 68499 45903
0 45905 5 1 1 45904
0 45906 7 1 2 4908 45905
0 45907 5 1 1 45906
0 45908 7 1 2 78184 45907
0 45909 5 1 1 45908
0 45910 7 1 2 45897 45909
0 45911 5 1 1 45910
0 45912 7 1 2 69607 45911
0 45913 5 1 1 45912
0 45914 7 1 2 89954 97575
0 45915 5 1 1 45914
0 45916 7 1 2 45913 45915
0 45917 5 1 1 45916
0 45918 7 1 2 72756 45917
0 45919 5 1 1 45918
0 45920 7 2 2 79684 97153
0 45921 7 1 2 81484 104189
0 45922 5 1 1 45921
0 45923 7 2 2 92355 83636
0 45924 7 1 2 95923 105574
0 45925 5 1 1 45924
0 45926 7 1 2 45922 45925
0 45927 5 1 1 45926
0 45928 7 1 2 105572 45927
0 45929 5 1 1 45928
0 45930 7 1 2 78708 84682
0 45931 5 1 1 45930
0 45932 7 2 2 64485 82267
0 45933 5 1 1 105576
0 45934 7 1 2 72757 105577
0 45935 5 1 1 45934
0 45936 7 1 2 70252 104236
0 45937 7 1 2 45935 45936
0 45938 5 1 1 45937
0 45939 7 1 2 45931 45938
0 45940 5 1 1 45939
0 45941 7 1 2 71860 45940
0 45942 5 1 1 45941
0 45943 7 1 2 83331 81421
0 45944 5 2 1 45943
0 45945 7 1 2 81177 96034
0 45946 5 1 1 45945
0 45947 7 1 2 105578 45946
0 45948 5 1 1 45947
0 45949 7 1 2 70253 45948
0 45950 5 1 1 45949
0 45951 7 1 2 37164 45950
0 45952 5 1 1 45951
0 45953 7 1 2 68703 45952
0 45954 5 1 1 45953
0 45955 7 1 2 45942 45954
0 45956 5 1 1 45955
0 45957 7 1 2 81346 45956
0 45958 5 1 1 45957
0 45959 7 1 2 79830 82802
0 45960 5 1 1 45959
0 45961 7 1 2 84942 45960
0 45962 5 1 1 45961
0 45963 7 1 2 67763 96901
0 45964 5 1 1 45963
0 45965 7 1 2 68500 45964
0 45966 7 1 2 45962 45965
0 45967 5 1 1 45966
0 45968 7 1 2 67764 104908
0 45969 5 1 1 45968
0 45970 7 1 2 45967 45969
0 45971 5 1 1 45970
0 45972 7 1 2 80193 45971
0 45973 5 1 1 45972
0 45974 7 1 2 45958 45973
0 45975 5 1 1 45974
0 45976 7 1 2 66891 45975
0 45977 5 1 1 45976
0 45978 7 1 2 45929 45977
0 45979 5 1 1 45978
0 45980 7 1 2 70519 45979
0 45981 5 1 1 45980
0 45982 7 1 2 87869 91119
0 45983 7 1 2 97254 45982
0 45984 5 1 1 45983
0 45985 7 1 2 100029 84589
0 45986 7 1 2 81347 45985
0 45987 5 1 1 45986
0 45988 7 1 2 45984 45987
0 45989 5 1 1 45988
0 45990 7 1 2 93805 45989
0 45991 5 1 1 45990
0 45992 7 1 2 64486 82302
0 45993 5 1 1 45992
0 45994 7 1 2 81178 94214
0 45995 5 1 1 45994
0 45996 7 1 2 45993 45995
0 45997 5 1 1 45996
0 45998 7 1 2 81348 45997
0 45999 5 1 1 45998
0 46000 7 1 2 96007 80194
0 46001 7 1 2 95790 46000
0 46002 5 1 1 46001
0 46003 7 1 2 45999 46002
0 46004 5 1 1 46003
0 46005 7 1 2 66892 46004
0 46006 5 1 1 46005
0 46007 7 1 2 88825 92133
0 46008 7 2 2 92403 86092
0 46009 7 1 2 84154 105580
0 46010 7 1 2 46007 46009
0 46011 5 1 1 46010
0 46012 7 1 2 46006 46011
0 46013 5 1 1 46012
0 46014 7 1 2 67765 46013
0 46015 5 1 1 46014
0 46016 7 1 2 45991 46015
0 46017 7 1 2 45981 46016
0 46018 7 1 2 45919 46017
0 46019 5 1 1 46018
0 46020 7 1 2 71167 46019
0 46021 5 1 1 46020
0 46022 7 1 2 66071 101721
0 46023 5 1 1 46022
0 46024 7 1 2 104074 46023
0 46025 5 1 1 46024
0 46026 7 1 2 67766 46025
0 46027 5 1 1 46026
0 46028 7 1 2 69965 105339
0 46029 5 1 1 46028
0 46030 7 1 2 46027 46029
0 46031 5 1 1 46030
0 46032 7 1 2 69608 46031
0 46033 5 1 1 46032
0 46034 7 1 2 89029 103662
0 46035 5 1 1 46034
0 46036 7 1 2 46033 46035
0 46037 5 1 1 46036
0 46038 7 1 2 81349 46037
0 46039 5 1 1 46038
0 46040 7 1 2 82141 86752
0 46041 5 1 1 46040
0 46042 7 1 2 19038 78038
0 46043 5 1 1 46042
0 46044 7 1 2 71861 10250
0 46045 7 1 2 46043 46044
0 46046 5 1 1 46045
0 46047 7 1 2 46041 46046
0 46048 5 1 1 46047
0 46049 7 1 2 75441 46048
0 46050 5 1 1 46049
0 46051 7 2 2 71862 84187
0 46052 7 1 2 87129 105582
0 46053 5 1 1 46052
0 46054 7 1 2 91434 105067
0 46055 5 1 1 46054
0 46056 7 1 2 102887 98915
0 46057 5 1 1 46056
0 46058 7 1 2 46055 46057
0 46059 5 1 1 46058
0 46060 7 1 2 68501 46059
0 46061 5 1 1 46060
0 46062 7 1 2 46053 46061
0 46063 7 1 2 46050 46062
0 46064 5 1 1 46063
0 46065 7 1 2 69609 46064
0 46066 5 1 1 46065
0 46067 7 2 2 88826 105225
0 46068 5 1 1 105584
0 46069 7 1 2 67767 75442
0 46070 7 1 2 105585 46069
0 46071 5 1 1 46070
0 46072 7 1 2 46066 46071
0 46073 5 1 1 46072
0 46074 7 1 2 80195 46073
0 46075 5 1 1 46074
0 46076 7 1 2 46039 46075
0 46077 5 1 1 46076
0 46078 7 1 2 66893 46077
0 46079 5 1 1 46078
0 46080 7 2 2 89023 78438
0 46081 7 1 2 80031 105573
0 46082 7 1 2 105586 46081
0 46083 5 1 1 46082
0 46084 7 1 2 72465 46083
0 46085 7 1 2 46079 46084
0 46086 7 1 2 46021 46085
0 46087 5 1 1 46086
0 46088 7 1 2 98321 104590
0 46089 5 1 1 46088
0 46090 7 1 2 79286 83731
0 46091 7 1 2 46089 46090
0 46092 5 2 1 46091
0 46093 7 1 2 64487 105341
0 46094 5 1 1 46093
0 46095 7 1 2 81010 46094
0 46096 5 1 1 46095
0 46097 7 1 2 77477 89040
0 46098 5 1 1 46097
0 46099 7 1 2 64858 11305
0 46100 7 1 2 46098 46099
0 46101 7 1 2 46096 46100
0 46102 5 1 1 46101
0 46103 7 1 2 105588 46102
0 46104 5 1 1 46103
0 46105 7 1 2 79152 46104
0 46106 5 1 1 46105
0 46107 7 1 2 83012 4164
0 46108 5 4 1 46107
0 46109 7 3 2 75443 105590
0 46110 5 1 1 105594
0 46111 7 1 2 64859 105595
0 46112 5 1 1 46111
0 46113 7 1 2 68704 94208
0 46114 5 1 1 46113
0 46115 7 1 2 46112 46114
0 46116 5 1 1 46115
0 46117 7 1 2 66072 95422
0 46118 7 1 2 46116 46117
0 46119 5 1 1 46118
0 46120 7 1 2 46106 46119
0 46121 5 1 1 46120
0 46122 7 1 2 74454 46121
0 46123 5 1 1 46122
0 46124 7 1 2 104075 104048
0 46125 5 1 1 46124
0 46126 7 1 2 83732 97705
0 46127 7 1 2 46125 46126
0 46128 5 1 1 46127
0 46129 7 1 2 67400 46128
0 46130 7 1 2 46123 46129
0 46131 5 1 1 46130
0 46132 7 1 2 73867 46131
0 46133 7 1 2 46087 46132
0 46134 5 1 1 46133
0 46135 7 1 2 82142 98836
0 46136 5 1 1 46135
0 46137 7 1 2 87631 95403
0 46138 5 1 1 46137
0 46139 7 1 2 46136 46138
0 46140 5 1 1 46139
0 46141 7 1 2 70520 46140
0 46142 5 1 1 46141
0 46143 7 2 2 83046 82143
0 46144 5 1 1 105597
0 46145 7 1 2 105579 46144
0 46146 5 1 1 46145
0 46147 7 1 2 80378 46146
0 46148 5 1 1 46147
0 46149 7 1 2 46142 46148
0 46150 5 1 1 46149
0 46151 7 1 2 77478 46150
0 46152 5 1 1 46151
0 46153 7 1 2 69966 105587
0 46154 5 1 1 46153
0 46155 7 1 2 85639 92550
0 46156 5 1 1 46155
0 46157 7 1 2 46154 46156
0 46158 7 1 2 46152 46157
0 46159 5 1 1 46158
0 46160 7 1 2 70254 46159
0 46161 5 1 1 46160
0 46162 7 1 2 101722 78516
0 46163 5 1 1 46162
0 46164 7 1 2 82144 105331
0 46165 5 1 1 46164
0 46166 7 1 2 83805 81485
0 46167 5 1 1 46166
0 46168 7 1 2 46165 46167
0 46169 5 1 1 46168
0 46170 7 1 2 68502 46169
0 46171 5 1 1 46170
0 46172 7 1 2 101710 98916
0 46173 5 1 1 46172
0 46174 7 1 2 46171 46173
0 46175 5 1 1 46174
0 46176 7 1 2 71168 46175
0 46177 5 1 1 46176
0 46178 7 1 2 46163 46177
0 46179 7 1 2 46161 46178
0 46180 5 1 1 46179
0 46181 7 1 2 88588 46180
0 46182 5 1 1 46181
0 46183 7 1 2 80379 87130
0 46184 5 1 1 46183
0 46185 7 1 2 102888 97542
0 46186 5 1 1 46185
0 46187 7 1 2 46184 46186
0 46188 5 1 1 46187
0 46189 7 1 2 69610 46188
0 46190 5 1 1 46189
0 46191 7 1 2 64860 90115
0 46192 7 1 2 94325 46191
0 46193 5 1 1 46192
0 46194 7 1 2 46068 46193
0 46195 5 1 1 46194
0 46196 7 1 2 75444 46195
0 46197 5 1 1 46196
0 46198 7 1 2 103471 104911
0 46199 5 1 1 46198
0 46200 7 1 2 77525 46199
0 46201 5 1 1 46200
0 46202 7 1 2 46197 46201
0 46203 7 1 2 46190 46202
0 46204 5 1 1 46203
0 46205 7 1 2 67768 46204
0 46206 5 1 1 46205
0 46207 7 2 2 81916 77185
0 46208 5 1 1 105599
0 46209 7 1 2 80459 87063
0 46210 5 1 1 46209
0 46211 7 1 2 46208 46210
0 46212 5 1 1 46211
0 46213 7 1 2 81422 46212
0 46214 5 1 1 46213
0 46215 7 1 2 46206 46214
0 46216 5 1 1 46215
0 46217 7 1 2 88233 46216
0 46218 5 1 1 46217
0 46219 7 1 2 46182 46218
0 46220 5 1 1 46219
0 46221 7 1 2 72466 46220
0 46222 5 1 1 46221
0 46223 7 1 2 99936 90407
0 46224 5 1 1 46223
0 46225 7 1 2 89884 105591
0 46226 5 1 1 46225
0 46227 7 1 2 46224 46226
0 46228 5 1 1 46227
0 46229 7 1 2 64861 46228
0 46230 5 1 1 46229
0 46231 7 1 2 101723 88589
0 46232 5 1 1 46231
0 46233 7 1 2 46232 45762
0 46234 5 1 1 46233
0 46235 7 1 2 64488 46234
0 46236 5 1 1 46235
0 46237 7 1 2 46230 46236
0 46238 5 1 1 46237
0 46239 7 1 2 97753 46238
0 46240 5 1 1 46239
0 46241 7 1 2 46222 46240
0 46242 5 1 1 46241
0 46243 7 1 2 90355 46242
0 46244 5 1 1 46243
0 46245 7 1 2 64862 93532
0 46246 7 1 2 89048 46245
0 46247 5 1 1 46246
0 46248 7 1 2 105589 46247
0 46249 5 1 1 46248
0 46250 7 1 2 88234 46249
0 46251 5 1 1 46250
0 46252 7 1 2 83007 78439
0 46253 5 1 1 46252
0 46254 7 1 2 66781 78497
0 46255 7 1 2 98662 46254
0 46256 7 1 2 98353 46255
0 46257 5 1 1 46256
0 46258 7 1 2 46253 46257
0 46259 5 1 1 46258
0 46260 7 1 2 64489 103409
0 46261 7 1 2 92694 46260
0 46262 7 1 2 46259 46261
0 46263 5 1 1 46262
0 46264 7 1 2 46251 46263
0 46265 5 1 1 46264
0 46266 7 1 2 67401 46265
0 46267 5 1 1 46266
0 46268 7 1 2 80901 89738
0 46269 5 1 1 46268
0 46270 7 1 2 89700 6243
0 46271 5 1 1 46270
0 46272 7 1 2 101257 46271
0 46273 5 1 1 46272
0 46274 7 1 2 46269 46273
0 46275 5 1 1 46274
0 46276 7 1 2 70255 46275
0 46277 5 1 1 46276
0 46278 7 1 2 104101 94527
0 46279 5 1 1 46278
0 46280 7 1 2 46277 46279
0 46281 5 1 1 46280
0 46282 7 1 2 68705 46281
0 46283 5 1 1 46282
0 46284 7 1 2 89635 79328
0 46285 7 1 2 102440 46284
0 46286 5 1 1 46285
0 46287 7 1 2 46283 46286
0 46288 5 1 1 46287
0 46289 7 1 2 98724 46288
0 46290 5 1 1 46289
0 46291 7 2 2 80738 98304
0 46292 5 1 1 105601
0 46293 7 1 2 100846 46292
0 46294 5 1 1 46293
0 46295 7 1 2 98616 88235
0 46296 7 1 2 99148 46295
0 46297 7 1 2 46294 46296
0 46298 5 1 1 46297
0 46299 7 1 2 79984 92003
0 46300 7 1 2 98410 46299
0 46301 7 1 2 98535 46300
0 46302 5 1 1 46301
0 46303 7 1 2 46298 46302
0 46304 7 1 2 46290 46303
0 46305 7 1 2 46267 46304
0 46306 5 1 1 46305
0 46307 7 1 2 105145 46306
0 46308 5 1 1 46307
0 46309 7 1 2 82462 46308
0 46310 7 1 2 46244 46309
0 46311 7 1 2 46134 46310
0 46312 5 1 1 46311
0 46313 7 1 2 74431 76094
0 46314 7 1 2 46312 46313
0 46315 7 1 2 45878 46314
0 46316 5 1 1 46315
0 46317 7 1 2 45579 46316
0 46318 7 1 2 45107 46317
0 46319 5 1 1 46318
0 46320 7 1 2 72064 46319
0 46321 5 1 1 46320
0 46322 7 3 2 67132 90294
0 46323 7 1 2 101508 101724
0 46324 5 1 1 46323
0 46325 7 1 2 100798 105456
0 46326 5 1 1 46325
0 46327 7 1 2 46324 46326
0 46328 5 1 1 46327
0 46329 7 1 2 105269 46328
0 46330 5 1 1 46329
0 46331 7 1 2 78517 105602
0 46332 5 1 1 46331
0 46333 7 1 2 100841 93350
0 46334 5 1 1 46333
0 46335 7 1 2 46332 46334
0 46336 5 1 1 46335
0 46337 7 1 2 64863 46336
0 46338 5 1 1 46337
0 46339 7 1 2 93751 104431
0 46340 5 1 1 46339
0 46341 7 1 2 82706 46340
0 46342 5 1 1 46341
0 46343 7 1 2 67769 46342
0 46344 5 1 1 46343
0 46345 7 1 2 85614 88002
0 46346 7 1 2 97975 46345
0 46347 5 1 1 46346
0 46348 7 1 2 46344 46347
0 46349 5 1 1 46348
0 46350 7 1 2 69967 46349
0 46351 5 1 1 46350
0 46352 7 1 2 67770 82699
0 46353 7 1 2 94285 46352
0 46354 5 1 1 46353
0 46355 7 1 2 46351 46354
0 46356 7 1 2 46338 46355
0 46357 5 1 1 46356
0 46358 7 1 2 67402 46357
0 46359 5 1 1 46358
0 46360 7 4 2 67771 96920
0 46361 7 1 2 66073 104162
0 46362 5 1 1 46361
0 46363 7 1 2 86071 46362
0 46364 5 1 1 46363
0 46365 7 1 2 78066 46364
0 46366 5 1 1 46365
0 46367 7 1 2 68503 46366
0 46368 5 1 1 46367
0 46369 7 1 2 77479 83030
0 46370 5 1 1 46369
0 46371 7 1 2 1450 46370
0 46372 7 1 2 46368 46371
0 46373 5 1 1 46372
0 46374 7 1 2 105606 46373
0 46375 5 1 1 46374
0 46376 7 1 2 46359 46375
0 46377 5 1 1 46376
0 46378 7 1 2 70875 46377
0 46379 5 1 1 46378
0 46380 7 1 2 46330 46379
0 46381 5 1 1 46380
0 46382 7 1 2 65653 46381
0 46383 5 1 1 46382
0 46384 7 2 2 98461 102070
0 46385 7 1 2 102027 105305
0 46386 7 1 2 105610 46385
0 46387 5 1 1 46386
0 46388 7 1 2 46383 46387
0 46389 5 1 1 46388
0 46390 7 1 2 105603 46389
0 46391 5 1 1 46390
0 46392 7 1 2 64864 101767
0 46393 5 1 1 46392
0 46394 7 1 2 84628 87259
0 46395 5 1 1 46394
0 46396 7 1 2 46393 46395
0 46397 5 1 1 46396
0 46398 7 1 2 96763 46397
0 46399 5 1 1 46398
0 46400 7 1 2 77480 101262
0 46401 5 1 1 46400
0 46402 7 1 2 86844 95781
0 46403 5 1 1 46402
0 46404 7 1 2 46401 46403
0 46405 5 1 1 46404
0 46406 7 1 2 97058 46405
0 46407 5 1 1 46406
0 46408 7 1 2 46399 46407
0 46409 5 1 1 46408
0 46410 7 1 2 68706 46409
0 46411 5 1 1 46410
0 46412 7 1 2 101139 103524
0 46413 5 1 1 46412
0 46414 7 1 2 46411 46413
0 46415 5 1 1 46414
0 46416 7 1 2 69254 46415
0 46417 5 1 1 46416
0 46418 7 2 2 68707 104703
0 46419 7 1 2 94353 105612
0 46420 5 1 1 46419
0 46421 7 1 2 98537 46420
0 46422 5 1 1 46421
0 46423 7 1 2 69968 46422
0 46424 5 1 1 46423
0 46425 7 1 2 82700 103443
0 46426 5 1 1 46425
0 46427 7 1 2 46424 46426
0 46428 5 1 1 46427
0 46429 7 1 2 98767 46428
0 46430 5 1 1 46429
0 46431 7 1 2 46417 46430
0 46432 5 1 1 46431
0 46433 7 1 2 70876 46432
0 46434 5 1 1 46433
0 46435 7 1 2 101509 103525
0 46436 5 1 1 46435
0 46437 7 2 2 77186 86845
0 46438 7 1 2 90005 105614
0 46439 5 1 1 46438
0 46440 7 1 2 46436 46439
0 46441 5 1 1 46440
0 46442 7 1 2 105270 46441
0 46443 5 1 1 46442
0 46444 7 1 2 46434 46443
0 46445 5 1 1 46444
0 46446 7 1 2 96370 46445
0 46447 5 1 1 46446
0 46448 7 4 2 69611 65690
0 46449 7 3 2 63980 105616
0 46450 7 1 2 95341 98768
0 46451 7 1 2 105620 46450
0 46452 5 1 1 46451
0 46453 7 1 2 94666 93325
0 46454 7 1 2 105611 46453
0 46455 5 1 1 46454
0 46456 7 1 2 46452 46455
0 46457 5 1 1 46456
0 46458 7 1 2 64195 46457
0 46459 5 1 1 46458
0 46460 7 1 2 96764 92990
0 46461 5 1 1 46460
0 46462 7 1 2 103671 46461
0 46463 5 1 1 46462
0 46464 7 1 2 97854 46463
0 46465 5 1 1 46464
0 46466 7 1 2 93060 99067
0 46467 5 3 1 46466
0 46468 7 1 2 46465 105623
0 46469 5 1 1 46468
0 46470 7 2 2 69255 46469
0 46471 5 1 1 105626
0 46472 7 1 2 88920 105627
0 46473 5 1 1 46472
0 46474 7 1 2 46459 46473
0 46475 5 2 1 46474
0 46476 7 1 2 69005 105628
0 46477 5 1 1 46476
0 46478 7 1 2 99464 101036
0 46479 5 3 1 46478
0 46480 7 1 2 46471 105630
0 46481 5 1 1 46480
0 46482 7 1 2 92153 46481
0 46483 5 1 1 46482
0 46484 7 1 2 46477 46483
0 46485 5 1 1 46484
0 46486 7 1 2 65654 46485
0 46487 5 1 1 46486
0 46488 7 1 2 46447 46487
0 46489 5 1 1 46488
0 46490 7 1 2 72178 46489
0 46491 5 1 1 46490
0 46492 7 3 2 89676 73831
0 46493 5 1 1 105633
0 46494 7 1 2 96286 17394
0 46495 5 1 1 46494
0 46496 7 1 2 88921 46495
0 46497 5 1 1 46496
0 46498 7 1 2 46493 46497
0 46499 5 1 1 46498
0 46500 7 1 2 63914 46499
0 46501 5 1 1 46500
0 46502 7 4 2 88590 91533
0 46503 7 1 2 68708 105636
0 46504 5 1 1 46503
0 46505 7 1 2 46501 46504
0 46506 5 1 1 46505
0 46507 7 1 2 83756 105450
0 46508 5 1 1 46507
0 46509 7 1 2 100040 104239
0 46510 5 3 1 46509
0 46511 7 2 2 64865 78384
0 46512 7 1 2 89248 105643
0 46513 5 1 1 46512
0 46514 7 1 2 105640 46513
0 46515 7 1 2 46508 46514
0 46516 5 1 1 46515
0 46517 7 1 2 71863 46516
0 46518 7 1 2 46506 46517
0 46519 5 1 1 46518
0 46520 7 4 2 88236 90318
0 46521 7 2 2 68709 105645
0 46522 7 1 2 76970 91735
0 46523 7 1 2 78461 46522
0 46524 7 1 2 45933 46523
0 46525 5 1 1 46524
0 46526 7 1 2 88735 105644
0 46527 5 1 1 46526
0 46528 7 1 2 105641 46527
0 46529 7 1 2 46525 46528
0 46530 5 1 1 46529
0 46531 7 1 2 105649 46530
0 46532 5 1 1 46531
0 46533 7 1 2 46519 46532
0 46534 5 1 1 46533
0 46535 7 1 2 70521 46534
0 46536 5 1 1 46535
0 46537 7 2 2 83047 80032
0 46538 5 1 1 105651
0 46539 7 1 2 105445 46538
0 46540 5 1 1 46539
0 46541 7 1 2 78462 46540
0 46542 5 1 1 46541
0 46543 7 1 2 78385 105598
0 46544 5 1 1 46543
0 46545 7 1 2 105642 46544
0 46546 7 1 2 46542 46545
0 46547 5 1 1 46546
0 46548 7 1 2 71864 105650
0 46549 7 1 2 46547 46548
0 46550 5 1 1 46549
0 46551 7 1 2 46536 46550
0 46552 5 1 1 46551
0 46553 7 1 2 67403 46552
0 46554 5 1 1 46553
0 46555 7 1 2 101754 89677
0 46556 5 1 1 46555
0 46557 7 1 2 65655 85185
0 46558 5 1 1 46557
0 46559 7 1 2 46556 46558
0 46560 5 1 1 46559
0 46561 7 1 2 88922 46560
0 46562 5 1 1 46561
0 46563 7 1 2 71865 105634
0 46564 5 1 1 46563
0 46565 7 1 2 46562 46564
0 46566 5 1 1 46565
0 46567 7 1 2 70522 46566
0 46568 5 1 1 46567
0 46569 7 1 2 91534 96632
0 46570 5 1 1 46569
0 46571 7 1 2 46568 46570
0 46572 5 1 1 46571
0 46573 7 1 2 63915 46572
0 46574 5 1 1 46573
0 46575 7 1 2 86683 105637
0 46576 5 1 1 46575
0 46577 7 1 2 46574 46576
0 46578 5 1 1 46577
0 46579 7 1 2 80885 80838
0 46580 7 1 2 97224 46579
0 46581 7 1 2 46578 46580
0 46582 5 1 1 46581
0 46583 7 1 2 46554 46582
0 46584 5 1 1 46583
0 46585 7 1 2 70256 46584
0 46586 5 1 1 46585
0 46587 7 1 2 82262 102071
0 46588 5 1 1 46587
0 46589 7 1 2 101258 78518
0 46590 5 1 1 46589
0 46591 7 1 2 46588 46590
0 46592 5 1 1 46591
0 46593 7 2 2 65188 96371
0 46594 7 4 2 65494 84599
0 46595 7 1 2 97205 105655
0 46596 7 1 2 105653 46595
0 46597 7 1 2 46592 46596
0 46598 5 1 1 46597
0 46599 7 1 2 46586 46598
0 46600 5 1 1 46599
0 46601 7 1 2 74432 46600
0 46602 5 1 1 46601
0 46603 7 1 2 46491 46602
0 46604 7 1 2 46391 46603
0 46605 5 1 1 46604
0 46606 7 1 2 66365 46605
0 46607 5 1 1 46606
0 46608 7 1 2 99410 79913
0 46609 5 1 1 46608
0 46610 7 1 2 99389 101857
0 46611 5 1 1 46610
0 46612 7 1 2 46609 46611
0 46613 5 1 1 46612
0 46614 7 1 2 71467 46613
0 46615 5 1 1 46614
0 46616 7 1 2 73565 99755
0 46617 7 1 2 105349 46616
0 46618 5 1 1 46617
0 46619 7 1 2 46615 46618
0 46620 5 1 1 46619
0 46621 7 1 2 77481 46620
0 46622 5 1 1 46621
0 46623 7 1 2 69256 97868
0 46624 5 1 1 46623
0 46625 7 1 2 14507 46624
0 46626 5 4 1 46625
0 46627 7 1 2 75445 104061
0 46628 5 1 1 46627
0 46629 7 1 2 94708 46628
0 46630 5 1 1 46629
0 46631 7 1 2 68710 46630
0 46632 5 1 1 46631
0 46633 7 1 2 101734 46632
0 46634 5 1 1 46633
0 46635 7 1 2 105659 46634
0 46636 5 1 1 46635
0 46637 7 1 2 82843 105660
0 46638 5 1 1 46637
0 46639 7 1 2 100381 100481
0 46640 5 1 1 46639
0 46641 7 1 2 46638 46640
0 46642 5 1 1 46641
0 46643 7 1 2 85640 46642
0 46644 5 1 1 46643
0 46645 7 1 2 73927 94475
0 46646 7 1 2 104422 46645
0 46647 5 1 1 46646
0 46648 7 1 2 46644 46647
0 46649 7 1 2 46636 46648
0 46650 5 1 1 46649
0 46651 7 1 2 72467 46650
0 46652 5 1 1 46651
0 46653 7 1 2 67404 98529
0 46654 7 1 2 100842 46653
0 46655 5 1 1 46654
0 46656 7 1 2 46652 46655
0 46657 5 1 1 46656
0 46658 7 1 2 69969 46657
0 46659 5 1 1 46658
0 46660 7 1 2 74433 98260
0 46661 5 1 1 46660
0 46662 7 1 2 67405 98525
0 46663 5 1 1 46662
0 46664 7 2 2 99761 46663
0 46665 5 1 1 105663
0 46666 7 1 2 46661 105664
0 46667 5 6 1 46666
0 46668 7 1 2 105420 105665
0 46669 5 1 1 46668
0 46670 7 2 2 72468 83551
0 46671 7 1 2 105671 105661
0 46672 5 1 1 46671
0 46673 7 1 2 102805 98168
0 46674 5 1 1 46673
0 46675 7 1 2 46672 46674
0 46676 5 1 1 46675
0 46677 7 1 2 83332 46676
0 46678 5 1 1 46677
0 46679 7 2 2 99451 92004
0 46680 7 1 2 104704 105673
0 46681 5 1 1 46680
0 46682 7 1 2 46678 46681
0 46683 5 1 1 46682
0 46684 7 1 2 80739 46683
0 46685 5 1 1 46684
0 46686 7 1 2 46669 46685
0 46687 7 1 2 46659 46686
0 46688 5 1 1 46687
0 46689 7 1 2 71468 46688
0 46690 5 1 1 46689
0 46691 7 1 2 46622 46690
0 46692 5 1 1 46691
0 46693 7 1 2 46692 105604
0 46694 5 1 1 46693
0 46695 7 1 2 81057 105674
0 46696 5 1 1 46695
0 46697 7 1 2 35588 46696
0 46698 5 1 1 46697
0 46699 7 1 2 73566 46698
0 46700 5 1 1 46699
0 46701 7 1 2 104102 105666
0 46702 5 1 1 46701
0 46703 7 1 2 46700 46702
0 46704 5 1 1 46703
0 46705 7 1 2 81769 46704
0 46706 5 1 1 46705
0 46707 7 2 2 100030 96651
0 46708 7 1 2 105667 105675
0 46709 5 1 1 46708
0 46710 7 1 2 46706 46709
0 46711 5 1 1 46710
0 46712 7 1 2 68711 46711
0 46713 5 1 1 46712
0 46714 7 2 2 80103 81184
0 46715 7 1 2 81770 105677
0 46716 5 3 1 46715
0 46717 7 1 2 79890 82661
0 46718 7 1 2 105679 46717
0 46719 5 1 1 46718
0 46720 7 1 2 99480 46719
0 46721 5 1 1 46720
0 46722 7 1 2 73567 102293
0 46723 7 1 2 102713 46722
0 46724 5 1 1 46723
0 46725 7 1 2 46721 46724
0 46726 5 1 1 46725
0 46727 7 1 2 77482 46726
0 46728 5 1 1 46727
0 46729 7 1 2 46713 46728
0 46730 5 1 1 46729
0 46731 7 1 2 71469 46730
0 46732 5 2 1 46731
0 46733 7 1 2 99481 83767
0 46734 5 1 1 46733
0 46735 7 1 2 72469 99667
0 46736 7 1 2 22891 46735
0 46737 5 1 1 46736
0 46738 7 1 2 46734 46737
0 46739 5 1 1 46738
0 46740 7 1 2 77483 46739
0 46741 5 1 1 46740
0 46742 7 1 2 99482 77187
0 46743 5 1 1 46742
0 46744 7 1 2 46741 46743
0 46745 5 2 1 46744
0 46746 7 1 2 81771 105684
0 46747 5 1 1 46746
0 46748 7 1 2 100501 98553
0 46749 5 1 1 46748
0 46750 7 1 2 46747 46749
0 46751 5 1 1 46750
0 46752 7 1 2 73568 46751
0 46753 5 1 1 46752
0 46754 7 1 2 105682 46753
0 46755 5 1 1 46754
0 46756 7 1 2 91359 9126
0 46757 5 1 1 46756
0 46758 7 1 2 72179 46757
0 46759 7 1 2 46755 46758
0 46760 5 1 1 46759
0 46761 7 1 2 46694 46760
0 46762 5 1 1 46761
0 46763 7 1 2 65656 46762
0 46764 5 1 1 46763
0 46765 7 1 2 85747 105685
0 46766 5 1 1 46765
0 46767 7 1 2 105683 46766
0 46768 5 1 1 46767
0 46769 7 1 2 96432 90295
0 46770 7 1 2 46768 46769
0 46771 5 1 1 46770
0 46772 7 1 2 46764 46771
0 46773 5 1 1 46772
0 46774 7 1 2 67772 46773
0 46775 5 1 1 46774
0 46776 7 1 2 16926 96287
0 46777 5 4 1 46776
0 46778 7 1 2 66366 105629
0 46779 5 1 1 46778
0 46780 7 1 2 65691 82463
0 46781 7 1 2 81111 96252
0 46782 7 1 2 46780 46781
0 46783 7 1 2 103588 46782
0 46784 5 1 1 46783
0 46785 7 1 2 46779 46784
0 46786 5 1 1 46785
0 46787 7 1 2 63916 46786
0 46788 5 1 1 46787
0 46789 7 1 2 97170 98158
0 46790 7 1 2 93426 46789
0 46791 7 1 2 104965 93654
0 46792 7 1 2 46790 46791
0 46793 5 1 1 46792
0 46794 7 1 2 46788 46793
0 46795 5 1 1 46794
0 46796 7 1 2 105686 46795
0 46797 5 1 1 46796
0 46798 7 1 2 69970 101768
0 46799 5 1 1 46798
0 46800 7 1 2 101352 46799
0 46801 5 1 1 46800
0 46802 7 1 2 81058 46801
0 46803 5 1 1 46802
0 46804 7 1 2 87518 105652
0 46805 5 1 1 46804
0 46806 7 1 2 46803 46805
0 46807 5 1 1 46806
0 46808 7 1 2 96483 46807
0 46809 5 1 1 46808
0 46810 7 2 2 81059 105605
0 46811 7 1 2 100374 105454
0 46812 7 1 2 105690 46811
0 46813 5 1 1 46812
0 46814 7 1 2 46809 46813
0 46815 5 1 1 46814
0 46816 7 1 2 68712 46815
0 46817 5 1 1 46816
0 46818 7 1 2 65657 105676
0 46819 7 1 2 105691 46818
0 46820 5 1 1 46819
0 46821 7 1 2 46817 46820
0 46822 5 1 1 46821
0 46823 7 1 2 74434 46822
0 46824 5 1 1 46823
0 46825 7 1 2 94718 96718
0 46826 5 1 1 46825
0 46827 7 1 2 98202 96582
0 46828 5 1 1 46827
0 46829 7 1 2 46826 46828
0 46830 5 1 1 46829
0 46831 7 1 2 88923 46830
0 46832 5 1 1 46831
0 46833 7 1 2 94719 105635
0 46834 5 1 1 46833
0 46835 7 1 2 46832 46834
0 46836 5 1 1 46835
0 46837 7 1 2 101831 46836
0 46838 5 1 1 46837
0 46839 7 1 2 90319 90975
0 46840 7 1 2 104573 46839
0 46841 5 1 1 46840
0 46842 7 1 2 46838 46841
0 46843 5 1 1 46842
0 46844 7 1 2 65495 46843
0 46845 5 1 1 46844
0 46846 7 1 2 94804 91535
0 46847 7 1 2 105563 46846
0 46848 5 1 1 46847
0 46849 7 1 2 46845 46848
0 46850 5 1 1 46849
0 46851 7 1 2 63917 46850
0 46852 5 1 1 46851
0 46853 7 1 2 82125 91536
0 46854 7 2 2 69006 84357
0 46855 7 1 2 87593 105692
0 46856 7 1 2 46853 46855
0 46857 5 1 1 46856
0 46858 7 1 2 46852 46857
0 46859 5 1 1 46858
0 46860 7 1 2 74176 46859
0 46861 5 1 1 46860
0 46862 7 1 2 46824 46861
0 46863 5 1 1 46862
0 46864 7 1 2 103289 46863
0 46865 5 1 1 46864
0 46866 7 1 2 46797 46865
0 46867 7 1 2 46775 46866
0 46868 7 1 2 46607 46867
0 46869 5 1 1 46868
0 46870 7 1 2 73234 46869
0 46871 5 1 1 46870
0 46872 7 1 2 99734 79886
0 46873 5 1 1 46872
0 46874 7 1 2 71699 100829
0 46875 7 2 2 104117 46874
0 46876 5 1 1 105694
0 46877 7 1 2 46873 46876
0 46878 5 1 1 46877
0 46879 7 1 2 82464 46878
0 46880 5 1 1 46879
0 46881 7 1 2 102878 84727
0 46882 5 1 1 46881
0 46883 7 1 2 71169 105695
0 46884 5 1 1 46883
0 46885 7 1 2 71866 81991
0 46886 7 1 2 74157 46885
0 46887 7 3 2 69971 80301
0 46888 7 1 2 103425 105696
0 46889 7 1 2 46886 46888
0 46890 5 1 1 46889
0 46891 7 1 2 46884 46890
0 46892 5 1 1 46891
0 46893 7 1 2 69612 46892
0 46894 5 1 1 46893
0 46895 7 1 2 46882 46894
0 46896 5 1 1 46895
0 46897 7 1 2 74435 46896
0 46898 5 1 1 46897
0 46899 7 1 2 46880 46898
0 46900 5 1 1 46899
0 46901 7 1 2 67773 46900
0 46902 5 1 1 46901
0 46903 7 1 2 101058 105600
0 46904 5 1 1 46903
0 46905 7 1 2 46902 46904
0 46906 5 1 1 46905
0 46907 7 1 2 72470 46906
0 46908 5 1 1 46907
0 46909 7 1 2 100005 92775
0 46910 5 1 1 46909
0 46911 7 1 2 80128 89443
0 46912 5 1 1 46911
0 46913 7 1 2 46910 46912
0 46914 5 2 1 46913
0 46915 7 1 2 64490 105699
0 46916 5 1 1 46915
0 46917 7 1 2 99811 104401
0 46918 5 1 1 46917
0 46919 7 1 2 46916 46918
0 46920 5 1 1 46919
0 46921 7 1 2 74436 46920
0 46922 5 1 1 46921
0 46923 7 1 2 92849 80843
0 46924 5 1 1 46923
0 46925 7 1 2 46922 46924
0 46926 5 1 1 46925
0 46927 7 1 2 35656 82091
0 46928 5 1 1 46927
0 46929 7 1 2 1352 46928
0 46930 7 1 2 46926 46929
0 46931 5 1 1 46930
0 46932 7 1 2 69613 105700
0 46933 5 1 1 46932
0 46934 7 1 2 42263 46933
0 46935 5 1 1 46934
0 46936 7 1 2 92531 93124
0 46937 5 1 1 46936
0 46938 7 1 2 84207 82553
0 46939 5 1 1 46938
0 46940 7 1 2 46937 46939
0 46941 5 1 1 46940
0 46942 7 1 2 46935 46941
0 46943 5 1 1 46942
0 46944 7 1 2 79478 105575
0 46945 5 1 1 46944
0 46946 7 1 2 99971 102072
0 46947 5 1 1 46946
0 46948 7 1 2 46945 46947
0 46949 5 1 1 46948
0 46950 7 1 2 69257 46949
0 46951 5 1 1 46950
0 46952 7 1 2 73928 85085
0 46953 7 1 2 98713 46952
0 46954 5 1 1 46953
0 46955 7 1 2 46951 46954
0 46956 5 1 1 46955
0 46957 7 1 2 104980 46956
0 46958 5 1 1 46957
0 46959 7 1 2 46943 46958
0 46960 7 1 2 46931 46959
0 46961 5 1 1 46960
0 46962 7 1 2 67406 46961
0 46963 5 1 1 46962
0 46964 7 1 2 67774 105668
0 46965 5 1 1 46964
0 46966 7 1 2 98644 98542
0 46967 5 1 1 46966
0 46968 7 1 2 46965 46967
0 46969 5 1 1 46968
0 46970 7 1 2 42588 105149
0 46971 5 1 1 46970
0 46972 7 1 2 101252 46971
0 46973 7 1 2 46969 46972
0 46974 5 1 1 46973
0 46975 7 1 2 46963 46974
0 46976 7 1 2 46908 46975
0 46977 5 1 1 46976
0 46978 7 1 2 68713 46977
0 46979 5 1 1 46978
0 46980 7 1 2 100123 103234
0 46981 5 1 1 46980
0 46982 7 1 2 100502 86128
0 46983 5 1 1 46982
0 46984 7 1 2 46981 46983
0 46985 5 1 1 46984
0 46986 7 1 2 72758 46985
0 46987 5 1 1 46986
0 46988 7 1 2 76608 82328
0 46989 5 1 1 46988
0 46990 7 1 2 8251 46989
0 46991 5 1 1 46990
0 46992 7 1 2 84218 87289
0 46993 5 1 1 46992
0 46994 7 1 2 46991 46993
0 46995 5 1 1 46994
0 46996 7 2 2 67775 46995
0 46997 7 1 2 78141 105701
0 46998 5 1 1 46997
0 46999 7 1 2 46987 46998
0 47000 5 1 1 46999
0 47001 7 1 2 67407 47000
0 47002 5 1 1 47001
0 47003 7 1 2 94260 104195
0 47004 5 1 1 47003
0 47005 7 1 2 101059 47004
0 47006 5 1 1 47005
0 47007 7 1 2 85544 105702
0 47008 5 1 1 47007
0 47009 7 1 2 47006 47008
0 47010 5 1 1 47009
0 47011 7 1 2 98289 47010
0 47012 5 1 1 47011
0 47013 7 1 2 47002 47012
0 47014 7 1 2 46979 47013
0 47015 5 2 1 47014
0 47016 7 2 2 72180 73868
0 47017 7 1 2 105703 105705
0 47018 5 1 1 47017
0 47019 7 1 2 67408 93533
0 47020 5 1 1 47019
0 47021 7 1 2 103672 47020
0 47022 5 3 1 47021
0 47023 7 1 2 70877 105707
0 47024 5 2 1 47023
0 47025 7 2 2 82506 98769
0 47026 7 1 2 77188 105712
0 47027 5 1 1 47026
0 47028 7 1 2 105710 47027
0 47029 5 1 1 47028
0 47030 7 1 2 101305 47029
0 47031 5 1 1 47030
0 47032 7 1 2 99158 105416
0 47033 7 1 2 92890 47032
0 47034 5 1 1 47033
0 47035 7 1 2 47031 47034
0 47036 5 1 1 47035
0 47037 7 1 2 93806 47036
0 47038 5 1 1 47037
0 47039 7 1 2 76502 89024
0 47040 7 1 2 105669 47039
0 47041 5 1 1 47040
0 47042 7 1 2 88385 101279
0 47043 5 1 1 47042
0 47044 7 2 2 99929 101474
0 47045 5 1 1 105714
0 47046 7 1 2 47043 47045
0 47047 5 1 1 47046
0 47048 7 1 2 98645 81060
0 47049 7 1 2 47047 47048
0 47050 5 1 1 47049
0 47051 7 1 2 47041 47050
0 47052 5 1 1 47051
0 47053 7 1 2 70257 47052
0 47054 5 1 1 47053
0 47055 7 1 2 103603 47054
0 47056 5 1 1 47055
0 47057 7 1 2 72759 47056
0 47058 5 1 1 47057
0 47059 7 1 2 105670 105715
0 47060 5 1 1 47059
0 47061 7 1 2 96952 98230
0 47062 5 1 1 47061
0 47063 7 1 2 65846 102327
0 47064 5 1 1 47063
0 47065 7 1 2 76238 47064
0 47066 7 1 2 47062 47065
0 47067 5 1 1 47066
0 47068 7 1 2 76337 81011
0 47069 5 1 1 47068
0 47070 7 2 2 80275 47069
0 47071 7 1 2 99456 18649
0 47072 7 1 2 105716 47071
0 47073 5 1 1 47072
0 47074 7 1 2 47067 47073
0 47075 5 1 1 47074
0 47076 7 1 2 89025 47075
0 47077 5 1 1 47076
0 47078 7 1 2 47060 47077
0 47079 5 1 1 47078
0 47080 7 1 2 70258 47079
0 47081 5 1 1 47080
0 47082 7 1 2 101483 104549
0 47083 5 1 1 47082
0 47084 7 1 2 47081 47083
0 47085 5 1 1 47084
0 47086 7 1 2 67776 47085
0 47087 5 1 1 47086
0 47088 7 1 2 47058 47087
0 47089 7 1 2 47038 47088
0 47090 5 1 1 47089
0 47091 7 1 2 96827 47090
0 47092 5 1 1 47091
0 47093 7 1 2 47018 47092
0 47094 5 1 1 47093
0 47095 7 1 2 68150 47094
0 47096 5 1 1 47095
0 47097 7 2 2 85754 96433
0 47098 5 1 1 105718
0 47099 7 1 2 96288 47098
0 47100 5 1 1 47099
0 47101 7 1 2 81969 47100
0 47102 5 1 1 47101
0 47103 7 1 2 83941 105687
0 47104 5 1 1 47103
0 47105 7 1 2 47102 47104
0 47106 5 1 1 47105
0 47107 7 1 2 98278 47106
0 47108 5 1 1 47107
0 47109 7 1 2 70259 95125
0 47110 5 1 1 47109
0 47111 7 2 2 77944 47110
0 47112 5 1 1 105720
0 47113 7 1 2 86072 89489
0 47114 5 1 1 47113
0 47115 7 1 2 105721 47114
0 47116 5 1 1 47115
0 47117 7 1 2 96434 47116
0 47118 5 1 1 47117
0 47119 7 1 2 86275 86073
0 47120 5 1 1 47119
0 47121 7 1 2 89487 47120
0 47122 5 1 1 47121
0 47123 7 1 2 96279 47122
0 47124 5 1 1 47123
0 47125 7 1 2 47118 47124
0 47126 5 1 1 47125
0 47127 7 1 2 72760 47126
0 47128 5 1 1 47127
0 47129 7 3 2 101289 77965
0 47130 5 2 1 105722
0 47131 7 1 2 96435 105723
0 47132 5 2 1 47131
0 47133 7 1 2 47128 105727
0 47134 5 1 1 47133
0 47135 7 1 2 98290 47134
0 47136 5 1 1 47135
0 47137 7 1 2 47108 47136
0 47138 5 1 1 47137
0 47139 7 1 2 70878 47138
0 47140 5 1 1 47139
0 47141 7 1 2 96785 104269
0 47142 5 3 1 47141
0 47143 7 1 2 85641 96280
0 47144 5 1 1 47143
0 47145 7 1 2 32059 105719
0 47146 5 1 1 47145
0 47147 7 1 2 47144 47146
0 47148 5 1 1 47147
0 47149 7 1 2 71700 47148
0 47150 5 1 1 47149
0 47151 7 1 2 82310 96907
0 47152 5 1 1 47151
0 47153 7 1 2 47150 47152
0 47154 5 1 1 47153
0 47155 7 1 2 105729 47154
0 47156 5 1 1 47155
0 47157 7 1 2 93752 105656
0 47158 5 1 1 47157
0 47159 7 1 2 76338 105688
0 47160 7 1 2 47158 47159
0 47161 5 1 1 47160
0 47162 7 1 2 76503 96436
0 47163 5 1 1 47162
0 47164 7 1 2 83682 96281
0 47165 5 1 1 47164
0 47166 7 1 2 47163 47165
0 47167 7 1 2 47161 47166
0 47168 5 1 1 47167
0 47169 7 1 2 72761 47168
0 47170 5 1 1 47169
0 47171 7 1 2 105728 47170
0 47172 5 1 1 47171
0 47173 7 1 2 67409 47172
0 47174 5 1 1 47173
0 47175 7 1 2 47156 47174
0 47176 5 1 1 47175
0 47177 7 1 2 98526 47176
0 47178 5 1 1 47177
0 47179 7 1 2 47140 47178
0 47180 5 1 1 47179
0 47181 7 1 2 88924 47180
0 47182 5 1 1 47181
0 47183 7 1 2 72762 47112
0 47184 5 1 1 47183
0 47185 7 1 2 105725 47184
0 47186 5 2 1 47185
0 47187 7 1 2 98511 105732
0 47188 5 1 1 47187
0 47189 7 1 2 65847 105730
0 47190 5 1 1 47189
0 47191 7 2 2 72471 84000
0 47192 7 1 2 70879 105734
0 47193 5 1 1 47192
0 47194 7 1 2 47190 47193
0 47195 5 2 1 47194
0 47196 7 1 2 81917 105736
0 47197 5 1 1 47196
0 47198 7 1 2 34041 47197
0 47199 5 1 1 47198
0 47200 7 1 2 80945 47199
0 47201 5 1 1 47200
0 47202 7 1 2 81918 98386
0 47203 5 1 1 47202
0 47204 7 1 2 30334 47203
0 47205 5 1 1 47204
0 47206 7 1 2 89235 47205
0 47207 5 1 1 47206
0 47208 7 2 2 84208 98482
0 47209 7 1 2 81142 105738
0 47210 5 1 1 47209
0 47211 7 1 2 47207 47210
0 47212 7 1 2 47201 47211
0 47213 7 1 2 47188 47212
0 47214 5 1 1 47213
0 47215 7 1 2 77189 47214
0 47216 5 1 1 47215
0 47217 7 1 2 72763 85802
0 47218 5 1 1 47217
0 47219 7 1 2 103594 82072
0 47220 7 2 2 47218 47219
0 47221 5 1 1 105740
0 47222 7 1 2 47216 47221
0 47223 5 1 1 47222
0 47224 7 1 2 72181 73832
0 47225 7 1 2 47223 47224
0 47226 5 1 1 47225
0 47227 7 1 2 47182 47226
0 47228 5 1 1 47227
0 47229 7 1 2 69258 47228
0 47230 5 1 1 47229
0 47231 7 1 2 98512 78395
0 47232 5 1 1 47231
0 47233 7 1 2 25728 47232
0 47234 5 2 1 47233
0 47235 7 1 2 95774 105742
0 47236 5 1 1 47235
0 47237 7 1 2 66367 95787
0 47238 5 2 1 47237
0 47239 7 1 2 96084 105744
0 47240 5 1 1 47239
0 47241 7 1 2 64866 47240
0 47242 5 1 1 47241
0 47243 7 1 2 102789 96883
0 47244 5 1 1 47243
0 47245 7 1 2 96089 47244
0 47246 5 1 1 47245
0 47247 7 1 2 67410 47246
0 47248 7 1 2 47242 47247
0 47249 5 1 1 47248
0 47250 7 1 2 47236 47249
0 47251 5 1 1 47250
0 47252 7 1 2 96828 47251
0 47253 5 1 1 47252
0 47254 7 1 2 73929 101156
0 47255 5 1 1 47254
0 47256 7 1 2 96786 47255
0 47257 5 1 1 47256
0 47258 7 1 2 70880 47257
0 47259 5 1 1 47258
0 47260 7 1 2 84209 105271
0 47261 5 1 1 47260
0 47262 7 1 2 47259 47261
0 47263 5 1 1 47262
0 47264 7 1 2 69972 47263
0 47265 5 1 1 47264
0 47266 7 1 2 77632 101095
0 47267 5 1 1 47266
0 47268 7 1 2 47265 47267
0 47269 5 1 1 47268
0 47270 7 1 2 87290 47269
0 47271 5 1 1 47270
0 47272 7 1 2 87780 105726
0 47273 5 2 1 47272
0 47274 7 1 2 99452 105746
0 47275 5 1 1 47274
0 47276 7 1 2 82311 105743
0 47277 5 1 1 47276
0 47278 7 1 2 99453 89236
0 47279 5 1 1 47278
0 47280 7 1 2 47277 47279
0 47281 5 1 1 47280
0 47282 7 1 2 78709 47281
0 47283 5 1 1 47282
0 47284 7 1 2 47275 47283
0 47285 7 1 2 47271 47284
0 47286 5 1 1 47285
0 47287 7 1 2 105706 47286
0 47288 5 1 1 47287
0 47289 7 1 2 47253 47288
0 47290 5 1 1 47289
0 47291 7 1 2 101007 47290
0 47292 5 1 1 47291
0 47293 7 1 2 47230 47292
0 47294 7 1 2 47096 47293
0 47295 5 1 1 47294
0 47296 7 1 2 63918 47295
0 47297 5 1 1 47296
0 47298 7 1 2 75033 87775
0 47299 5 1 1 47298
0 47300 7 2 2 73569 79510
0 47301 7 1 2 81671 105748
0 47302 5 1 1 47301
0 47303 7 1 2 104009 47302
0 47304 5 1 1 47303
0 47305 7 1 2 81772 47304
0 47306 5 1 1 47305
0 47307 7 1 2 66368 82660
0 47308 5 1 1 47307
0 47309 7 1 2 67777 47308
0 47310 7 1 2 47306 47309
0 47311 5 1 1 47310
0 47312 7 1 2 72764 103002
0 47313 5 1 1 47312
0 47314 7 1 2 68151 47313
0 47315 7 1 2 47311 47314
0 47316 5 1 1 47315
0 47317 7 1 2 47299 47316
0 47318 5 1 1 47317
0 47319 7 1 2 99483 47318
0 47320 5 1 1 47319
0 47321 7 1 2 69259 98387
0 47322 5 1 1 47321
0 47323 7 1 2 99469 47322
0 47324 5 3 1 47323
0 47325 7 1 2 81919 105750
0 47326 5 1 1 47325
0 47327 7 3 2 80645 99756
0 47328 5 1 1 105753
0 47329 7 1 2 47326 47328
0 47330 5 1 1 47329
0 47331 7 3 2 90047 90161
0 47332 7 1 2 72765 105756
0 47333 7 1 2 47330 47332
0 47334 5 1 1 47333
0 47335 7 1 2 98034 104832
0 47336 7 1 2 105724 47335
0 47337 5 1 1 47336
0 47338 7 1 2 47334 47337
0 47339 7 1 2 47320 47338
0 47340 5 1 1 47339
0 47341 7 1 2 96484 47340
0 47342 5 1 1 47341
0 47343 7 1 2 79948 94286
0 47344 5 1 1 47343
0 47345 7 1 2 80167 47344
0 47346 5 1 1 47345
0 47347 7 1 2 72766 47346
0 47348 5 1 1 47347
0 47349 7 1 2 82154 47348
0 47350 5 1 1 47349
0 47351 7 1 2 99484 105646
0 47352 7 1 2 47350 47351
0 47353 5 1 1 47352
0 47354 7 1 2 89281 77622
0 47355 5 1 1 47354
0 47356 7 1 2 86074 47355
0 47357 5 1 1 47356
0 47358 7 1 2 104234 47357
0 47359 5 1 1 47358
0 47360 7 1 2 70260 47359
0 47361 5 1 1 47360
0 47362 7 1 2 87466 82210
0 47363 5 1 1 47362
0 47364 7 1 2 47361 47363
0 47365 5 1 1 47364
0 47366 7 2 2 102485 99060
0 47367 7 1 2 90290 99195
0 47368 7 1 2 105759 47367
0 47369 7 1 2 47365 47368
0 47370 5 1 1 47369
0 47371 7 1 2 47353 47370
0 47372 7 1 2 47342 47371
0 47373 5 1 1 47372
0 47374 7 1 2 77484 47373
0 47375 5 1 1 47374
0 47376 7 1 2 68152 105704
0 47377 5 1 1 47376
0 47378 7 1 2 69260 105741
0 47379 5 1 1 47378
0 47380 7 1 2 69261 105737
0 47381 5 1 1 47380
0 47382 7 1 2 35165 47381
0 47383 5 1 1 47382
0 47384 7 1 2 81920 47383
0 47385 5 1 1 47384
0 47386 7 1 2 72767 105754
0 47387 5 1 1 47386
0 47388 7 1 2 47385 47387
0 47389 5 1 1 47388
0 47390 7 1 2 70261 47389
0 47391 5 1 1 47390
0 47392 7 1 2 85461 99312
0 47393 5 1 1 47392
0 47394 7 1 2 47391 47393
0 47395 5 1 1 47394
0 47396 7 1 2 78710 47395
0 47397 5 1 1 47396
0 47398 7 1 2 69262 105733
0 47399 5 1 1 47398
0 47400 7 1 2 82335 89062
0 47401 5 1 1 47400
0 47402 7 1 2 104371 47401
0 47403 5 1 1 47402
0 47404 7 1 2 47399 47403
0 47405 5 1 1 47404
0 47406 7 1 2 98513 47405
0 47407 5 1 1 47406
0 47408 7 1 2 96963 105747
0 47409 5 1 1 47408
0 47410 7 1 2 96921 95126
0 47411 7 1 2 105072 47410
0 47412 5 1 1 47411
0 47413 7 1 2 47409 47412
0 47414 5 1 1 47413
0 47415 7 1 2 70881 47414
0 47416 5 1 1 47415
0 47417 7 1 2 95127 103853
0 47418 5 1 1 47417
0 47419 7 1 2 100166 105739
0 47420 5 1 1 47419
0 47421 7 1 2 47418 47420
0 47422 5 1 1 47421
0 47423 7 1 2 82286 47422
0 47424 5 1 1 47423
0 47425 7 1 2 99592 105068
0 47426 7 1 2 95128 47425
0 47427 5 1 1 47426
0 47428 7 1 2 47424 47427
0 47429 7 1 2 47416 47428
0 47430 7 1 2 47407 47429
0 47431 7 1 2 47397 47430
0 47432 5 1 1 47431
0 47433 7 1 2 77190 47432
0 47434 5 1 1 47433
0 47435 7 1 2 47379 47434
0 47436 7 1 2 47377 47435
0 47437 5 1 1 47436
0 47438 7 1 2 105638 47437
0 47439 5 1 1 47438
0 47440 7 1 2 47375 47439
0 47441 7 1 2 47297 47440
0 47442 7 1 2 46871 47441
0 47443 5 1 1 47442
0 47444 7 1 2 65607 47443
0 47445 5 1 1 47444
0 47446 7 1 2 67133 98000
0 47447 7 1 2 105382 47446
0 47448 5 1 1 47447
0 47449 7 1 2 81921 99079
0 47450 7 1 2 84620 47449
0 47451 7 1 2 97855 47450
0 47452 5 1 1 47451
0 47453 7 1 2 47448 47452
0 47454 5 1 1 47453
0 47455 7 1 2 64196 47454
0 47456 5 1 1 47455
0 47457 7 1 2 99422 97139
0 47458 5 1 1 47457
0 47459 7 1 2 81922 101091
0 47460 5 1 1 47459
0 47461 7 1 2 47458 47460
0 47462 5 1 1 47461
0 47463 7 1 2 77485 47462
0 47464 5 1 1 47463
0 47465 7 1 2 77995 103865
0 47466 5 1 1 47465
0 47467 7 1 2 47464 47466
0 47468 5 1 1 47467
0 47469 7 1 2 102794 47468
0 47470 5 1 1 47469
0 47471 7 1 2 47456 47470
0 47472 5 1 1 47471
0 47473 7 1 2 66593 47472
0 47474 5 1 1 47473
0 47475 7 1 2 100503 102519
0 47476 5 1 1 47475
0 47477 7 1 2 99473 30122
0 47478 5 1 1 47477
0 47479 7 1 2 82582 86453
0 47480 7 1 2 47478 47479
0 47481 5 1 1 47480
0 47482 7 1 2 47476 47481
0 47483 5 1 1 47482
0 47484 7 1 2 84621 47483
0 47485 5 1 1 47484
0 47486 7 1 2 47474 47485
0 47487 5 1 1 47486
0 47488 7 1 2 65189 47487
0 47489 5 1 1 47488
0 47490 7 2 2 86446 82583
0 47491 7 1 2 98554 105761
0 47492 5 1 1 47491
0 47493 7 1 2 82507 47492
0 47494 5 1 1 47493
0 47495 7 1 2 98159 105762
0 47496 5 1 1 47495
0 47497 7 1 2 98279 104495
0 47498 5 1 1 47497
0 47499 7 1 2 82465 47498
0 47500 7 1 2 47496 47499
0 47501 5 1 1 47500
0 47502 7 1 2 74437 84622
0 47503 7 1 2 47501 47502
0 47504 7 1 2 47494 47503
0 47505 5 1 1 47504
0 47506 7 1 2 47489 47505
0 47507 5 1 1 47506
0 47508 7 1 2 63919 47507
0 47509 5 1 1 47508
0 47510 7 1 2 102005 103632
0 47511 7 1 2 103646 75520
0 47512 7 1 2 47510 47511
0 47513 5 1 1 47512
0 47514 7 1 2 47509 47513
0 47515 5 1 1 47514
0 47516 7 1 2 73869 47515
0 47517 5 1 1 47516
0 47518 7 4 2 98841 84325
0 47519 7 1 2 77383 105763
0 47520 7 1 2 98121 47519
0 47521 5 1 1 47520
0 47522 7 2 2 68153 104000
0 47523 5 1 1 105767
0 47524 7 1 2 38629 47523
0 47525 5 1 1 47524
0 47526 7 1 2 73984 95355
0 47527 7 1 2 47525 47526
0 47528 5 1 1 47527
0 47529 7 1 2 47521 47528
0 47530 5 1 1 47529
0 47531 7 1 2 80740 47530
0 47532 5 1 1 47531
0 47533 7 1 2 78665 95356
0 47534 7 1 2 105768 47533
0 47535 5 1 1 47534
0 47536 7 1 2 47532 47535
0 47537 5 1 1 47536
0 47538 7 1 2 67134 47537
0 47539 5 1 1 47538
0 47540 7 1 2 92825 102446
0 47541 7 1 2 101904 47540
0 47542 7 1 2 96020 47541
0 47543 5 1 1 47542
0 47544 7 1 2 81923 87705
0 47545 5 3 1 47544
0 47546 7 1 2 103223 105769
0 47547 5 1 1 47546
0 47548 7 1 2 99485 84299
0 47549 7 1 2 47547 47548
0 47550 5 1 1 47549
0 47551 7 1 2 47543 47550
0 47552 5 1 1 47551
0 47553 7 1 2 77486 47552
0 47554 5 1 1 47553
0 47555 7 1 2 82329 103866
0 47556 7 1 2 78002 47555
0 47557 7 1 2 89063 47556
0 47558 5 1 1 47557
0 47559 7 1 2 47554 47558
0 47560 5 1 1 47559
0 47561 7 1 2 88591 47560
0 47562 5 1 1 47561
0 47563 7 1 2 47539 47562
0 47564 5 1 1 47563
0 47565 7 1 2 91537 47564
0 47566 5 1 1 47565
0 47567 7 2 2 72768 98627
0 47568 7 2 2 77677 105772
0 47569 7 1 2 92465 84966
0 47570 7 2 2 105774 47569
0 47571 7 3 2 75512 91174
0 47572 7 2 2 84530 91558
0 47573 7 1 2 105778 105781
0 47574 7 1 2 105776 47573
0 47575 5 1 1 47574
0 47576 7 1 2 47566 47575
0 47577 7 1 2 47517 47576
0 47578 5 1 1 47577
0 47579 7 1 2 65608 47578
0 47580 5 1 1 47579
0 47581 7 1 2 94999 84232
0 47582 7 1 2 105157 47581
0 47583 7 1 2 105777 47582
0 47584 5 1 1 47583
0 47585 7 1 2 47580 47584
0 47586 5 1 1 47585
0 47587 7 1 2 76609 47586
0 47588 5 1 1 47587
0 47589 7 1 2 103841 85423
0 47590 5 1 1 47589
0 47591 7 1 2 93114 98770
0 47592 5 1 1 47591
0 47593 7 1 2 47590 47592
0 47594 5 1 1 47593
0 47595 7 1 2 73870 47594
0 47596 5 1 1 47595
0 47597 7 1 2 98771 90425
0 47598 7 1 2 105760 47597
0 47599 5 1 1 47598
0 47600 7 2 2 70689 93326
0 47601 7 1 2 85419 91559
0 47602 7 1 2 103868 47601
0 47603 7 1 2 105783 47602
0 47604 5 1 1 47603
0 47605 7 1 2 47599 47604
0 47606 7 1 2 47596 47605
0 47607 5 1 1 47606
0 47608 7 1 2 77384 47607
0 47609 5 1 1 47608
0 47610 7 2 2 97856 99162
0 47611 7 1 2 84358 105785
0 47612 7 1 2 96372 47611
0 47613 5 1 1 47612
0 47614 7 1 2 47609 47613
0 47615 5 1 1 47614
0 47616 7 1 2 65609 47615
0 47617 5 1 1 47616
0 47618 7 3 2 84233 96253
0 47619 7 2 2 98462 105787
0 47620 7 2 2 96315 92440
0 47621 7 1 2 99310 105792
0 47622 7 1 2 105790 47621
0 47623 5 1 1 47622
0 47624 7 1 2 47617 47623
0 47625 5 1 1 47624
0 47626 7 1 2 82330 47625
0 47627 5 1 1 47626
0 47628 7 1 2 67778 79528
0 47629 7 1 2 82258 47628
0 47630 7 1 2 99486 47629
0 47631 7 1 2 105654 47630
0 47632 5 1 1 47631
0 47633 7 1 2 47627 47632
0 47634 5 1 1 47633
0 47635 7 1 2 72182 47634
0 47636 5 1 1 47635
0 47637 7 1 2 99267 95530
0 47638 7 1 2 96418 47637
0 47639 5 1 1 47638
0 47640 7 1 2 70882 99299
0 47641 7 1 2 93662 47640
0 47642 7 1 2 91538 47641
0 47643 5 1 1 47642
0 47644 7 1 2 47639 47643
0 47645 5 1 1 47644
0 47646 7 1 2 63920 47645
0 47647 5 1 1 47646
0 47648 7 2 2 69007 96254
0 47649 7 1 2 65692 93265
0 47650 7 2 2 105794 47649
0 47651 7 1 2 100880 103869
0 47652 7 1 2 105796 47651
0 47653 5 1 1 47652
0 47654 7 1 2 47647 47653
0 47655 5 1 1 47654
0 47656 7 1 2 80741 47655
0 47657 5 1 1 47656
0 47658 7 1 2 72769 97968
0 47659 7 1 2 101426 47658
0 47660 7 1 2 96373 47659
0 47661 5 1 1 47660
0 47662 7 1 2 47657 47661
0 47663 5 1 1 47662
0 47664 7 1 2 64197 47663
0 47665 5 1 1 47664
0 47666 7 1 2 103177 40088
0 47667 5 1 1 47666
0 47668 7 1 2 77487 47667
0 47669 5 1 1 47668
0 47670 7 1 2 77996 78440
0 47671 5 2 1 47670
0 47672 7 1 2 47669 105798
0 47673 5 1 1 47672
0 47674 7 3 2 65693 67411
0 47675 5 1 1 105800
0 47676 7 1 2 102486 105801
0 47677 7 1 2 105504 47676
0 47678 7 1 2 47673 47677
0 47679 5 1 1 47678
0 47680 7 1 2 47665 47679
0 47681 5 1 1 47680
0 47682 7 1 2 76010 47681
0 47683 5 1 1 47682
0 47684 7 1 2 47636 47683
0 47685 5 1 1 47684
0 47686 7 1 2 73985 47685
0 47687 5 1 1 47686
0 47688 7 1 2 104034 94139
0 47689 7 1 2 105788 47688
0 47690 7 1 2 99335 47689
0 47691 5 1 1 47690
0 47692 7 1 2 47687 47691
0 47693 5 1 1 47692
0 47694 7 1 2 73235 47693
0 47695 5 1 1 47694
0 47696 7 2 2 80742 104785
0 47697 7 1 2 102240 105803
0 47698 5 1 1 47697
0 47699 7 1 2 76504 87291
0 47700 5 2 1 47699
0 47701 7 2 2 67779 102321
0 47702 7 1 2 96301 105807
0 47703 7 1 2 105805 47702
0 47704 5 1 1 47703
0 47705 7 1 2 47698 47704
0 47706 5 1 1 47705
0 47707 7 1 2 77385 47706
0 47708 5 1 1 47707
0 47709 7 1 2 93127 105657
0 47710 7 1 2 105786 47709
0 47711 5 1 1 47710
0 47712 7 1 2 47708 47711
0 47713 5 1 1 47712
0 47714 7 1 2 63921 47713
0 47715 5 1 1 47714
0 47716 7 2 2 99033 91488
0 47717 7 1 2 93427 105809
0 47718 7 1 2 105309 47717
0 47719 5 1 1 47718
0 47720 7 1 2 47715 47719
0 47721 5 1 1 47720
0 47722 7 1 2 73871 47721
0 47723 5 1 1 47722
0 47724 7 1 2 88592 105806
0 47725 5 1 1 47724
0 47726 7 1 2 96113 47725
0 47727 5 1 1 47726
0 47728 7 1 2 95215 47727
0 47729 5 1 1 47728
0 47730 7 1 2 100727 92970
0 47731 7 1 2 89771 47730
0 47732 5 1 1 47731
0 47733 7 1 2 47729 47732
0 47734 5 1 1 47733
0 47735 7 1 2 105292 47734
0 47736 5 1 1 47735
0 47737 7 1 2 104329 105764
0 47738 7 1 2 105804 47737
0 47739 5 1 1 47738
0 47740 7 1 2 47736 47739
0 47741 5 1 1 47740
0 47742 7 1 2 91539 47741
0 47743 5 1 1 47742
0 47744 7 1 2 91777 93327
0 47745 7 1 2 94144 47744
0 47746 7 1 2 105782 105810
0 47747 7 1 2 47745 47746
0 47748 5 1 1 47747
0 47749 7 1 2 47743 47748
0 47750 7 1 2 47723 47749
0 47751 5 1 1 47750
0 47752 7 1 2 65610 47751
0 47753 5 1 1 47752
0 47754 7 1 2 65190 91286
0 47755 7 1 2 103842 47754
0 47756 7 3 2 66782 89548
0 47757 7 1 2 94108 105789
0 47758 7 1 2 105811 47757
0 47759 7 1 2 47755 47758
0 47760 5 1 1 47759
0 47761 7 1 2 47753 47760
0 47762 7 1 2 47695 47761
0 47763 5 1 1 47762
0 47764 7 1 2 87039 47763
0 47765 5 1 1 47764
0 47766 7 1 2 47588 47765
0 47767 7 1 2 47445 47766
0 47768 5 1 1 47767
0 47769 7 1 2 66894 47768
0 47770 5 1 1 47769
0 47771 7 1 2 75446 94752
0 47772 5 1 1 47771
0 47773 7 1 2 88843 86623
0 47774 7 1 2 47772 47773
0 47775 5 1 1 47774
0 47776 7 1 2 73236 47775
0 47777 5 1 1 47776
0 47778 7 1 2 77126 75937
0 47779 5 1 1 47778
0 47780 7 1 2 83048 104649
0 47781 7 1 2 47779 47780
0 47782 5 1 1 47781
0 47783 7 1 2 47777 47782
0 47784 5 1 1 47783
0 47785 7 1 2 71170 47784
0 47786 5 1 1 47785
0 47787 7 1 2 103444 84395
0 47788 5 1 1 47787
0 47789 7 1 2 47786 47788
0 47790 5 1 1 47789
0 47791 7 1 2 69973 47790
0 47792 5 1 1 47791
0 47793 7 2 2 81773 75987
0 47794 7 1 2 73570 105814
0 47795 5 4 1 47794
0 47796 7 1 2 96678 105816
0 47797 5 1 1 47796
0 47798 7 1 2 74565 100764
0 47799 7 1 2 47797 47798
0 47800 5 1 1 47799
0 47801 7 1 2 47792 47800
0 47802 5 1 1 47801
0 47803 7 1 2 72770 47802
0 47804 5 1 1 47803
0 47805 7 1 2 86635 105817
0 47806 5 3 1 47805
0 47807 7 1 2 75447 105820
0 47808 5 1 1 47807
0 47809 7 1 2 85755 82082
0 47810 5 1 1 47809
0 47811 7 1 2 47808 47810
0 47812 5 1 1 47811
0 47813 7 1 2 69974 47812
0 47814 5 1 1 47813
0 47815 7 1 2 92713 87005
0 47816 5 1 1 47815
0 47817 7 1 2 47814 47816
0 47818 5 1 1 47817
0 47819 7 1 2 78441 47818
0 47820 5 1 1 47819
0 47821 7 1 2 100010 97535
0 47822 5 2 1 47821
0 47823 7 1 2 69975 105823
0 47824 5 1 1 47823
0 47825 7 1 2 71171 99562
0 47826 5 1 1 47825
0 47827 7 1 2 47824 47826
0 47828 5 1 1 47827
0 47829 7 1 2 73571 47828
0 47830 5 1 1 47829
0 47831 7 1 2 69976 77089
0 47832 5 2 1 47831
0 47833 7 1 2 66074 105825
0 47834 5 1 1 47833
0 47835 7 1 2 88870 47834
0 47836 5 1 1 47835
0 47837 7 1 2 71172 89203
0 47838 5 1 1 47837
0 47839 7 1 2 47836 47838
0 47840 5 1 1 47839
0 47841 7 1 2 65191 47840
0 47842 5 1 1 47841
0 47843 7 1 2 47830 47842
0 47844 5 1 1 47843
0 47845 7 1 2 93019 47844
0 47846 5 2 1 47845
0 47847 7 1 2 47820 105827
0 47848 7 1 2 47804 47847
0 47849 5 1 1 47848
0 47850 7 1 2 85545 47849
0 47851 5 1 1 47850
0 47852 7 1 2 88709 77074
0 47853 7 1 2 96021 47852
0 47854 7 1 2 102714 47853
0 47855 5 1 1 47854
0 47856 7 1 2 47851 47855
0 47857 5 1 1 47856
0 47858 7 1 2 67412 47857
0 47859 5 1 1 47858
0 47860 7 1 2 74407 99068
0 47861 5 2 1 47860
0 47862 7 4 2 85546 78488
0 47863 7 1 2 72472 105831
0 47864 5 1 1 47863
0 47865 7 1 2 105829 47864
0 47866 5 1 1 47865
0 47867 7 1 2 104232 47866
0 47868 5 1 1 47867
0 47869 7 1 2 87152 79511
0 47870 5 1 1 47869
0 47871 7 1 2 101293 47870
0 47872 5 1 1 47871
0 47873 7 2 2 83049 94476
0 47874 5 2 1 105835
0 47875 7 1 2 79495 105836
0 47876 5 1 1 47875
0 47877 7 1 2 100863 105837
0 47878 5 1 1 47877
0 47879 7 1 2 68714 47878
0 47880 5 1 1 47879
0 47881 7 1 2 79786 95188
0 47882 5 1 1 47881
0 47883 7 1 2 105838 47882
0 47884 5 1 1 47883
0 47885 7 1 2 75448 47884
0 47886 5 1 1 47885
0 47887 7 1 2 81924 450
0 47888 7 1 2 91628 47887
0 47889 5 1 1 47888
0 47890 7 1 2 84177 84210
0 47891 5 1 1 47890
0 47892 7 1 2 47889 47891
0 47893 7 1 2 47886 47892
0 47894 7 1 2 47880 47893
0 47895 5 1 1 47894
0 47896 7 1 2 68154 47895
0 47897 5 1 1 47896
0 47898 7 1 2 47876 47897
0 47899 5 1 1 47898
0 47900 7 1 2 72771 47899
0 47901 5 1 1 47900
0 47902 7 1 2 47872 47901
0 47903 5 1 1 47902
0 47904 7 1 2 69977 47903
0 47905 5 1 1 47904
0 47906 7 1 2 101294 83867
0 47907 5 1 1 47906
0 47908 7 1 2 101266 103487
0 47909 5 1 1 47908
0 47910 7 1 2 68715 47909
0 47911 5 1 1 47910
0 47912 7 1 2 66369 103438
0 47913 5 1 1 47912
0 47914 7 1 2 47911 47913
0 47915 5 1 1 47914
0 47916 7 1 2 78417 47915
0 47917 5 1 1 47916
0 47918 7 1 2 47907 47917
0 47919 5 1 1 47918
0 47920 7 1 2 68155 47919
0 47921 5 1 1 47920
0 47922 7 1 2 78418 101822
0 47923 5 1 1 47922
0 47924 7 1 2 66075 94553
0 47925 5 1 1 47924
0 47926 7 2 2 81598 88736
0 47927 5 1 1 105839
0 47928 7 1 2 47925 105840
0 47929 5 1 1 47928
0 47930 7 1 2 47923 47929
0 47931 5 1 1 47930
0 47932 7 1 2 71470 47931
0 47933 5 1 1 47932
0 47934 7 1 2 81925 104799
0 47935 5 1 1 47934
0 47936 7 1 2 72772 97564
0 47937 5 1 1 47936
0 47938 7 1 2 47935 47937
0 47939 5 1 1 47938
0 47940 7 1 2 80946 47939
0 47941 5 1 1 47940
0 47942 7 1 2 81313 83757
0 47943 5 1 1 47942
0 47944 7 1 2 47941 47943
0 47945 5 1 1 47944
0 47946 7 1 2 69978 47945
0 47947 5 1 1 47946
0 47948 7 1 2 47933 47947
0 47949 5 1 1 47948
0 47950 7 1 2 73237 47949
0 47951 5 1 1 47950
0 47952 7 1 2 105828 47951
0 47953 7 1 2 47921 47952
0 47954 7 1 2 47905 47953
0 47955 5 1 1 47954
0 47956 7 1 2 99390 47955
0 47957 5 1 1 47956
0 47958 7 1 2 47868 47957
0 47959 7 1 2 47859 47958
0 47960 5 1 1 47959
0 47961 7 1 2 69614 47960
0 47962 5 1 1 47961
0 47963 7 1 2 89217 75021
0 47964 5 1 1 47963
0 47965 7 1 2 75449 74977
0 47966 5 2 1 47965
0 47967 7 1 2 105815 105841
0 47968 5 1 1 47967
0 47969 7 1 2 47964 47968
0 47970 5 1 1 47969
0 47971 7 1 2 73572 47970
0 47972 5 1 1 47971
0 47973 7 1 2 81774 78898
0 47974 5 1 1 47973
0 47975 7 1 2 86468 47974
0 47976 5 2 1 47975
0 47977 7 1 2 75022 105843
0 47978 5 1 1 47977
0 47979 7 2 2 47972 47978
0 47980 5 3 1 105845
0 47981 7 1 2 101047 105847
0 47982 5 1 1 47981
0 47983 7 2 2 74075 90864
0 47984 5 1 1 105850
0 47985 7 1 2 105848 105851
0 47986 5 1 1 47985
0 47987 7 1 2 64491 105846
0 47988 5 1 1 47987
0 47989 7 1 2 69615 103458
0 47990 5 1 1 47989
0 47991 7 1 2 78463 47990
0 47992 7 1 2 47988 47991
0 47993 5 1 1 47992
0 47994 7 2 2 81775 92260
0 47995 5 4 1 105852
0 47996 7 1 2 75290 95458
0 47997 7 1 2 105853 47996
0 47998 5 1 1 47997
0 47999 7 1 2 93514 105849
0 48000 5 1 1 47999
0 48001 7 1 2 47998 48000
0 48002 7 1 2 47993 48001
0 48003 5 1 1 48002
0 48004 7 1 2 70883 48003
0 48005 5 1 1 48004
0 48006 7 1 2 47986 48005
0 48007 5 1 1 48006
0 48008 7 1 2 69263 48007
0 48009 5 1 1 48008
0 48010 7 1 2 47982 48009
0 48011 5 1 1 48010
0 48012 7 1 2 67413 48011
0 48013 5 1 1 48012
0 48014 7 1 2 77488 102054
0 48015 5 3 1 48014
0 48016 7 1 2 10768 105858
0 48017 5 1 1 48016
0 48018 7 1 2 67414 48017
0 48019 5 1 1 48018
0 48020 7 1 2 35185 48019
0 48021 5 2 1 48020
0 48022 7 1 2 84558 105861
0 48023 5 1 1 48022
0 48024 7 1 2 95640 100382
0 48025 7 1 2 97178 48024
0 48026 5 1 1 48025
0 48027 7 1 2 48023 48026
0 48028 5 1 1 48027
0 48029 7 1 2 99738 48028
0 48030 5 1 1 48029
0 48031 7 1 2 99608 94512
0 48032 5 1 1 48031
0 48033 7 1 2 77809 87168
0 48034 5 1 1 48033
0 48035 7 1 2 48032 48034
0 48036 5 1 1 48035
0 48037 7 1 2 70884 98108
0 48038 5 1 1 48037
0 48039 7 1 2 95388 102471
0 48040 5 1 1 48039
0 48041 7 1 2 48038 48040
0 48042 5 1 1 48041
0 48043 7 1 2 69264 48042
0 48044 5 1 1 48043
0 48045 7 1 2 85462 99080
0 48046 7 1 2 97216 48045
0 48047 5 1 1 48046
0 48048 7 1 2 48044 48047
0 48049 5 1 1 48048
0 48050 7 1 2 48036 48049
0 48051 5 1 1 48050
0 48052 7 1 2 99783 104001
0 48053 5 1 1 48052
0 48054 7 1 2 102782 105023
0 48055 5 1 1 48054
0 48056 7 1 2 48053 48055
0 48057 5 1 1 48056
0 48058 7 1 2 97268 48057
0 48059 5 1 1 48058
0 48060 7 1 2 79071 95372
0 48061 7 1 2 84514 48060
0 48062 7 1 2 99519 48061
0 48063 5 1 1 48062
0 48064 7 1 2 48059 48063
0 48065 7 1 2 48051 48064
0 48066 7 1 2 48030 48065
0 48067 5 1 1 48066
0 48068 7 1 2 68716 48067
0 48069 5 1 1 48068
0 48070 7 1 2 103225 103227
0 48071 5 1 1 48070
0 48072 7 3 2 98291 96210
0 48073 7 1 2 48071 105863
0 48074 5 1 1 48073
0 48075 7 1 2 81061 102600
0 48076 5 1 1 48075
0 48077 7 1 2 34081 48076
0 48078 5 1 1 48077
0 48079 7 1 2 82651 48078
0 48080 5 1 1 48079
0 48081 7 1 2 48074 48080
0 48082 7 1 2 48069 48081
0 48083 7 1 2 48013 48082
0 48084 5 1 1 48083
0 48085 7 1 2 64867 48084
0 48086 5 1 1 48085
0 48087 7 1 2 67780 105821
0 48088 5 1 1 48087
0 48089 7 1 2 85656 85045
0 48090 5 1 1 48089
0 48091 7 1 2 48088 48090
0 48092 5 1 1 48091
0 48093 7 1 2 71173 48092
0 48094 5 1 1 48093
0 48095 7 1 2 93201 85795
0 48096 5 1 1 48095
0 48097 7 1 2 48094 48096
0 48098 5 2 1 48097
0 48099 7 2 2 83333 105866
0 48100 5 1 1 105868
0 48101 7 1 2 97532 90239
0 48102 5 1 1 48101
0 48103 7 1 2 48100 48102
0 48104 5 1 1 48103
0 48105 7 1 2 72473 76339
0 48106 7 1 2 48104 48105
0 48107 5 1 1 48106
0 48108 7 1 2 72773 92776
0 48109 7 1 2 100418 48108
0 48110 7 1 2 105822 48109
0 48111 5 1 1 48110
0 48112 7 1 2 48107 48111
0 48113 5 1 1 48112
0 48114 7 1 2 70885 48113
0 48115 5 1 1 48114
0 48116 7 1 2 97916 105869
0 48117 5 1 1 48116
0 48118 7 1 2 48115 48117
0 48119 5 1 1 48118
0 48120 7 1 2 64492 48119
0 48121 5 1 1 48120
0 48122 7 1 2 38587 105818
0 48123 5 2 1 48122
0 48124 7 1 2 96765 105870
0 48125 5 1 1 48124
0 48126 7 2 2 87028 104497
0 48127 7 1 2 101157 105872
0 48128 5 1 1 48127
0 48129 7 1 2 48125 48128
0 48130 5 1 1 48129
0 48131 7 1 2 70886 48130
0 48132 5 1 1 48131
0 48133 7 1 2 102591 87481
0 48134 5 1 1 48133
0 48135 7 1 2 48132 48134
0 48136 5 1 1 48135
0 48137 7 1 2 101498 48136
0 48138 5 1 1 48137
0 48139 7 2 2 100640 84515
0 48140 5 1 1 105874
0 48141 7 1 2 67781 105871
0 48142 5 1 1 48141
0 48143 7 1 2 81970 105873
0 48144 5 1 1 48143
0 48145 7 1 2 48142 48144
0 48146 5 1 1 48145
0 48147 7 1 2 69979 48146
0 48148 5 1 1 48147
0 48149 7 1 2 48140 48148
0 48150 5 1 1 48149
0 48151 7 1 2 98592 48150
0 48152 5 1 1 48151
0 48153 7 1 2 65848 48152
0 48154 5 1 1 48153
0 48155 7 1 2 72474 87482
0 48156 7 1 2 102529 48155
0 48157 5 1 1 48156
0 48158 7 1 2 101934 104270
0 48159 5 2 1 48158
0 48160 7 1 2 85748 105876
0 48161 5 1 1 48160
0 48162 7 1 2 70887 48161
0 48163 7 1 2 48157 48162
0 48164 5 1 1 48163
0 48165 7 1 2 64493 48164
0 48166 5 1 1 48165
0 48167 7 1 2 82727 81423
0 48168 7 1 2 103565 48167
0 48169 7 1 2 101240 48168
0 48170 5 1 1 48169
0 48171 7 1 2 48166 48170
0 48172 5 1 1 48171
0 48173 7 1 2 71174 48172
0 48174 7 1 2 48154 48173
0 48175 5 1 1 48174
0 48176 7 1 2 48138 48175
0 48177 5 1 1 48176
0 48178 7 1 2 70262 48177
0 48179 5 1 1 48178
0 48180 7 1 2 48121 48179
0 48181 5 1 1 48180
0 48182 7 1 2 69265 48181
0 48183 5 1 1 48182
0 48184 7 1 2 75450 105867
0 48185 5 1 1 48184
0 48186 7 3 2 74566 82652
0 48187 5 1 1 105878
0 48188 7 1 2 105406 105879
0 48189 5 1 1 48188
0 48190 7 1 2 48185 48189
0 48191 5 1 1 48190
0 48192 7 1 2 69980 48191
0 48193 5 1 1 48192
0 48194 7 2 2 86898 81404
0 48195 7 1 2 77810 76710
0 48196 7 1 2 105881 48195
0 48197 5 1 1 48196
0 48198 7 1 2 48193 48197
0 48199 5 1 1 48198
0 48200 7 1 2 64494 102302
0 48201 7 1 2 48199 48200
0 48202 5 1 1 48201
0 48203 7 1 2 96922 104817
0 48204 5 2 1 48203
0 48205 7 1 2 99411 82653
0 48206 5 1 1 48205
0 48207 7 1 2 105883 48206
0 48208 5 1 1 48207
0 48209 7 1 2 76664 48208
0 48210 5 1 1 48209
0 48211 7 1 2 85547 80236
0 48212 7 1 2 100984 48211
0 48213 5 1 1 48212
0 48214 7 1 2 48210 48213
0 48215 5 1 1 48214
0 48216 7 1 2 69616 48215
0 48217 5 1 1 48216
0 48218 7 1 2 80814 82419
0 48219 5 1 1 48218
0 48220 7 1 2 104815 104412
0 48221 5 1 1 48220
0 48222 7 1 2 48219 48221
0 48223 5 1 1 48222
0 48224 7 1 2 69266 48223
0 48225 5 1 1 48224
0 48226 7 1 2 96868 100387
0 48227 7 1 2 100823 48226
0 48228 5 1 1 48227
0 48229 7 1 2 48225 48228
0 48230 5 1 1 48229
0 48231 7 1 2 67415 48230
0 48232 5 1 1 48231
0 48233 7 1 2 48217 48232
0 48234 5 1 1 48233
0 48235 7 1 2 83758 48234
0 48236 5 1 1 48235
0 48237 7 4 2 2667 105508
0 48238 7 1 2 100014 86822
0 48239 5 1 1 48238
0 48240 7 1 2 64495 103526
0 48241 5 1 1 48240
0 48242 7 1 2 48239 48241
0 48243 5 1 1 48242
0 48244 7 1 2 105885 48243
0 48245 5 1 1 48244
0 48246 7 1 2 75034 86837
0 48247 5 1 1 48246
0 48248 7 1 2 47927 48247
0 48249 5 1 1 48248
0 48250 7 1 2 69981 48249
0 48251 5 1 1 48250
0 48252 7 1 2 78419 101263
0 48253 5 1 1 48252
0 48254 7 1 2 48251 48253
0 48255 5 1 1 48254
0 48256 7 1 2 68717 104111
0 48257 7 1 2 48255 48256
0 48258 5 1 1 48257
0 48259 7 1 2 48245 48258
0 48260 5 1 1 48259
0 48261 7 1 2 67416 48260
0 48262 5 1 1 48261
0 48263 7 1 2 82798 101759
0 48264 5 1 1 48263
0 48265 7 1 2 71175 48264
0 48266 5 1 1 48265
0 48267 7 1 2 101232 38648
0 48268 7 1 2 48266 48267
0 48269 5 1 1 48268
0 48270 7 1 2 69982 48269
0 48271 5 1 1 48270
0 48272 7 1 2 91136 103857
0 48273 5 1 1 48272
0 48274 7 1 2 80947 104531
0 48275 5 1 1 48274
0 48276 7 1 2 48273 48275
0 48277 7 1 2 48271 48276
0 48278 5 1 1 48277
0 48279 7 1 2 105316 48278
0 48280 5 1 1 48279
0 48281 7 1 2 48262 48280
0 48282 7 1 2 48236 48281
0 48283 5 1 1 48282
0 48284 7 1 2 76095 48283
0 48285 5 1 1 48284
0 48286 7 1 2 81926 95864
0 48287 5 1 1 48286
0 48288 7 1 2 64496 105826
0 48289 5 1 1 48288
0 48290 7 1 2 88871 48289
0 48291 5 1 1 48290
0 48292 7 1 2 48287 48291
0 48293 5 1 1 48292
0 48294 7 1 2 65192 48293
0 48295 5 1 1 48294
0 48296 7 1 2 69983 100012
0 48297 5 1 1 48296
0 48298 7 1 2 69617 89204
0 48299 5 1 1 48298
0 48300 7 1 2 48297 48299
0 48301 5 1 1 48300
0 48302 7 1 2 73573 48301
0 48303 5 1 1 48302
0 48304 7 1 2 48295 48303
0 48305 5 1 1 48304
0 48306 7 1 2 66076 48305
0 48307 5 1 1 48306
0 48308 7 1 2 105770 105680
0 48309 5 1 1 48308
0 48310 7 1 2 78386 48309
0 48311 5 1 1 48310
0 48312 7 1 2 48307 48311
0 48313 5 1 1 48312
0 48314 7 1 2 102601 48313
0 48315 5 1 1 48314
0 48316 7 1 2 82636 104522
0 48317 5 1 1 48316
0 48318 7 1 2 71176 99487
0 48319 7 1 2 101772 48318
0 48320 5 1 1 48319
0 48321 7 1 2 48317 48320
0 48322 5 1 1 48321
0 48323 7 1 2 69984 48322
0 48324 5 1 1 48323
0 48325 7 2 2 87222 105771
0 48326 5 1 1 105889
0 48327 7 1 2 104523 48326
0 48328 5 1 1 48327
0 48329 7 1 2 48324 48328
0 48330 5 1 1 48329
0 48331 7 1 2 93020 48330
0 48332 5 1 1 48331
0 48333 7 1 2 48315 48332
0 48334 7 1 2 48285 48333
0 48335 7 1 2 48202 48334
0 48336 7 1 2 48183 48335
0 48337 7 1 2 48086 48336
0 48338 7 1 2 47962 48337
0 48339 5 1 1 48338
0 48340 7 1 2 96330 48339
0 48341 5 1 1 48340
0 48342 7 1 2 99034 96512
0 48343 7 1 2 96022 48342
0 48344 7 1 2 85424 99333
0 48345 7 1 2 105779 48344
0 48346 7 1 2 48343 48345
0 48347 5 1 1 48346
0 48348 7 1 2 48341 48347
0 48349 5 1 1 48348
0 48350 7 1 2 67135 48349
0 48351 5 1 1 48350
0 48352 7 1 2 95086 82405
0 48353 5 1 1 48352
0 48354 7 1 2 80743 101475
0 48355 5 1 1 48354
0 48356 7 1 2 48353 48355
0 48357 5 1 1 48356
0 48358 7 1 2 67782 48357
0 48359 5 1 1 48358
0 48360 7 1 2 88681 87776
0 48361 5 1 1 48360
0 48362 7 1 2 48359 48361
0 48363 5 1 1 48362
0 48364 7 1 2 71177 48363
0 48365 5 1 1 48364
0 48366 7 2 2 80380 85086
0 48367 7 1 2 105226 105891
0 48368 5 1 1 48367
0 48369 7 1 2 48365 48368
0 48370 5 1 1 48369
0 48371 7 1 2 69618 48370
0 48372 5 1 1 48371
0 48373 7 2 2 80839 88353
0 48374 7 1 2 105892 105893
0 48375 5 1 1 48374
0 48376 7 1 2 48372 48375
0 48377 5 1 1 48376
0 48378 7 1 2 99391 48377
0 48379 5 1 1 48378
0 48380 7 1 2 68504 103032
0 48381 5 1 1 48380
0 48382 7 1 2 103493 48381
0 48383 5 1 1 48382
0 48384 7 1 2 100514 48383
0 48385 5 1 1 48384
0 48386 7 1 2 99423 103269
0 48387 7 1 2 104705 48386
0 48388 5 1 1 48387
0 48389 7 1 2 48385 48388
0 48390 5 1 1 48389
0 48391 7 1 2 67783 48390
0 48392 5 1 1 48391
0 48393 7 1 2 68505 87185
0 48394 5 1 1 48393
0 48395 7 1 2 82855 48394
0 48396 5 6 1 48395
0 48397 7 1 2 82466 98543
0 48398 7 3 2 105895 48397
0 48399 5 1 1 105901
0 48400 7 1 2 76610 105902
0 48401 5 1 1 48400
0 48402 7 1 2 48392 48401
0 48403 5 1 1 48402
0 48404 7 1 2 67417 48403
0 48405 5 1 1 48404
0 48406 7 1 2 101204 101915
0 48407 7 1 2 105896 48406
0 48408 5 1 1 48407
0 48409 7 1 2 48405 48408
0 48410 5 1 1 48409
0 48411 7 1 2 66594 48410
0 48412 5 1 1 48411
0 48413 7 2 2 72774 104432
0 48414 5 1 1 105904
0 48415 7 1 2 93521 48414
0 48416 5 1 1 48415
0 48417 7 1 2 70888 48416
0 48418 5 1 1 48417
0 48419 7 1 2 47984 48418
0 48420 5 1 1 48419
0 48421 7 1 2 69267 48420
0 48422 5 1 1 48421
0 48423 7 1 2 101049 48422
0 48424 5 1 1 48423
0 48425 7 1 2 101476 48424
0 48426 5 1 1 48425
0 48427 7 2 2 85463 92787
0 48428 5 1 1 105906
0 48429 7 1 2 69268 104803
0 48430 5 1 1 48429
0 48431 7 1 2 48428 48430
0 48432 5 4 1 48431
0 48433 7 1 2 104800 105908
0 48434 5 1 1 48433
0 48435 7 1 2 69269 104809
0 48436 5 1 1 48435
0 48437 7 1 2 25661 48436
0 48438 5 2 1 48437
0 48439 7 1 2 105082 105912
0 48440 5 1 1 48439
0 48441 7 1 2 48434 48440
0 48442 5 1 1 48441
0 48443 7 1 2 80646 48442
0 48444 5 1 1 48443
0 48445 7 1 2 48426 48444
0 48446 5 1 1 48445
0 48447 7 1 2 67418 48446
0 48448 5 1 1 48447
0 48449 7 1 2 48412 48448
0 48450 7 1 2 48379 48449
0 48451 5 1 1 48450
0 48452 7 1 2 65193 48451
0 48453 5 1 1 48452
0 48454 7 1 2 80545 104779
0 48455 5 1 1 48454
0 48456 7 4 2 85548 81062
0 48457 7 2 2 70523 96035
0 48458 7 1 2 105914 105918
0 48459 5 1 1 48458
0 48460 7 1 2 48455 48459
0 48461 5 1 1 48460
0 48462 7 1 2 74863 48461
0 48463 5 1 1 48462
0 48464 7 1 2 90838 43176
0 48465 5 1 1 48464
0 48466 7 1 2 80546 48465
0 48467 5 1 1 48466
0 48468 7 1 2 93885 96075
0 48469 5 1 1 48468
0 48470 7 1 2 48467 48469
0 48471 5 1 1 48470
0 48472 7 1 2 104112 48471
0 48473 5 1 1 48472
0 48474 7 1 2 82856 86760
0 48475 5 2 1 48474
0 48476 7 1 2 93357 105920
0 48477 5 1 1 48476
0 48478 7 1 2 105489 105832
0 48479 5 1 1 48478
0 48480 7 1 2 48477 48479
0 48481 5 1 1 48480
0 48482 7 1 2 64497 48481
0 48483 5 1 1 48482
0 48484 7 1 2 48473 48483
0 48485 5 1 1 48484
0 48486 7 1 2 74567 48485
0 48487 5 1 1 48486
0 48488 7 1 2 48463 48487
0 48489 5 1 1 48488
0 48490 7 1 2 79865 48489
0 48491 5 1 1 48490
0 48492 7 2 2 74076 95272
0 48493 5 1 1 105922
0 48494 7 1 2 104807 48493
0 48495 5 1 1 48494
0 48496 7 1 2 64498 48495
0 48497 5 1 1 48496
0 48498 7 1 2 103798 104796
0 48499 5 2 1 48498
0 48500 7 1 2 93061 105924
0 48501 5 1 1 48500
0 48502 7 1 2 48497 48501
0 48503 5 1 1 48502
0 48504 7 1 2 89070 48503
0 48505 5 1 1 48504
0 48506 7 1 2 94840 105905
0 48507 5 1 1 48506
0 48508 7 1 2 87459 104775
0 48509 5 1 1 48508
0 48510 7 1 2 48507 48509
0 48511 5 1 1 48510
0 48512 7 1 2 73574 48511
0 48513 5 1 1 48512
0 48514 7 1 2 48505 48513
0 48515 5 1 1 48514
0 48516 7 1 2 69270 48515
0 48517 5 1 1 48516
0 48518 7 1 2 69619 105925
0 48519 5 1 1 48518
0 48520 7 1 2 71867 78500
0 48521 5 1 1 48520
0 48522 7 1 2 48519 48521
0 48523 5 1 1 48522
0 48524 7 1 2 89071 48523
0 48525 5 1 1 48524
0 48526 7 1 2 88851 101037
0 48527 5 1 1 48526
0 48528 7 1 2 48525 48527
0 48529 5 1 1 48528
0 48530 7 1 2 85464 48529
0 48531 5 1 1 48530
0 48532 7 1 2 48517 48531
0 48533 5 1 1 48532
0 48534 7 1 2 97411 48533
0 48535 5 1 1 48534
0 48536 7 1 2 72775 78055
0 48537 5 1 1 48536
0 48538 7 1 2 90839 48537
0 48539 5 1 1 48538
0 48540 7 1 2 105909 48539
0 48541 5 1 1 48540
0 48542 7 1 2 100515 82087
0 48543 5 1 1 48542
0 48544 7 1 2 48541 48543
0 48545 5 1 1 48544
0 48546 7 1 2 84856 48545
0 48547 5 1 1 48546
0 48548 7 1 2 99930 105833
0 48549 5 1 1 48548
0 48550 7 1 2 99553 86141
0 48551 7 1 2 104805 48550
0 48552 5 1 1 48551
0 48553 7 1 2 48549 48552
0 48554 5 1 1 48553
0 48555 7 1 2 105083 48554
0 48556 5 1 1 48555
0 48557 7 1 2 83449 82057
0 48558 5 1 1 48557
0 48559 7 1 2 79937 83296
0 48560 5 1 1 48559
0 48561 7 1 2 48558 48560
0 48562 5 1 1 48561
0 48563 7 1 2 105913 48562
0 48564 5 1 1 48563
0 48565 7 1 2 85087 86653
0 48566 7 1 2 104695 48565
0 48567 5 1 1 48566
0 48568 7 1 2 48564 48567
0 48569 7 1 2 48556 48568
0 48570 7 1 2 48547 48569
0 48571 7 1 2 86311 18568
0 48572 5 1 1 48571
0 48573 7 1 2 105910 48572
0 48574 5 1 1 48573
0 48575 7 1 2 92656 83465
0 48576 5 1 1 48575
0 48577 7 1 2 30387 48576
0 48578 5 1 1 48577
0 48579 7 1 2 104113 48578
0 48580 5 1 1 48579
0 48581 7 1 2 83450 74200
0 48582 7 1 2 74347 48581
0 48583 5 1 1 48582
0 48584 7 1 2 48580 48583
0 48585 7 1 2 48574 48584
0 48586 5 1 1 48585
0 48587 7 1 2 104801 48586
0 48588 5 1 1 48587
0 48589 7 1 2 93358 105592
0 48590 5 1 1 48589
0 48591 7 1 2 80744 105834
0 48592 5 1 1 48591
0 48593 7 1 2 48590 48592
0 48594 5 1 1 48593
0 48595 7 1 2 105084 48594
0 48596 5 1 1 48595
0 48597 7 1 2 65496 105185
0 48598 5 1 1 48597
0 48599 7 1 2 16212 48598
0 48600 5 1 1 48599
0 48601 7 1 2 105911 48600
0 48602 5 1 1 48601
0 48603 7 1 2 48596 48602
0 48604 5 1 1 48603
0 48605 7 1 2 75451 48604
0 48606 5 1 1 48605
0 48607 7 1 2 48588 48606
0 48608 7 1 2 48570 48607
0 48609 7 1 2 48535 48608
0 48610 7 1 2 48491 48609
0 48611 5 1 1 48610
0 48612 7 1 2 67419 48611
0 48613 5 1 1 48612
0 48614 7 1 2 77921 105897
0 48615 5 1 1 48614
0 48616 7 1 2 76505 105593
0 48617 5 1 1 48616
0 48618 7 1 2 48615 48617
0 48619 5 1 1 48618
0 48620 7 1 2 70263 48619
0 48621 5 1 1 48620
0 48622 7 1 2 78711 87186
0 48623 5 1 1 48622
0 48624 7 1 2 93687 83160
0 48625 7 1 2 95199 48624
0 48626 5 1 1 48625
0 48627 7 1 2 48623 48626
0 48628 5 1 1 48627
0 48629 7 1 2 76506 48628
0 48630 5 1 1 48629
0 48631 7 1 2 48621 48630
0 48632 5 1 1 48631
0 48633 7 1 2 78519 48632
0 48634 5 1 1 48633
0 48635 7 1 2 90006 104901
0 48636 5 1 1 48635
0 48637 7 1 2 73575 94261
0 48638 7 1 2 101038 48637
0 48639 5 1 1 48638
0 48640 7 1 2 48636 48639
0 48641 5 1 1 48640
0 48642 7 1 2 97412 48641
0 48643 5 1 1 48642
0 48644 7 1 2 86684 73986
0 48645 5 1 1 48644
0 48646 7 1 2 46110 48645
0 48647 5 1 1 48646
0 48648 7 1 2 78489 82058
0 48649 7 1 2 48647 48648
0 48650 5 1 1 48649
0 48651 7 1 2 48643 48650
0 48652 7 1 2 48634 48651
0 48653 5 1 1 48652
0 48654 7 1 2 99392 48653
0 48655 5 1 1 48654
0 48656 7 1 2 48613 48655
0 48657 7 1 2 48453 48656
0 48658 5 1 1 48657
0 48659 7 1 2 73238 48658
0 48660 5 1 1 48659
0 48661 7 1 2 99465 78490
0 48662 5 2 1 48661
0 48663 7 1 2 70889 98411
0 48664 5 1 1 48663
0 48665 7 1 2 103706 48664
0 48666 5 1 1 48665
0 48667 7 1 2 69271 48666
0 48668 5 1 1 48667
0 48669 7 1 2 105926 48668
0 48670 5 5 1 48669
0 48671 7 2 2 98936 105928
0 48672 5 1 1 105933
0 48673 7 1 2 71471 48672
0 48674 5 1 1 48673
0 48675 7 1 2 97206 98821
0 48676 5 1 1 48675
0 48677 7 1 2 86276 105431
0 48678 5 1 1 48677
0 48679 7 1 2 48676 48678
0 48680 5 1 1 48679
0 48681 7 1 2 69272 48680
0 48682 5 1 1 48681
0 48683 7 1 2 101042 97207
0 48684 5 1 1 48683
0 48685 7 1 2 48682 48684
0 48686 5 1 1 48685
0 48687 7 1 2 84857 48686
0 48688 5 1 1 48687
0 48689 7 1 2 66783 102806
0 48690 7 2 2 105886 48689
0 48691 5 1 1 105935
0 48692 7 1 2 66370 48691
0 48693 7 1 2 48688 48692
0 48694 5 1 1 48693
0 48695 7 1 2 69985 48694
0 48696 7 1 2 48674 48695
0 48697 5 1 1 48696
0 48698 7 1 2 76711 97225
0 48699 5 1 1 48698
0 48700 7 1 2 66784 97754
0 48701 5 1 1 48700
0 48702 7 1 2 48699 48701
0 48703 5 1 1 48702
0 48704 7 1 2 70890 48703
0 48705 5 1 1 48704
0 48706 7 1 2 78491 102454
0 48707 5 1 1 48706
0 48708 7 1 2 48705 48707
0 48709 5 1 1 48708
0 48710 7 1 2 69273 48709
0 48711 5 1 1 48710
0 48712 7 1 2 101043 102447
0 48713 5 1 1 48712
0 48714 7 1 2 48711 48713
0 48715 5 1 1 48714
0 48716 7 1 2 102143 48715
0 48717 5 1 1 48716
0 48718 7 1 2 65497 102148
0 48719 5 1 1 48718
0 48720 7 1 2 66371 94935
0 48721 5 1 1 48720
0 48722 7 1 2 73576 99501
0 48723 5 1 1 48722
0 48724 7 1 2 103464 48723
0 48725 7 1 2 48721 48724
0 48726 5 1 1 48725
0 48727 7 1 2 80647 48726
0 48728 5 1 1 48727
0 48729 7 1 2 48719 48728
0 48730 5 1 1 48729
0 48731 7 1 2 98378 78492
0 48732 5 1 1 48731
0 48733 7 1 2 98394 48732
0 48734 5 1 1 48733
0 48735 7 1 2 70891 48734
0 48736 5 1 1 48735
0 48737 7 1 2 103707 48736
0 48738 5 1 1 48737
0 48739 7 1 2 69274 48738
0 48740 5 1 1 48739
0 48741 7 1 2 48740 105927
0 48742 5 1 1 48741
0 48743 7 1 2 48730 48742
0 48744 5 1 1 48743
0 48745 7 1 2 71472 103254
0 48746 5 1 1 48745
0 48747 7 1 2 100710 103862
0 48748 7 1 2 48746 48747
0 48749 5 1 1 48748
0 48750 7 1 2 97371 104956
0 48751 5 1 1 48750
0 48752 7 1 2 97208 48751
0 48753 7 1 2 105887 48752
0 48754 5 1 1 48753
0 48755 7 1 2 48749 48754
0 48756 5 1 1 48755
0 48757 7 1 2 84858 48756
0 48758 5 1 1 48757
0 48759 7 2 2 81287 79512
0 48760 7 1 2 105936 105937
0 48761 5 1 1 48760
0 48762 7 1 2 64499 48761
0 48763 7 1 2 48758 48762
0 48764 7 1 2 48744 48763
0 48765 7 1 2 48717 48764
0 48766 7 1 2 48697 48765
0 48767 5 1 1 48766
0 48768 7 1 2 99695 98198
0 48769 5 1 1 48768
0 48770 7 1 2 96964 94349
0 48771 5 1 1 48770
0 48772 7 1 2 48769 48771
0 48773 5 1 1 48772
0 48774 7 1 2 98822 48773
0 48775 5 1 1 48774
0 48776 7 1 2 85465 98191
0 48777 7 1 2 82219 95515
0 48778 7 1 2 48776 48777
0 48779 5 1 1 48778
0 48780 7 1 2 97741 103514
0 48781 7 1 2 92184 48780
0 48782 5 1 1 48781
0 48783 7 1 2 48779 48782
0 48784 7 1 2 48775 48783
0 48785 5 1 1 48784
0 48786 7 1 2 82997 48785
0 48787 5 1 1 48786
0 48788 7 2 2 77526 97059
0 48789 5 1 1 105939
0 48790 7 1 2 98395 48789
0 48791 5 1 1 48790
0 48792 7 1 2 85549 48791
0 48793 5 1 1 48792
0 48794 7 1 2 100113 93359
0 48795 5 1 1 48794
0 48796 7 1 2 105830 48795
0 48797 7 1 2 48793 48796
0 48798 5 1 1 48797
0 48799 7 1 2 80823 48798
0 48800 5 1 1 48799
0 48801 7 1 2 48787 48800
0 48802 5 1 1 48801
0 48803 7 1 2 76507 48802
0 48804 5 1 1 48803
0 48805 7 1 2 76239 105934
0 48806 5 1 1 48805
0 48807 7 1 2 69620 48806
0 48808 7 1 2 48804 48807
0 48809 5 1 1 48808
0 48810 7 1 2 48767 48809
0 48811 5 1 1 48810
0 48812 7 1 2 87187 102149
0 48813 5 1 1 48812
0 48814 7 2 2 68506 97515
0 48815 5 1 1 105941
0 48816 7 1 2 97413 105942
0 48817 5 1 1 48816
0 48818 7 1 2 48813 48817
0 48819 5 1 1 48818
0 48820 7 1 2 99757 48819
0 48821 5 1 1 48820
0 48822 7 2 2 99412 84859
0 48823 5 1 1 105943
0 48824 7 1 2 68718 105944
0 48825 7 1 2 103281 48824
0 48826 5 1 1 48825
0 48827 7 1 2 48821 48826
0 48828 5 1 1 48827
0 48829 7 1 2 69621 48828
0 48830 5 1 1 48829
0 48831 7 1 2 71473 102900
0 48832 5 1 1 48831
0 48833 7 1 2 101694 48832
0 48834 5 1 1 48833
0 48835 7 1 2 69622 48834
0 48836 5 1 1 48835
0 48837 7 1 2 83781 79915
0 48838 5 1 1 48837
0 48839 7 1 2 48836 48838
0 48840 5 1 1 48839
0 48841 7 1 2 80648 48840
0 48842 5 1 1 48841
0 48843 7 1 2 79251 89955
0 48844 5 1 1 48843
0 48845 7 1 2 48842 48844
0 48846 5 1 1 48845
0 48847 7 1 2 105751 48846
0 48848 5 1 1 48847
0 48849 7 1 2 98514 92788
0 48850 5 1 1 48849
0 48851 7 1 2 70892 104198
0 48852 5 1 1 48851
0 48853 7 1 2 48850 48852
0 48854 5 1 1 48853
0 48855 7 1 2 69275 48854
0 48856 5 1 1 48855
0 48857 7 2 2 67420 105907
0 48858 5 1 1 105945
0 48859 7 1 2 48856 48858
0 48860 5 1 1 48859
0 48861 7 1 2 87236 48860
0 48862 5 1 1 48861
0 48863 7 1 2 102150 105514
0 48864 5 1 1 48863
0 48865 7 1 2 48862 48864
0 48866 5 1 1 48865
0 48867 7 1 2 80745 48866
0 48868 5 1 1 48867
0 48869 7 1 2 99668 98199
0 48870 5 1 1 48869
0 48871 7 3 2 68719 99413
0 48872 5 1 1 105947
0 48873 7 1 2 83793 105948
0 48874 5 1 1 48873
0 48875 7 1 2 48870 48874
0 48876 5 1 1 48875
0 48877 7 1 2 79287 95189
0 48878 7 1 2 48876 48877
0 48879 5 1 1 48878
0 48880 7 1 2 48868 48879
0 48881 7 1 2 48848 48880
0 48882 7 1 2 48830 48881
0 48883 5 1 1 48882
0 48884 7 1 2 83759 48883
0 48885 5 1 1 48884
0 48886 7 1 2 48811 48885
0 48887 5 1 1 48886
0 48888 7 1 2 68156 48887
0 48889 5 1 1 48888
0 48890 7 1 2 67784 103036
0 48891 7 1 2 100516 48890
0 48892 5 1 1 48891
0 48893 7 1 2 48399 48892
0 48894 5 1 1 48893
0 48895 7 1 2 67421 48894
0 48896 5 1 1 48895
0 48897 7 1 2 105864 105898
0 48898 5 1 1 48897
0 48899 7 1 2 48896 48898
0 48900 5 1 1 48899
0 48901 7 1 2 81302 48900
0 48902 5 1 1 48901
0 48903 7 1 2 48889 48902
0 48904 7 1 2 48660 48903
0 48905 5 1 1 48904
0 48906 7 1 2 98128 48905
0 48907 5 1 1 48906
0 48908 7 1 2 48351 48907
0 48909 5 1 1 48908
0 48910 7 1 2 76810 48909
0 48911 5 1 1 48910
0 48912 7 1 2 63809 48911
0 48913 7 1 2 47770 48912
0 48914 5 1 1 48913
0 48915 7 1 2 71178 100045
0 48916 5 1 1 48915
0 48917 7 1 2 104098 48916
0 48918 5 1 1 48917
0 48919 7 1 2 69623 48918
0 48920 5 1 1 48919
0 48921 7 2 2 77090 104852
0 48922 7 1 2 82013 105950
0 48923 5 1 1 48922
0 48924 7 1 2 48920 48923
0 48925 5 1 1 48924
0 48926 7 1 2 70524 48925
0 48927 5 1 1 48926
0 48928 7 1 2 100054 23234
0 48929 5 1 1 48928
0 48930 7 1 2 100052 48929
0 48931 5 1 1 48930
0 48932 7 1 2 77191 48931
0 48933 5 1 1 48932
0 48934 7 1 2 48927 48933
0 48935 5 1 1 48934
0 48936 7 1 2 64198 48935
0 48937 5 1 1 48936
0 48938 7 1 2 82662 105890
0 48939 5 1 1 48938
0 48940 7 1 2 64500 48939
0 48941 5 1 1 48940
0 48942 7 2 2 81776 93753
0 48943 7 1 2 105556 105952
0 48944 5 1 1 48943
0 48945 7 1 2 48941 48944
0 48946 5 1 1 48945
0 48947 7 1 2 98344 48946
0 48948 5 1 1 48947
0 48949 7 1 2 48937 48948
0 48950 5 1 1 48949
0 48951 7 2 2 94830 48950
0 48952 5 1 1 105954
0 48953 7 1 2 78076 105955
0 48954 5 1 1 48953
0 48955 7 1 2 100517 103258
0 48956 5 1 1 48955
0 48957 7 2 2 74692 101017
0 48958 7 1 2 73577 95277
0 48959 7 1 2 105956 48958
0 48960 5 1 1 48959
0 48961 7 1 2 48956 48960
0 48962 5 1 1 48961
0 48963 7 1 2 80746 48962
0 48964 5 1 1 48963
0 48965 7 3 2 70525 102907
0 48966 5 2 1 105958
0 48967 7 1 2 71868 105959
0 48968 5 1 1 48967
0 48969 7 1 2 88386 100757
0 48970 7 1 2 100518 48969
0 48971 7 1 2 48968 48970
0 48972 5 1 1 48971
0 48973 7 1 2 48964 48972
0 48974 5 1 1 48973
0 48975 7 2 2 72183 48974
0 48976 5 1 1 105963
0 48977 7 1 2 75157 105964
0 48978 5 1 1 48977
0 48979 7 1 2 48954 48978
0 48980 5 1 1 48979
0 48981 7 1 2 67422 48980
0 48982 5 1 1 48981
0 48983 7 1 2 66785 103259
0 48984 5 1 1 48983
0 48985 7 1 2 103469 48984
0 48986 5 1 1 48985
0 48987 7 1 2 70526 48986
0 48988 5 1 1 48987
0 48989 7 1 2 82998 103260
0 48990 5 1 1 48989
0 48991 7 1 2 94930 48990
0 48992 5 1 1 48991
0 48993 7 1 2 65498 48992
0 48994 5 1 1 48993
0 48995 7 1 2 48988 48994
0 48996 5 1 1 48995
0 48997 7 1 2 98242 96302
0 48998 7 2 2 48996 48997
0 48999 7 1 2 94781 89867
0 49000 7 1 2 105965 48999
0 49001 5 1 1 49000
0 49002 7 1 2 48982 49001
0 49003 5 1 1 49002
0 49004 7 1 2 68157 49003
0 49005 5 1 1 49004
0 49006 7 1 2 95377 97479
0 49007 7 2 2 87661 49006
0 49008 7 3 2 65611 93734
0 49009 7 1 2 105967 105969
0 49010 5 2 1 49009
0 49011 7 2 2 85444 82571
0 49012 7 1 2 94753 78089
0 49013 5 1 1 49012
0 49014 7 1 2 95709 78118
0 49015 5 1 1 49014
0 49016 7 1 2 49013 49015
0 49017 5 1 1 49016
0 49018 7 1 2 105974 49017
0 49019 5 2 1 49018
0 49020 7 3 2 81927 78090
0 49021 5 2 1 105978
0 49022 7 1 2 104633 78119
0 49023 5 1 1 49022
0 49024 7 1 2 105981 49023
0 49025 5 1 1 49024
0 49026 7 1 2 68507 49025
0 49027 5 1 1 49026
0 49028 7 1 2 87188 87873
0 49029 5 1 1 49028
0 49030 7 1 2 49027 49029
0 49031 5 1 1 49030
0 49032 7 1 2 73239 49031
0 49033 5 1 1 49032
0 49034 7 2 2 89355 86009
0 49035 7 1 2 79044 105983
0 49036 5 1 1 49035
0 49037 7 1 2 49033 49036
0 49038 5 1 1 49037
0 49039 7 1 2 101018 49038
0 49040 5 1 1 49039
0 49041 7 2 2 79739 101008
0 49042 7 2 2 85642 78091
0 49043 5 1 1 105987
0 49044 7 1 2 83976 77733
0 49045 7 1 2 75158 49044
0 49046 5 1 1 49045
0 49047 7 1 2 49043 49046
0 49048 5 1 1 49047
0 49049 7 1 2 105985 49048
0 49050 5 1 1 49049
0 49051 7 1 2 49040 49050
0 49052 5 1 1 49051
0 49053 7 1 2 70893 49052
0 49054 5 1 1 49053
0 49055 7 1 2 105976 49054
0 49056 5 1 1 49055
0 49057 7 1 2 67423 49056
0 49058 5 1 1 49057
0 49059 7 1 2 105972 49058
0 49060 5 1 1 49059
0 49061 7 1 2 75452 49060
0 49062 5 1 1 49061
0 49063 7 1 2 75180 86757
0 49064 5 1 1 49063
0 49065 7 1 2 85756 78092
0 49066 5 1 1 49065
0 49067 7 1 2 49064 49066
0 49068 5 1 1 49067
0 49069 7 1 2 76665 49068
0 49070 5 1 1 49069
0 49071 7 1 2 69986 103475
0 49072 5 1 1 49071
0 49073 7 1 2 83552 83586
0 49074 5 1 1 49073
0 49075 7 1 2 49072 49074
0 49076 5 2 1 49075
0 49077 7 1 2 76125 105989
0 49078 5 1 1 49077
0 49079 7 1 2 49070 49078
0 49080 5 1 1 49079
0 49081 7 1 2 101019 49080
0 49082 5 1 1 49081
0 49083 7 1 2 68508 85377
0 49084 7 1 2 100905 49083
0 49085 5 1 1 49084
0 49086 7 1 2 98345 91950
0 49087 7 1 2 104413 49086
0 49088 5 1 1 49087
0 49089 7 1 2 49085 49088
0 49090 5 2 1 49089
0 49091 7 1 2 97710 105991
0 49092 5 1 1 49091
0 49093 7 1 2 49082 49092
0 49094 5 1 1 49093
0 49095 7 1 2 67424 49094
0 49096 5 1 1 49095
0 49097 7 1 2 104291 78093
0 49098 5 1 1 49097
0 49099 7 1 2 97595 105539
0 49100 5 1 1 49099
0 49101 7 1 2 49098 49100
0 49102 5 1 1 49101
0 49103 7 1 2 104945 49102
0 49104 5 1 1 49103
0 49105 7 1 2 49096 49104
0 49106 5 1 1 49105
0 49107 7 1 2 70894 49106
0 49108 5 1 1 49107
0 49109 7 1 2 71179 88837
0 49110 5 1 1 49109
0 49111 7 1 2 105567 49110
0 49112 5 1 1 49111
0 49113 7 1 2 70527 49112
0 49114 5 1 1 49113
0 49115 7 1 2 76666 97558
0 49116 5 1 1 49115
0 49117 7 1 2 49114 49116
0 49118 5 1 1 49117
0 49119 7 1 2 69624 49118
0 49120 5 1 1 49119
0 49121 7 1 2 105697 105951
0 49122 5 1 1 49121
0 49123 7 1 2 49120 49122
0 49124 5 1 1 49123
0 49125 7 1 2 65849 97439
0 49126 7 2 2 49124 49125
0 49127 7 1 2 105993 105970
0 49128 5 1 1 49127
0 49129 7 1 2 49108 49128
0 49130 5 1 1 49129
0 49131 7 1 2 73240 49130
0 49132 5 1 1 49131
0 49133 7 1 2 82610 98203
0 49134 7 1 2 99414 49133
0 49135 7 2 2 100074 49134
0 49136 7 1 2 69625 85188
0 49137 7 1 2 105995 49136
0 49138 5 1 1 49137
0 49139 7 1 2 49132 49138
0 49140 7 1 2 49062 49139
0 49141 7 1 2 49005 49140
0 49142 5 1 1 49141
0 49143 7 1 2 72776 49142
0 49144 5 1 1 49143
0 49145 7 2 2 68158 105170
0 49146 7 1 2 92386 105997
0 49147 5 1 1 49146
0 49148 7 1 2 102107 98861
0 49149 5 1 1 49148
0 49150 7 1 2 49147 49149
0 49151 5 2 1 49150
0 49152 7 1 2 75181 105999
0 49153 5 1 1 49152
0 49154 7 1 2 65850 78094
0 49155 7 1 2 104229 49154
0 49156 5 1 1 49155
0 49157 7 1 2 49153 49156
0 49158 5 1 1 49157
0 49159 7 1 2 77192 49158
0 49160 5 1 1 49159
0 49161 7 1 2 72184 77075
0 49162 7 2 2 105998 49161
0 49163 7 1 2 79093 87965
0 49164 7 1 2 106001 49163
0 49165 5 1 1 49164
0 49166 7 1 2 49160 49165
0 49167 5 1 1 49166
0 49168 7 1 2 69276 49167
0 49169 5 1 1 49168
0 49170 7 1 2 100383 104618
0 49171 7 2 2 104221 49170
0 49172 7 1 2 103983 84234
0 49173 7 1 2 106003 49172
0 49174 5 1 1 49173
0 49175 7 1 2 72475 49174
0 49176 7 1 2 49169 49175
0 49177 5 1 1 49176
0 49178 7 1 2 79288 95153
0 49179 5 1 1 49178
0 49180 7 1 2 82654 81215
0 49181 5 2 1 49180
0 49182 7 1 2 69987 18576
0 49183 7 1 2 106005 49182
0 49184 5 1 1 49183
0 49185 7 1 2 64868 97808
0 49186 5 1 1 49185
0 49187 7 1 2 74568 49186
0 49188 7 1 2 49184 49187
0 49189 5 1 1 49188
0 49190 7 1 2 49179 49189
0 49191 5 1 1 49190
0 49192 7 1 2 101714 49191
0 49193 5 1 1 49192
0 49194 7 1 2 80063 101127
0 49195 5 1 1 49194
0 49196 7 1 2 82574 49195
0 49197 5 1 1 49196
0 49198 7 1 2 86823 49197
0 49199 5 1 1 49198
0 49200 7 1 2 49193 49199
0 49201 5 1 1 49200
0 49202 7 1 2 85466 49201
0 49203 5 1 1 49202
0 49204 7 1 2 69626 92342
0 49205 7 1 2 83910 49204
0 49206 5 1 1 49205
0 49207 7 1 2 19272 49206
0 49208 5 1 1 49207
0 49209 7 1 2 103028 49208
0 49210 5 1 1 49209
0 49211 7 1 2 49203 49210
0 49212 5 1 1 49211
0 49213 7 2 2 67136 49212
0 49214 7 1 2 78077 106007
0 49215 5 1 1 49214
0 49216 7 1 2 98749 93879
0 49217 5 1 1 49216
0 49218 7 1 2 78021 98734
0 49219 5 1 1 49218
0 49220 7 1 2 49217 49219
0 49221 5 1 1 49220
0 49222 7 1 2 80948 49221
0 49223 5 1 1 49222
0 49224 7 1 2 93886 98738
0 49225 5 1 1 49224
0 49226 7 1 2 102220 79787
0 49227 5 1 1 49226
0 49228 7 1 2 49225 49227
0 49229 5 1 1 49228
0 49230 7 1 2 74569 49229
0 49231 5 1 1 49230
0 49232 7 1 2 49223 49231
0 49233 5 1 1 49232
0 49234 7 1 2 82728 49233
0 49235 5 1 1 49234
0 49236 7 1 2 77678 100519
0 49237 7 1 2 103372 49236
0 49238 5 1 1 49237
0 49239 7 1 2 49235 49238
0 49240 5 2 1 49239
0 49241 7 1 2 75182 106009
0 49242 5 1 1 49241
0 49243 7 1 2 67425 49242
0 49244 7 1 2 49215 49243
0 49245 5 1 1 49244
0 49246 7 1 2 67785 49245
0 49247 7 1 2 49177 49246
0 49248 5 1 1 49247
0 49249 7 1 2 74693 101128
0 49250 5 2 1 49249
0 49251 7 1 2 87371 106011
0 49252 5 1 1 49251
0 49253 7 1 2 71869 49252
0 49254 5 1 1 49253
0 49255 7 1 2 66786 100935
0 49256 5 1 1 49255
0 49257 7 1 2 102480 92096
0 49258 5 1 1 49257
0 49259 7 1 2 49256 49258
0 49260 7 1 2 49254 49259
0 49261 5 1 1 49260
0 49262 7 1 2 70528 49261
0 49263 5 1 1 49262
0 49264 7 1 2 95846 78938
0 49265 5 2 1 49264
0 49266 7 1 2 97543 106013
0 49267 5 1 1 49266
0 49268 7 1 2 79425 95847
0 49269 5 2 1 49268
0 49270 7 1 2 80554 106015
0 49271 5 1 1 49270
0 49272 7 1 2 49267 49271
0 49273 7 1 2 49263 49272
0 49274 5 1 1 49273
0 49275 7 1 2 67786 49274
0 49276 5 1 1 49275
0 49277 7 1 2 97944 105199
0 49278 5 1 1 49277
0 49279 7 1 2 49276 49278
0 49280 5 2 1 49279
0 49281 7 1 2 75183 106017
0 49282 5 1 1 49281
0 49283 7 1 2 86530 76014
0 49284 7 1 2 84516 49283
0 49285 5 1 1 49284
0 49286 7 1 2 49282 49285
0 49287 5 1 1 49286
0 49288 7 1 2 85550 49287
0 49289 5 1 1 49288
0 49290 7 1 2 100547 96023
0 49291 5 1 1 49290
0 49292 7 2 2 64199 84300
0 49293 7 2 2 68509 106019
0 49294 5 1 1 106021
0 49295 7 1 2 49291 49294
0 49296 5 1 1 49295
0 49297 7 1 2 81777 49296
0 49298 5 1 1 49297
0 49299 7 1 2 31357 106020
0 49300 5 1 1 49299
0 49301 7 1 2 49298 49300
0 49302 5 1 1 49301
0 49303 7 1 2 65194 49302
0 49304 5 1 1 49303
0 49305 7 1 2 67787 87040
0 49306 5 1 1 49305
0 49307 7 1 2 87824 49306
0 49308 5 1 1 49307
0 49309 7 1 2 69988 49308
0 49310 5 1 1 49309
0 49311 7 1 2 84260 82145
0 49312 5 1 1 49311
0 49313 7 1 2 49310 49312
0 49314 5 1 1 49313
0 49315 7 1 2 64200 85757
0 49316 7 1 2 49314 49315
0 49317 5 1 1 49316
0 49318 7 1 2 49304 49317
0 49319 5 1 1 49318
0 49320 7 2 2 94831 49319
0 49321 7 1 2 78078 106023
0 49322 5 1 1 49321
0 49323 7 1 2 87817 92642
0 49324 5 1 1 49323
0 49325 7 1 2 85657 49324
0 49326 5 1 1 49325
0 49327 7 1 2 69989 104958
0 49328 5 1 1 49327
0 49329 7 1 2 49326 49328
0 49330 5 1 1 49329
0 49331 7 2 2 94832 49330
0 49332 7 1 2 97493 106025
0 49333 5 1 1 49332
0 49334 7 1 2 80747 101129
0 49335 5 1 1 49334
0 49336 7 1 2 68720 104502
0 49337 5 1 1 49336
0 49338 7 1 2 49335 49337
0 49339 5 1 1 49338
0 49340 7 1 2 102055 49339
0 49341 5 1 1 49340
0 49342 7 1 2 92673 76755
0 49343 7 1 2 104507 49342
0 49344 5 1 1 49343
0 49345 7 1 2 49341 49344
0 49346 5 1 1 49345
0 49347 7 2 2 72185 49346
0 49348 7 1 2 75159 106027
0 49349 5 1 1 49348
0 49350 7 1 2 49333 49349
0 49351 5 1 1 49350
0 49352 7 1 2 75453 49351
0 49353 5 1 1 49352
0 49354 7 1 2 49322 49353
0 49355 7 1 2 49289 49354
0 49356 5 1 1 49355
0 49357 7 1 2 67426 49356
0 49358 5 1 1 49357
0 49359 7 1 2 101130 105474
0 49360 7 2 2 105596 49359
0 49361 7 2 2 70643 93103
0 49362 7 1 2 106029 106031
0 49363 5 1 1 49362
0 49364 7 2 2 64869 74744
0 49365 5 1 1 106033
0 49366 7 1 2 106012 49365
0 49367 5 1 1 49366
0 49368 7 1 2 80381 49367
0 49369 5 1 1 49368
0 49370 7 1 2 74800 86654
0 49371 5 1 1 49370
0 49372 7 1 2 88799 83800
0 49373 5 1 1 49372
0 49374 7 1 2 49371 49373
0 49375 7 1 2 49369 49374
0 49376 5 1 1 49375
0 49377 7 1 2 70529 49376
0 49378 5 1 1 49377
0 49379 7 1 2 86758 106014
0 49380 5 1 1 49379
0 49381 7 1 2 49378 49380
0 49382 5 1 1 49381
0 49383 7 1 2 67788 49382
0 49384 5 1 1 49383
0 49385 7 1 2 104222 105200
0 49386 5 1 1 49385
0 49387 7 1 2 49384 49386
0 49388 5 2 1 49387
0 49389 7 1 2 75184 106035
0 49390 5 1 1 49389
0 49391 7 2 2 76006 86010
0 49392 7 1 2 90241 106037
0 49393 5 1 1 49392
0 49394 7 1 2 49390 49393
0 49395 5 1 1 49394
0 49396 7 1 2 99393 49395
0 49397 5 1 1 49396
0 49398 7 1 2 49363 49397
0 49399 7 1 2 49358 49398
0 49400 5 1 1 49399
0 49401 7 1 2 81063 49400
0 49402 5 1 1 49401
0 49403 7 1 2 101399 92643
0 49404 5 2 1 49403
0 49405 7 1 2 104574 75185
0 49406 5 1 1 49405
0 49407 7 1 2 82844 89356
0 49408 7 1 2 78079 49407
0 49409 7 1 2 80064 49408
0 49410 5 1 1 49409
0 49411 7 1 2 49406 49410
0 49412 5 1 1 49411
0 49413 7 1 2 83031 49412
0 49414 5 1 1 49413
0 49415 7 1 2 10577 104982
0 49416 5 1 1 49415
0 49417 7 2 2 94513 49416
0 49418 7 1 2 76015 106041
0 49419 5 1 1 49418
0 49420 7 1 2 49414 49419
0 49421 5 1 1 49420
0 49422 7 1 2 64201 49421
0 49423 5 1 1 49422
0 49424 7 2 2 83297 89357
0 49425 7 1 2 84967 106043
0 49426 7 1 2 105971 49425
0 49427 5 1 1 49426
0 49428 7 1 2 49423 49427
0 49429 5 1 1 49428
0 49430 7 1 2 67427 49429
0 49431 5 1 1 49430
0 49432 7 1 2 100551 90982
0 49433 7 2 2 104575 49432
0 49434 7 2 2 94782 89143
0 49435 7 1 2 106045 106047
0 49436 5 1 1 49435
0 49437 7 1 2 49431 49436
0 49438 5 1 1 49437
0 49439 7 1 2 70895 49438
0 49440 5 1 1 49439
0 49441 7 1 2 75454 80205
0 49442 7 1 2 102748 49441
0 49443 7 2 2 104576 49442
0 49444 7 1 2 106049 106048
0 49445 5 1 1 49444
0 49446 7 1 2 49440 49445
0 49447 5 1 1 49446
0 49448 7 1 2 106039 49447
0 49449 5 1 1 49448
0 49450 7 1 2 84308 10766
0 49451 5 1 1 49450
0 49452 7 1 2 23435 79426
0 49453 7 2 2 49451 49452
0 49454 7 1 2 81778 104984
0 49455 5 1 1 49454
0 49456 7 1 2 82862 49455
0 49457 5 1 1 49456
0 49458 7 1 2 66077 49457
0 49459 5 1 1 49458
0 49460 7 1 2 85749 78387
0 49461 5 1 1 49460
0 49462 7 1 2 49459 49461
0 49463 5 1 1 49462
0 49464 7 1 2 67428 94833
0 49465 7 2 2 49463 49464
0 49466 5 1 1 106053
0 49467 7 1 2 78080 106054
0 49468 5 1 1 49467
0 49469 7 1 2 99454 97827
0 49470 7 1 2 104706 49469
0 49471 5 1 1 49470
0 49472 7 1 2 97925 30320
0 49473 5 1 1 49472
0 49474 7 1 2 77193 49473
0 49475 5 1 1 49474
0 49476 7 1 2 103597 49475
0 49477 5 1 1 49476
0 49478 7 1 2 78022 80237
0 49479 7 1 2 49477 49478
0 49480 5 1 1 49479
0 49481 7 1 2 49471 49480
0 49482 5 1 1 49481
0 49483 7 2 2 72186 49482
0 49484 5 1 1 106055
0 49485 7 1 2 75160 106056
0 49486 5 1 1 49485
0 49487 7 1 2 49468 49486
0 49488 5 1 1 49487
0 49489 7 1 2 106051 49488
0 49490 5 1 1 49489
0 49491 7 1 2 49449 49490
0 49492 7 1 2 49402 49491
0 49493 7 1 2 49248 49492
0 49494 7 1 2 49144 49493
0 49495 5 1 1 49494
0 49496 7 1 2 71474 49495
0 49497 5 1 1 49496
0 49498 7 1 2 68510 96457
0 49499 5 1 1 49498
0 49500 7 1 2 104485 49499
0 49501 5 1 1 49500
0 49502 7 2 2 84380 49501
0 49503 5 1 1 106057
0 49504 7 1 2 75161 106058
0 49505 5 1 1 49504
0 49506 7 1 2 95907 76126
0 49507 5 1 1 49506
0 49508 7 1 2 77755 106038
0 49509 5 2 1 49508
0 49510 7 1 2 49507 106059
0 49511 5 1 1 49510
0 49512 7 1 2 73578 49511
0 49513 5 1 1 49512
0 49514 7 1 2 49505 49513
0 49515 5 1 1 49514
0 49516 7 1 2 85551 49515
0 49517 5 1 1 49516
0 49518 7 2 2 67137 87483
0 49519 7 2 2 103202 106061
0 49520 7 1 2 97494 106063
0 49521 5 1 1 49520
0 49522 7 1 2 49517 49521
0 49523 5 1 1 49522
0 49524 7 1 2 92895 49523
0 49525 5 1 1 49524
0 49526 7 2 2 97592 84649
0 49527 7 1 2 73241 99900
0 49528 7 1 2 106065 49527
0 49529 5 1 1 49528
0 49530 7 1 2 106060 49529
0 49531 5 1 1 49530
0 49532 7 1 2 73579 49531
0 49533 5 1 1 49532
0 49534 7 1 2 87484 78095
0 49535 5 1 1 49534
0 49536 7 1 2 70644 77734
0 49537 7 1 2 77502 49536
0 49538 7 1 2 104168 49537
0 49539 5 1 1 49538
0 49540 7 1 2 49535 49539
0 49541 5 1 1 49540
0 49542 7 1 2 73242 49541
0 49543 5 1 1 49542
0 49544 7 1 2 49533 49543
0 49545 5 1 1 49544
0 49546 7 1 2 101020 49545
0 49547 5 1 1 49546
0 49548 7 2 2 82611 83114
0 49549 5 2 1 106067
0 49550 7 1 2 96825 106069
0 49551 5 1 1 49550
0 49552 7 2 2 68721 98204
0 49553 7 2 2 49551 106071
0 49554 7 2 2 84326 95563
0 49555 7 1 2 106073 106075
0 49556 5 1 1 49555
0 49557 7 1 2 49547 49556
0 49558 5 1 1 49557
0 49559 7 1 2 70896 49558
0 49560 5 1 1 49559
0 49561 7 2 2 95641 74077
0 49562 7 1 2 77510 105984
0 49563 5 1 1 49562
0 49564 7 2 2 74801 106066
0 49565 5 1 1 106079
0 49566 7 1 2 49563 49565
0 49567 5 1 1 49566
0 49568 7 1 2 65499 49567
0 49569 5 1 1 49568
0 49570 7 1 2 73243 105988
0 49571 5 1 1 49570
0 49572 7 1 2 49569 49571
0 49573 5 1 1 49572
0 49574 7 1 2 68722 49573
0 49575 5 1 1 49574
0 49576 7 1 2 82710 105979
0 49577 5 1 1 49576
0 49578 7 1 2 49575 49577
0 49579 5 1 1 49578
0 49580 7 1 2 106077 49579
0 49581 5 1 1 49580
0 49582 7 1 2 49560 49581
0 49583 5 1 1 49582
0 49584 7 1 2 72777 49583
0 49585 5 1 1 49584
0 49586 7 1 2 49525 49585
0 49587 5 1 1 49586
0 49588 7 1 2 67429 49587
0 49589 5 1 1 49588
0 49590 7 1 2 92896 105899
0 49591 5 1 1 49590
0 49592 7 1 2 68511 95317
0 49593 7 1 2 103719 49592
0 49594 5 1 1 49593
0 49595 7 1 2 49591 49594
0 49596 5 2 1 49595
0 49597 7 1 2 75186 106081
0 49598 5 1 1 49597
0 49599 7 2 2 65612 89128
0 49600 7 2 2 98205 106083
0 49601 7 1 2 105073 106085
0 49602 5 1 1 49601
0 49603 7 1 2 49598 49602
0 49604 5 1 1 49603
0 49605 7 1 2 71701 49604
0 49606 5 1 1 49605
0 49607 7 2 2 71180 105458
0 49608 7 1 2 106087 106084
0 49609 5 1 1 49608
0 49610 7 1 2 49606 49609
0 49611 5 1 1 49610
0 49612 7 1 2 103203 49611
0 49613 5 1 1 49612
0 49614 7 1 2 80206 98206
0 49615 7 1 2 76979 49614
0 49616 7 2 2 69008 96728
0 49617 7 1 2 92956 106089
0 49618 7 1 2 49615 49617
0 49619 5 1 1 49618
0 49620 7 1 2 49613 49619
0 49621 5 1 1 49620
0 49622 7 1 2 96923 49621
0 49623 5 1 1 49622
0 49624 7 1 2 49589 49623
0 49625 5 1 1 49624
0 49626 7 1 2 70264 49625
0 49627 5 1 1 49626
0 49628 7 1 2 84860 97571
0 49629 5 1 1 49628
0 49630 7 1 2 105982 49629
0 49631 5 1 1 49630
0 49632 7 1 2 85467 49631
0 49633 5 1 1 49632
0 49634 7 2 2 88767 95651
0 49635 7 1 2 106091 106032
0 49636 5 1 1 49635
0 49637 7 1 2 49633 49636
0 49638 5 1 1 49637
0 49639 7 1 2 74802 49638
0 49640 5 1 1 49639
0 49641 7 1 2 99424 91610
0 49642 7 1 2 97495 49641
0 49643 5 1 1 49642
0 49644 7 1 2 49640 49643
0 49645 5 1 1 49644
0 49646 7 1 2 100419 49645
0 49647 5 1 1 49646
0 49648 7 1 2 84343 83911
0 49649 7 1 2 104683 49648
0 49650 7 1 2 97597 49649
0 49651 5 1 1 49650
0 49652 7 1 2 49647 49651
0 49653 5 1 1 49652
0 49654 7 1 2 92897 49653
0 49655 5 1 1 49654
0 49656 7 1 2 74745 97598
0 49657 5 1 1 49656
0 49658 7 1 2 68723 106080
0 49659 5 1 1 49658
0 49660 7 1 2 49657 49659
0 49661 5 1 1 49660
0 49662 7 1 2 65500 49661
0 49663 5 1 1 49662
0 49664 7 1 2 86631 78096
0 49665 5 1 1 49664
0 49666 7 1 2 49663 49665
0 49667 5 1 1 49666
0 49668 7 1 2 101021 49667
0 49669 5 1 1 49668
0 49670 7 2 2 96822 106072
0 49671 7 1 2 106093 106076
0 49672 5 1 1 49671
0 49673 7 1 2 49669 49672
0 49674 5 1 1 49673
0 49675 7 1 2 70897 49674
0 49676 5 1 1 49675
0 49677 7 1 2 105977 49676
0 49678 5 1 1 49677
0 49679 7 1 2 67430 49678
0 49680 5 1 1 49679
0 49681 7 1 2 105973 49680
0 49682 5 1 1 49681
0 49683 7 1 2 71702 49682
0 49684 5 1 1 49683
0 49685 7 1 2 86974 96679
0 49686 5 2 1 49685
0 49687 7 1 2 85468 106095
0 49688 5 1 1 49687
0 49689 7 1 2 91955 103515
0 49690 5 1 1 49689
0 49691 7 1 2 49688 49690
0 49692 5 1 1 49691
0 49693 7 2 2 97209 49692
0 49694 7 1 2 106097 106086
0 49695 5 1 1 49694
0 49696 7 1 2 49684 49695
0 49697 5 1 1 49696
0 49698 7 1 2 72778 49697
0 49699 5 1 1 49698
0 49700 7 1 2 49655 49699
0 49701 7 1 2 49627 49700
0 49702 5 1 1 49701
0 49703 7 1 2 69990 49702
0 49704 5 1 1 49703
0 49705 7 1 2 94220 89780
0 49706 5 2 1 49705
0 49707 7 1 2 86472 106099
0 49708 5 1 1 49707
0 49709 7 1 2 80033 104791
0 49710 5 1 1 49709
0 49711 7 1 2 103877 83760
0 49712 5 1 1 49711
0 49713 7 1 2 49710 49712
0 49714 5 1 1 49713
0 49715 7 1 2 49708 49714
0 49716 5 1 1 49715
0 49717 7 1 2 77091 96869
0 49718 7 1 2 99142 49717
0 49719 7 1 2 106096 49718
0 49720 5 1 1 49719
0 49721 7 1 2 49716 49720
0 49722 5 2 1 49721
0 49723 7 1 2 78097 106101
0 49724 5 1 1 49723
0 49725 7 1 2 101022 98917
0 49726 5 1 1 49725
0 49727 7 1 2 69277 87189
0 49728 7 1 2 98544 49727
0 49729 5 1 1 49728
0 49730 7 1 2 49726 49729
0 49731 5 1 1 49730
0 49732 7 1 2 68512 49731
0 49733 5 1 1 49732
0 49734 7 1 2 69278 86838
0 49735 7 1 2 105613 49734
0 49736 5 1 1 49735
0 49737 7 1 2 49733 49736
0 49738 5 1 1 49737
0 49739 7 2 2 95005 49738
0 49740 7 1 2 92065 94140
0 49741 7 1 2 106103 49740
0 49742 5 1 1 49741
0 49743 7 1 2 49724 49742
0 49744 5 1 1 49743
0 49745 7 1 2 67431 49744
0 49746 5 1 1 49745
0 49747 7 1 2 87808 92368
0 49748 7 1 2 98628 49747
0 49749 7 2 2 105900 49748
0 49750 7 1 2 84359 89868
0 49751 7 1 2 86508 49750
0 49752 7 1 2 106105 49751
0 49753 5 1 1 49752
0 49754 7 1 2 49746 49753
0 49755 5 1 1 49754
0 49756 7 1 2 70898 49755
0 49757 5 1 1 49756
0 49758 7 2 2 67432 74078
0 49759 7 2 2 95642 106107
0 49760 7 1 2 87897 89758
0 49761 7 1 2 76790 49760
0 49762 7 1 2 96636 49761
0 49763 5 1 1 49762
0 49764 7 1 2 103105 75187
0 49765 5 1 1 49764
0 49766 7 2 2 86899 89358
0 49767 7 1 2 76138 106111
0 49768 5 1 1 49767
0 49769 7 1 2 49765 49768
0 49770 5 1 1 49769
0 49771 7 2 2 67789 75291
0 49772 7 1 2 64870 106113
0 49773 7 1 2 49770 49772
0 49774 5 1 1 49773
0 49775 7 1 2 49763 49774
0 49776 5 1 1 49775
0 49777 7 1 2 106109 49776
0 49778 5 1 1 49777
0 49779 7 1 2 49757 49778
0 49780 7 1 2 49704 49779
0 49781 7 1 2 49497 49780
0 49782 5 1 1 49781
0 49783 7 1 2 73872 49782
0 49784 5 1 1 49783
0 49785 7 1 2 69009 95643
0 49786 7 1 2 105966 49785
0 49787 5 1 1 49786
0 49788 7 1 2 63922 48952
0 49789 5 1 1 49788
0 49790 7 1 2 69010 48976
0 49791 5 1 1 49790
0 49792 7 1 2 67433 49791
0 49793 7 1 2 49789 49792
0 49794 5 1 1 49793
0 49795 7 1 2 49787 49794
0 49796 5 1 1 49795
0 49797 7 1 2 68159 49796
0 49798 5 1 1 49797
0 49799 7 1 2 94754 88237
0 49800 5 1 1 49799
0 49801 7 1 2 88827 92616
0 49802 5 1 1 49801
0 49803 7 1 2 49800 49802
0 49804 5 1 1 49803
0 49805 7 1 2 105975 49804
0 49806 5 2 1 49805
0 49807 7 1 2 104634 92617
0 49808 5 1 1 49807
0 49809 7 1 2 89701 49808
0 49810 5 1 1 49809
0 49811 7 1 2 68513 49810
0 49812 5 1 1 49811
0 49813 7 1 2 87190 90956
0 49814 5 1 1 49813
0 49815 7 1 2 49812 49814
0 49816 5 1 1 49815
0 49817 7 1 2 73244 49816
0 49818 5 1 1 49817
0 49819 7 1 2 95070 89365
0 49820 5 1 1 49819
0 49821 7 1 2 49818 49820
0 49822 5 1 1 49821
0 49823 7 1 2 101023 49822
0 49824 5 1 1 49823
0 49825 7 2 2 85643 88238
0 49826 5 2 1 106117
0 49827 7 1 2 101588 88593
0 49828 5 1 1 49827
0 49829 7 1 2 106119 49828
0 49830 5 1 1 49829
0 49831 7 1 2 49830 105986
0 49832 5 1 1 49831
0 49833 7 1 2 49824 49832
0 49834 5 1 1 49833
0 49835 7 1 2 70899 49834
0 49836 5 1 1 49835
0 49837 7 1 2 106115 49836
0 49838 5 1 1 49837
0 49839 7 1 2 67434 49838
0 49840 5 1 1 49839
0 49841 7 1 2 93104 105968
0 49842 5 2 1 49841
0 49843 7 1 2 49840 106121
0 49844 5 1 1 49843
0 49845 7 1 2 75455 49844
0 49846 5 1 1 49845
0 49847 7 1 2 95007 105996
0 49848 5 1 1 49847
0 49849 7 1 2 72187 83013
0 49850 5 1 1 49849
0 49851 7 1 2 68514 89296
0 49852 7 1 2 49850 49851
0 49853 5 1 1 49852
0 49854 7 1 2 89702 49853
0 49855 5 1 1 49854
0 49856 7 1 2 76667 49855
0 49857 5 1 1 49856
0 49858 7 1 2 89810 105990
0 49859 5 1 1 49858
0 49860 7 1 2 49857 49859
0 49861 5 1 1 49860
0 49862 7 1 2 101024 49861
0 49863 5 1 1 49862
0 49864 7 1 2 90615 105992
0 49865 5 1 1 49864
0 49866 7 1 2 49863 49865
0 49867 5 1 1 49866
0 49868 7 1 2 67435 49867
0 49869 5 1 1 49868
0 49870 7 1 2 87339 77735
0 49871 7 1 2 87601 49870
0 49872 5 1 1 49871
0 49873 7 1 2 86075 93304
0 49874 5 1 1 49873
0 49875 7 1 2 49872 49874
0 49876 5 1 1 49875
0 49877 7 1 2 104946 49876
0 49878 5 1 1 49877
0 49879 7 1 2 49869 49878
0 49880 5 1 1 49879
0 49881 7 1 2 70900 49880
0 49882 5 1 1 49881
0 49883 7 1 2 93105 105994
0 49884 5 1 1 49883
0 49885 7 1 2 49882 49884
0 49886 5 1 1 49885
0 49887 7 1 2 73245 49886
0 49888 5 1 1 49887
0 49889 7 1 2 49848 49888
0 49890 7 1 2 49846 49889
0 49891 7 1 2 49798 49890
0 49892 5 1 1 49891
0 49893 7 1 2 72779 49892
0 49894 5 1 1 49893
0 49895 7 1 2 88594 106000
0 49896 5 1 1 49895
0 49897 7 1 2 104230 93431
0 49898 5 1 1 49897
0 49899 7 1 2 49896 49898
0 49900 5 1 1 49899
0 49901 7 1 2 77194 49900
0 49902 5 1 1 49901
0 49903 7 1 2 92071 106002
0 49904 5 1 1 49903
0 49905 7 1 2 49902 49904
0 49906 5 1 1 49905
0 49907 7 1 2 69279 49906
0 49908 5 1 1 49907
0 49909 7 1 2 84327 100932
0 49910 7 1 2 106004 49909
0 49911 5 1 1 49910
0 49912 7 1 2 72476 49911
0 49913 7 1 2 49908 49912
0 49914 5 1 1 49913
0 49915 7 1 2 63923 106008
0 49916 5 1 1 49915
0 49917 7 1 2 88595 106010
0 49918 5 1 1 49917
0 49919 7 1 2 67436 49918
0 49920 7 1 2 49916 49919
0 49921 5 1 1 49920
0 49922 7 1 2 67790 49921
0 49923 7 1 2 49914 49922
0 49924 5 1 1 49923
0 49925 7 1 2 88596 106018
0 49926 5 1 1 49925
0 49927 7 1 2 75808 93175
0 49928 7 1 2 86968 49927
0 49929 5 1 1 49928
0 49930 7 1 2 49926 49929
0 49931 5 1 1 49930
0 49932 7 1 2 85552 49931
0 49933 5 1 1 49932
0 49934 7 1 2 63924 106024
0 49935 5 1 1 49934
0 49936 7 1 2 84235 106026
0 49937 5 1 1 49936
0 49938 7 1 2 69011 106028
0 49939 5 1 1 49938
0 49940 7 1 2 49937 49939
0 49941 5 1 1 49940
0 49942 7 1 2 75456 49941
0 49943 5 1 1 49942
0 49944 7 1 2 49935 49943
0 49945 7 1 2 49933 49944
0 49946 5 1 1 49945
0 49947 7 1 2 67437 49946
0 49948 5 1 1 49947
0 49949 7 1 2 93735 106030
0 49950 5 1 1 49949
0 49951 7 1 2 104959 90846
0 49952 5 1 1 49951
0 49953 7 1 2 88597 106036
0 49954 5 1 1 49953
0 49955 7 1 2 49952 49954
0 49956 5 1 1 49955
0 49957 7 1 2 99394 49956
0 49958 5 1 1 49957
0 49959 7 1 2 49950 49958
0 49960 7 1 2 49948 49959
0 49961 5 1 1 49960
0 49962 7 1 2 81064 49961
0 49963 5 1 1 49962
0 49964 7 1 2 80065 94702
0 49965 5 1 1 49964
0 49966 7 1 2 81065 92701
0 49967 5 1 1 49966
0 49968 7 1 2 49965 49967
0 49969 5 1 1 49968
0 49970 7 1 2 70265 49969
0 49971 5 1 1 49970
0 49972 7 1 2 104577 90964
0 49973 5 1 1 49972
0 49974 7 1 2 49971 49973
0 49975 5 1 1 49974
0 49976 7 1 2 80649 49975
0 49977 5 1 1 49976
0 49978 7 1 2 89990 106042
0 49979 5 1 1 49978
0 49980 7 1 2 49977 49979
0 49981 5 1 1 49980
0 49982 7 1 2 64202 49981
0 49983 5 1 1 49982
0 49984 7 2 2 84968 93106
0 49985 7 1 2 106044 106123
0 49986 5 1 1 49985
0 49987 7 1 2 49983 49986
0 49988 5 1 1 49987
0 49989 7 1 2 67438 49988
0 49990 5 1 1 49989
0 49991 7 2 2 70530 93736
0 49992 7 1 2 106125 106046
0 49993 5 1 1 49992
0 49994 7 1 2 49990 49993
0 49995 5 1 1 49994
0 49996 7 1 2 70901 49995
0 49997 5 1 1 49996
0 49998 7 1 2 106126 106050
0 49999 5 1 1 49998
0 50000 7 1 2 49997 49999
0 50001 5 1 1 50000
0 50002 7 1 2 106040 50001
0 50003 5 1 1 50002
0 50004 7 1 2 63925 49466
0 50005 5 1 1 50004
0 50006 7 1 2 69012 49484
0 50007 5 1 1 50006
0 50008 7 1 2 106052 50007
0 50009 7 1 2 50005 50008
0 50010 5 1 1 50009
0 50011 7 1 2 50003 50010
0 50012 7 1 2 49963 50011
0 50013 7 1 2 49924 50012
0 50014 7 1 2 49894 50013
0 50015 5 1 1 50014
0 50016 7 1 2 71475 50015
0 50017 5 1 1 50016
0 50018 7 1 2 84236 106064
0 50019 5 1 1 50018
0 50020 7 1 2 73580 104519
0 50021 5 1 1 50020
0 50022 7 1 2 49503 50021
0 50023 5 1 1 50022
0 50024 7 1 2 69013 50023
0 50025 5 1 1 50024
0 50026 7 1 2 83488 95974
0 50027 5 1 1 50026
0 50028 7 1 2 50025 50027
0 50029 5 1 1 50028
0 50030 7 1 2 85553 50029
0 50031 5 1 1 50030
0 50032 7 1 2 50019 50031
0 50033 5 1 1 50032
0 50034 7 1 2 92898 50033
0 50035 5 1 1 50034
0 50036 7 1 2 104517 96045
0 50037 5 1 1 50036
0 50038 7 1 2 75648 95975
0 50039 5 1 1 50038
0 50040 7 1 2 50037 50039
0 50041 5 1 1 50040
0 50042 7 1 2 73581 50041
0 50043 5 1 1 50042
0 50044 7 1 2 79200 88598
0 50045 7 1 2 104169 50044
0 50046 5 1 1 50045
0 50047 7 1 2 63926 106062
0 50048 5 1 1 50047
0 50049 7 1 2 50046 50048
0 50050 5 1 1 50049
0 50051 7 1 2 73246 50050
0 50052 5 1 1 50051
0 50053 7 1 2 50043 50052
0 50054 5 1 1 50053
0 50055 7 1 2 101025 50054
0 50056 5 1 1 50055
0 50057 7 3 2 69627 84237
0 50058 7 1 2 106074 106127
0 50059 5 1 1 50058
0 50060 7 1 2 50056 50059
0 50061 5 1 1 50060
0 50062 7 1 2 70902 50061
0 50063 5 1 1 50062
0 50064 7 1 2 82612 90641
0 50065 5 1 1 50064
0 50066 7 1 2 74803 89719
0 50067 5 1 1 50066
0 50068 7 1 2 50065 50067
0 50069 5 1 1 50068
0 50070 7 1 2 65501 50069
0 50071 5 1 1 50070
0 50072 7 1 2 73247 106118
0 50073 5 1 1 50072
0 50074 7 1 2 50071 50073
0 50075 5 1 1 50074
0 50076 7 1 2 68724 50075
0 50077 5 1 1 50076
0 50078 7 1 2 87216 92684
0 50079 5 1 1 50078
0 50080 7 1 2 50077 50079
0 50081 5 1 1 50080
0 50082 7 1 2 50081 106078
0 50083 5 1 1 50082
0 50084 7 1 2 50063 50083
0 50085 5 1 1 50084
0 50086 7 1 2 72780 50085
0 50087 5 1 1 50086
0 50088 7 1 2 50035 50087
0 50089 5 1 1 50088
0 50090 7 1 2 67439 50089
0 50091 5 1 1 50090
0 50092 7 1 2 88599 106082
0 50093 5 1 1 50092
0 50094 7 1 2 93185 105074
0 50095 5 1 1 50094
0 50096 7 1 2 50093 50095
0 50097 5 1 1 50096
0 50098 7 1 2 71703 50097
0 50099 5 1 1 50098
0 50100 7 1 2 89869 106088
0 50101 5 1 1 50100
0 50102 7 1 2 50099 50101
0 50103 5 1 1 50102
0 50104 7 1 2 103204 50103
0 50105 5 1 1 50104
0 50106 7 1 2 77527 89763
0 50107 7 1 2 98623 105424
0 50108 7 1 2 50106 50107
0 50109 5 1 1 50108
0 50110 7 1 2 50105 50109
0 50111 5 1 1 50110
0 50112 7 1 2 96924 50111
0 50113 5 1 1 50112
0 50114 7 1 2 50091 50113
0 50115 5 1 1 50114
0 50116 7 1 2 70266 50115
0 50117 5 1 1 50116
0 50118 7 1 2 89703 90023
0 50119 5 1 1 50118
0 50120 7 1 2 85469 50119
0 50121 5 1 1 50120
0 50122 7 1 2 93737 106092
0 50123 5 1 1 50122
0 50124 7 1 2 50121 50123
0 50125 5 1 1 50124
0 50126 7 1 2 74804 50125
0 50127 5 1 1 50126
0 50128 7 1 2 85470 77503
0 50129 7 1 2 106112 50128
0 50130 5 1 1 50129
0 50131 7 1 2 50127 50130
0 50132 5 1 1 50131
0 50133 7 1 2 100420 50132
0 50134 5 1 1 50133
0 50135 7 5 2 93107 97480
0 50136 5 1 1 106130
0 50137 7 1 2 74746 100119
0 50138 7 1 2 106131 50137
0 50139 5 1 1 50138
0 50140 7 1 2 50134 50139
0 50141 5 1 1 50140
0 50142 7 1 2 92899 50141
0 50143 5 1 1 50142
0 50144 7 1 2 76791 89731
0 50145 5 1 1 50144
0 50146 7 1 2 93847 91611
0 50147 5 1 1 50146
0 50148 7 1 2 50145 50147
0 50149 5 1 1 50148
0 50150 7 1 2 65502 50149
0 50151 5 1 1 50150
0 50152 7 1 2 81928 98654
0 50153 5 1 1 50152
0 50154 7 1 2 50151 50153
0 50155 5 1 1 50154
0 50156 7 1 2 101026 50155
0 50157 5 1 1 50156
0 50158 7 1 2 106128 106094
0 50159 5 1 1 50158
0 50160 7 1 2 50157 50159
0 50161 5 1 1 50160
0 50162 7 1 2 70903 50161
0 50163 5 1 1 50162
0 50164 7 1 2 106116 50163
0 50165 5 1 1 50164
0 50166 7 1 2 67440 50165
0 50167 5 1 1 50166
0 50168 7 1 2 106122 50167
0 50169 5 1 1 50168
0 50170 7 1 2 71704 50169
0 50171 5 1 1 50170
0 50172 7 1 2 93186 106098
0 50173 5 1 1 50172
0 50174 7 1 2 50171 50173
0 50175 5 1 1 50174
0 50176 7 1 2 72781 50175
0 50177 5 1 1 50176
0 50178 7 1 2 50143 50177
0 50179 7 1 2 50117 50178
0 50180 5 1 1 50179
0 50181 7 1 2 69991 50180
0 50182 5 1 1 50181
0 50183 7 1 2 96016 106104
0 50184 5 1 1 50183
0 50185 7 1 2 88239 106102
0 50186 5 1 1 50185
0 50187 7 1 2 50184 50186
0 50188 5 1 1 50187
0 50189 7 1 2 67441 50188
0 50190 5 1 1 50189
0 50191 7 1 2 77833 104389
0 50192 7 1 2 106106 50191
0 50193 5 1 1 50192
0 50194 7 1 2 50190 50193
0 50195 5 1 1 50194
0 50196 7 1 2 70904 50195
0 50197 5 1 1 50196
0 50198 7 1 2 103406 105882
0 50199 5 1 1 50198
0 50200 7 1 2 79740 81424
0 50201 7 1 2 102441 50200
0 50202 5 1 1 50201
0 50203 7 1 2 50199 50202
0 50204 5 1 1 50203
0 50205 7 1 2 88240 50204
0 50206 5 1 1 50205
0 50207 7 1 2 103410 90560
0 50208 7 1 2 103106 50207
0 50209 5 1 1 50208
0 50210 7 1 2 50206 50209
0 50211 5 1 1 50210
0 50212 7 1 2 106110 50211
0 50213 5 1 1 50212
0 50214 7 1 2 50197 50213
0 50215 7 1 2 50182 50214
0 50216 7 1 2 50017 50215
0 50217 5 1 1 50216
0 50218 7 1 2 89585 50217
0 50219 5 1 1 50218
0 50220 7 2 2 85658 82032
0 50221 5 1 1 106135
0 50222 7 1 2 66595 103728
0 50223 5 1 1 50222
0 50224 7 1 2 70267 96682
0 50225 7 1 2 50223 50224
0 50226 5 1 1 50225
0 50227 7 1 2 37337 50226
0 50228 5 1 1 50227
0 50229 7 1 2 68725 50228
0 50230 5 1 1 50229
0 50231 7 1 2 50221 50230
0 50232 5 1 1 50231
0 50233 7 1 2 69992 50232
0 50234 5 1 1 50233
0 50235 7 1 2 104219 50234
0 50236 5 1 1 50235
0 50237 7 1 2 101009 50236
0 50238 5 1 1 50237
0 50239 7 1 2 89213 13896
0 50240 5 1 1 50239
0 50241 7 1 2 68160 50240
0 50242 5 1 1 50241
0 50243 7 1 2 69993 97603
0 50244 5 1 1 50243
0 50245 7 1 2 50242 50244
0 50246 5 1 1 50245
0 50247 7 1 2 73582 50246
0 50248 5 1 1 50247
0 50249 7 1 2 78939 95913
0 50250 5 1 1 50249
0 50251 7 1 2 81929 50250
0 50252 5 1 1 50251
0 50253 7 1 2 99011 50252
0 50254 7 1 2 50248 50253
0 50255 5 1 1 50254
0 50256 7 1 2 81066 50255
0 50257 5 1 1 50256
0 50258 7 1 2 82637 87085
0 50259 5 1 1 50258
0 50260 7 1 2 2101 50259
0 50261 5 1 1 50260
0 50262 7 1 2 101131 50261
0 50263 5 1 1 50262
0 50264 7 1 2 101161 101769
0 50265 5 1 1 50264
0 50266 7 1 2 103456 105487
0 50267 5 1 1 50266
0 50268 7 1 2 50265 50267
0 50269 7 1 2 50263 50268
0 50270 5 1 1 50269
0 50271 7 1 2 68726 50270
0 50272 5 1 1 50271
0 50273 7 1 2 81067 106016
0 50274 5 1 1 50273
0 50275 7 1 2 93506 105018
0 50276 5 1 1 50275
0 50277 7 1 2 50274 50276
0 50278 5 1 1 50277
0 50279 7 1 2 82655 50278
0 50280 5 1 1 50279
0 50281 7 1 2 101308 104392
0 50282 5 1 1 50281
0 50283 7 1 2 101499 106136
0 50284 5 1 1 50283
0 50285 7 1 2 50282 50284
0 50286 7 1 2 50280 50285
0 50287 7 1 2 50272 50286
0 50288 7 1 2 50257 50287
0 50289 5 1 1 50288
0 50290 7 1 2 69280 50289
0 50291 5 1 1 50290
0 50292 7 1 2 93560 76972
0 50293 7 1 2 105880 50292
0 50294 5 1 1 50293
0 50295 7 1 2 50291 50294
0 50296 7 1 2 50238 50295
0 50297 5 1 1 50296
0 50298 7 1 2 67791 50297
0 50299 5 1 1 50298
0 50300 7 1 2 81779 7127
0 50301 5 1 1 50300
0 50302 7 1 2 89214 50301
0 50303 5 1 1 50302
0 50304 7 1 2 68161 50303
0 50305 5 1 1 50304
0 50306 7 1 2 99499 50305
0 50307 5 1 1 50306
0 50308 7 1 2 73583 50307
0 50309 5 1 1 50308
0 50310 7 1 2 74908 86655
0 50311 5 1 1 50310
0 50312 7 1 2 91750 50311
0 50313 5 1 1 50312
0 50314 7 1 2 73248 50313
0 50315 5 1 1 50314
0 50316 7 1 2 50309 50315
0 50317 5 1 1 50316
0 50318 7 1 2 71181 50317
0 50319 5 1 1 50318
0 50320 7 1 2 66078 103445
0 50321 5 1 1 50320
0 50322 7 1 2 101773 50321
0 50323 5 1 1 50322
0 50324 7 1 2 69994 50323
0 50325 5 1 1 50324
0 50326 7 1 2 81930 79856
0 50327 5 2 1 50326
0 50328 7 1 2 104056 106137
0 50329 5 1 1 50328
0 50330 7 1 2 71182 50329
0 50331 5 1 1 50330
0 50332 7 1 2 102879 105557
0 50333 5 2 1 50332
0 50334 7 1 2 50331 106139
0 50335 7 1 2 50325 50334
0 50336 5 1 1 50335
0 50337 7 1 2 68162 50336
0 50338 5 1 1 50337
0 50339 7 1 2 50319 50338
0 50340 5 1 1 50339
0 50341 7 1 2 69628 50340
0 50342 5 1 1 50341
0 50343 7 1 2 64501 103446
0 50344 5 1 1 50343
0 50345 7 1 2 101774 50344
0 50346 5 1 1 50345
0 50347 7 1 2 69995 50346
0 50348 5 1 1 50347
0 50349 7 1 2 106140 50348
0 50350 5 1 1 50349
0 50351 7 1 2 98944 50350
0 50352 5 1 1 50351
0 50353 7 1 2 50342 50352
0 50354 5 1 1 50353
0 50355 7 1 2 93351 50354
0 50356 5 1 1 50355
0 50357 7 1 2 50299 50356
0 50358 5 1 1 50357
0 50359 7 1 2 71476 50358
0 50360 5 1 1 50359
0 50361 7 1 2 73249 87093
0 50362 7 1 2 86710 50361
0 50363 5 1 1 50362
0 50364 7 1 2 75649 95318
0 50365 7 1 2 99581 50364
0 50366 5 1 1 50365
0 50367 7 1 2 50363 50366
0 50368 5 1 1 50367
0 50369 7 1 2 73584 50368
0 50370 5 1 1 50369
0 50371 7 1 2 82146 105844
0 50372 5 1 1 50371
0 50373 7 1 2 72782 89956
0 50374 5 1 1 50373
0 50375 7 1 2 50372 50374
0 50376 5 1 1 50375
0 50377 7 1 2 73250 50376
0 50378 5 1 1 50377
0 50379 7 1 2 50370 50378
0 50380 5 1 1 50379
0 50381 7 1 2 77195 50380
0 50382 5 1 1 50381
0 50383 7 1 2 73251 103441
0 50384 5 1 1 50383
0 50385 7 1 2 69996 908
0 50386 7 1 2 85813 50385
0 50387 7 1 2 92900 50386
0 50388 7 1 2 50384 50387
0 50389 5 1 1 50388
0 50390 7 1 2 50382 50389
0 50391 5 1 1 50390
0 50392 7 1 2 69281 50391
0 50393 5 1 1 50392
0 50394 7 1 2 83506 77528
0 50395 7 1 2 92809 50394
0 50396 7 1 2 81633 76827
0 50397 7 1 2 50395 50396
0 50398 5 1 1 50397
0 50399 7 1 2 50393 50398
0 50400 7 1 2 50360 50399
0 50401 5 1 1 50400
0 50402 7 1 2 98049 50401
0 50403 5 1 1 50402
0 50404 7 2 2 85615 87385
0 50405 5 1 1 106141
0 50406 7 1 2 78520 106142
0 50407 5 1 1 50406
0 50408 7 1 2 86277 87191
0 50409 5 1 1 50408
0 50410 7 1 2 74694 88682
0 50411 5 1 1 50410
0 50412 7 1 2 48815 50411
0 50413 7 1 2 50409 50412
0 50414 5 1 1 50413
0 50415 7 1 2 93179 50414
0 50416 5 1 1 50415
0 50417 7 1 2 50407 50416
0 50418 5 1 1 50417
0 50419 7 1 2 76508 50418
0 50420 5 1 1 50419
0 50421 7 1 2 82083 99143
0 50422 7 1 2 105921 50421
0 50423 5 1 1 50422
0 50424 7 1 2 50420 50423
0 50425 5 1 1 50424
0 50426 7 1 2 76340 102795
0 50427 7 1 2 96386 50426
0 50428 7 1 2 50425 50427
0 50429 5 1 1 50428
0 50430 7 1 2 50403 50429
0 50431 5 1 1 50430
0 50432 7 1 2 98515 50431
0 50433 5 1 1 50432
0 50434 7 1 2 50219 50433
0 50435 7 1 2 49784 50434
0 50436 5 1 1 50435
0 50437 7 1 2 71959 50436
0 50438 5 1 1 50437
0 50439 7 1 2 75162 73873
0 50440 5 1 1 50439
0 50441 7 1 2 44419 50440
0 50442 5 1 1 50441
0 50443 7 1 2 95319 103205
0 50444 5 1 1 50443
0 50445 7 3 2 68163 82554
0 50446 7 1 2 82359 106143
0 50447 5 1 1 50446
0 50448 7 1 2 50444 50447
0 50449 5 1 1 50448
0 50450 7 1 2 69282 50449
0 50451 5 1 1 50450
0 50452 7 1 2 102355 106022
0 50453 5 1 1 50452
0 50454 7 1 2 50451 50453
0 50455 5 1 1 50454
0 50456 7 1 2 70531 50455
0 50457 5 1 1 50456
0 50458 7 1 2 72783 105302
0 50459 7 1 2 101684 50458
0 50460 5 1 1 50459
0 50461 7 1 2 50457 50460
0 50462 5 1 1 50461
0 50463 7 1 2 81068 50462
0 50464 5 1 1 50463
0 50465 7 1 2 100520 98931
0 50466 5 1 1 50465
0 50467 7 1 2 50464 50466
0 50468 5 1 1 50467
0 50469 7 1 2 67442 50468
0 50470 5 1 1 50469
0 50471 7 1 2 82360 104880
0 50472 5 1 1 50471
0 50473 7 1 2 20945 50472
0 50474 5 1 1 50473
0 50475 7 1 2 71183 50474
0 50476 5 1 1 50475
0 50477 7 1 2 76828 103796
0 50478 5 1 1 50477
0 50479 7 1 2 50476 50478
0 50480 5 1 1 50479
0 50481 7 1 2 70532 50480
0 50482 5 1 1 50481
0 50483 7 1 2 87809 76712
0 50484 7 1 2 90116 50483
0 50485 5 1 1 50484
0 50486 7 1 2 50482 50485
0 50487 5 1 1 50486
0 50488 7 1 2 69629 50487
0 50489 5 1 1 50488
0 50490 7 1 2 92957 104697
0 50491 5 1 1 50490
0 50492 7 1 2 50489 50491
0 50493 5 1 1 50492
0 50494 7 1 2 99395 50493
0 50495 5 1 1 50494
0 50496 7 1 2 50470 50495
0 50497 5 1 1 50496
0 50498 7 1 2 75457 50497
0 50499 5 1 1 50498
0 50500 7 1 2 80129 103275
0 50501 5 1 1 50500
0 50502 7 1 2 73252 90837
0 50503 5 1 1 50502
0 50504 7 1 2 50501 50503
0 50505 5 1 1 50504
0 50506 7 1 2 64502 50505
0 50507 5 1 1 50506
0 50508 7 1 2 69630 93679
0 50509 7 1 2 103276 50508
0 50510 5 1 1 50509
0 50511 7 1 2 50507 50510
0 50512 5 1 1 50511
0 50513 7 1 2 67443 50512
0 50514 5 1 1 50513
0 50515 7 1 2 92356 98160
0 50516 7 1 2 100482 50515
0 50517 5 1 1 50516
0 50518 7 1 2 50514 50517
0 50519 5 1 1 50518
0 50520 7 1 2 70905 50519
0 50521 5 1 1 50520
0 50522 7 2 2 87810 97210
0 50523 7 1 2 92816 106146
0 50524 5 1 1 50523
0 50525 7 1 2 50521 50524
0 50526 5 1 1 50525
0 50527 7 1 2 69283 50526
0 50528 5 1 1 50527
0 50529 7 1 2 100494 106147
0 50530 5 1 1 50529
0 50531 7 1 2 50528 50530
0 50532 5 1 1 50531
0 50533 7 1 2 84861 50532
0 50534 5 1 1 50533
0 50535 7 2 2 79705 83094
0 50536 5 2 1 106148
0 50537 7 1 2 50405 106150
0 50538 5 1 1 50537
0 50539 7 1 2 105865 50538
0 50540 5 1 1 50539
0 50541 7 2 2 87714 98918
0 50542 7 1 2 97887 106152
0 50543 5 1 1 50542
0 50544 7 1 2 97828 85026
0 50545 5 1 1 50544
0 50546 7 1 2 81780 92637
0 50547 5 1 1 50546
0 50548 7 1 2 50545 50547
0 50549 5 1 1 50548
0 50550 7 1 2 73585 50549
0 50551 5 1 1 50550
0 50552 7 1 2 72784 106149
0 50553 5 1 1 50552
0 50554 7 1 2 50551 50553
0 50555 5 1 1 50554
0 50556 7 1 2 70906 81069
0 50557 7 1 2 50555 50556
0 50558 5 1 1 50557
0 50559 7 1 2 50543 50558
0 50560 5 1 1 50559
0 50561 7 1 2 69284 50560
0 50562 5 1 1 50561
0 50563 7 1 2 100495 106153
0 50564 5 1 1 50563
0 50565 7 1 2 50562 50564
0 50566 5 1 1 50565
0 50567 7 1 2 67444 50566
0 50568 5 1 1 50567
0 50569 7 1 2 50540 50568
0 50570 7 1 2 50534 50569
0 50571 7 1 2 50499 50570
0 50572 5 1 1 50571
0 50573 7 1 2 72188 50572
0 50574 5 1 1 50573
0 50575 7 1 2 96898 94736
0 50576 7 1 2 96108 50575
0 50577 7 1 2 103772 50576
0 50578 5 1 1 50577
0 50579 7 1 2 50574 50578
0 50580 5 1 1 50579
0 50581 7 1 2 50442 50580
0 50582 5 1 1 50581
0 50583 7 1 2 96657 97060
0 50584 5 1 1 50583
0 50585 7 1 2 82276 98109
0 50586 5 1 1 50585
0 50587 7 1 2 50584 50586
0 50588 5 1 1 50587
0 50589 7 1 2 77489 50588
0 50590 5 1 1 50589
0 50591 7 1 2 72785 96658
0 50592 5 1 1 50591
0 50593 7 1 2 82277 97269
0 50594 5 1 1 50593
0 50595 7 1 2 50592 50594
0 50596 5 1 1 50595
0 50597 7 1 2 97742 50596
0 50598 5 1 1 50597
0 50599 7 1 2 50590 50598
0 50600 5 1 1 50599
0 50601 7 1 2 68727 50600
0 50602 5 1 1 50601
0 50603 7 1 2 101331 105708
0 50604 5 1 1 50603
0 50605 7 1 2 97130 94354
0 50606 7 1 2 92891 50605
0 50607 5 1 1 50606
0 50608 7 1 2 50604 50607
0 50609 7 1 2 50602 50608
0 50610 5 1 1 50609
0 50611 7 1 2 82467 50610
0 50612 5 1 1 50611
0 50613 7 1 2 73253 104858
0 50614 5 1 1 50613
0 50615 7 1 2 66079 10521
0 50616 5 1 1 50615
0 50617 7 1 2 105333 50616
0 50618 5 1 1 50617
0 50619 7 1 2 50614 50618
0 50620 5 1 1 50619
0 50621 7 1 2 68515 50620
0 50622 5 1 1 50621
0 50623 7 1 2 74747 105824
0 50624 5 1 1 50623
0 50625 7 1 2 50622 50624
0 50626 5 1 1 50625
0 50627 7 1 2 69631 50626
0 50628 5 1 1 50627
0 50629 7 1 2 71705 99010
0 50630 5 1 1 50629
0 50631 7 1 2 96661 50630
0 50632 5 1 1 50631
0 50633 7 1 2 100765 50632
0 50634 5 1 1 50633
0 50635 7 1 2 50628 50634
0 50636 5 1 1 50635
0 50637 7 1 2 105713 50636
0 50638 5 1 1 50637
0 50639 7 1 2 50612 50638
0 50640 5 1 1 50639
0 50641 7 1 2 74438 98050
0 50642 7 1 2 50640 50641
0 50643 5 1 1 50642
0 50644 7 1 2 50582 50643
0 50645 5 1 1 50644
0 50646 7 1 2 71960 50645
0 50647 5 1 1 50646
0 50648 7 2 2 72189 88900
0 50649 7 1 2 92441 93649
0 50650 7 1 2 106154 50649
0 50651 7 1 2 103744 50650
0 50652 5 1 1 50651
0 50653 7 1 2 102330 90253
0 50654 7 1 2 103331 50653
0 50655 5 1 1 50654
0 50656 7 1 2 50652 50655
0 50657 5 1 1 50656
0 50658 7 1 2 63927 50657
0 50659 5 1 1 50658
0 50660 7 1 2 86459 105485
0 50661 5 1 1 50660
0 50662 7 1 2 83478 96831
0 50663 5 1 1 50662
0 50664 7 1 2 50661 50663
0 50665 5 1 1 50664
0 50666 7 1 2 101873 98772
0 50667 7 1 2 50665 50666
0 50668 5 1 1 50667
0 50669 7 1 2 50659 50668
0 50670 5 1 1 50669
0 50671 7 1 2 66080 50670
0 50672 5 1 1 50671
0 50673 7 1 2 86460 96340
0 50674 5 2 1 50673
0 50675 7 1 2 83479 98129
0 50676 5 1 1 50675
0 50677 7 1 2 106156 50676
0 50678 5 2 1 50677
0 50679 7 1 2 73785 106157
0 50680 5 1 1 50679
0 50681 7 1 2 82468 50680
0 50682 7 2 2 106158 50681
0 50683 7 1 2 96766 91636
0 50684 7 1 2 106160 50683
0 50685 5 1 1 50684
0 50686 7 1 2 50672 50685
0 50687 5 1 1 50686
0 50688 7 1 2 64503 50687
0 50689 5 1 1 50688
0 50690 7 1 2 98412 106161
0 50691 5 1 1 50690
0 50692 7 1 2 99415 78493
0 50693 7 1 2 106159 50692
0 50694 5 1 1 50693
0 50695 7 1 2 50691 50694
0 50696 5 1 1 50695
0 50697 7 1 2 92495 50696
0 50698 5 1 1 50697
0 50699 7 1 2 50689 50698
0 50700 5 1 1 50699
0 50701 7 1 2 65613 50700
0 50702 5 1 1 50701
0 50703 7 1 2 105624 105711
0 50704 5 1 1 50703
0 50705 7 1 2 69285 50704
0 50706 5 1 1 50705
0 50707 7 1 2 105631 50706
0 50708 5 1 1 50707
0 50709 7 2 2 102985 50708
0 50710 7 1 2 92066 90320
0 50711 7 1 2 106162 50710
0 50712 5 1 1 50711
0 50713 7 1 2 67445 20712
0 50714 5 1 1 50713
0 50715 7 1 2 98379 101039
0 50716 5 1 1 50715
0 50717 7 1 2 50714 50716
0 50718 5 1 1 50717
0 50719 7 1 2 70907 50718
0 50720 5 1 1 50719
0 50721 7 1 2 105625 50720
0 50722 5 1 1 50721
0 50723 7 1 2 69286 50722
0 50724 5 1 1 50723
0 50725 7 1 2 105632 50724
0 50726 5 2 1 50725
0 50727 7 1 2 83480 96485
0 50728 7 1 2 106164 50727
0 50729 5 1 1 50728
0 50730 7 1 2 50712 50729
0 50731 5 1 1 50730
0 50732 7 1 2 76811 50731
0 50733 5 1 1 50732
0 50734 7 1 2 50702 50733
0 50735 5 1 1 50734
0 50736 7 1 2 73987 50735
0 50737 5 1 1 50736
0 50738 7 1 2 98045 106163
0 50739 5 1 1 50738
0 50740 7 1 2 79771 105378
0 50741 5 1 1 50740
0 50742 7 1 2 96353 105262
0 50743 5 1 1 50742
0 50744 7 1 2 50741 50743
0 50745 5 1 1 50744
0 50746 7 1 2 89728 50745
0 50747 7 1 2 106165 50746
0 50748 5 1 1 50747
0 50749 7 1 2 50739 50748
0 50750 5 1 1 50749
0 50751 7 1 2 71961 50750
0 50752 5 1 1 50751
0 50753 7 2 2 77776 92442
0 50754 7 2 2 91717 87440
0 50755 7 1 2 95320 106168
0 50756 7 1 2 106166 50755
0 50757 7 1 2 105791 50756
0 50758 5 1 1 50757
0 50759 7 1 2 50752 50758
0 50760 5 1 1 50759
0 50761 7 1 2 87041 50760
0 50762 5 1 1 50761
0 50763 7 1 2 75669 82684
0 50764 7 1 2 91287 50763
0 50765 7 1 2 103633 50764
0 50766 7 1 2 98892 50765
0 50767 5 1 1 50766
0 50768 7 1 2 50762 50767
0 50769 7 1 2 50737 50768
0 50770 7 1 2 50647 50769
0 50771 5 1 1 50770
0 50772 7 1 2 64871 50771
0 50773 5 1 1 50772
0 50774 7 1 2 75852 97683
0 50775 7 1 2 102820 50774
0 50776 5 1 1 50775
0 50777 7 1 2 98445 90865
0 50778 7 1 2 77701 50777
0 50779 5 1 1 50778
0 50780 7 1 2 50776 50779
0 50781 5 1 1 50780
0 50782 7 1 2 96652 50781
0 50783 5 1 1 50782
0 50784 7 2 2 82278 98617
0 50785 7 1 2 100384 104893
0 50786 7 1 2 106170 50785
0 50787 5 1 1 50786
0 50788 7 1 2 50783 50787
0 50789 5 1 1 50788
0 50790 7 1 2 69287 50789
0 50791 5 1 1 50790
0 50792 7 1 2 73254 101761
0 50793 5 1 1 50792
0 50794 7 1 2 66787 97761
0 50795 5 1 1 50794
0 50796 7 1 2 50793 50795
0 50797 5 1 1 50796
0 50798 7 1 2 105862 50797
0 50799 5 1 1 50798
0 50800 7 1 2 99466 102442
0 50801 7 1 2 97689 50800
0 50802 5 1 1 50801
0 50803 7 1 2 50799 50802
0 50804 7 1 2 50791 50803
0 50805 5 2 1 50804
0 50806 7 1 2 88241 106172
0 50807 5 1 1 50806
0 50808 7 1 2 28153 12538
0 50809 5 1 1 50808
0 50810 7 1 2 99396 50809
0 50811 5 1 1 50810
0 50812 7 1 2 48823 50811
0 50813 5 1 1 50812
0 50814 7 1 2 68164 50813
0 50815 5 1 1 50814
0 50816 7 1 2 95910 105755
0 50817 5 1 1 50816
0 50818 7 1 2 50815 50817
0 50819 5 1 1 50818
0 50820 7 1 2 78521 50819
0 50821 5 1 1 50820
0 50822 7 1 2 100521 95911
0 50823 5 1 1 50822
0 50824 7 1 2 100504 86900
0 50825 5 1 1 50824
0 50826 7 1 2 50823 50825
0 50827 5 1 1 50826
0 50828 7 1 2 70533 50827
0 50829 5 1 1 50828
0 50830 7 1 2 80547 81216
0 50831 7 1 2 93693 50830
0 50832 5 1 1 50831
0 50833 7 1 2 50829 50832
0 50834 5 1 1 50833
0 50835 7 1 2 96767 50834
0 50836 5 1 1 50835
0 50837 7 1 2 50821 50836
0 50838 5 1 1 50837
0 50839 7 2 2 72190 50838
0 50840 7 1 2 69014 106174
0 50841 5 1 1 50840
0 50842 7 1 2 50807 50841
0 50843 5 1 1 50842
0 50844 7 1 2 68728 50843
0 50845 5 1 1 50844
0 50846 7 1 2 95037 103846
0 50847 5 1 1 50846
0 50848 7 1 2 103673 38421
0 50849 5 1 1 50848
0 50850 7 1 2 98088 50849
0 50851 5 1 1 50850
0 50852 7 1 2 50847 50851
0 50853 5 1 1 50852
0 50854 7 1 2 82469 50853
0 50855 5 1 1 50854
0 50856 7 3 2 67446 82508
0 50857 7 1 2 95038 106176
0 50858 7 1 2 78522 50857
0 50859 5 1 1 50858
0 50860 7 1 2 50855 50859
0 50861 5 1 1 50860
0 50862 7 1 2 80748 74439
0 50863 7 1 2 50861 50862
0 50864 5 1 1 50863
0 50865 7 1 2 74695 89239
0 50866 5 1 1 50865
0 50867 7 1 2 2993 105854
0 50868 7 1 2 50866 50867
0 50869 5 1 1 50868
0 50870 7 1 2 100522 50869
0 50871 5 1 1 50870
0 50872 7 1 2 87388 95914
0 50873 5 1 1 50872
0 50874 7 1 2 101087 105915
0 50875 7 1 2 50873 50874
0 50876 5 1 1 50875
0 50877 7 1 2 50871 50876
0 50878 5 1 1 50877
0 50879 7 1 2 67447 50878
0 50880 5 1 1 50879
0 50881 7 1 2 4236 96463
0 50882 5 1 1 50881
0 50883 7 1 2 82656 102315
0 50884 7 1 2 78523 50883
0 50885 7 1 2 50882 50884
0 50886 5 1 1 50885
0 50887 7 1 2 50880 50886
0 50888 7 1 2 50864 50887
0 50889 5 2 1 50888
0 50890 7 1 2 88600 106179
0 50891 5 1 1 50890
0 50892 7 1 2 83050 96604
0 50893 5 1 1 50892
0 50894 7 1 2 106006 50893
0 50895 5 1 1 50894
0 50896 7 1 2 105929 50895
0 50897 5 1 1 50896
0 50898 7 1 2 82638 97131
0 50899 7 1 2 78003 50898
0 50900 5 1 1 50899
0 50901 7 1 2 69632 85809
0 50902 7 1 2 99488 50901
0 50903 5 1 1 50902
0 50904 7 1 2 50900 50903
0 50905 5 1 1 50904
0 50906 7 1 2 83761 50905
0 50907 5 1 1 50906
0 50908 7 1 2 50897 50907
0 50909 5 1 1 50908
0 50910 7 2 2 67138 50909
0 50911 7 1 2 63928 106181
0 50912 5 1 1 50911
0 50913 7 1 2 50891 50912
0 50914 7 1 2 50845 50913
0 50915 5 1 1 50914
0 50916 7 1 2 69997 50915
0 50917 5 1 1 50916
0 50918 7 1 2 83466 105752
0 50919 5 1 1 50918
0 50920 7 1 2 100912 102448
0 50921 5 1 1 50920
0 50922 7 1 2 105884 48872
0 50923 5 1 1 50922
0 50924 7 1 2 84862 50923
0 50925 5 1 1 50924
0 50926 7 1 2 50921 50925
0 50927 7 1 2 50919 50926
0 50928 5 1 1 50927
0 50929 7 1 2 74570 50928
0 50930 5 1 1 50929
0 50931 7 1 2 86986 105949
0 50932 5 1 1 50931
0 50933 7 1 2 50930 50932
0 50934 5 1 1 50933
0 50935 7 1 2 68165 90983
0 50936 7 2 2 50934 50935
0 50937 7 1 2 89129 106183
0 50938 5 1 1 50937
0 50939 7 2 2 68166 103447
0 50940 7 1 2 85471 104547
0 50941 5 1 1 50940
0 50942 7 1 2 69633 99471
0 50943 5 1 1 50942
0 50944 7 1 2 50941 50943
0 50945 5 1 1 50944
0 50946 7 1 2 106185 50945
0 50947 5 1 1 50946
0 50948 7 1 2 65503 104986
0 50949 5 1 1 50948
0 50950 7 1 2 87145 50949
0 50951 5 1 1 50950
0 50952 7 1 2 65195 50951
0 50953 5 1 1 50952
0 50954 7 1 2 88855 50953
0 50955 5 1 1 50954
0 50956 7 1 2 82470 98593
0 50957 7 1 2 50955 50956
0 50958 5 1 1 50957
0 50959 7 1 2 50947 50958
0 50960 5 2 1 50959
0 50961 7 1 2 88242 106187
0 50962 5 1 1 50961
0 50963 7 1 2 50938 50962
0 50964 5 1 1 50963
0 50965 7 1 2 83762 50964
0 50966 5 1 1 50965
0 50967 7 1 2 85027 101264
0 50968 5 1 1 50967
0 50969 7 1 2 105855 50968
0 50970 5 1 1 50969
0 50971 7 2 2 68729 50970
0 50972 5 1 1 106189
0 50973 7 2 2 86222 97772
0 50974 7 1 2 83567 106191
0 50975 5 1 1 50974
0 50976 7 1 2 50972 50975
0 50977 5 1 1 50976
0 50978 7 1 2 69634 50977
0 50979 5 1 1 50978
0 50980 7 1 2 9310 50979
0 50981 5 1 1 50980
0 50982 7 1 2 104109 50981
0 50983 5 1 1 50982
0 50984 7 1 2 22765 78780
0 50985 5 1 1 50984
0 50986 7 1 2 94658 50985
0 50987 5 1 1 50986
0 50988 7 1 2 9308 50987
0 50989 5 1 1 50988
0 50990 7 1 2 105888 50989
0 50991 5 1 1 50990
0 50992 7 1 2 100124 106190
0 50993 5 1 1 50992
0 50994 7 1 2 50991 50993
0 50995 5 1 1 50994
0 50996 7 1 2 67448 50995
0 50997 5 1 1 50996
0 50998 7 1 2 80238 81217
0 50999 5 1 1 50998
0 51000 7 1 2 84244 79926
0 51001 5 1 1 51000
0 51002 7 1 2 50999 51001
0 51003 5 1 1 51002
0 51004 7 1 2 81931 51003
0 51005 7 1 2 105930 51004
0 51006 5 1 1 51005
0 51007 7 1 2 50997 51006
0 51008 7 1 2 50983 51007
0 51009 5 2 1 51008
0 51010 7 1 2 88243 106193
0 51011 5 1 1 51010
0 51012 7 3 2 99416 80749
0 51013 5 1 1 106195
0 51014 7 1 2 99758 87192
0 51015 5 1 1 51014
0 51016 7 1 2 51013 51015
0 51017 5 1 1 51016
0 51018 7 1 2 68516 51017
0 51019 5 1 1 51018
0 51020 7 1 2 82471 102131
0 51021 7 1 2 88683 51020
0 51022 5 1 1 51021
0 51023 7 1 2 51019 51022
0 51024 5 1 1 51023
0 51025 7 2 2 104848 51024
0 51026 7 1 2 69015 106198
0 51027 5 1 1 51026
0 51028 7 1 2 89697 105931
0 51029 5 1 1 51028
0 51030 7 1 2 51027 51029
0 51031 5 1 1 51030
0 51032 7 1 2 95858 51031
0 51033 5 1 1 51032
0 51034 7 1 2 83362 98919
0 51035 5 1 1 51034
0 51036 7 1 2 104881 86013
0 51037 5 1 1 51036
0 51038 7 1 2 51035 51037
0 51039 5 1 1 51038
0 51040 7 1 2 68517 51039
0 51041 5 1 1 51040
0 51042 7 1 2 87822 105490
0 51043 5 1 1 51042
0 51044 7 1 2 51041 51043
0 51045 5 1 1 51044
0 51046 7 1 2 93694 51045
0 51047 5 1 1 51046
0 51048 7 1 2 67792 103749
0 51049 7 1 2 103682 51048
0 51050 5 1 1 51049
0 51051 7 1 2 51047 51050
0 51052 5 1 1 51051
0 51053 7 1 2 64504 51052
0 51054 5 1 1 51053
0 51055 7 1 2 83363 105903
0 51056 5 1 1 51055
0 51057 7 1 2 51054 51056
0 51058 5 1 1 51057
0 51059 7 2 2 102749 51058
0 51060 7 1 2 69016 106200
0 51061 5 1 1 51060
0 51062 7 1 2 51033 51061
0 51063 7 1 2 51011 51062
0 51064 7 1 2 50966 51063
0 51065 7 1 2 50917 51064
0 51066 5 1 1 51065
0 51067 7 1 2 89586 51066
0 51068 5 1 1 51067
0 51069 7 1 2 78098 106173
0 51070 5 1 1 51069
0 51071 7 1 2 75163 106175
0 51072 5 1 1 51071
0 51073 7 1 2 51070 51072
0 51074 5 1 1 51073
0 51075 7 1 2 68730 51074
0 51076 5 1 1 51075
0 51077 7 1 2 75188 106180
0 51078 5 1 1 51077
0 51079 7 1 2 78081 106182
0 51080 5 1 1 51079
0 51081 7 1 2 51078 51080
0 51082 7 1 2 51076 51081
0 51083 5 1 1 51082
0 51084 7 1 2 69998 51083
0 51085 5 1 1 51084
0 51086 7 1 2 78099 106188
0 51087 5 1 1 51086
0 51088 7 1 2 70645 89870
0 51089 7 1 2 106184 51088
0 51090 5 1 1 51089
0 51091 7 1 2 51087 51090
0 51092 5 1 1 51091
0 51093 7 1 2 83763 51092
0 51094 5 1 1 51093
0 51095 7 1 2 78100 106194
0 51096 5 1 1 51095
0 51097 7 1 2 75164 106199
0 51098 5 1 1 51097
0 51099 7 1 2 105932 105980
0 51100 5 1 1 51099
0 51101 7 1 2 51098 51100
0 51102 5 1 1 51101
0 51103 7 1 2 95859 51102
0 51104 5 1 1 51103
0 51105 7 1 2 75165 106201
0 51106 5 1 1 51105
0 51107 7 1 2 51104 51106
0 51108 7 1 2 51096 51107
0 51109 7 1 2 51094 51108
0 51110 7 1 2 51085 51109
0 51111 5 1 1 51110
0 51112 7 1 2 73874 51111
0 51113 5 1 1 51112
0 51114 7 1 2 51068 51113
0 51115 5 1 1 51114
0 51116 7 1 2 71962 51115
0 51117 5 1 1 51116
0 51118 7 1 2 65504 90291
0 51119 7 2 2 91294 51118
0 51120 7 2 2 64505 106202
0 51121 7 1 2 93266 101870
0 51122 7 2 2 105775 51121
0 51123 7 1 2 64203 106206
0 51124 7 1 2 106204 51123
0 51125 5 1 1 51124
0 51126 7 1 2 51117 51125
0 51127 7 1 2 50773 51126
0 51128 5 1 1 51127
0 51129 7 1 2 66372 51128
0 51130 5 1 1 51129
0 51131 7 1 2 105306 106203
0 51132 7 1 2 106207 51131
0 51133 5 1 1 51132
0 51134 7 1 2 68892 51133
0 51135 7 1 2 51130 51134
0 51136 7 1 2 50438 51135
0 51137 5 1 1 51136
0 51138 7 1 2 67007 51137
0 51139 7 1 2 48914 51138
0 51140 5 1 1 51139
0 51141 7 1 2 71870 100914
0 51142 5 1 1 51141
0 51143 7 1 2 71477 93462
0 51144 7 1 2 51142 51143
0 51145 5 1 1 51144
0 51146 7 1 2 70534 88713
0 51147 7 1 2 89948 51146
0 51148 7 1 2 51145 51147
0 51149 5 1 1 51148
0 51150 7 1 2 81613 103386
0 51151 5 2 1 51150
0 51152 7 1 2 72786 106208
0 51153 7 1 2 51149 51152
0 51154 5 1 1 51153
0 51155 7 1 2 87205 103391
0 51156 5 1 1 51155
0 51157 7 1 2 76240 94429
0 51158 5 1 1 51157
0 51159 7 1 2 67793 51158
0 51160 7 1 2 51156 51159
0 51161 5 1 1 51160
0 51162 7 1 2 69635 51161
0 51163 7 1 2 51154 51162
0 51164 5 1 1 51163
0 51165 7 1 2 81012 51164
0 51166 5 1 1 51165
0 51167 7 1 2 71478 100915
0 51168 5 1 1 51167
0 51169 7 1 2 83313 51168
0 51170 5 1 1 51169
0 51171 7 1 2 80650 51170
0 51172 5 1 1 51171
0 51173 7 1 2 95071 81649
0 51174 5 1 1 51173
0 51175 7 1 2 77271 51174
0 51176 7 1 2 51172 51175
0 51177 5 1 1 51176
0 51178 7 1 2 88601 98853
0 51179 7 1 2 51177 51178
0 51180 7 1 2 51166 51179
0 51181 5 1 1 51180
0 51182 7 1 2 80130 89249
0 51183 7 1 2 99961 51182
0 51184 7 1 2 89841 51183
0 51185 5 1 1 51184
0 51186 7 1 2 51181 51185
0 51187 5 1 1 51186
0 51188 7 1 2 91910 51187
0 51189 5 1 1 51188
0 51190 7 1 2 92240 84650
0 51191 7 1 2 94373 51190
0 51192 5 2 1 51191
0 51193 7 5 2 94016 96699
0 51194 7 3 2 105151 106212
0 51195 7 1 2 87075 1223
0 51196 5 7 1 51195
0 51197 7 1 2 66373 106220
0 51198 7 1 2 106217 51197
0 51199 5 1 1 51198
0 51200 7 1 2 106210 51199
0 51201 5 1 1 51200
0 51202 7 1 2 66596 51201
0 51203 5 1 1 51202
0 51204 7 1 2 93830 100646
0 51205 5 1 1 51204
0 51206 7 1 2 91315 51205
0 51207 5 1 1 51206
0 51208 7 1 2 51203 51207
0 51209 5 1 1 51208
0 51210 7 1 2 64872 51209
0 51211 5 1 1 51210
0 51212 7 1 2 99824 103024
0 51213 5 1 1 51212
0 51214 7 1 2 65196 51213
0 51215 5 1 1 51214
0 51216 7 1 2 66597 94903
0 51217 5 1 1 51216
0 51218 7 1 2 51215 51217
0 51219 5 1 1 51218
0 51220 7 1 2 91316 51219
0 51221 5 1 1 51220
0 51222 7 1 2 51211 51221
0 51223 5 1 1 51222
0 51224 7 1 2 73586 51223
0 51225 5 1 1 51224
0 51226 7 2 2 91310 88925
0 51227 7 2 2 70535 106227
0 51228 7 2 2 67139 87107
0 51229 7 1 2 87206 106231
0 51230 7 1 2 106229 51229
0 51231 5 1 1 51230
0 51232 7 1 2 51225 51231
0 51233 5 1 1 51232
0 51234 7 1 2 68167 51233
0 51235 5 1 1 51234
0 51236 7 1 2 73255 84166
0 51237 7 1 2 92241 51236
0 51238 7 1 2 100046 51237
0 51239 7 1 2 106230 51238
0 51240 5 1 1 51239
0 51241 7 1 2 51235 51240
0 51242 5 1 1 51241
0 51243 7 1 2 67794 51242
0 51244 5 1 1 51243
0 51245 7 6 2 80750 87706
0 51246 7 1 2 94247 106233
0 51247 5 1 1 51246
0 51248 7 2 2 75458 105531
0 51249 5 1 1 106239
0 51250 7 1 2 51247 51249
0 51251 5 1 1 51250
0 51252 7 1 2 72787 51251
0 51253 5 1 1 51252
0 51254 7 3 2 91706 106234
0 51255 7 1 2 94340 106241
0 51256 5 1 1 51255
0 51257 7 1 2 51253 51256
0 51258 5 1 1 51257
0 51259 7 1 2 68168 51258
0 51260 5 1 1 51259
0 51261 7 3 2 71963 84683
0 51262 7 1 2 96613 91190
0 51263 7 1 2 106244 51262
0 51264 5 1 1 51263
0 51265 7 1 2 81495 105856
0 51266 5 1 1 51265
0 51267 7 1 2 88994 51266
0 51268 5 1 1 51267
0 51269 7 1 2 71479 51268
0 51270 7 1 2 51264 51269
0 51271 7 1 2 51260 51270
0 51272 5 1 1 51271
0 51273 7 1 2 69636 87825
0 51274 7 1 2 87819 51273
0 51275 5 1 1 51274
0 51276 7 1 2 80751 84946
0 51277 7 1 2 88080 51276
0 51278 7 1 2 95876 51277
0 51279 7 1 2 51275 51278
0 51280 5 1 1 51279
0 51281 7 1 2 63981 66895
0 51282 7 1 2 81781 51281
0 51283 7 1 2 92232 51282
0 51284 7 1 2 84517 51283
0 51285 5 1 1 51284
0 51286 7 1 2 66374 51285
0 51287 7 1 2 51280 51286
0 51288 5 1 1 51287
0 51289 7 1 2 51272 51288
0 51290 5 1 1 51289
0 51291 7 1 2 73256 75491
0 51292 5 1 1 51291
0 51293 7 1 2 81486 88995
0 51294 7 1 2 51292 51293
0 51295 5 1 1 51294
0 51296 7 1 2 51290 51295
0 51297 5 1 1 51296
0 51298 7 1 2 88244 51297
0 51299 5 1 1 51298
0 51300 7 3 2 74748 106221
0 51301 7 1 2 91416 106247
0 51302 5 1 1 51301
0 51303 7 1 2 63982 80104
0 51304 7 1 2 96614 51303
0 51305 7 1 2 91262 51304
0 51306 5 1 1 51305
0 51307 7 1 2 51302 51306
0 51308 5 1 1 51307
0 51309 7 1 2 67795 51308
0 51310 5 1 1 51309
0 51311 7 1 2 100568 82159
0 51312 7 1 2 98874 51311
0 51313 5 1 1 51312
0 51314 7 1 2 51310 51313
0 51315 5 1 1 51314
0 51316 7 1 2 66598 51315
0 51317 5 1 1 51316
0 51318 7 1 2 65197 77679
0 51319 5 1 1 51318
0 51320 7 1 2 69637 51319
0 51321 5 1 1 51320
0 51322 7 1 2 88996 98920
0 51323 7 1 2 51321 51322
0 51324 5 1 1 51323
0 51325 7 1 2 51317 51324
0 51326 5 1 1 51325
0 51327 7 1 2 93166 51326
0 51328 5 1 1 51327
0 51329 7 1 2 70536 100353
0 51330 7 1 2 91290 90296
0 51331 7 1 2 51329 51330
0 51332 5 1 1 51331
0 51333 7 1 2 79579 91405
0 51334 7 1 2 95000 95611
0 51335 7 1 2 91395 51334
0 51336 7 1 2 51333 51335
0 51337 5 1 1 51336
0 51338 7 1 2 51332 51337
0 51339 5 1 1 51338
0 51340 7 1 2 71871 51339
0 51341 5 1 1 51340
0 51342 7 1 2 74498 88448
0 51343 5 2 1 51342
0 51344 7 1 2 66375 106250
0 51345 5 1 1 51344
0 51346 7 1 2 81225 51345
0 51347 5 1 1 51346
0 51348 7 1 2 91375 98921
0 51349 7 1 2 51347 51348
0 51350 5 1 1 51349
0 51351 7 1 2 51341 51350
0 51352 7 1 2 51328 51351
0 51353 7 1 2 51299 51352
0 51354 5 1 1 51353
0 51355 7 1 2 69999 51354
0 51356 5 1 1 51355
0 51357 7 1 2 92134 91573
0 51358 7 1 2 105581 51357
0 51359 5 1 1 51358
0 51360 7 1 2 91579 51359
0 51361 5 1 1 51360
0 51362 7 1 2 83236 51361
0 51363 5 1 1 51362
0 51364 7 1 2 88997 90780
0 51365 5 1 1 51364
0 51366 7 1 2 80250 94248
0 51367 7 1 2 90677 51366
0 51368 5 1 1 51367
0 51369 7 1 2 51365 51368
0 51370 5 2 1 51369
0 51371 7 1 2 76096 106252
0 51372 5 1 1 51371
0 51373 7 1 2 91376 105414
0 51374 5 1 1 51373
0 51375 7 1 2 51372 51374
0 51376 5 1 1 51375
0 51377 7 1 2 64873 51376
0 51378 5 1 1 51377
0 51379 7 1 2 51363 51378
0 51380 5 1 1 51379
0 51381 7 1 2 67796 51380
0 51382 5 1 1 51381
0 51383 7 1 2 81614 105107
0 51384 7 1 2 96049 51383
0 51385 7 1 2 91654 51384
0 51386 5 1 1 51385
0 51387 7 1 2 51382 51386
0 51388 5 1 1 51387
0 51389 7 1 2 80752 51388
0 51390 5 1 1 51389
0 51391 7 1 2 81487 85997
0 51392 7 1 2 92245 51391
0 51393 7 1 2 102604 51392
0 51394 5 1 1 51393
0 51395 7 1 2 51390 51394
0 51396 7 1 2 51356 51395
0 51397 7 1 2 51244 51396
0 51398 5 1 1 51397
0 51399 7 1 2 71184 51398
0 51400 5 1 1 51399
0 51401 7 1 2 72788 106240
0 51402 5 1 1 51401
0 51403 7 1 2 100364 90377
0 51404 7 1 2 106242 51403
0 51405 5 1 1 51404
0 51406 7 1 2 51402 51405
0 51407 5 1 1 51406
0 51408 7 1 2 68169 51407
0 51409 5 1 1 51408
0 51410 7 2 2 91884 90535
0 51411 7 1 2 93371 96615
0 51412 7 1 2 106254 51411
0 51413 5 1 1 51412
0 51414 7 1 2 51409 51413
0 51415 5 1 1 51414
0 51416 7 1 2 88245 51415
0 51417 5 1 1 51416
0 51418 7 1 2 101865 90789
0 51419 5 1 1 51418
0 51420 7 1 2 94052 106248
0 51421 5 1 1 51420
0 51422 7 1 2 51419 51421
0 51423 5 1 1 51422
0 51424 7 1 2 101748 84623
0 51425 7 1 2 51423 51424
0 51426 5 1 1 51425
0 51427 7 1 2 51417 51426
0 51428 5 1 1 51427
0 51429 7 1 2 71480 51428
0 51430 5 1 1 51429
0 51431 7 1 2 91377 105364
0 51432 5 1 1 51431
0 51433 7 1 2 66376 75166
0 51434 7 1 2 87671 51433
0 51435 7 1 2 94086 96224
0 51436 7 1 2 51434 51435
0 51437 5 1 1 51436
0 51438 7 1 2 51432 51437
0 51439 5 1 1 51438
0 51440 7 1 2 98922 51439
0 51441 5 1 1 51440
0 51442 7 1 2 51430 51441
0 51443 5 1 1 51442
0 51444 7 1 2 70000 51443
0 51445 5 1 1 51444
0 51446 7 1 2 64874 82084
0 51447 5 1 1 51446
0 51448 7 1 2 87057 51447
0 51449 5 1 1 51448
0 51450 7 1 2 91378 51449
0 51451 5 1 1 51450
0 51452 7 2 2 75167 94093
0 51453 7 1 2 87672 96225
0 51454 7 1 2 106256 51453
0 51455 5 1 1 51454
0 51456 7 1 2 51451 51455
0 51457 5 1 1 51456
0 51458 7 1 2 71481 51457
0 51459 5 1 1 51458
0 51460 7 1 2 92166 97157
0 51461 7 1 2 105165 51460
0 51462 5 2 1 51461
0 51463 7 1 2 51459 106258
0 51464 5 1 1 51463
0 51465 7 1 2 98923 51464
0 51466 5 1 1 51465
0 51467 7 1 2 51445 51466
0 51468 5 1 1 51467
0 51469 7 1 2 69638 51468
0 51470 5 1 1 51469
0 51471 7 1 2 77777 90426
0 51472 7 1 2 86118 51471
0 51473 7 1 2 96248 51472
0 51474 7 1 2 105105 51473
0 51475 5 1 1 51474
0 51476 7 1 2 51470 51475
0 51477 7 1 2 51400 51476
0 51478 5 1 1 51477
0 51479 7 1 2 85953 51478
0 51480 5 1 1 51479
0 51481 7 1 2 51189 51480
0 51482 5 1 1 51481
0 51483 7 1 2 69288 51482
0 51484 5 1 1 51483
0 51485 7 2 2 93848 89359
0 51486 5 1 1 106260
0 51487 7 1 2 93935 106261
0 51488 5 1 1 51487
0 51489 7 1 2 104062 88602
0 51490 5 1 1 51489
0 51491 7 1 2 98533 51490
0 51492 5 1 1 51491
0 51493 7 1 2 75292 51492
0 51494 5 1 1 51493
0 51495 7 1 2 51488 51494
0 51496 5 3 1 51495
0 51497 7 1 2 92280 76973
0 51498 7 1 2 92595 92603
0 51499 7 1 2 51497 51498
0 51500 7 1 2 106262 51499
0 51501 5 1 1 51500
0 51502 7 1 2 51484 51501
0 51503 5 1 1 51502
0 51504 7 1 2 67449 51503
0 51505 5 1 1 51504
0 51506 7 2 2 75050 75223
0 51507 5 1 1 106265
0 51508 7 1 2 87707 78549
0 51509 5 1 1 51508
0 51510 7 1 2 51507 51509
0 51511 5 1 1 51510
0 51512 7 1 2 75938 51511
0 51513 5 1 1 51512
0 51514 7 1 2 65198 75195
0 51515 7 2 2 93964 51514
0 51516 5 1 1 106267
0 51517 7 1 2 78666 106268
0 51518 5 1 1 51517
0 51519 7 1 2 51513 51518
0 51520 5 1 1 51519
0 51521 7 1 2 64875 51520
0 51522 5 1 1 51521
0 51523 7 1 2 63929 89817
0 51524 7 1 2 103374 51523
0 51525 5 1 1 51524
0 51526 7 1 2 51522 51525
0 51527 5 2 1 51526
0 51528 7 1 2 105142 106269
0 51529 5 1 1 51528
0 51530 7 3 2 70729 66377
0 51531 7 1 2 77680 106271
0 51532 7 1 2 101597 51531
0 51533 7 1 2 90796 91922
0 51534 7 1 2 51532 51533
0 51535 5 1 1 51534
0 51536 7 1 2 51529 51535
0 51537 5 1 1 51536
0 51538 7 1 2 80753 51537
0 51539 5 1 1 51538
0 51540 7 1 2 67008 90321
0 51541 7 2 2 78101 51540
0 51542 7 1 2 64876 89968
0 51543 5 1 1 51542
0 51544 7 1 2 104996 51543
0 51545 5 1 1 51544
0 51546 7 1 2 106274 51545
0 51547 5 1 1 51546
0 51548 7 4 2 63930 70690
0 51549 7 1 2 86223 75825
0 51550 7 1 2 106276 51549
0 51551 7 2 2 91711 106272
0 51552 7 1 2 95001 106280
0 51553 7 1 2 51550 51552
0 51554 5 1 1 51553
0 51555 7 1 2 51547 51554
0 51556 5 1 1 51555
0 51557 7 1 2 73988 51556
0 51558 5 1 1 51557
0 51559 7 1 2 93295 106275
0 51560 5 1 1 51559
0 51561 7 1 2 75939 75526
0 51562 7 1 2 77022 51561
0 51563 7 1 2 106257 51562
0 51564 5 1 1 51563
0 51565 7 1 2 51560 51564
0 51566 5 1 1 51565
0 51567 7 1 2 82331 51566
0 51568 5 1 1 51567
0 51569 7 1 2 51558 51568
0 51570 5 1 1 51569
0 51571 7 1 2 78185 51570
0 51572 5 1 1 51571
0 51573 7 1 2 87750 87516
0 51574 7 1 2 102172 51573
0 51575 7 1 2 106281 51574
0 51576 7 1 2 94120 51575
0 51577 5 1 1 51576
0 51578 7 1 2 51572 51577
0 51579 7 1 2 51539 51578
0 51580 5 1 1 51579
0 51581 7 1 2 101557 98698
0 51582 7 1 2 51580 51581
0 51583 5 1 1 51582
0 51584 7 1 2 51505 51583
0 51585 5 1 1 51584
0 51586 7 1 2 65851 51585
0 51587 5 1 1 51586
0 51588 7 1 2 79857 96185
0 51589 5 1 1 51588
0 51590 7 1 2 86142 75762
0 51591 7 1 2 78335 51590
0 51592 5 1 1 51591
0 51593 7 1 2 51589 51592
0 51594 5 1 1 51593
0 51595 7 1 2 65505 51594
0 51596 5 1 1 51595
0 51597 7 1 2 79772 95929
0 51598 5 1 1 51597
0 51599 7 1 2 51596 51598
0 51600 5 1 1 51599
0 51601 7 1 2 81405 51600
0 51602 5 1 1 51601
0 51603 7 1 2 64506 105961
0 51604 5 2 1 51603
0 51605 7 1 2 104668 106282
0 51606 5 1 1 51605
0 51607 7 1 2 51602 51606
0 51608 5 1 1 51607
0 51609 7 1 2 71482 51608
0 51610 5 1 1 51609
0 51611 7 1 2 64507 45637
0 51612 5 2 1 51611
0 51613 7 1 2 70001 106284
0 51614 5 1 1 51613
0 51615 7 1 2 70537 94963
0 51616 5 1 1 51615
0 51617 7 1 2 51614 51616
0 51618 5 1 1 51617
0 51619 7 1 2 72789 51618
0 51620 5 1 1 51619
0 51621 7 1 2 82147 86155
0 51622 5 1 1 51621
0 51623 7 1 2 51620 51622
0 51624 5 1 1 51623
0 51625 7 1 2 78270 51624
0 51626 5 1 1 51625
0 51627 7 1 2 51610 51626
0 51628 5 1 1 51627
0 51629 7 1 2 68170 51628
0 51630 5 1 1 51629
0 51631 7 1 2 94966 102996
0 51632 5 1 1 51631
0 51633 7 1 2 70002 51632
0 51634 5 1 1 51633
0 51635 7 1 2 69639 103000
0 51636 5 1 1 51635
0 51637 7 1 2 51634 51636
0 51638 5 1 1 51637
0 51639 7 1 2 72790 51638
0 51640 5 1 1 51639
0 51641 7 1 2 86174 92193
0 51642 5 1 1 51641
0 51643 7 1 2 51640 51642
0 51644 5 1 1 51643
0 51645 7 1 2 70538 51644
0 51646 5 1 1 51645
0 51647 7 2 2 1927 51646
0 51648 5 1 1 106286
0 51649 7 1 2 78271 51648
0 51650 5 1 1 51649
0 51651 7 1 2 51630 51650
0 51652 5 1 1 51651
0 51653 7 1 2 71185 51652
0 51654 5 1 1 51653
0 51655 7 1 2 69640 98659
0 51656 7 2 2 102161 51655
0 51657 5 1 1 106288
0 51658 7 1 2 91023 106289
0 51659 5 1 1 51658
0 51660 7 1 2 51654 51659
0 51661 5 1 1 51660
0 51662 7 1 2 88246 51661
0 51663 5 1 1 51662
0 51664 7 1 2 103829 96568
0 51665 5 1 1 51664
0 51666 7 1 2 70539 104733
0 51667 5 1 1 51666
0 51668 7 1 2 51665 51667
0 51669 5 1 1 51668
0 51670 7 1 2 68518 51669
0 51671 5 1 1 51670
0 51672 7 1 2 85771 106070
0 51673 5 1 1 51672
0 51674 7 1 2 70268 51673
0 51675 5 1 1 51674
0 51676 7 1 2 38619 51675
0 51677 5 2 1 51676
0 51678 7 1 2 91109 106290
0 51679 5 1 1 51678
0 51680 7 1 2 51671 51679
0 51681 5 1 1 51680
0 51682 7 1 2 71483 51681
0 51683 5 1 1 51682
0 51684 7 2 2 96729 90083
0 51685 7 1 2 101665 88778
0 51686 5 2 1 51685
0 51687 7 1 2 106292 106294
0 51688 5 1 1 51687
0 51689 7 1 2 51683 51688
0 51690 5 1 1 51689
0 51691 7 1 2 72791 51690
0 51692 5 1 1 51691
0 51693 7 1 2 79125 105875
0 51694 5 1 1 51693
0 51695 7 1 2 64508 105370
0 51696 5 1 1 51695
0 51697 7 1 2 83794 92194
0 51698 5 1 1 51697
0 51699 7 1 2 51696 51698
0 51700 5 1 1 51699
0 51701 7 1 2 104742 51700
0 51702 5 1 1 51701
0 51703 7 1 2 51694 51702
0 51704 7 1 2 51692 51703
0 51705 5 1 1 51704
0 51706 7 1 2 70003 51705
0 51707 5 1 1 51706
0 51708 7 1 2 84086 106293
0 51709 5 1 1 51708
0 51710 7 1 2 94568 95741
0 51711 7 1 2 101866 51710
0 51712 5 1 1 51711
0 51713 7 1 2 51709 51712
0 51714 5 1 1 51713
0 51715 7 1 2 73587 51714
0 51716 5 1 1 51715
0 51717 7 1 2 104727 87949
0 51718 5 1 1 51717
0 51719 7 1 2 51716 51718
0 51720 5 1 1 51719
0 51721 7 1 2 64877 51720
0 51722 5 1 1 51721
0 51723 7 1 2 71484 87365
0 51724 7 1 2 95841 51723
0 51725 5 1 1 51724
0 51726 7 1 2 51722 51725
0 51727 5 1 1 51726
0 51728 7 1 2 67797 51727
0 51729 5 1 1 51728
0 51730 7 1 2 99740 82160
0 51731 7 1 2 91110 51730
0 51732 5 1 1 51731
0 51733 7 1 2 51729 51732
0 51734 5 1 1 51733
0 51735 7 1 2 74696 51734
0 51736 5 1 1 51735
0 51737 7 1 2 98327 103625
0 51738 7 2 2 71485 80302
0 51739 7 1 2 94921 106296
0 51740 7 1 2 51737 51739
0 51741 5 1 1 51740
0 51742 7 1 2 51736 51741
0 51743 7 1 2 51707 51742
0 51744 5 1 1 51743
0 51745 7 1 2 71186 51744
0 51746 5 1 1 51745
0 51747 7 1 2 90084 86147
0 51748 5 1 1 51747
0 51749 7 1 2 104744 51748
0 51750 5 1 1 51749
0 51751 7 1 2 75023 51750
0 51752 5 1 1 51751
0 51753 7 1 2 95056 95988
0 51754 5 1 1 51753
0 51755 7 1 2 51752 51754
0 51756 5 1 1 51755
0 51757 7 1 2 64878 51756
0 51758 5 1 1 51757
0 51759 7 1 2 96616 78272
0 51760 5 1 1 51759
0 51761 7 2 2 66599 89931
0 51762 7 1 2 95943 83489
0 51763 7 1 2 106298 51762
0 51764 5 1 1 51763
0 51765 7 1 2 51760 51764
0 51766 5 1 1 51765
0 51767 7 1 2 66378 51766
0 51768 5 1 1 51767
0 51769 7 1 2 71187 51768
0 51770 7 1 2 51758 51769
0 51771 5 1 1 51770
0 51772 7 1 2 103389 31990
0 51773 7 1 2 85728 51772
0 51774 5 3 1 51773
0 51775 7 1 2 85177 106300
0 51776 5 1 1 51775
0 51777 7 1 2 104745 51776
0 51778 5 1 1 51777
0 51779 7 1 2 74978 51778
0 51780 5 1 1 51779
0 51781 7 1 2 84058 75988
0 51782 7 1 2 94578 51781
0 51783 5 1 1 51782
0 51784 7 1 2 66081 51783
0 51785 7 1 2 51780 51784
0 51786 5 1 1 51785
0 51787 7 1 2 51771 51786
0 51788 5 1 1 51787
0 51789 7 1 2 99849 78273
0 51790 7 1 2 102848 51789
0 51791 5 1 1 51790
0 51792 7 1 2 51788 51791
0 51793 5 1 1 51792
0 51794 7 1 2 69641 51793
0 51795 5 1 1 51794
0 51796 7 1 2 86161 104754
0 51797 5 1 1 51796
0 51798 7 1 2 104746 51797
0 51799 5 1 1 51798
0 51800 7 1 2 64509 51799
0 51801 5 1 1 51800
0 51802 7 1 2 94579 104032
0 51803 5 1 1 51802
0 51804 7 1 2 51801 51803
0 51805 5 1 1 51804
0 51806 7 1 2 105195 51805
0 51807 5 1 1 51806
0 51808 7 2 2 84059 79479
0 51809 7 1 2 76430 106303
0 51810 7 1 2 102849 51809
0 51811 5 1 1 51810
0 51812 7 1 2 51807 51811
0 51813 7 1 2 51795 51812
0 51814 5 1 1 51813
0 51815 7 1 2 67798 51814
0 51816 5 1 1 51815
0 51817 7 1 2 68171 93195
0 51818 7 1 2 97544 104452
0 51819 7 1 2 51817 51818
0 51820 5 1 1 51819
0 51821 7 1 2 51816 51820
0 51822 7 1 2 51746 51821
0 51823 5 1 1 51822
0 51824 7 1 2 88603 51823
0 51825 5 1 1 51824
0 51826 7 1 2 51663 51825
0 51827 5 2 1 51826
0 51828 7 1 2 67450 106305
0 51829 5 1 1 51828
0 51830 7 1 2 65852 51829
0 51831 5 1 1 51830
0 51832 7 1 2 103005 104748
0 51833 5 1 1 51832
0 51834 7 1 2 103488 93859
0 51835 5 2 1 51834
0 51836 7 1 2 66379 81070
0 51837 7 1 2 106307 51836
0 51838 5 1 1 51837
0 51839 7 1 2 51833 51838
0 51840 5 1 1 51839
0 51841 7 1 2 73257 51840
0 51842 5 1 1 51841
0 51843 7 1 2 82639 81615
0 51844 5 1 1 51843
0 51845 7 1 2 68172 94904
0 51846 5 1 1 51845
0 51847 7 1 2 51844 51846
0 51848 5 1 1 51847
0 51849 7 1 2 101500 51848
0 51850 5 1 1 51849
0 51851 7 1 2 51842 51850
0 51852 5 1 1 51851
0 51853 7 1 2 72792 51852
0 51854 5 1 1 51853
0 51855 7 1 2 88752 84985
0 51856 7 1 2 84518 51855
0 51857 5 1 1 51856
0 51858 7 1 2 51854 51857
0 51859 5 1 1 51858
0 51860 7 1 2 88604 51859
0 51861 5 1 1 51860
0 51862 7 1 2 75459 103218
0 51863 5 1 1 51862
0 51864 7 1 2 106100 51863
0 51865 5 1 1 51864
0 51866 7 1 2 81071 51865
0 51867 5 1 1 51866
0 51868 7 2 2 88003 77050
0 51869 7 1 2 87175 106309
0 51870 5 1 1 51869
0 51871 7 1 2 51867 51870
0 51872 5 1 1 51871
0 51873 7 1 2 72793 51872
0 51874 5 1 1 51873
0 51875 7 2 2 68173 105749
0 51876 5 1 1 106311
0 51877 7 1 2 83298 96076
0 51878 7 1 2 106312 51877
0 51879 5 1 1 51878
0 51880 7 1 2 51874 51879
0 51881 5 1 1 51880
0 51882 7 1 2 88605 51881
0 51883 5 1 1 51882
0 51884 7 2 2 86257 89842
0 51885 5 1 1 106313
0 51886 7 1 2 93522 103709
0 51887 5 1 1 51886
0 51888 7 1 2 106314 51887
0 51889 5 1 1 51888
0 51890 7 1 2 51883 51889
0 51891 5 1 1 51890
0 51892 7 1 2 64879 51891
0 51893 5 1 1 51892
0 51894 7 1 2 67451 51893
0 51895 7 1 2 51861 51894
0 51896 5 1 1 51895
0 51897 7 1 2 85178 51896
0 51898 5 1 1 51897
0 51899 7 1 2 70908 51898
0 51900 5 1 1 51899
0 51901 7 1 2 97414 98678
0 51902 5 2 1 51901
0 51903 7 1 2 88606 95119
0 51904 5 1 1 51903
0 51905 7 1 2 106315 51904
0 51906 5 1 1 51905
0 51907 7 1 2 70269 51906
0 51908 5 1 1 51907
0 51909 7 1 2 76611 79169
0 51910 5 1 1 51909
0 51911 7 1 2 97415 82876
0 51912 5 1 1 51911
0 51913 7 1 2 51910 51912
0 51914 5 1 1 51913
0 51915 7 1 2 88247 51914
0 51916 5 1 1 51915
0 51917 7 1 2 80034 90151
0 51918 5 1 1 51917
0 51919 7 1 2 51916 51918
0 51920 7 1 2 51908 51919
0 51921 5 1 1 51920
0 51922 7 1 2 81782 51921
0 51923 5 1 1 51922
0 51924 7 1 2 94648 102986
0 51925 7 1 2 103169 51924
0 51926 5 1 1 51925
0 51927 7 1 2 51923 51926
0 51928 5 1 1 51927
0 51929 7 1 2 73588 51928
0 51930 5 1 1 51929
0 51931 7 1 2 86701 90492
0 51932 7 1 2 103261 51931
0 51933 5 1 1 51932
0 51934 7 1 2 51930 51933
0 51935 5 1 1 51934
0 51936 7 1 2 68174 51935
0 51937 5 1 1 51936
0 51938 7 2 2 69017 91137
0 51939 7 1 2 87340 78113
0 51940 7 1 2 106317 51939
0 51941 5 1 1 51940
0 51942 7 1 2 16782 51941
0 51943 5 1 1 51942
0 51944 7 1 2 75085 51943
0 51945 5 1 1 51944
0 51946 7 1 2 100065 92045
0 51947 5 1 1 51946
0 51948 7 1 2 51945 51947
0 51949 5 1 1 51948
0 51950 7 1 2 70004 51949
0 51951 5 1 1 51950
0 51952 7 1 2 78324 90274
0 51953 7 1 2 104503 51952
0 51954 5 1 1 51953
0 51955 7 1 2 51951 51954
0 51956 7 1 2 51937 51955
0 51957 5 1 1 51956
0 51958 7 1 2 67799 51957
0 51959 5 1 1 51958
0 51960 7 1 2 96730 90643
0 51961 5 1 1 51960
0 51962 7 1 2 77756 90267
0 51963 7 1 2 94168 51962
0 51964 5 1 1 51963
0 51965 7 1 2 51961 51964
0 51966 5 1 1 51965
0 51967 7 1 2 68519 51966
0 51968 5 1 1 51967
0 51969 7 1 2 87341 92618
0 51970 5 1 1 51969
0 51971 7 1 2 94447 51970
0 51972 5 1 1 51971
0 51973 7 1 2 71486 51972
0 51974 5 1 1 51973
0 51975 7 1 2 94484 90965
0 51976 5 1 1 51975
0 51977 7 1 2 51974 51976
0 51978 5 1 1 51977
0 51979 7 1 2 79927 51978
0 51980 5 1 1 51979
0 51981 7 1 2 51968 51980
0 51982 5 1 1 51981
0 51983 7 1 2 70270 51982
0 51984 5 1 1 51983
0 51985 7 1 2 75086 96458
0 51986 7 1 2 89879 51985
0 51987 5 1 1 51986
0 51988 7 1 2 51984 51987
0 51989 5 1 1 51988
0 51990 7 1 2 92674 51989
0 51991 5 1 1 51990
0 51992 7 1 2 51959 51991
0 51993 5 1 1 51992
0 51994 7 1 2 71188 51993
0 51995 5 1 1 51994
0 51996 7 2 2 82393 88607
0 51997 7 1 2 76341 106319
0 51998 5 1 1 51997
0 51999 7 1 2 106316 51998
0 52000 5 1 1 51999
0 52001 7 1 2 68175 52000
0 52002 5 1 1 52001
0 52003 7 1 2 93196 88608
0 52004 5 1 1 52003
0 52005 7 1 2 52002 52004
0 52006 5 1 1 52005
0 52007 7 1 2 85750 52006
0 52008 5 1 1 52007
0 52009 7 1 2 70005 81370
0 52010 5 1 1 52009
0 52011 7 1 2 87131 88609
0 52012 7 1 2 79996 52011
0 52013 7 1 2 52010 52012
0 52014 5 1 1 52013
0 52015 7 1 2 52008 52014
0 52016 5 1 1 52015
0 52017 7 1 2 70271 52016
0 52018 5 1 1 52017
0 52019 7 1 2 71487 87132
0 52020 7 1 2 90740 52019
0 52021 7 1 2 24491 52020
0 52022 5 1 1 52021
0 52023 7 1 2 52018 52022
0 52024 5 1 1 52023
0 52025 7 1 2 90866 52024
0 52026 5 1 1 52025
0 52027 7 1 2 72477 52026
0 52028 7 1 2 51995 52027
0 52029 5 1 1 52028
0 52030 7 1 2 51900 52029
0 52031 5 1 1 52030
0 52032 7 1 2 87086 105230
0 52033 5 1 1 52032
0 52034 7 1 2 97755 79262
0 52035 5 1 1 52034
0 52036 7 1 2 52033 52035
0 52037 5 1 1 52036
0 52038 7 1 2 85708 52037
0 52039 5 1 1 52038
0 52040 7 1 2 98280 98924
0 52041 7 1 2 94116 52040
0 52042 5 1 1 52041
0 52043 7 1 2 52039 52042
0 52044 5 1 1 52043
0 52045 7 1 2 88610 52044
0 52046 5 1 1 52045
0 52047 7 1 2 82657 16079
0 52048 5 1 1 52047
0 52049 7 2 2 79858 52048
0 52050 5 1 1 106321
0 52051 7 1 2 71189 52050
0 52052 5 1 1 52051
0 52053 7 1 2 106283 52052
0 52054 5 1 1 52053
0 52055 7 1 2 78390 52054
0 52056 5 1 1 52055
0 52057 7 1 2 66380 52056
0 52058 5 1 1 52057
0 52059 7 2 2 82640 91435
0 52060 5 1 1 106323
0 52061 7 1 2 66082 106324
0 52062 5 1 1 52061
0 52063 7 1 2 52058 52062
0 52064 5 1 1 52063
0 52065 7 1 2 73258 52064
0 52066 5 1 1 52065
0 52067 7 1 2 79289 80001
0 52068 5 1 1 52067
0 52069 7 1 2 52066 52068
0 52070 5 1 1 52069
0 52071 7 1 2 72794 52070
0 52072 5 1 1 52071
0 52073 7 1 2 95216 106322
0 52074 5 1 1 52073
0 52075 7 1 2 67452 52074
0 52076 7 1 2 52072 52075
0 52077 5 1 1 52076
0 52078 7 1 2 70540 103262
0 52079 5 1 1 52078
0 52080 7 2 2 103489 52079
0 52081 5 1 1 106325
0 52082 7 1 2 66381 52081
0 52083 5 1 1 52082
0 52084 7 1 2 101591 103494
0 52085 5 1 1 52084
0 52086 7 1 2 75293 52085
0 52087 5 1 1 52086
0 52088 7 1 2 78839 52087
0 52089 7 1 2 52083 52088
0 52090 5 1 1 52089
0 52091 7 1 2 71190 52090
0 52092 5 1 1 52091
0 52093 7 1 2 86278 99831
0 52094 5 1 1 52093
0 52095 7 2 2 76342 81314
0 52096 5 1 1 106327
0 52097 7 1 2 66083 106328
0 52098 5 1 1 52097
0 52099 7 1 2 52094 52098
0 52100 5 1 1 52099
0 52101 7 1 2 70541 52100
0 52102 5 2 1 52101
0 52103 7 1 2 66382 103485
0 52104 5 1 1 52103
0 52105 7 1 2 81273 52104
0 52106 5 1 1 52105
0 52107 7 1 2 69642 52106
0 52108 5 1 1 52107
0 52109 7 1 2 106329 52108
0 52110 7 1 2 52092 52109
0 52111 5 1 1 52110
0 52112 7 1 2 68176 52111
0 52113 5 1 1 52112
0 52114 7 2 2 87133 79938
0 52115 5 2 1 106331
0 52116 7 1 2 101889 103495
0 52117 5 1 1 52116
0 52118 7 1 2 64880 52117
0 52119 5 1 1 52118
0 52120 7 1 2 81783 100702
0 52121 5 1 1 52120
0 52122 7 1 2 52119 52121
0 52123 5 2 1 52122
0 52124 7 1 2 77490 106335
0 52125 5 1 1 52124
0 52126 7 1 2 106333 52125
0 52127 5 1 1 52126
0 52128 7 1 2 74571 52127
0 52129 5 1 1 52128
0 52130 7 1 2 76612 79822
0 52131 5 1 1 52130
0 52132 7 1 2 1592 52131
0 52133 5 1 1 52132
0 52134 7 1 2 26299 52133
0 52135 7 1 2 52129 52134
0 52136 7 1 2 52113 52135
0 52137 5 1 1 52136
0 52138 7 1 2 67800 52137
0 52139 5 1 1 52138
0 52140 7 1 2 88359 44895
0 52141 5 1 1 52140
0 52142 7 1 2 76629 52141
0 52143 5 1 1 52142
0 52144 7 1 2 69643 106332
0 52145 5 1 1 52144
0 52146 7 1 2 52143 52145
0 52147 5 1 1 52146
0 52148 7 1 2 68177 52147
0 52149 5 1 1 52148
0 52150 7 1 2 72478 52149
0 52151 7 1 2 52139 52150
0 52152 5 1 1 52151
0 52153 7 1 2 88248 52152
0 52154 7 1 2 52077 52153
0 52155 5 1 1 52154
0 52156 7 1 2 52046 52155
0 52157 5 1 1 52156
0 52158 7 1 2 78274 52157
0 52159 5 1 1 52158
0 52160 7 1 2 77834 98831
0 52161 7 1 2 87978 52160
0 52162 5 1 1 52161
0 52163 7 1 2 91043 52162
0 52164 5 1 1 52163
0 52165 7 1 2 81072 52164
0 52166 5 1 1 52165
0 52167 7 1 2 80131 84612
0 52168 7 1 2 86479 95810
0 52169 7 1 2 52167 52168
0 52170 5 1 1 52169
0 52171 7 1 2 52166 52170
0 52172 5 1 1 52171
0 52173 7 1 2 72795 52172
0 52174 5 1 1 52173
0 52175 7 1 2 94096 94625
0 52176 5 1 1 52175
0 52177 7 1 2 90632 52176
0 52178 5 1 1 52177
0 52179 7 1 2 65506 52178
0 52180 5 1 1 52179
0 52181 7 1 2 75294 89732
0 52182 5 1 1 52181
0 52183 7 1 2 51486 52182
0 52184 5 1 1 52183
0 52185 7 1 2 104755 52184
0 52186 5 1 1 52185
0 52187 7 1 2 78275 97020
0 52188 5 1 1 52187
0 52189 7 1 2 52186 52188
0 52190 7 1 2 52180 52189
0 52191 5 1 1 52190
0 52192 7 1 2 95217 52191
0 52193 5 1 1 52192
0 52194 7 1 2 52174 52193
0 52195 5 1 1 52194
0 52196 7 1 2 67453 52195
0 52197 5 1 1 52196
0 52198 7 1 2 103736 97226
0 52199 7 1 2 91121 52198
0 52200 5 1 1 52199
0 52201 7 1 2 52197 52200
0 52202 5 1 1 52201
0 52203 7 1 2 64881 52202
0 52204 5 1 1 52203
0 52205 7 1 2 104063 85179
0 52206 5 1 1 52205
0 52207 7 1 2 78281 52206
0 52208 5 1 1 52207
0 52209 7 1 2 88249 52208
0 52210 5 1 1 52209
0 52211 7 1 2 94497 90623
0 52212 5 1 1 52211
0 52213 7 1 2 52210 52212
0 52214 5 1 1 52213
0 52215 7 1 2 75295 52214
0 52216 5 1 1 52215
0 52217 7 1 2 79597 93849
0 52218 7 1 2 89623 52217
0 52219 5 1 1 52218
0 52220 7 1 2 52216 52219
0 52221 5 1 1 52220
0 52222 7 1 2 67454 93518
0 52223 7 1 2 52221 52222
0 52224 5 1 1 52223
0 52225 7 1 2 52204 52224
0 52226 5 1 1 52225
0 52227 7 1 2 75024 52226
0 52228 5 1 1 52227
0 52229 7 1 2 89641 103980
0 52230 5 1 1 52229
0 52231 7 1 2 81089 89909
0 52232 5 1 1 52231
0 52233 7 1 2 52230 52232
0 52234 5 1 1 52233
0 52235 7 1 2 85709 52234
0 52236 5 1 1 52235
0 52237 7 1 2 85831 79452
0 52238 7 1 2 98903 52237
0 52239 7 1 2 94528 52238
0 52240 5 1 1 52239
0 52241 7 1 2 52236 52240
0 52242 5 1 1 52241
0 52243 7 1 2 75940 52242
0 52244 5 1 1 52243
0 52245 7 1 2 71488 95989
0 52246 5 1 1 52245
0 52247 7 1 2 38347 52246
0 52248 5 1 1 52247
0 52249 7 1 2 101524 90551
0 52250 7 1 2 52248 52249
0 52251 5 1 1 52250
0 52252 7 1 2 52244 52251
0 52253 5 1 1 52252
0 52254 7 1 2 96768 52253
0 52255 5 1 1 52254
0 52256 7 1 2 101106 92716
0 52257 5 1 1 52256
0 52258 7 1 2 97743 90493
0 52259 5 1 1 52258
0 52260 7 1 2 52257 52259
0 52261 5 1 1 52260
0 52262 7 1 2 73259 52261
0 52263 5 1 1 52262
0 52264 7 2 2 97744 80260
0 52265 7 1 2 88611 106337
0 52266 5 1 1 52265
0 52267 7 1 2 52263 52266
0 52268 5 1 1 52267
0 52269 7 1 2 80754 52268
0 52270 5 1 1 52269
0 52271 7 2 2 99177 84600
0 52272 7 1 2 87913 76713
0 52273 7 1 2 106339 52272
0 52274 5 1 1 52273
0 52275 7 1 2 52270 52274
0 52276 5 1 1 52275
0 52277 7 1 2 78276 52276
0 52278 5 1 1 52277
0 52279 7 1 2 87169 84155
0 52280 7 2 2 67009 102750
0 52281 7 1 2 103349 106341
0 52282 7 1 2 52279 52281
0 52283 5 1 1 52282
0 52284 7 1 2 52278 52283
0 52285 5 1 1 52284
0 52286 7 1 2 73589 52285
0 52287 5 1 1 52286
0 52288 7 2 2 97416 79355
0 52289 7 1 2 82765 106343
0 52290 5 1 1 52289
0 52291 7 2 2 84492 74252
0 52292 7 1 2 79290 87418
0 52293 7 1 2 106345 52292
0 52294 5 1 1 52293
0 52295 7 1 2 52290 52294
0 52296 5 1 1 52295
0 52297 7 1 2 71191 52296
0 52298 5 1 1 52297
0 52299 7 1 2 92782 90683
0 52300 7 1 2 87974 52299
0 52301 5 1 1 52300
0 52302 7 1 2 52298 52301
0 52303 5 1 1 52302
0 52304 7 1 2 98035 52303
0 52305 5 1 1 52304
0 52306 7 2 2 63931 97440
0 52307 7 1 2 89594 106347
0 52308 7 1 2 81547 52307
0 52309 5 1 1 52308
0 52310 7 1 2 52305 52309
0 52311 5 1 1 52310
0 52312 7 1 2 85710 52311
0 52313 5 1 1 52312
0 52314 7 1 2 86296 88612
0 52315 5 1 1 52314
0 52316 7 1 2 89849 52315
0 52317 5 1 1 52316
0 52318 7 1 2 67455 75025
0 52319 7 1 2 90085 52318
0 52320 7 1 2 104330 52319
0 52321 7 1 2 52317 52320
0 52322 5 1 1 52321
0 52323 7 1 2 52313 52322
0 52324 7 1 2 52287 52323
0 52325 5 1 1 52324
0 52326 7 1 2 67801 52325
0 52327 5 1 1 52326
0 52328 7 1 2 52255 52327
0 52329 5 1 1 52328
0 52330 7 1 2 74697 52329
0 52331 5 1 1 52330
0 52332 7 1 2 52228 52331
0 52333 7 1 2 52159 52332
0 52334 7 1 2 52031 52333
0 52335 5 1 1 52334
0 52336 7 1 2 51831 52335
0 52337 5 1 1 52336
0 52338 7 1 2 69289 52337
0 52339 5 1 1 52338
0 52340 7 1 2 99455 106306
0 52341 5 1 1 52340
0 52342 7 1 2 78186 106270
0 52343 5 1 1 52342
0 52344 7 1 2 77702 77841
0 52345 7 1 2 90166 52344
0 52346 5 1 1 52345
0 52347 7 1 2 52343 52346
0 52348 5 1 1 52347
0 52349 7 1 2 80755 52348
0 52350 5 1 1 52349
0 52351 7 1 2 102125 75838
0 52352 7 1 2 104437 52351
0 52353 5 1 1 52352
0 52354 7 1 2 52350 52353
0 52355 5 1 1 52354
0 52356 7 1 2 98703 52355
0 52357 5 1 1 52356
0 52358 7 1 2 64204 52357
0 52359 7 1 2 52341 52358
0 52360 5 1 1 52359
0 52361 7 1 2 52339 52360
0 52362 5 1 1 52361
0 52363 7 1 2 105543 106196
0 52364 5 1 1 52363
0 52365 7 1 2 70006 89049
0 52366 5 1 1 52365
0 52367 7 5 2 68520 96569
0 52368 7 1 2 64882 106349
0 52369 5 1 1 52368
0 52370 7 1 2 52366 52369
0 52371 5 4 1 52370
0 52372 7 1 2 99759 106354
0 52373 5 1 1 52372
0 52374 7 1 2 52364 52373
0 52375 5 1 1 52374
0 52376 7 1 2 71192 52375
0 52377 5 1 1 52376
0 52378 7 1 2 69644 105541
0 52379 7 1 2 106197 52378
0 52380 5 1 1 52379
0 52381 7 1 2 52377 52380
0 52382 5 1 1 52381
0 52383 7 1 2 95572 52382
0 52384 5 1 1 52383
0 52385 7 1 2 86123 48187
0 52386 5 1 1 52385
0 52387 7 2 2 86829 52386
0 52388 5 1 1 106358
0 52389 7 1 2 96769 52388
0 52390 5 1 1 52389
0 52391 7 2 2 97061 102908
0 52392 7 1 2 70542 106360
0 52393 5 1 1 52392
0 52394 7 1 2 52390 52393
0 52395 5 1 1 52394
0 52396 7 1 2 70909 52395
0 52397 5 1 1 52396
0 52398 7 1 2 80909 105272
0 52399 5 1 1 52398
0 52400 7 1 2 52397 52399
0 52401 5 1 1 52400
0 52402 7 1 2 69290 52401
0 52403 5 1 1 52402
0 52404 7 1 2 80910 104479
0 52405 5 1 1 52404
0 52406 7 1 2 52403 52405
0 52407 5 1 1 52406
0 52408 7 1 2 81073 52407
0 52409 5 1 1 52408
0 52410 7 1 2 67802 106359
0 52411 5 1 1 52410
0 52412 7 1 2 72796 105962
0 52413 5 1 1 52412
0 52414 7 1 2 103619 52413
0 52415 7 1 2 52411 52414
0 52416 5 1 1 52415
0 52417 7 1 2 52409 52416
0 52418 5 1 1 52417
0 52419 7 1 2 85180 52418
0 52420 5 1 1 52419
0 52421 7 1 2 52384 52420
0 52422 5 1 1 52421
0 52423 7 1 2 88613 52422
0 52424 5 1 1 52423
0 52425 7 1 2 98816 45283
0 52426 5 1 1 52425
0 52427 7 1 2 70007 52426
0 52428 5 1 1 52427
0 52429 7 1 2 97284 98058
0 52430 5 1 1 52429
0 52431 7 1 2 52428 52430
0 52432 5 1 1 52431
0 52433 7 1 2 73590 52432
0 52434 5 1 1 52433
0 52435 7 1 2 74698 74079
0 52436 7 1 2 92357 52435
0 52437 5 1 1 52436
0 52438 7 1 2 52434 52437
0 52439 5 1 1 52438
0 52440 7 1 2 81784 52439
0 52441 5 1 1 52440
0 52442 7 1 2 100047 105923
0 52443 5 1 1 52442
0 52444 7 1 2 81559 95252
0 52445 5 1 1 52444
0 52446 7 1 2 52443 52445
0 52447 5 1 1 52446
0 52448 7 1 2 70543 52447
0 52449 5 1 1 52448
0 52450 7 1 2 52441 52449
0 52451 5 1 1 52450
0 52452 7 1 2 69291 52451
0 52453 5 1 1 52452
0 52454 7 1 2 101044 106301
0 52455 5 1 1 52454
0 52456 7 1 2 52453 52455
0 52457 5 1 1 52456
0 52458 7 1 2 78277 52457
0 52459 5 1 1 52458
0 52460 7 2 2 84863 100031
0 52461 7 1 2 102056 104850
0 52462 7 1 2 106362 52461
0 52463 5 1 1 52462
0 52464 7 1 2 52459 52463
0 52465 5 1 1 52464
0 52466 7 1 2 67456 88250
0 52467 7 1 2 52465 52466
0 52468 5 1 1 52467
0 52469 7 1 2 52424 52468
0 52470 5 1 1 52469
0 52471 7 1 2 76097 52470
0 52472 5 1 1 52471
0 52473 7 1 2 85711 101389
0 52474 5 2 1 52473
0 52475 7 1 2 106326 106364
0 52476 5 3 1 52475
0 52477 7 1 2 98292 106366
0 52478 5 1 1 52477
0 52479 7 2 2 95089 86317
0 52480 5 1 1 106369
0 52481 7 1 2 86313 106370
0 52482 5 2 1 52481
0 52483 7 1 2 98281 106371
0 52484 5 1 1 52483
0 52485 7 1 2 52478 52484
0 52486 5 1 1 52485
0 52487 7 1 2 88614 52486
0 52488 5 1 1 52487
0 52489 7 1 2 97745 98639
0 52490 5 2 1 52489
0 52491 7 1 2 98243 104103
0 52492 5 1 1 52491
0 52493 7 1 2 106373 52492
0 52494 5 1 1 52493
0 52495 7 1 2 89843 52494
0 52496 5 1 1 52495
0 52497 7 1 2 52488 52496
0 52498 5 1 1 52497
0 52499 7 1 2 82472 52498
0 52500 5 1 1 52499
0 52501 7 1 2 83334 89844
0 52502 5 1 1 52501
0 52503 7 1 2 89130 105658
0 52504 5 1 1 52503
0 52505 7 1 2 52502 52504
0 52506 5 1 1 52505
0 52507 7 1 2 68521 52506
0 52508 5 1 1 52507
0 52509 7 1 2 96731 91919
0 52510 5 1 1 52509
0 52511 7 1 2 52508 52510
0 52512 5 1 1 52511
0 52513 7 1 2 65199 52512
0 52514 5 1 1 52513
0 52515 7 1 2 89839 52480
0 52516 5 1 1 52515
0 52517 7 1 2 52514 52516
0 52518 5 1 1 52517
0 52519 7 1 2 71193 106177
0 52520 7 1 2 52518 52519
0 52521 5 1 1 52520
0 52522 7 1 2 52500 52521
0 52523 5 1 1 52522
0 52524 7 1 2 74440 90086
0 52525 7 1 2 52523 52524
0 52526 5 1 1 52525
0 52527 7 1 2 97746 93191
0 52528 5 1 1 52527
0 52529 7 1 2 98244 90957
0 52530 7 1 2 106350 52529
0 52531 5 1 1 52530
0 52532 7 1 2 52528 52531
0 52533 5 1 1 52532
0 52534 7 1 2 82473 91024
0 52535 7 1 2 52533 52534
0 52536 5 1 1 52535
0 52537 7 1 2 52526 52536
0 52538 5 1 1 52537
0 52539 7 1 2 93021 52538
0 52540 5 1 1 52539
0 52541 7 1 2 52472 52540
0 52542 7 1 2 52362 52541
0 52543 5 1 1 52542
0 52544 7 1 2 89587 52543
0 52545 5 1 1 52544
0 52546 7 1 2 90678 91771
0 52547 5 1 1 52546
0 52548 7 1 2 88032 106273
0 52549 7 1 2 95861 52548
0 52550 7 1 2 106213 52549
0 52551 5 1 1 52550
0 52552 7 1 2 52547 52551
0 52553 5 1 1 52552
0 52554 7 1 2 70544 52553
0 52555 5 1 1 52554
0 52556 7 1 2 70691 100778
0 52557 7 2 2 70730 88710
0 52558 7 4 2 72191 79315
0 52559 7 1 2 95657 106377
0 52560 7 1 2 106375 52559
0 52561 7 1 2 52556 52560
0 52562 5 1 1 52561
0 52563 7 1 2 52555 52562
0 52564 5 1 1 52563
0 52565 7 1 2 96965 52564
0 52566 5 1 1 52565
0 52567 7 1 2 79170 104382
0 52568 7 1 2 93547 52567
0 52569 7 1 2 106214 52568
0 52570 7 1 2 100992 52569
0 52571 5 1 1 52570
0 52572 7 1 2 52566 52571
0 52573 5 1 1 52572
0 52574 7 1 2 64883 52573
0 52575 5 1 1 52574
0 52576 7 1 2 102958 93650
0 52577 7 1 2 90421 96200
0 52578 7 1 2 98102 52577
0 52579 7 1 2 52576 52578
0 52580 5 1 1 52579
0 52581 7 1 2 52575 52580
0 52582 5 1 1 52581
0 52583 7 1 2 73591 52582
0 52584 5 1 1 52583
0 52585 7 2 2 69292 79291
0 52586 7 1 2 97490 106381
0 52587 7 1 2 106228 52586
0 52588 5 1 1 52587
0 52589 7 1 2 52584 52588
0 52590 5 1 1 52589
0 52591 7 1 2 68178 52590
0 52592 5 1 1 52591
0 52593 7 1 2 78725 91890
0 52594 5 1 1 52593
0 52595 7 1 2 91580 52594
0 52596 5 1 1 52595
0 52597 7 1 2 64510 52596
0 52598 5 1 1 52597
0 52599 7 1 2 92155 99049
0 52600 5 1 1 52599
0 52601 7 1 2 91363 84381
0 52602 5 1 1 52601
0 52603 7 1 2 52600 52602
0 52604 5 1 1 52603
0 52605 7 1 2 87708 52604
0 52606 5 1 1 52605
0 52607 7 1 2 52598 52606
0 52608 5 1 1 52607
0 52609 7 1 2 96966 52608
0 52610 5 1 1 52609
0 52611 7 2 2 100302 88926
0 52612 5 1 1 106383
0 52613 7 1 2 21317 52612
0 52614 5 1 1 52613
0 52615 7 1 2 87237 52614
0 52616 5 1 1 52615
0 52617 7 1 2 97722 96513
0 52618 7 1 2 93994 52617
0 52619 5 1 1 52618
0 52620 7 1 2 52616 52619
0 52621 5 1 1 52620
0 52622 7 1 2 106132 52621
0 52623 5 1 1 52622
0 52624 7 1 2 52610 52623
0 52625 5 1 1 52624
0 52626 7 1 2 70008 52625
0 52627 5 1 1 52626
0 52628 7 4 2 92558 96356
0 52629 7 1 2 98594 77784
0 52630 7 1 2 106385 52629
0 52631 5 1 1 52630
0 52632 7 1 2 52627 52631
0 52633 5 1 1 52632
0 52634 7 1 2 80756 52633
0 52635 5 1 1 52634
0 52636 7 1 2 90540 105248
0 52637 5 1 1 52636
0 52638 7 1 2 96925 79037
0 52639 7 1 2 97016 52638
0 52640 5 1 1 52639
0 52641 7 1 2 52637 52640
0 52642 5 1 1 52641
0 52643 7 1 2 74699 52642
0 52644 5 1 1 52643
0 52645 7 2 2 72479 92826
0 52646 5 1 1 106389
0 52647 7 1 2 106378 106390
0 52648 5 1 1 52647
0 52649 7 2 2 63932 98149
0 52650 7 1 2 66788 97441
0 52651 7 2 2 106391 52650
0 52652 5 1 1 106393
0 52653 7 1 2 52648 52652
0 52654 5 1 1 52653
0 52655 7 1 2 70009 52654
0 52656 5 1 1 52655
0 52657 7 1 2 52644 52656
0 52658 5 1 1 52657
0 52659 7 1 2 73260 52658
0 52660 5 1 1 52659
0 52661 7 3 2 98150 102449
0 52662 5 1 1 106395
0 52663 7 1 2 75296 89482
0 52664 7 1 2 106396 52663
0 52665 5 1 1 52664
0 52666 7 1 2 52660 52665
0 52667 5 1 1 52666
0 52668 7 1 2 73592 52667
0 52669 5 1 1 52668
0 52670 7 1 2 96926 81170
0 52671 5 1 1 52670
0 52672 7 2 2 96967 86148
0 52673 5 1 1 106398
0 52674 7 1 2 73261 106399
0 52675 5 1 1 52674
0 52676 7 1 2 52671 52675
0 52677 5 1 1 52676
0 52678 7 1 2 88251 52677
0 52679 5 1 1 52678
0 52680 7 1 2 99035 93379
0 52681 7 1 2 84629 52680
0 52682 7 1 2 106379 52681
0 52683 5 1 1 52682
0 52684 7 1 2 52679 52683
0 52685 7 1 2 52669 52684
0 52686 5 1 1 52685
0 52687 7 1 2 88998 52686
0 52688 5 1 1 52687
0 52689 7 1 2 96968 106222
0 52690 5 1 1 52689
0 52691 7 1 2 100993 92827
0 52692 5 1 1 52691
0 52693 7 1 2 52690 52692
0 52694 5 1 1 52693
0 52695 7 1 2 72192 78667
0 52696 7 1 2 96700 52695
0 52697 7 1 2 94599 90503
0 52698 7 1 2 52696 52697
0 52699 7 1 2 52694 52698
0 52700 5 1 1 52699
0 52701 7 1 2 52688 52700
0 52702 7 1 2 52635 52701
0 52703 5 1 1 52702
0 52704 7 1 2 71489 52703
0 52705 5 1 1 52704
0 52706 7 1 2 91379 95877
0 52707 5 1 1 52706
0 52708 7 2 2 92135 106251
0 52709 7 1 2 91655 106400
0 52710 5 1 1 52709
0 52711 7 1 2 52707 52710
0 52712 5 1 1 52711
0 52713 7 1 2 96969 52712
0 52714 5 1 1 52713
0 52715 7 1 2 70731 91650
0 52716 7 2 2 69293 88033
0 52717 7 1 2 97458 106402
0 52718 7 1 2 52715 52717
0 52719 7 1 2 88444 52718
0 52720 5 1 1 52719
0 52721 7 1 2 52714 52720
0 52722 5 1 1 52721
0 52723 7 1 2 66383 52722
0 52724 5 1 1 52723
0 52725 7 4 2 97132 77778
0 52726 7 2 2 90309 105617
0 52727 7 1 2 97496 106408
0 52728 7 1 2 106404 52727
0 52729 5 1 1 52728
0 52730 7 1 2 52724 52729
0 52731 5 1 1 52730
0 52732 7 1 2 64884 52731
0 52733 5 1 1 52732
0 52734 7 2 2 99337 106386
0 52735 7 1 2 69645 75989
0 52736 5 1 1 52735
0 52737 7 1 2 105102 52736
0 52738 7 1 2 106410 52737
0 52739 5 1 1 52738
0 52740 7 1 2 52733 52739
0 52741 5 1 1 52740
0 52742 7 1 2 80757 52741
0 52743 5 1 1 52742
0 52744 7 2 2 63983 106133
0 52745 7 1 2 102081 94110
0 52746 7 1 2 106412 52745
0 52747 5 1 1 52746
0 52748 7 1 2 52743 52747
0 52749 7 1 2 52705 52748
0 52750 7 1 2 52592 52749
0 52751 5 1 1 52750
0 52752 7 1 2 85954 52751
0 52753 5 1 1 52752
0 52754 7 3 2 74201 88081
0 52755 5 1 1 106414
0 52756 7 1 2 84864 79171
0 52757 7 1 2 88999 52756
0 52758 5 1 1 52757
0 52759 7 1 2 52755 52758
0 52760 5 1 1 52759
0 52761 7 1 2 73593 52760
0 52762 5 1 1 52761
0 52763 7 1 2 98885 105523
0 52764 5 1 1 52763
0 52765 7 1 2 52762 52764
0 52766 5 1 1 52765
0 52767 7 1 2 65200 52766
0 52768 5 1 1 52767
0 52769 7 1 2 97618 106415
0 52770 5 1 1 52769
0 52771 7 1 2 52768 52770
0 52772 5 1 1 52771
0 52773 7 1 2 68179 52772
0 52774 5 1 1 52773
0 52775 7 1 2 106291 106416
0 52776 5 1 1 52775
0 52777 7 1 2 52774 52776
0 52778 5 1 1 52777
0 52779 7 1 2 88615 52778
0 52780 5 1 1 52779
0 52781 7 1 2 73262 97777
0 52782 5 1 1 52781
0 52783 7 1 2 104177 96491
0 52784 7 1 2 52782 52783
0 52785 5 1 1 52784
0 52786 7 1 2 99099 52785
0 52787 5 1 1 52786
0 52788 7 2 2 94169 88054
0 52789 7 1 2 87016 94783
0 52790 7 1 2 90526 52789
0 52791 7 1 2 106417 52790
0 52792 5 1 1 52791
0 52793 7 1 2 52787 52792
0 52794 5 1 1 52793
0 52795 7 1 2 73594 52794
0 52796 5 1 1 52795
0 52797 7 1 2 92650 93674
0 52798 7 1 2 106409 52797
0 52799 5 1 1 52798
0 52800 7 1 2 52796 52799
0 52801 5 1 1 52800
0 52802 7 1 2 88252 52801
0 52803 5 1 1 52802
0 52804 7 1 2 52780 52803
0 52805 5 1 1 52804
0 52806 7 1 2 72480 52805
0 52807 5 1 1 52806
0 52808 7 1 2 88354 89733
0 52809 5 1 1 52808
0 52810 7 1 2 51885 52809
0 52811 5 1 1 52810
0 52812 7 1 2 73263 52811
0 52813 5 1 1 52812
0 52814 7 1 2 83490 95968
0 52815 5 1 1 52814
0 52816 7 1 2 52813 52815
0 52817 5 1 1 52816
0 52818 7 3 2 64205 71964
0 52819 7 1 2 91175 106419
0 52820 7 1 2 105427 52819
0 52821 7 1 2 52817 52820
0 52822 5 1 1 52821
0 52823 7 1 2 52807 52822
0 52824 5 1 1 52823
0 52825 7 1 2 70010 52824
0 52826 5 1 1 52825
0 52827 7 1 2 96927 87348
0 52828 5 1 1 52827
0 52829 7 1 2 85378 98103
0 52830 5 1 1 52829
0 52831 7 1 2 52828 52830
0 52832 5 1 1 52831
0 52833 7 1 2 73595 52832
0 52834 5 1 1 52833
0 52835 7 1 2 52673 52834
0 52836 5 1 1 52835
0 52837 7 1 2 81218 52836
0 52838 5 1 1 52837
0 52839 7 1 2 102098 92011
0 52840 7 1 2 104390 52839
0 52841 5 1 1 52840
0 52842 7 1 2 52838 52841
0 52843 5 1 1 52842
0 52844 7 1 2 98855 52843
0 52845 5 1 1 52844
0 52846 7 1 2 52826 52845
0 52847 5 1 1 52846
0 52848 7 1 2 71490 52847
0 52849 5 1 1 52848
0 52850 7 1 2 82332 88253
0 52851 5 2 1 52850
0 52852 7 2 2 84865 90174
0 52853 5 1 1 106424
0 52854 7 1 2 106422 52853
0 52855 5 2 1 52854
0 52856 7 2 2 67457 105160
0 52857 7 1 2 106426 106428
0 52858 5 1 1 52857
0 52859 7 1 2 94236 98629
0 52860 7 1 2 91406 52859
0 52861 7 2 2 98868 52860
0 52862 5 1 1 106430
0 52863 7 1 2 52858 52862
0 52864 5 1 1 52863
0 52865 7 1 2 66600 52864
0 52866 5 1 1 52865
0 52867 7 1 2 52646 52662
0 52868 5 1 1 52867
0 52869 7 1 2 106218 52868
0 52870 5 1 1 52869
0 52871 7 1 2 52866 52870
0 52872 5 1 1 52871
0 52873 7 1 2 73596 52872
0 52874 5 1 1 52873
0 52875 7 1 2 94784 91176
0 52876 7 1 2 106215 52875
0 52877 7 1 2 106171 52876
0 52878 5 1 1 52877
0 52879 7 1 2 52874 52878
0 52880 5 1 1 52879
0 52881 7 1 2 68180 52880
0 52882 5 1 1 52881
0 52883 7 1 2 96928 94485
0 52884 5 1 1 52883
0 52885 7 1 2 96970 96562
0 52886 5 1 1 52885
0 52887 7 1 2 52884 52886
0 52888 5 1 1 52887
0 52889 7 1 2 106219 52888
0 52890 5 1 1 52889
0 52891 7 1 2 83121 93672
0 52892 7 1 2 96255 52891
0 52893 7 1 2 91843 106348
0 52894 7 1 2 52892 52893
0 52895 5 1 1 52894
0 52896 7 1 2 52890 52895
0 52897 5 1 1 52896
0 52898 7 1 2 73989 52897
0 52899 5 1 1 52898
0 52900 7 2 2 93314 106090
0 52901 7 1 2 98181 94017
0 52902 7 1 2 97317 52901
0 52903 7 1 2 106432 52902
0 52904 5 1 1 52903
0 52905 7 1 2 52899 52904
0 52906 7 1 2 52882 52905
0 52907 5 1 1 52906
0 52908 7 1 2 66384 52907
0 52909 5 1 1 52908
0 52910 7 1 2 90175 96996
0 52911 5 1 1 52910
0 52912 7 1 2 50136 52911
0 52913 5 1 1 52912
0 52914 7 2 2 97723 91177
0 52915 7 3 2 90375 106434
0 52916 7 1 2 94659 78668
0 52917 7 1 2 106436 52916
0 52918 7 1 2 52913 52917
0 52919 5 1 1 52918
0 52920 7 1 2 52909 52919
0 52921 5 1 1 52920
0 52922 7 1 2 64885 52921
0 52923 5 1 1 52922
0 52924 7 1 2 96997 106310
0 52925 5 1 1 52924
0 52926 7 1 2 96929 91144
0 52927 5 1 1 52926
0 52928 7 1 2 52925 52927
0 52929 5 1 1 52928
0 52930 7 1 2 88616 52929
0 52931 5 1 1 52930
0 52932 7 2 2 63933 95644
0 52933 7 1 2 89646 98161
0 52934 7 1 2 106439 52933
0 52935 5 1 1 52934
0 52936 7 1 2 52931 52935
0 52937 5 1 1 52936
0 52938 7 1 2 82641 106437
0 52939 7 1 2 52937 52938
0 52940 5 1 1 52939
0 52941 7 1 2 52923 52940
0 52942 7 1 2 52849 52941
0 52943 5 1 1 52942
0 52944 7 1 2 85335 52943
0 52945 5 1 1 52944
0 52946 7 1 2 52753 52945
0 52947 5 1 1 52946
0 52948 7 1 2 71194 52947
0 52949 5 1 1 52948
0 52950 7 1 2 98036 86427
0 52951 7 1 2 89366 52950
0 52952 7 1 2 94789 52951
0 52953 5 1 1 52952
0 52954 7 1 2 104684 93856
0 52955 5 1 1 52954
0 52956 7 1 2 84328 99240
0 52957 5 1 1 52956
0 52958 7 1 2 52955 52957
0 52959 5 1 1 52958
0 52960 7 1 2 92981 90565
0 52961 7 1 2 52959 52960
0 52962 5 1 1 52961
0 52963 7 1 2 52953 52962
0 52964 5 1 1 52963
0 52965 7 1 2 65507 52964
0 52966 5 1 1 52965
0 52967 7 1 2 89156 92982
0 52968 7 1 2 106405 52967
0 52969 7 1 2 106387 52968
0 52970 5 1 1 52969
0 52971 7 1 2 52966 52970
0 52972 5 1 1 52971
0 52973 7 1 2 83192 52972
0 52974 5 1 1 52973
0 52975 7 1 2 73264 87460
0 52976 7 1 2 105161 52975
0 52977 5 1 1 52976
0 52978 7 1 2 68181 93315
0 52979 7 1 2 106418 52978
0 52980 5 1 1 52979
0 52981 7 1 2 52977 52980
0 52982 5 1 1 52981
0 52983 7 1 2 67458 52982
0 52984 5 1 1 52983
0 52985 7 1 2 99533 89207
0 52986 5 2 1 52985
0 52987 7 5 2 98037 93575
0 52988 7 1 2 94600 106443
0 52989 7 1 2 106441 52988
0 52990 5 1 1 52989
0 52991 7 1 2 52984 52990
0 52992 5 1 1 52991
0 52993 7 1 2 88254 52992
0 52994 5 1 1 52993
0 52995 7 2 2 97198 93576
0 52996 7 3 2 105152 106448
0 52997 5 1 1 106450
0 52998 7 1 2 106429 106442
0 52999 5 1 1 52998
0 53000 7 1 2 52997 52999
0 53001 5 1 1 53000
0 53002 7 1 2 90129 53001
0 53003 5 1 1 53002
0 53004 7 1 2 52994 53003
0 53005 5 1 1 53004
0 53006 7 1 2 65201 53005
0 53007 5 1 1 53006
0 53008 7 1 2 91696 94343
0 53009 7 1 2 106444 53008
0 53010 5 1 1 53009
0 53011 7 1 2 97133 105162
0 53012 5 1 1 53011
0 53013 7 1 2 53010 53012
0 53014 5 1 1 53013
0 53015 7 1 2 88255 53014
0 53016 5 1 1 53015
0 53017 7 2 2 90322 106406
0 53018 7 1 2 64511 78082
0 53019 7 2 2 106453 53018
0 53020 5 1 1 106455
0 53021 7 1 2 70272 106456
0 53022 5 1 1 53021
0 53023 7 1 2 53016 53022
0 53024 5 1 1 53023
0 53025 7 1 2 81785 53024
0 53026 5 1 1 53025
0 53027 7 1 2 73265 106431
0 53028 5 1 1 53027
0 53029 7 1 2 53026 53028
0 53030 5 1 1 53029
0 53031 7 1 2 66601 53030
0 53032 5 1 1 53031
0 53033 7 1 2 53007 53032
0 53034 5 1 1 53033
0 53035 7 1 2 73597 53034
0 53036 5 1 1 53035
0 53037 7 1 2 94660 84245
0 53038 5 1 1 53037
0 53039 7 1 2 82033 88355
0 53040 5 1 1 53039
0 53041 7 1 2 53038 53040
0 53042 5 1 1 53041
0 53043 7 1 2 96930 53042
0 53044 5 1 1 53043
0 53045 7 1 2 96971 88362
0 53046 5 1 1 53045
0 53047 7 1 2 53044 53046
0 53048 5 1 1 53047
0 53049 7 1 2 98856 53048
0 53050 5 1 1 53049
0 53051 7 1 2 86224 99328
0 53052 7 1 2 84023 53051
0 53053 7 1 2 106205 53052
0 53054 5 1 1 53053
0 53055 7 1 2 53050 53054
0 53056 7 1 2 53036 53055
0 53057 5 1 1 53056
0 53058 7 1 2 85336 53057
0 53059 5 1 1 53058
0 53060 7 1 2 80758 106253
0 53061 5 1 1 53060
0 53062 7 1 2 106211 53061
0 53063 5 1 1 53062
0 53064 7 1 2 96972 53063
0 53065 5 1 1 53064
0 53066 7 1 2 106263 106451
0 53067 5 1 1 53066
0 53068 7 1 2 53065 53067
0 53069 5 1 1 53068
0 53070 7 1 2 73266 53069
0 53071 5 1 1 53070
0 53072 7 1 2 87709 106411
0 53073 5 1 1 53072
0 53074 7 1 2 70273 96998
0 53075 7 1 2 97252 53074
0 53076 7 1 2 92156 53075
0 53077 5 1 1 53076
0 53078 7 1 2 53073 53077
0 53079 5 1 1 53078
0 53080 7 1 2 80759 53079
0 53081 5 1 1 53080
0 53082 7 1 2 73598 106394
0 53083 5 1 1 53082
0 53084 7 1 2 6839 7312
0 53085 5 1 1 53084
0 53086 7 1 2 85712 53085
0 53087 5 1 1 53086
0 53088 7 1 2 85751 92795
0 53089 5 1 1 53088
0 53090 7 1 2 53087 53089
0 53091 5 1 1 53090
0 53092 7 1 2 96931 53091
0 53093 5 1 1 53092
0 53094 7 1 2 53083 53093
0 53095 5 1 1 53094
0 53096 7 1 2 89000 53095
0 53097 5 1 1 53096
0 53098 7 1 2 53081 53097
0 53099 5 1 1 53098
0 53100 7 1 2 68182 53099
0 53101 5 1 1 53100
0 53102 7 1 2 86170 79605
0 53103 7 1 2 105812 53102
0 53104 7 1 2 106413 53103
0 53105 5 1 1 53104
0 53106 7 1 2 53101 53105
0 53107 7 1 2 53071 53106
0 53108 5 1 1 53107
0 53109 7 1 2 85955 53108
0 53110 5 1 1 53109
0 53111 7 1 2 71195 53110
0 53112 7 1 2 53059 53111
0 53113 5 1 1 53112
0 53114 7 1 2 104438 90212
0 53115 5 1 1 53114
0 53116 7 1 2 80760 95742
0 53117 7 1 2 96871 53116
0 53118 7 1 2 105146 53117
0 53119 5 1 1 53118
0 53120 7 1 2 53115 53119
0 53121 5 1 1 53120
0 53122 7 1 2 88256 53121
0 53123 5 1 1 53122
0 53124 7 1 2 81786 96797
0 53125 5 1 1 53124
0 53126 7 1 2 77681 89372
0 53127 7 2 2 53125 53126
0 53128 7 1 2 89001 106457
0 53129 5 1 1 53128
0 53130 7 1 2 104081 92450
0 53131 7 1 2 106435 53130
0 53132 5 1 1 53131
0 53133 7 1 2 53129 53132
0 53134 5 1 1 53133
0 53135 7 1 2 89314 53134
0 53136 5 1 1 53135
0 53137 7 1 2 53123 53136
0 53138 5 1 1 53137
0 53139 7 1 2 69646 53138
0 53140 5 1 1 53139
0 53141 7 1 2 91697 95257
0 53142 7 2 2 93714 91560
0 53143 7 1 2 76863 106459
0 53144 7 1 2 53141 53143
0 53145 7 1 2 106235 53144
0 53146 5 1 1 53145
0 53147 7 1 2 53140 53146
0 53148 5 1 1 53147
0 53149 7 1 2 67459 53148
0 53150 5 1 1 53149
0 53151 7 5 2 85956 94440
0 53152 7 1 2 74572 106461
0 53153 5 1 1 53152
0 53154 7 1 2 75488 89315
0 53155 5 1 1 53154
0 53156 7 1 2 53153 53155
0 53157 5 1 1 53156
0 53158 7 1 2 68183 106452
0 53159 7 1 2 53157 53158
0 53160 5 1 1 53159
0 53161 7 1 2 66084 53160
0 53162 7 1 2 53150 53161
0 53163 5 1 1 53162
0 53164 7 1 2 53113 53163
0 53165 5 1 1 53164
0 53166 7 1 2 52974 53165
0 53167 5 1 1 53166
0 53168 7 1 2 97417 53167
0 53169 5 1 1 53168
0 53170 7 1 2 87207 98595
0 53171 5 1 1 53170
0 53172 7 1 2 77922 98475
0 53173 5 1 1 53172
0 53174 7 1 2 53171 53173
0 53175 5 1 1 53174
0 53176 7 1 2 68184 53175
0 53177 5 1 1 53176
0 53178 7 1 2 100933 103567
0 53179 5 1 1 53178
0 53180 7 1 2 53177 53179
0 53181 5 1 1 53180
0 53182 7 1 2 97017 53181
0 53183 5 1 1 53182
0 53184 7 1 2 64886 105842
0 53185 5 1 1 53184
0 53186 7 1 2 102605 53185
0 53187 5 2 1 53186
0 53188 7 2 2 97442 106466
0 53189 7 1 2 64512 84651
0 53190 7 1 2 106468 53189
0 53191 5 1 1 53190
0 53192 7 1 2 53183 53191
0 53193 5 1 1 53192
0 53194 7 1 2 65508 53193
0 53195 5 1 1 53194
0 53196 7 1 2 100790 88815
0 53197 5 1 1 53196
0 53198 7 2 2 76965 99178
0 53199 5 1 1 106470
0 53200 7 1 2 53197 53199
0 53201 5 1 1 53200
0 53202 7 1 2 92796 53201
0 53203 5 1 1 53202
0 53204 7 1 2 88356 93850
0 53205 7 1 2 106469 53204
0 53206 5 1 1 53205
0 53207 7 1 2 53203 53206
0 53208 7 1 2 53195 53207
0 53209 5 1 1 53208
0 53210 7 1 2 73599 53209
0 53211 5 1 1 53210
0 53212 7 1 2 69647 79045
0 53213 7 1 2 106340 53212
0 53214 5 1 1 53213
0 53215 7 1 2 79968 98596
0 53216 7 1 2 89845 53215
0 53217 5 1 1 53216
0 53218 7 1 2 53214 53217
0 53219 5 1 1 53218
0 53220 7 1 2 74700 53219
0 53221 5 1 1 53220
0 53222 7 1 2 101061 90494
0 53223 7 1 2 103584 53222
0 53224 5 1 1 53223
0 53225 7 1 2 53221 53224
0 53226 7 1 2 53211 53225
0 53227 5 1 1 53226
0 53228 7 1 2 69294 53227
0 53229 5 1 1 53228
0 53230 7 1 2 70011 103392
0 53231 5 1 1 53230
0 53232 7 1 2 80651 88445
0 53233 5 1 1 53232
0 53234 7 1 2 53231 53233
0 53235 5 1 1 53234
0 53236 7 1 2 99300 84329
0 53237 7 1 2 104535 53236
0 53238 7 1 2 53235 53237
0 53239 5 1 1 53238
0 53240 7 1 2 53229 53239
0 53241 5 1 1 53240
0 53242 7 1 2 88082 53241
0 53243 5 1 1 53242
0 53244 7 1 2 67460 105085
0 53245 7 1 2 93555 53244
0 53246 7 1 2 106264 53245
0 53247 5 1 1 53246
0 53248 7 1 2 53243 53247
0 53249 5 1 1 53248
0 53250 7 1 2 89435 53249
0 53251 5 1 1 53250
0 53252 7 1 2 90048 98618
0 53253 5 1 1 53252
0 53254 7 1 2 80168 87490
0 53255 5 1 1 53254
0 53256 7 1 2 80180 86830
0 53257 7 1 2 53255 53256
0 53258 5 1 1 53257
0 53259 7 1 2 98597 53258
0 53260 5 1 1 53259
0 53261 7 1 2 53253 53260
0 53262 5 1 1 53261
0 53263 7 1 2 88257 53262
0 53264 5 1 1 53263
0 53265 7 4 2 67461 80761
0 53266 7 1 2 90495 106472
0 53267 7 1 2 90163 53266
0 53268 5 1 1 53267
0 53269 7 1 2 53264 53268
0 53270 5 1 1 53269
0 53271 7 1 2 66085 53270
0 53272 5 1 1 53271
0 53273 7 1 2 64887 75489
0 53274 5 1 1 53273
0 53275 7 2 2 103490 53274
0 53276 5 1 1 106476
0 53277 7 1 2 102042 89880
0 53278 7 1 2 53276 53277
0 53279 5 1 1 53278
0 53280 7 1 2 53272 53279
0 53281 5 1 1 53280
0 53282 7 1 2 89002 53281
0 53283 5 1 1 53282
0 53284 7 1 2 104199 106223
0 53285 5 1 1 53284
0 53286 7 1 2 77516 100996
0 53287 5 1 1 53286
0 53288 7 1 2 53285 53287
0 53289 5 1 1 53288
0 53290 7 1 2 94772 53289
0 53291 5 1 1 53290
0 53292 7 1 2 87710 21795
0 53293 7 1 2 5614 42398
0 53294 5 1 1 53293
0 53295 7 1 2 94441 53294
0 53296 7 1 2 53292 53295
0 53297 5 1 1 53296
0 53298 7 1 2 53291 53297
0 53299 5 1 1 53298
0 53300 7 1 2 68185 53299
0 53301 5 1 1 53300
0 53302 7 1 2 91155 78726
0 53303 7 1 2 82018 53302
0 53304 7 1 2 106473 53303
0 53305 5 1 1 53304
0 53306 7 1 2 53301 53305
0 53307 5 1 1 53306
0 53308 7 1 2 91792 53307
0 53309 5 1 1 53308
0 53310 7 1 2 53283 53309
0 53311 5 1 1 53310
0 53312 7 1 2 69295 53311
0 53313 5 1 1 53312
0 53314 7 1 2 75990 91380
0 53315 5 1 1 53314
0 53316 7 1 2 91516 91935
0 53317 7 1 2 106401 53316
0 53318 5 1 1 53317
0 53319 7 1 2 53315 53318
0 53320 5 1 1 53319
0 53321 7 1 2 70012 53320
0 53322 5 1 1 53321
0 53323 7 2 2 69018 92031
0 53324 7 1 2 91422 106478
0 53325 5 1 1 53324
0 53326 7 1 2 53322 53325
0 53327 5 1 1 53326
0 53328 7 1 2 66086 53327
0 53329 5 1 1 53328
0 53330 7 1 2 106259 53329
0 53331 5 1 1 53330
0 53332 7 1 2 69648 53331
0 53333 5 1 1 53332
0 53334 7 1 2 74573 74317
0 53335 7 1 2 90552 53334
0 53336 7 1 2 95686 53335
0 53337 5 1 1 53336
0 53338 7 1 2 53333 53337
0 53339 5 1 1 53338
0 53340 7 1 2 80762 53339
0 53341 5 1 1 53340
0 53342 7 1 2 69649 91801
0 53343 7 1 2 80136 106216
0 53344 7 1 2 53342 53343
0 53345 7 1 2 106249 53344
0 53346 5 1 1 53345
0 53347 7 1 2 53341 53346
0 53348 5 1 1 53347
0 53349 7 1 2 96973 53348
0 53350 5 1 1 53349
0 53351 7 1 2 53313 53350
0 53352 5 1 1 53351
0 53353 7 1 2 85957 53352
0 53354 5 1 1 53353
0 53355 7 1 2 96932 75460
0 53356 7 1 2 96259 53355
0 53357 5 1 1 53356
0 53358 7 1 2 99525 93561
0 53359 7 1 2 87208 53358
0 53360 5 1 1 53359
0 53361 7 1 2 53357 53360
0 53362 5 1 1 53361
0 53363 7 1 2 70545 53362
0 53364 5 1 1 53363
0 53365 7 1 2 104685 97533
0 53366 7 1 2 105938 53365
0 53367 5 1 1 53366
0 53368 7 1 2 53364 53367
0 53369 5 1 1 53368
0 53370 7 1 2 99110 53369
0 53371 5 1 1 53370
0 53372 7 1 2 67803 53371
0 53373 7 1 2 53354 53372
0 53374 7 1 2 53251 53373
0 53375 7 1 2 53169 53374
0 53376 7 1 2 52949 53375
0 53377 5 1 1 53376
0 53378 7 2 2 72065 94436
0 53379 7 2 2 84360 87751
0 53380 7 1 2 104762 106482
0 53381 7 1 2 106480 53380
0 53382 5 1 1 53381
0 53383 7 1 2 85337 89711
0 53384 5 1 1 53383
0 53385 7 1 2 99683 94442
0 53386 5 1 1 53385
0 53387 7 1 2 53384 53386
0 53388 5 1 1 53387
0 53389 7 1 2 68186 101027
0 53390 7 1 2 53388 53389
0 53391 5 1 1 53390
0 53392 7 1 2 53382 53391
0 53393 5 1 1 53392
0 53394 7 1 2 71491 53393
0 53395 5 1 1 53394
0 53396 7 2 2 104410 106462
0 53397 7 1 2 101136 106484
0 53398 5 1 1 53397
0 53399 7 1 2 53395 53398
0 53400 5 1 1 53399
0 53401 7 1 2 88083 53400
0 53402 5 1 1 53401
0 53403 7 1 2 69650 101112
0 53404 5 1 1 53403
0 53405 7 1 2 76509 105412
0 53406 5 1 1 53405
0 53407 7 1 2 53404 53406
0 53408 5 3 1 53407
0 53409 7 1 2 89408 106486
0 53410 5 1 1 53409
0 53411 7 1 2 81124 93381
0 53412 5 1 1 53411
0 53413 7 1 2 53410 53412
0 53414 5 1 1 53413
0 53415 7 1 2 81787 89003
0 53416 7 1 2 53414 53415
0 53417 5 1 1 53416
0 53418 7 1 2 53402 53417
0 53419 5 1 1 53418
0 53420 7 1 2 73600 53419
0 53421 5 1 1 53420
0 53422 7 1 2 99233 84196
0 53423 7 2 2 93108 91899
0 53424 7 2 2 75763 91178
0 53425 7 1 2 106489 106491
0 53426 7 1 2 53422 53425
0 53427 7 1 2 94174 53426
0 53428 5 1 1 53427
0 53429 7 1 2 53421 53428
0 53430 5 1 1 53429
0 53431 7 1 2 67462 53430
0 53432 5 1 1 53431
0 53433 7 1 2 76714 103968
0 53434 7 1 2 102786 91646
0 53435 7 1 2 105472 106460
0 53436 7 1 2 53434 53435
0 53437 7 1 2 53433 53436
0 53438 5 1 1 53437
0 53439 7 1 2 53432 53438
0 53440 5 1 1 53439
0 53441 7 1 2 74701 53440
0 53442 5 1 1 53441
0 53443 7 1 2 101689 92427
0 53444 5 2 1 53443
0 53445 7 1 2 89409 106493
0 53446 5 1 1 53445
0 53447 7 2 2 101923 81074
0 53448 5 1 1 106495
0 53449 7 1 2 79480 90504
0 53450 5 1 1 53449
0 53451 7 1 2 53448 53450
0 53452 5 1 1 53451
0 53453 7 1 2 75297 89334
0 53454 7 1 2 53452 53453
0 53455 5 1 1 53454
0 53456 7 1 2 53446 53455
0 53457 5 1 1 53456
0 53458 7 1 2 69296 53457
0 53459 5 1 1 53458
0 53460 7 1 2 78130 80138
0 53461 7 1 2 89402 53460
0 53462 5 1 1 53461
0 53463 7 1 2 53459 53462
0 53464 5 1 1 53463
0 53465 7 1 2 88084 53464
0 53466 5 1 1 53465
0 53467 7 1 2 63984 79392
0 53468 7 2 2 75298 89549
0 53469 7 1 2 95468 106497
0 53470 7 1 2 53467 53469
0 53471 7 1 2 106487 53470
0 53472 5 1 1 53471
0 53473 7 1 2 53466 53472
0 53474 5 1 1 53473
0 53475 7 1 2 67463 53474
0 53476 5 1 1 53475
0 53477 7 1 2 95743 97199
0 53478 7 1 2 91390 53477
0 53479 7 2 2 79580 93625
0 53480 7 1 2 97319 105536
0 53481 7 1 2 106499 53480
0 53482 7 1 2 53478 53481
0 53483 5 1 1 53482
0 53484 7 1 2 53476 53483
0 53485 5 1 1 53484
0 53486 7 1 2 84866 53485
0 53487 5 1 1 53486
0 53488 7 1 2 76396 103317
0 53489 7 2 2 105647 53488
0 53490 7 1 2 71196 103585
0 53491 5 1 1 53490
0 53492 7 1 2 89917 91436
0 53493 5 1 1 53492
0 53494 7 1 2 4772 79294
0 53495 5 1 1 53494
0 53496 7 1 2 76098 53495
0 53497 5 1 1 53496
0 53498 7 1 2 53493 53497
0 53499 7 1 2 53491 53498
0 53500 5 1 1 53499
0 53501 7 1 2 106501 53500
0 53502 5 1 1 53501
0 53503 7 1 2 92089 79868
0 53504 5 1 1 53503
0 53505 7 1 2 81075 53504
0 53506 5 1 1 53505
0 53507 7 1 2 77878 104408
0 53508 5 1 1 53507
0 53509 7 1 2 81076 104393
0 53510 5 1 1 53509
0 53511 7 1 2 101494 53510
0 53512 5 1 1 53511
0 53513 7 1 2 71492 53512
0 53514 5 1 1 53513
0 53515 7 1 2 53508 53514
0 53516 7 1 2 53506 53515
0 53517 5 1 1 53516
0 53518 7 1 2 69297 53517
0 53519 5 1 1 53518
0 53520 7 1 2 74574 103532
0 53521 5 1 1 53520
0 53522 7 1 2 53519 53521
0 53523 5 1 1 53522
0 53524 7 1 2 91232 53523
0 53525 5 1 1 53524
0 53526 7 1 2 53502 53525
0 53527 5 1 1 53526
0 53528 7 1 2 101104 53527
0 53529 5 1 1 53528
0 53530 7 1 2 53487 53529
0 53531 5 1 1 53530
0 53532 7 1 2 73601 53531
0 53533 5 1 1 53532
0 53534 7 1 2 91233 105086
0 53535 5 1 1 53534
0 53536 7 1 2 91211 106344
0 53537 5 1 1 53536
0 53538 7 1 2 53535 53537
0 53539 5 1 1 53538
0 53540 7 1 2 66087 53539
0 53541 5 1 1 53540
0 53542 7 2 2 91623 105384
0 53543 7 1 2 79382 96147
0 53544 7 1 2 106503 53543
0 53545 5 1 1 53544
0 53546 7 1 2 53541 53545
0 53547 5 1 1 53546
0 53548 7 1 2 73267 53547
0 53549 5 1 1 53548
0 53550 7 1 2 82538 99108
0 53551 5 1 1 53550
0 53552 7 1 2 69298 53551
0 53553 7 1 2 53549 53552
0 53554 5 1 1 53553
0 53555 7 1 2 100939 91221
0 53556 5 1 1 53555
0 53557 7 1 2 95234 91322
0 53558 7 1 2 99254 53557
0 53559 7 1 2 99112 53558
0 53560 5 1 1 53559
0 53561 7 1 2 64206 53560
0 53562 7 1 2 53556 53561
0 53563 5 1 1 53562
0 53564 7 1 2 67464 53563
0 53565 7 1 2 53554 53564
0 53566 5 1 1 53565
0 53567 7 1 2 98245 89901
0 53568 7 2 2 93738 91900
0 53569 7 1 2 105153 106505
0 53570 7 1 2 53567 53569
0 53571 7 1 2 99962 53570
0 53572 5 1 1 53571
0 53573 7 1 2 53566 53572
0 53574 5 1 1 53573
0 53575 7 1 2 70546 53574
0 53576 5 1 1 53575
0 53577 7 1 2 74103 93626
0 53578 7 1 2 85616 53577
0 53579 7 1 2 100667 105038
0 53580 7 1 2 106490 53579
0 53581 7 1 2 53578 53580
0 53582 5 1 1 53581
0 53583 7 1 2 53576 53582
0 53584 5 1 1 53583
0 53585 7 1 2 75461 53584
0 53586 5 1 1 53585
0 53587 7 1 2 67465 106496
0 53588 5 1 1 53587
0 53589 7 1 2 71197 106471
0 53590 5 1 1 53589
0 53591 7 1 2 53588 53590
0 53592 5 1 1 53591
0 53593 7 1 2 91234 53592
0 53594 5 1 1 53593
0 53595 7 1 2 92596 99169
0 53596 7 1 2 91302 53595
0 53597 5 1 1 53596
0 53598 7 1 2 53594 53597
0 53599 5 1 1 53598
0 53600 7 1 2 74702 53599
0 53601 5 1 1 53600
0 53602 7 1 2 91651 105467
0 53603 7 2 2 98038 92136
0 53604 7 1 2 106500 106507
0 53605 7 1 2 53602 53604
0 53606 5 1 1 53605
0 53607 7 1 2 102751 91364
0 53608 7 1 2 106494 53607
0 53609 5 1 1 53608
0 53610 7 1 2 53606 53609
0 53611 5 1 1 53610
0 53612 7 1 2 85958 53611
0 53613 5 1 1 53612
0 53614 7 1 2 53601 53613
0 53615 5 1 1 53614
0 53616 7 1 2 69299 53615
0 53617 5 1 1 53616
0 53618 7 1 2 99329 74104
0 53619 7 1 2 92283 53618
0 53620 7 1 2 106498 53619
0 53621 7 1 2 106488 53620
0 53622 5 1 1 53621
0 53623 7 1 2 53617 53622
0 53624 5 1 1 53623
0 53625 7 1 2 85713 53624
0 53626 5 1 1 53625
0 53627 7 1 2 70013 92947
0 53628 7 1 2 83305 53627
0 53629 5 1 1 53628
0 53630 7 1 2 64888 99872
0 53631 5 1 1 53630
0 53632 7 1 2 106463 53631
0 53633 7 1 2 53629 53632
0 53634 5 1 1 53633
0 53635 7 1 2 80652 90857
0 53636 7 1 2 99505 53635
0 53637 5 1 1 53636
0 53638 7 1 2 53634 53637
0 53639 5 1 1 53638
0 53640 7 1 2 101028 53639
0 53641 5 1 1 53640
0 53642 7 1 2 64889 92090
0 53643 7 1 2 102585 53642
0 53644 5 1 1 53643
0 53645 7 1 2 103582 53644
0 53646 7 1 2 106485 53645
0 53647 5 1 1 53646
0 53648 7 1 2 53641 53647
0 53649 5 1 1 53648
0 53650 7 1 2 88085 53649
0 53651 5 1 1 53650
0 53652 7 1 2 101690 92432
0 53653 5 1 1 53652
0 53654 7 1 2 106502 53653
0 53655 5 1 1 53654
0 53656 7 1 2 53651 53655
0 53657 5 1 1 53656
0 53658 7 1 2 67466 53657
0 53659 5 1 1 53658
0 53660 7 3 2 67467 101029
0 53661 7 1 2 91222 106509
0 53662 5 1 1 53661
0 53663 7 1 2 98476 89902
0 53664 7 1 2 93631 106068
0 53665 7 1 2 106506 53664
0 53666 7 1 2 53663 53665
0 53667 5 1 1 53666
0 53668 7 1 2 53662 53667
0 53669 5 1 1 53668
0 53670 7 1 2 90049 53669
0 53671 5 1 1 53670
0 53672 7 1 2 72797 53671
0 53673 7 1 2 53659 53672
0 53674 7 1 2 53626 53673
0 53675 7 1 2 53586 53674
0 53676 7 1 2 53533 53675
0 53677 7 1 2 53442 53676
0 53678 5 1 1 53677
0 53679 7 1 2 70910 53678
0 53680 7 1 2 53377 53679
0 53681 5 1 1 53680
0 53682 7 2 2 98773 90213
0 53683 7 1 2 101532 106427
0 53684 5 1 1 53683
0 53685 7 3 2 72193 93739
0 53686 7 1 2 83350 84986
0 53687 7 1 2 106514 53686
0 53688 5 1 1 53687
0 53689 7 1 2 53684 53688
0 53690 5 1 1 53689
0 53691 7 1 2 70014 53690
0 53692 5 1 1 53691
0 53693 7 1 2 100444 99238
0 53694 7 1 2 105243 53693
0 53695 5 1 1 53694
0 53696 7 1 2 53692 53695
0 53697 5 1 1 53696
0 53698 7 1 2 69651 53697
0 53699 5 1 1 53698
0 53700 7 1 2 91138 76715
0 53701 7 1 2 94791 53700
0 53702 7 1 2 101168 53701
0 53703 5 1 1 53702
0 53704 7 1 2 53699 53703
0 53705 5 1 1 53704
0 53706 7 1 2 73602 53705
0 53707 5 1 1 53706
0 53708 7 1 2 66789 77504
0 53709 7 1 2 77757 53708
0 53710 7 2 2 64207 88004
0 53711 7 1 2 99255 106517
0 53712 7 1 2 53709 53711
0 53713 5 1 1 53712
0 53714 7 1 2 53707 53713
0 53715 5 1 1 53714
0 53716 7 1 2 66602 53715
0 53717 5 1 1 53716
0 53718 7 1 2 93610 77794
0 53719 7 1 2 88005 53718
0 53720 7 1 2 100641 91612
0 53721 7 1 2 53719 53720
0 53722 5 1 1 53721
0 53723 7 1 2 53717 53722
0 53724 5 1 1 53723
0 53725 7 1 2 106512 53724
0 53726 5 1 1 53725
0 53727 7 1 2 97134 81077
0 53728 7 1 2 75682 53727
0 53729 5 1 1 53728
0 53730 7 1 2 95284 84075
0 53731 7 1 2 106508 53730
0 53732 5 1 1 53731
0 53733 7 1 2 53729 53732
0 53734 5 1 1 53733
0 53735 7 1 2 63810 53734
0 53736 5 1 1 53735
0 53737 7 2 2 87419 97331
0 53738 7 1 2 98039 91640
0 53739 7 1 2 106519 53738
0 53740 5 1 1 53739
0 53741 7 1 2 53736 53740
0 53742 5 1 1 53741
0 53743 7 1 2 73875 53742
0 53744 5 1 1 53743
0 53745 7 3 2 98040 103322
0 53746 7 1 2 96214 106521
0 53747 5 1 1 53746
0 53748 7 1 2 53020 53747
0 53749 5 1 1 53748
0 53750 7 1 2 63811 53749
0 53751 5 1 1 53750
0 53752 7 1 2 97724 106134
0 53753 7 1 2 90386 53752
0 53754 5 1 1 53753
0 53755 7 1 2 53751 53754
0 53756 5 1 1 53755
0 53757 7 1 2 71198 53756
0 53758 5 1 1 53757
0 53759 7 1 2 94100 91426
0 53760 7 1 2 99241 98910
0 53761 7 1 2 53759 53760
0 53762 5 1 1 53761
0 53763 7 1 2 53758 53762
0 53764 7 1 2 53744 53763
0 53765 5 1 1 53764
0 53766 7 1 2 76241 53765
0 53767 5 1 1 53766
0 53768 7 1 2 101743 79393
0 53769 7 1 2 106454 53768
0 53770 5 1 1 53769
0 53771 7 2 2 75670 95586
0 53772 7 1 2 99242 106304
0 53773 7 1 2 106524 53772
0 53774 7 1 2 73876 53773
0 53775 5 1 1 53774
0 53776 7 1 2 53770 53775
0 53777 7 1 2 53767 53776
0 53778 5 1 1 53777
0 53779 7 1 2 70911 53778
0 53780 5 1 1 53779
0 53781 7 1 2 75861 96354
0 53782 5 1 1 53781
0 53783 7 2 2 91540 84032
0 53784 5 1 1 106526
0 53785 7 1 2 53782 53784
0 53786 5 1 1 53785
0 53787 7 1 2 82509 90898
0 53788 7 1 2 76943 53787
0 53789 7 1 2 106407 53788
0 53790 7 1 2 53786 53789
0 53791 5 1 1 53790
0 53792 7 1 2 53780 53791
0 53793 5 1 1 53792
0 53794 7 1 2 84421 53793
0 53795 5 1 1 53794
0 53796 7 1 2 95622 104619
0 53797 7 1 2 98966 53796
0 53798 7 1 2 91698 84496
0 53799 7 1 2 97320 53798
0 53800 7 1 2 53797 53799
0 53801 5 1 1 53800
0 53802 7 1 2 53795 53801
0 53803 5 1 1 53802
0 53804 7 1 2 101220 53803
0 53805 5 1 1 53804
0 53806 7 1 2 53726 53805
0 53807 7 1 2 53681 53806
0 53808 7 2 2 79394 106302
0 53809 7 1 2 103981 106528
0 53810 5 1 1 53809
0 53811 7 1 2 102850 78550
0 53812 5 1 1 53811
0 53813 7 1 2 14883 53812
0 53814 5 2 1 53813
0 53815 7 1 2 81090 106530
0 53816 5 1 1 53815
0 53817 7 3 2 76859 89131
0 53818 7 1 2 84412 106532
0 53819 7 1 2 106236 53818
0 53820 5 1 1 53819
0 53821 7 1 2 53816 53820
0 53822 5 1 1 53821
0 53823 7 1 2 79153 53822
0 53824 5 1 1 53823
0 53825 7 1 2 53810 53824
0 53826 5 1 1 53825
0 53827 7 1 2 67804 53826
0 53828 5 1 1 53827
0 53829 7 1 2 92675 76864
0 53830 7 1 2 97577 53829
0 53831 7 1 2 102851 53830
0 53832 5 1 1 53831
0 53833 7 1 2 53828 53832
0 53834 5 1 1 53833
0 53835 7 1 2 99593 53834
0 53836 5 1 1 53835
0 53837 7 2 2 79154 78551
0 53838 7 2 2 75462 106474
0 53839 7 1 2 64208 106537
0 53840 5 2 1 53839
0 53841 7 1 2 96933 96570
0 53842 5 1 1 53841
0 53843 7 1 2 106539 53842
0 53844 5 2 1 53843
0 53845 7 1 2 68522 106541
0 53846 5 1 1 53845
0 53847 7 1 2 96974 105346
0 53848 5 1 1 53847
0 53849 7 1 2 53846 53848
0 53850 5 1 1 53849
0 53851 7 1 2 92676 53850
0 53852 5 1 1 53851
0 53853 7 1 2 96975 82148
0 53854 7 1 2 106237 53853
0 53855 5 1 1 53854
0 53856 7 1 2 53852 53855
0 53857 5 1 1 53856
0 53858 7 1 2 106535 53857
0 53859 5 1 1 53858
0 53860 7 1 2 83335 85374
0 53861 7 1 2 86987 53860
0 53862 5 1 1 53861
0 53863 7 1 2 89036 86125
0 53864 5 1 1 53863
0 53865 7 1 2 76812 93715
0 53866 7 1 2 53864 53865
0 53867 5 1 1 53866
0 53868 7 1 2 53862 53867
0 53869 5 2 1 53868
0 53870 7 1 2 65202 106543
0 53871 5 1 1 53870
0 53872 7 3 2 84361 79795
0 53873 7 1 2 87477 106545
0 53874 5 1 1 53873
0 53875 7 1 2 53871 53874
0 53876 5 1 1 53875
0 53877 7 1 2 67805 53876
0 53878 5 1 1 53877
0 53879 7 1 2 97275 105960
0 53880 5 1 1 53879
0 53881 7 1 2 53878 53880
0 53882 5 1 1 53881
0 53883 7 1 2 72481 53882
0 53884 5 1 1 53883
0 53885 7 1 2 95417 98555
0 53886 7 1 2 104070 53885
0 53887 5 1 1 53886
0 53888 7 1 2 53884 53887
0 53889 5 1 1 53888
0 53890 7 1 2 75224 53889
0 53891 5 1 1 53890
0 53892 7 1 2 53859 53891
0 53893 5 1 1 53892
0 53894 7 1 2 69652 53893
0 53895 5 1 1 53894
0 53896 7 1 2 67468 92810
0 53897 7 1 2 79356 53896
0 53898 7 1 2 106529 53897
0 53899 5 1 1 53898
0 53900 7 1 2 53895 53899
0 53901 5 1 1 53900
0 53902 7 1 2 71199 53901
0 53903 5 1 1 53902
0 53904 7 2 2 94277 76771
0 53905 5 1 1 106548
0 53906 7 1 2 106546 106549
0 53907 5 1 1 53906
0 53908 7 1 2 75225 106544
0 53909 5 1 1 53908
0 53910 7 1 2 53907 53909
0 53911 5 1 1 53910
0 53912 7 1 2 65203 53911
0 53913 5 1 1 53912
0 53914 7 1 2 75196 94450
0 53915 5 2 1 53914
0 53916 7 1 2 85617 76772
0 53917 5 1 1 53916
0 53918 7 1 2 106550 53917
0 53919 5 1 1 53918
0 53920 7 1 2 66603 53919
0 53921 5 2 1 53920
0 53922 7 1 2 79078 90053
0 53923 5 1 1 53922
0 53924 7 1 2 106552 53923
0 53925 5 1 1 53924
0 53926 7 1 2 106547 53925
0 53927 5 1 1 53926
0 53928 7 1 2 53913 53927
0 53929 5 1 1 53928
0 53930 7 1 2 72798 53929
0 53931 5 1 1 53930
0 53932 7 1 2 98098 92996
0 53933 7 1 2 106531 53932
0 53934 5 1 1 53933
0 53935 7 1 2 53931 53934
0 53936 5 1 1 53935
0 53937 7 1 2 81078 53936
0 53938 5 1 1 53937
0 53939 7 6 2 93740 76860
0 53940 7 1 2 80763 79115
0 53941 7 2 2 101879 53940
0 53942 5 1 1 106560
0 53943 7 1 2 68523 106561
0 53944 5 1 1 53943
0 53945 7 1 2 83977 78887
0 53946 5 1 1 53945
0 53947 7 1 2 53944 53946
0 53948 5 1 1 53947
0 53949 7 1 2 75463 53948
0 53950 5 1 1 53949
0 53951 7 1 2 94958 53942
0 53952 5 1 1 53951
0 53953 7 1 2 74575 53952
0 53954 5 1 1 53953
0 53955 7 1 2 53950 53954
0 53956 5 1 1 53955
0 53957 7 1 2 72799 53956
0 53958 5 1 1 53957
0 53959 7 1 2 79116 94141
0 53960 7 1 2 106243 53959
0 53961 5 1 1 53960
0 53962 7 1 2 53958 53961
0 53963 5 1 1 53962
0 53964 7 1 2 66088 53963
0 53965 5 1 1 53964
0 53966 7 1 2 66896 83051
0 53967 7 1 2 92677 96057
0 53968 7 1 2 86011 53967
0 53969 7 1 2 53966 53968
0 53970 5 1 1 53969
0 53971 7 1 2 53965 53970
0 53972 5 1 1 53971
0 53973 7 1 2 106554 53972
0 53974 5 1 1 53973
0 53975 7 1 2 53938 53974
0 53976 5 1 1 53975
0 53977 7 1 2 67469 53976
0 53978 5 1 1 53977
0 53979 7 1 2 99554 81079
0 53980 7 1 2 87765 53979
0 53981 7 1 2 106361 53980
0 53982 5 1 1 53981
0 53983 7 1 2 53978 53982
0 53984 7 1 2 53903 53983
0 53985 5 1 1 53984
0 53986 7 1 2 70912 53985
0 53987 5 1 1 53986
0 53988 7 1 2 53836 53987
0 53989 5 1 1 53988
0 53990 7 1 2 76099 53989
0 53991 5 1 1 53990
0 53992 7 1 2 96571 76735
0 53993 5 1 1 53992
0 53994 7 2 2 84867 75774
0 53995 7 1 2 90259 106562
0 53996 5 1 1 53995
0 53997 7 1 2 53993 53996
0 53998 5 1 1 53997
0 53999 7 1 2 92759 53998
0 54000 5 1 1 53999
0 54001 7 1 2 77835 78352
0 54002 7 1 2 92213 54001
0 54003 7 1 2 104064 54002
0 54004 5 1 1 54003
0 54005 7 1 2 54000 54004
0 54006 5 1 1 54005
0 54007 7 1 2 71493 54006
0 54008 5 1 1 54007
0 54009 7 2 2 84868 84509
0 54010 7 1 2 90031 84437
0 54011 7 1 2 84559 54010
0 54012 7 1 2 106564 54011
0 54013 5 1 1 54012
0 54014 7 1 2 54008 54013
0 54015 5 1 1 54014
0 54016 7 1 2 70015 54015
0 54017 5 1 1 54016
0 54018 7 2 2 67140 87914
0 54019 7 1 2 84422 106566
0 54020 7 1 2 106565 54019
0 54021 7 1 2 101350 54020
0 54022 5 1 1 54021
0 54023 7 1 2 54017 54022
0 54024 5 2 1 54023
0 54025 7 1 2 106108 106568
0 54026 5 1 1 54025
0 54027 7 1 2 81986 86380
0 54028 5 1 1 54027
0 54029 7 2 2 66604 82333
0 54030 7 1 2 101225 87292
0 54031 7 1 2 106570 54030
0 54032 5 1 1 54031
0 54033 7 1 2 54028 54032
0 54034 5 1 1 54033
0 54035 7 1 2 97418 54034
0 54036 5 1 1 54035
0 54037 7 1 2 76613 79985
0 54038 7 1 2 95162 54037
0 54039 5 1 1 54038
0 54040 7 1 2 54036 54039
0 54041 5 1 1 54040
0 54042 7 1 2 68187 54041
0 54043 5 1 1 54042
0 54044 7 1 2 88731 80139
0 54045 5 1 1 54044
0 54046 7 1 2 54043 54045
0 54047 5 1 1 54046
0 54048 7 1 2 72482 54047
0 54049 5 1 1 54048
0 54050 7 1 2 97747 94175
0 54051 7 1 2 106467 54050
0 54052 5 1 1 54051
0 54053 7 1 2 54049 54052
0 54054 5 1 1 54053
0 54055 7 1 2 73603 54054
0 54056 5 1 1 54055
0 54057 7 1 2 74703 106338
0 54058 5 1 1 54057
0 54059 7 1 2 81987 103279
0 54060 7 1 2 101342 54059
0 54061 5 1 1 54060
0 54062 7 1 2 54058 54061
0 54063 5 1 1 54062
0 54064 7 1 2 73268 54063
0 54065 5 1 1 54064
0 54066 7 1 2 92525 98104
0 54067 5 1 1 54066
0 54068 7 1 2 54065 54067
0 54069 5 1 1 54068
0 54070 7 1 2 84869 54069
0 54071 5 1 1 54070
0 54072 7 1 2 54056 54071
0 54073 5 1 1 54072
0 54074 7 1 2 74121 54073
0 54075 5 1 1 54074
0 54076 7 1 2 76100 106355
0 54077 5 1 1 54076
0 54078 7 1 2 97362 104872
0 54079 5 1 1 54078
0 54080 7 1 2 99850 106351
0 54081 5 1 1 54080
0 54082 7 1 2 54079 54081
0 54083 7 1 2 54077 54082
0 54084 5 1 1 54083
0 54085 7 1 2 87609 98630
0 54086 7 1 2 54084 54085
0 54087 5 1 1 54086
0 54088 7 1 2 67806 54087
0 54089 7 1 2 54075 54088
0 54090 5 1 1 54089
0 54091 7 1 2 89050 99170
0 54092 5 1 1 54091
0 54093 7 1 2 72483 77545
0 54094 7 1 2 106352 54093
0 54095 5 1 1 54094
0 54096 7 1 2 54092 54095
0 54097 5 1 1 54096
0 54098 7 1 2 71200 54097
0 54099 5 1 1 54098
0 54100 7 1 2 80653 78899
0 54101 5 1 1 54100
0 54102 7 1 2 86114 54101
0 54103 5 1 1 54102
0 54104 7 1 2 104581 54103
0 54105 5 1 1 54104
0 54106 7 1 2 54099 54105
0 54107 5 1 1 54106
0 54108 7 1 2 76736 54107
0 54109 5 1 1 54108
0 54110 7 1 2 80840 98192
0 54111 7 1 2 96804 54110
0 54112 5 1 1 54111
0 54113 7 1 2 106374 54112
0 54114 5 1 1 54113
0 54115 7 1 2 74979 54114
0 54116 5 1 1 54115
0 54117 7 1 2 67470 100553
0 54118 7 1 2 92005 54117
0 54119 5 1 1 54118
0 54120 7 1 2 54116 54119
0 54121 5 1 1 54120
0 54122 7 1 2 84870 74122
0 54123 7 1 2 54121 54122
0 54124 5 1 1 54123
0 54125 7 1 2 72800 54124
0 54126 7 1 2 54109 54125
0 54127 5 1 1 54126
0 54128 7 1 2 70913 54127
0 54129 7 1 2 54090 54128
0 54130 5 1 1 54129
0 54131 7 1 2 54026 54130
0 54132 5 1 1 54131
0 54133 7 1 2 69300 54132
0 54134 5 1 1 54133
0 54135 7 1 2 77491 99866
0 54136 5 1 1 54135
0 54137 7 1 2 90361 54136
0 54138 5 1 1 54137
0 54139 7 2 2 85554 54138
0 54140 7 1 2 98774 77740
0 54141 7 1 2 106572 54140
0 54142 5 1 1 54141
0 54143 7 1 2 95645 98454
0 54144 7 1 2 99256 54143
0 54145 7 1 2 95156 54144
0 54146 5 1 1 54145
0 54147 7 1 2 54142 54146
0 54148 5 1 1 54147
0 54149 7 1 2 75464 54148
0 54150 5 1 1 54149
0 54151 7 1 2 70016 105371
0 54152 5 1 1 54151
0 54153 7 1 2 8126 54152
0 54154 5 1 1 54153
0 54155 7 1 2 105916 54154
0 54156 5 1 1 54155
0 54157 7 1 2 74576 106573
0 54158 5 1 1 54157
0 54159 7 1 2 79969 100523
0 54160 5 1 1 54159
0 54161 7 1 2 54158 54160
0 54162 5 1 1 54161
0 54163 7 1 2 67807 54162
0 54164 5 1 1 54163
0 54165 7 1 2 54156 54164
0 54166 5 1 1 54165
0 54167 7 1 2 102752 54166
0 54168 5 1 1 54167
0 54169 7 1 2 84273 105280
0 54170 5 1 1 54169
0 54171 7 1 2 95526 97481
0 54172 7 1 2 93497 54171
0 54173 5 1 1 54172
0 54174 7 1 2 54170 54173
0 54175 5 1 1 54174
0 54176 7 1 2 64890 54175
0 54177 5 1 1 54176
0 54178 7 1 2 95342 102753
0 54179 7 1 2 102527 54178
0 54180 5 1 1 54179
0 54181 7 1 2 54177 54180
0 54182 5 1 1 54181
0 54183 7 1 2 64209 54182
0 54184 5 1 1 54183
0 54185 7 1 2 99963 74080
0 54186 5 1 1 54185
0 54187 7 1 2 80169 98714
0 54188 5 1 1 54187
0 54189 7 1 2 54186 54188
0 54190 5 1 1 54189
0 54191 7 1 2 102322 84624
0 54192 7 1 2 54190 54191
0 54193 5 1 1 54192
0 54194 7 1 2 54184 54193
0 54195 5 1 1 54194
0 54196 7 1 2 87711 54195
0 54197 5 1 1 54196
0 54198 7 1 2 54168 54197
0 54199 5 1 1 54198
0 54200 7 1 2 77738 54199
0 54201 5 1 1 54200
0 54202 7 1 2 54150 54201
0 54203 5 1 1 54202
0 54204 7 1 2 80764 54203
0 54205 5 1 1 54204
0 54206 7 1 2 70914 103907
0 54207 7 1 2 106569 54206
0 54208 5 1 1 54207
0 54209 7 1 2 95326 95390
0 54210 7 1 2 105773 54209
0 54211 7 1 2 104439 54210
0 54212 5 1 1 54211
0 54213 7 1 2 54208 54212
0 54214 5 1 1 54213
0 54215 7 1 2 64210 54214
0 54216 5 1 1 54215
0 54217 7 1 2 54205 54216
0 54218 7 1 2 54134 54217
0 54219 5 1 1 54218
0 54220 7 1 2 74041 54219
0 54221 5 1 1 54220
0 54222 7 1 2 66385 106367
0 54223 5 1 1 54222
0 54224 7 1 2 85714 92920
0 54225 5 1 1 54224
0 54226 7 1 2 93860 54225
0 54227 5 1 1 54226
0 54228 7 1 2 64891 54227
0 54229 5 1 1 54228
0 54230 7 1 2 87264 54229
0 54231 7 1 2 54223 54230
0 54232 5 1 1 54231
0 54233 7 1 2 106555 54232
0 54234 5 1 1 54233
0 54235 7 1 2 84046 88007
0 54236 7 1 2 106363 54235
0 54237 5 1 1 54236
0 54238 7 1 2 54234 54237
0 54239 5 1 1 54238
0 54240 7 1 2 67808 54239
0 54241 5 1 1 54240
0 54242 7 1 2 84105 106556
0 54243 7 1 2 86988 54242
0 54244 5 1 1 54243
0 54245 7 1 2 54241 54244
0 54246 5 1 1 54245
0 54247 7 1 2 71201 54246
0 54248 5 1 1 54247
0 54249 7 1 2 73604 99827
0 54250 5 1 1 54249
0 54251 7 1 2 106330 54250
0 54252 5 1 1 54251
0 54253 7 2 2 67809 106557
0 54254 7 1 2 54252 106574
0 54255 5 1 1 54254
0 54256 7 1 2 54248 54255
0 54257 5 1 1 54256
0 54258 7 1 2 68188 54257
0 54259 5 1 1 54258
0 54260 7 1 2 76052 97829
0 54261 5 1 1 54260
0 54262 7 1 2 80085 87072
0 54263 5 1 1 54262
0 54264 7 1 2 54261 54263
0 54265 5 1 1 54264
0 54266 7 1 2 70017 54265
0 54267 5 1 1 54266
0 54268 7 1 2 70274 99510
0 54269 5 1 1 54268
0 54270 7 1 2 54267 54269
0 54271 5 1 1 54270
0 54272 7 1 2 73605 54271
0 54273 5 1 1 54272
0 54274 7 1 2 76242 106285
0 54275 5 1 1 54274
0 54276 7 1 2 54273 54275
0 54277 5 1 1 54276
0 54278 7 1 2 71202 54277
0 54279 5 1 1 54278
0 54280 7 1 2 69653 106336
0 54281 5 1 1 54280
0 54282 7 1 2 106334 54281
0 54283 5 1 1 54282
0 54284 7 1 2 74577 54283
0 54285 5 1 1 54284
0 54286 7 1 2 54279 54285
0 54287 5 1 1 54286
0 54288 7 1 2 106575 54287
0 54289 5 1 1 54288
0 54290 7 1 2 54259 54289
0 54291 5 1 1 54290
0 54292 7 1 2 70915 54291
0 54293 5 1 1 54292
0 54294 7 1 2 94741 106423
0 54295 5 1 1 54294
0 54296 7 1 2 93296 54295
0 54297 5 1 1 54296
0 54298 7 1 2 68189 87293
0 54299 5 1 1 54298
0 54300 7 1 2 88258 54299
0 54301 5 1 1 54300
0 54302 7 1 2 96617 88617
0 54303 5 1 1 54302
0 54304 7 1 2 54301 54303
0 54305 5 1 1 54304
0 54306 7 1 2 66386 54305
0 54307 5 1 1 54306
0 54308 7 1 2 65204 90094
0 54309 5 1 1 54308
0 54310 7 1 2 54307 54309
0 54311 5 1 1 54310
0 54312 7 1 2 64892 54311
0 54313 5 1 1 54312
0 54314 7 1 2 104994 88259
0 54315 5 1 1 54314
0 54316 7 1 2 54313 54315
0 54317 5 1 1 54316
0 54318 7 1 2 73990 54317
0 54319 5 1 1 54318
0 54320 7 1 2 54297 54319
0 54321 5 1 1 54320
0 54322 7 1 2 84531 95497
0 54323 7 1 2 54321 54322
0 54324 5 1 1 54323
0 54325 7 1 2 72484 54324
0 54326 7 1 2 54293 54325
0 54327 5 1 1 54326
0 54328 7 1 2 103431 19059
0 54329 5 1 1 54328
0 54330 7 1 2 82149 54329
0 54331 5 1 1 54330
0 54332 7 1 2 86279 80271
0 54333 5 1 1 54332
0 54334 7 1 2 52096 54333
0 54335 5 1 1 54334
0 54336 7 1 2 70547 54335
0 54337 5 1 1 54336
0 54338 7 1 2 93230 54337
0 54339 5 1 1 54338
0 54340 7 1 2 72801 54339
0 54341 5 1 1 54340
0 54342 7 1 2 54331 54341
0 54343 5 1 1 54342
0 54344 7 1 2 68190 54343
0 54345 5 1 1 54344
0 54346 7 1 2 106287 54345
0 54347 5 1 1 54346
0 54348 7 1 2 71203 54347
0 54349 5 1 1 54348
0 54350 7 1 2 51657 54349
0 54351 5 1 1 54350
0 54352 7 1 2 85555 54351
0 54353 5 1 1 54352
0 54354 7 1 2 79902 104498
0 54355 5 1 1 54354
0 54356 7 1 2 81538 54355
0 54357 5 1 1 54356
0 54358 7 1 2 79072 102909
0 54359 5 1 1 54358
0 54360 7 1 2 52060 54359
0 54361 5 1 1 54360
0 54362 7 1 2 72802 54361
0 54363 5 1 1 54362
0 54364 7 1 2 54357 54363
0 54365 5 1 1 54364
0 54366 7 1 2 73269 54365
0 54367 5 1 1 54366
0 54368 7 1 2 76343 87485
0 54369 5 1 1 54368
0 54370 7 1 2 78151 54369
0 54371 5 1 1 54370
0 54372 7 1 2 42418 54371
0 54373 5 1 1 54372
0 54374 7 1 2 64513 54373
0 54375 5 1 1 54374
0 54376 7 1 2 54367 54375
0 54377 5 1 1 54376
0 54378 7 1 2 66089 54377
0 54379 5 1 1 54378
0 54380 7 1 2 89268 87478
0 54381 5 1 1 54380
0 54382 7 1 2 54379 54381
0 54383 5 1 1 54382
0 54384 7 1 2 82474 54383
0 54385 5 1 1 54384
0 54386 7 1 2 54353 54385
0 54387 5 1 1 54386
0 54388 7 1 2 76773 54387
0 54389 5 1 1 54388
0 54390 7 1 2 81788 104011
0 54391 5 1 1 54390
0 54392 7 1 2 95087 73991
0 54393 5 1 1 54392
0 54394 7 1 2 54391 54393
0 54395 5 1 1 54394
0 54396 7 1 2 103750 54395
0 54397 5 1 1 54396
0 54398 7 1 2 100505 103421
0 54399 5 1 1 54398
0 54400 7 1 2 54397 54399
0 54401 5 1 1 54400
0 54402 7 1 2 67810 54401
0 54403 5 1 1 54402
0 54404 7 1 2 76243 87530
0 54405 5 1 1 54404
0 54406 7 1 2 81588 104689
0 54407 5 1 1 54406
0 54408 7 1 2 54405 54407
0 54409 5 1 1 54408
0 54410 7 1 2 95343 93352
0 54411 7 1 2 54409 54410
0 54412 5 1 1 54411
0 54413 7 1 2 54403 54412
0 54414 5 1 1 54413
0 54415 7 1 2 76774 54414
0 54416 5 1 1 54415
0 54417 7 1 2 81488 84390
0 54418 5 1 1 54417
0 54419 7 1 2 74980 93519
0 54420 5 1 1 54419
0 54421 7 1 2 54418 54420
0 54422 5 1 1 54421
0 54423 7 1 2 70916 54422
0 54424 5 1 1 54423
0 54425 7 1 2 85094 98163
0 54426 5 1 1 54425
0 54427 7 1 2 54424 54426
0 54428 5 1 1 54427
0 54429 7 1 2 100032 54428
0 54430 5 1 1 54429
0 54431 7 1 2 68524 82220
0 54432 7 1 2 100927 54431
0 54433 7 1 2 98166 54432
0 54434 5 1 1 54433
0 54435 7 1 2 54430 54434
0 54436 5 1 1 54435
0 54437 7 1 2 84871 74265
0 54438 7 1 2 54436 54437
0 54439 5 1 1 54438
0 54440 7 1 2 54416 54439
0 54441 5 1 1 54440
0 54442 7 1 2 65205 54441
0 54443 5 1 1 54442
0 54444 7 1 2 67471 54443
0 54445 7 1 2 54389 54444
0 54446 5 1 1 54445
0 54447 7 1 2 78888 54446
0 54448 7 1 2 54327 54447
0 54449 5 1 1 54448
0 54450 7 1 2 71494 106553
0 54451 5 1 1 54450
0 54452 7 1 2 78552 105347
0 54453 5 2 1 54452
0 54454 7 1 2 66387 106576
0 54455 5 1 1 54454
0 54456 7 1 2 105096 54455
0 54457 7 1 2 54451 54456
0 54458 5 1 1 54457
0 54459 7 1 2 78997 75809
0 54460 7 1 2 103808 54459
0 54461 5 1 1 54460
0 54462 7 1 2 79403 54461
0 54463 5 1 1 54462
0 54464 7 1 2 70548 54463
0 54465 5 1 1 54464
0 54466 7 1 2 99507 83670
0 54467 5 1 1 54466
0 54468 7 1 2 95889 80976
0 54469 5 1 1 54468
0 54470 7 1 2 54467 54469
0 54471 5 1 1 54470
0 54472 7 1 2 106536 54471
0 54473 5 1 1 54472
0 54474 7 1 2 54465 54473
0 54475 5 1 1 54474
0 54476 7 1 2 68525 54475
0 54477 5 1 1 54476
0 54478 7 1 2 72194 76892
0 54479 7 1 2 80798 54478
0 54480 7 1 2 95946 54479
0 54481 5 1 1 54480
0 54482 7 1 2 79404 54481
0 54483 5 1 1 54482
0 54484 7 1 2 75991 54483
0 54485 5 1 1 54484
0 54486 7 1 2 54477 54485
0 54487 7 1 2 54458 54486
0 54488 5 1 1 54487
0 54489 7 1 2 96934 54488
0 54490 5 1 1 54489
0 54491 7 1 2 53905 106551
0 54492 5 1 1 54491
0 54493 7 1 2 96935 54492
0 54494 5 1 1 54493
0 54495 7 1 2 96976 78553
0 54496 7 1 2 94278 54495
0 54497 5 1 1 54496
0 54498 7 1 2 54494 54497
0 54499 5 1 1 54498
0 54500 7 1 2 102336 54499
0 54501 5 1 1 54500
0 54502 7 1 2 98193 103060
0 54503 7 1 2 95677 54502
0 54504 7 1 2 94989 54503
0 54505 5 1 1 54504
0 54506 7 1 2 94649 102754
0 54507 7 1 2 100369 54506
0 54508 7 1 2 79606 54507
0 54509 5 1 1 54508
0 54510 7 1 2 54505 54509
0 54511 5 1 1 54510
0 54512 7 1 2 70549 54511
0 54513 5 1 1 54512
0 54514 7 1 2 99534 86145
0 54515 5 1 1 54514
0 54516 7 1 2 83224 102755
0 54517 7 1 2 84614 54516
0 54518 7 1 2 54515 54517
0 54519 5 1 1 54518
0 54520 7 1 2 54513 54519
0 54521 5 1 1 54520
0 54522 7 1 2 73270 54521
0 54523 5 1 1 54522
0 54524 7 1 2 54501 54523
0 54525 5 1 1 54524
0 54526 7 1 2 65206 54525
0 54527 5 1 1 54526
0 54528 7 1 2 91073 92076
0 54529 7 1 2 101188 54528
0 54530 7 1 2 101871 54529
0 54531 5 1 1 54530
0 54532 7 1 2 13451 1045
0 54533 5 1 1 54532
0 54534 7 1 2 74981 98099
0 54535 7 1 2 54533 54534
0 54536 5 1 1 54535
0 54537 7 1 2 54531 54536
0 54538 5 1 1 54537
0 54539 7 1 2 65509 54538
0 54540 5 1 1 54539
0 54541 7 3 2 84330 78998
0 54542 7 1 2 84713 78353
0 54543 7 1 2 91082 54542
0 54544 7 1 2 106578 54543
0 54545 5 1 1 54544
0 54546 7 1 2 54540 54545
0 54547 5 1 1 54546
0 54548 7 1 2 98182 54547
0 54549 5 1 1 54548
0 54550 7 1 2 54527 54549
0 54551 7 1 2 54490 54550
0 54552 5 1 1 54551
0 54553 7 1 2 70018 54552
0 54554 5 1 1 54553
0 54555 7 1 2 86702 93309
0 54556 7 1 2 86101 54555
0 54557 5 1 1 54556
0 54558 7 2 2 66897 84872
0 54559 7 1 2 79871 104067
0 54560 7 1 2 106581 54559
0 54561 5 1 1 54560
0 54562 7 1 2 54557 54561
0 54563 5 1 1 54562
0 54564 7 1 2 75226 54563
0 54565 5 1 1 54564
0 54566 7 1 2 100233 102955
0 54567 7 1 2 80949 54566
0 54568 7 1 2 106481 54567
0 54569 5 1 1 54568
0 54570 7 1 2 54565 54569
0 54571 5 1 1 54570
0 54572 7 1 2 67472 54571
0 54573 5 1 1 54572
0 54574 7 1 2 97545 78554
0 54575 5 1 1 54574
0 54576 7 2 2 70550 75227
0 54577 5 1 1 106583
0 54578 7 1 2 54575 54577
0 54579 5 1 1 54578
0 54580 7 1 2 75465 54579
0 54581 5 1 1 54580
0 54582 7 1 2 54581 106577
0 54583 5 1 1 54582
0 54584 7 1 2 75593 104655
0 54585 7 1 2 54583 54584
0 54586 5 1 1 54585
0 54587 7 1 2 54573 54586
0 54588 5 1 1 54587
0 54589 7 1 2 64893 54588
0 54590 5 1 1 54589
0 54591 7 1 2 96936 106308
0 54592 5 1 1 54591
0 54593 7 1 2 96977 86156
0 54594 5 1 1 54593
0 54595 7 1 2 54592 54594
0 54596 5 1 1 54595
0 54597 7 1 2 87766 54596
0 54598 5 1 1 54597
0 54599 7 1 2 96937 79402
0 54600 5 1 1 54599
0 54601 7 1 2 54598 54600
0 54602 5 1 1 54601
0 54603 7 1 2 71495 54602
0 54604 5 1 1 54603
0 54605 7 1 2 54590 54604
0 54606 5 1 1 54605
0 54607 7 1 2 68191 54606
0 54608 5 1 1 54607
0 54609 7 1 2 75197 103997
0 54610 7 1 2 106458 54609
0 54611 5 1 1 54610
0 54612 7 1 2 99555 98194
0 54613 7 1 2 78555 54612
0 54614 5 1 1 54613
0 54615 7 1 2 54611 54614
0 54616 5 1 1 54615
0 54617 7 1 2 79532 54616
0 54618 5 1 1 54617
0 54619 7 1 2 54608 54618
0 54620 7 1 2 54554 54619
0 54621 5 1 1 54620
0 54622 7 1 2 67811 54621
0 54623 5 1 1 54622
0 54624 7 1 2 104068 86198
0 54625 7 1 2 74266 54624
0 54626 7 1 2 87541 54625
0 54627 5 1 1 54626
0 54628 7 1 2 87930 76861
0 54629 7 1 2 96618 54628
0 54630 7 1 2 97189 54629
0 54631 5 1 1 54630
0 54632 7 1 2 54627 54631
0 54633 5 1 1 54632
0 54634 7 1 2 100033 54633
0 54635 5 1 1 54634
0 54636 7 1 2 70551 87980
0 54637 5 1 1 54636
0 54638 7 1 2 79405 54637
0 54639 5 1 1 54638
0 54640 7 1 2 79970 54639
0 54641 5 1 1 54640
0 54642 7 1 2 106365 106477
0 54643 5 1 1 54642
0 54644 7 1 2 75228 54643
0 54645 5 1 1 54644
0 54646 7 1 2 64894 80928
0 54647 5 1 1 54646
0 54648 7 1 2 70019 83782
0 54649 5 1 1 54648
0 54650 7 1 2 94437 74299
0 54651 7 1 2 54649 54650
0 54652 7 1 2 54647 54651
0 54653 5 1 1 54652
0 54654 7 1 2 54645 54653
0 54655 5 1 1 54654
0 54656 7 1 2 75941 54655
0 54657 5 1 1 54656
0 54658 7 1 2 78325 75883
0 54659 7 1 2 94486 54658
0 54660 7 1 2 98043 54659
0 54661 5 1 1 54660
0 54662 7 1 2 54657 54661
0 54663 5 1 1 54662
0 54664 7 1 2 79155 54663
0 54665 5 1 1 54664
0 54666 7 1 2 54641 54665
0 54667 5 1 1 54666
0 54668 7 1 2 69301 54667
0 54669 5 1 1 54668
0 54670 7 1 2 54635 54669
0 54671 5 1 1 54670
0 54672 7 1 2 96770 54671
0 54673 5 1 1 54672
0 54674 7 1 2 69302 76171
0 54675 7 1 2 98604 54674
0 54676 7 1 2 95752 90624
0 54677 7 1 2 54675 54676
0 54678 5 1 1 54677
0 54679 7 1 2 54673 54678
0 54680 7 1 2 54623 54679
0 54681 5 1 1 54680
0 54682 7 1 2 70917 54681
0 54683 5 1 1 54682
0 54684 7 2 2 93222 105097
0 54685 7 1 2 105678 106585
0 54686 5 1 1 54685
0 54687 7 1 2 97419 77682
0 54688 7 1 2 97273 54687
0 54689 5 1 1 54688
0 54690 7 1 2 93223 75583
0 54691 7 1 2 79796 54690
0 54692 5 1 1 54691
0 54693 7 1 2 54689 54692
0 54694 5 1 1 54693
0 54695 7 1 2 66605 54694
0 54696 5 1 1 54695
0 54697 7 1 2 54686 54696
0 54698 5 1 1 54697
0 54699 7 1 2 94889 54698
0 54700 5 1 1 54699
0 54701 7 3 2 78556 105544
0 54702 7 1 2 95602 92501
0 54703 7 1 2 106587 54702
0 54704 5 1 1 54703
0 54705 7 1 2 54700 54704
0 54706 5 1 1 54705
0 54707 7 1 2 65510 54706
0 54708 5 1 1 54707
0 54709 7 1 2 100048 95557
0 54710 5 1 1 54709
0 54711 7 1 2 66790 106588
0 54712 5 1 1 54711
0 54713 7 1 2 54710 54712
0 54714 5 1 1 54713
0 54715 7 1 2 106586 54714
0 54716 5 1 1 54715
0 54717 7 1 2 54708 54716
0 54718 5 1 1 54717
0 54719 7 1 2 105808 54718
0 54720 5 1 1 54719
0 54721 7 1 2 54683 54720
0 54722 5 1 1 54721
0 54723 7 1 2 81080 54722
0 54724 5 1 1 54723
0 54725 7 1 2 83441 87386
0 54726 5 1 1 54725
0 54727 7 1 2 43994 54726
0 54728 5 1 1 54727
0 54729 7 1 2 71496 54728
0 54730 5 1 1 54729
0 54731 7 1 2 70020 106295
0 54732 5 1 1 54731
0 54733 7 1 2 54730 54732
0 54734 5 1 1 54733
0 54735 7 1 2 70552 54734
0 54736 5 1 1 54735
0 54737 7 1 2 106209 54736
0 54738 5 1 1 54737
0 54739 7 1 2 100530 54738
0 54740 5 1 1 54739
0 54741 7 1 2 79674 105819
0 54742 5 1 1 54741
0 54743 7 1 2 99397 105615
0 54744 7 1 2 54742 54743
0 54745 5 1 1 54744
0 54746 7 1 2 54740 54745
0 54747 5 1 1 54746
0 54748 7 1 2 72803 54747
0 54749 5 1 1 54748
0 54750 7 1 2 76033 98775
0 54751 7 1 2 86824 54750
0 54752 7 1 2 100524 54751
0 54753 5 1 1 54752
0 54754 7 1 2 54749 54753
0 54755 5 1 1 54754
0 54756 7 1 2 75229 54755
0 54757 5 1 1 54756
0 54758 7 1 2 101001 95558
0 54759 5 1 1 54758
0 54760 7 1 2 95890 104710
0 54761 7 1 2 106533 54760
0 54762 5 1 1 54761
0 54763 7 1 2 54759 54762
0 54764 5 1 1 54763
0 54765 7 1 2 66388 54764
0 54766 5 1 1 54765
0 54767 7 2 2 65511 95344
0 54768 7 1 2 86225 101153
0 54769 7 1 2 106534 54768
0 54770 7 1 2 106590 54769
0 54771 5 1 1 54770
0 54772 7 1 2 54766 54771
0 54773 5 1 1 54772
0 54774 7 1 2 69303 54773
0 54775 5 1 1 54774
0 54776 7 1 2 95345 94905
0 54777 7 1 2 106129 106342
0 54778 7 1 2 54776 54777
0 54779 5 1 1 54778
0 54780 7 1 2 54775 54779
0 54781 5 1 1 54780
0 54782 7 1 2 87712 54781
0 54783 5 1 1 54782
0 54784 7 1 2 74704 79186
0 54785 5 1 1 54784
0 54786 7 1 2 51876 54785
0 54787 5 1 1 54786
0 54788 7 1 2 81789 54787
0 54789 5 1 1 54788
0 54790 7 1 2 83474 86601
0 54791 5 1 1 54790
0 54792 7 1 2 54789 54791
0 54793 5 1 1 54792
0 54794 7 1 2 100531 54793
0 54795 5 1 1 54794
0 54796 7 1 2 70553 79187
0 54797 5 1 1 54796
0 54798 7 1 2 86975 54797
0 54799 5 1 1 54798
0 54800 7 1 2 101069 87087
0 54801 7 1 2 54799 54800
0 54802 5 1 1 54801
0 54803 7 1 2 54795 54802
0 54804 5 1 1 54803
0 54805 7 1 2 75230 54804
0 54806 5 1 1 54805
0 54807 7 1 2 77887 78808
0 54808 7 1 2 78557 54807
0 54809 7 1 2 103620 54808
0 54810 5 1 1 54809
0 54811 7 1 2 54806 54810
0 54812 7 1 2 54783 54811
0 54813 5 1 1 54812
0 54814 7 1 2 67812 54813
0 54815 5 1 1 54814
0 54816 7 1 2 104679 104528
0 54817 5 1 1 54816
0 54818 7 1 2 78114 88880
0 54819 7 1 2 100355 54818
0 54820 5 1 1 54819
0 54821 7 1 2 54817 54820
0 54822 5 1 1 54821
0 54823 7 1 2 63934 54822
0 54824 5 1 1 54823
0 54825 7 1 2 83299 98463
0 54826 7 1 2 84601 54825
0 54827 7 1 2 84443 54826
0 54828 5 1 1 54827
0 54829 7 1 2 54824 54828
0 54830 5 1 1 54829
0 54831 7 1 2 79539 92586
0 54832 7 1 2 54830 54831
0 54833 5 1 1 54832
0 54834 7 1 2 54815 54833
0 54835 5 1 1 54834
0 54836 7 1 2 64895 54835
0 54837 5 1 1 54836
0 54838 7 1 2 80765 106589
0 54839 5 1 1 54838
0 54840 7 1 2 75231 106372
0 54841 5 1 1 54840
0 54842 7 1 2 54839 54841
0 54843 5 1 1 54842
0 54844 7 1 2 100532 54843
0 54845 5 1 1 54844
0 54846 7 1 2 75232 106368
0 54847 5 1 1 54846
0 54848 7 1 2 76775 106356
0 54849 5 1 1 54848
0 54850 7 1 2 54847 54849
0 54851 5 1 1 54850
0 54852 7 1 2 103621 54851
0 54853 5 1 1 54852
0 54854 7 1 2 54845 54853
0 54855 5 1 1 54854
0 54856 7 1 2 93022 54855
0 54857 5 1 1 54856
0 54858 7 1 2 54837 54857
0 54859 7 1 2 54757 54858
0 54860 5 1 1 54859
0 54861 7 1 2 79156 54860
0 54862 5 1 1 54861
0 54863 7 1 2 97443 95587
0 54864 7 1 2 103761 54863
0 54865 7 1 2 96164 54864
0 54866 7 1 2 93023 54865
0 54867 5 1 1 54866
0 54868 7 1 2 54862 54867
0 54869 7 1 2 54724 54868
0 54870 7 1 2 54449 54869
0 54871 7 1 2 54221 54870
0 54872 7 1 2 53991 54871
0 54873 5 1 1 54872
0 54874 7 1 2 73877 54873
0 54875 5 1 1 54874
0 54876 7 1 2 64896 100655
0 54877 5 1 1 54876
0 54878 7 1 2 78847 104050
0 54879 7 1 2 54877 54878
0 54880 5 1 1 54879
0 54881 7 1 2 79292 106297
0 54882 5 1 1 54881
0 54883 7 1 2 54880 54882
0 54884 5 1 1 54883
0 54885 7 1 2 66606 54884
0 54886 5 1 1 54885
0 54887 7 1 2 80086 80035
0 54888 7 1 2 106224 54887
0 54889 5 1 1 54888
0 54890 7 1 2 54886 54889
0 54891 5 1 1 54890
0 54892 7 1 2 73271 54891
0 54893 5 1 1 54892
0 54894 7 1 2 92404 79263
0 54895 7 1 2 106225 54894
0 54896 5 1 1 54895
0 54897 7 1 2 54893 54896
0 54898 5 1 1 54897
0 54899 7 1 2 85959 54898
0 54900 5 1 1 54899
0 54901 7 1 2 64897 78971
0 54902 5 1 1 54901
0 54903 7 1 2 79265 54902
0 54904 5 1 1 54903
0 54905 7 1 2 81790 93722
0 54906 7 1 2 54904 54905
0 54907 5 1 1 54906
0 54908 7 1 2 54900 54907
0 54909 5 1 1 54908
0 54910 7 1 2 88618 54909
0 54911 5 1 1 54910
0 54912 7 1 2 85960 97363
0 54913 7 1 2 93192 54912
0 54914 7 1 2 97818 54913
0 54915 5 1 1 54914
0 54916 7 1 2 54911 54915
0 54917 5 1 1 54916
0 54918 7 1 2 67813 54917
0 54919 5 1 1 54918
0 54920 7 1 2 89642 84438
0 54921 5 1 1 54920
0 54922 7 1 2 92678 75826
0 54923 7 1 2 90684 54922
0 54924 5 1 1 54923
0 54925 7 1 2 54921 54924
0 54926 5 1 1 54925
0 54927 7 1 2 84873 54926
0 54928 5 1 1 54927
0 54929 7 1 2 80902 94983
0 54930 7 1 2 96166 54929
0 54931 5 1 1 54930
0 54932 7 1 2 54928 54931
0 54933 5 1 1 54932
0 54934 7 1 2 65207 54933
0 54935 5 1 1 54934
0 54936 7 2 2 84684 94443
0 54937 5 1 1 106592
0 54938 7 1 2 96036 78115
0 54939 7 1 2 106318 54938
0 54940 5 1 1 54939
0 54941 7 1 2 54937 54940
0 54942 5 1 1 54941
0 54943 7 1 2 99684 54942
0 54944 5 1 1 54943
0 54945 7 1 2 54935 54944
0 54946 5 1 1 54945
0 54947 7 1 2 71706 54946
0 54948 5 1 1 54947
0 54949 7 1 2 70275 99685
0 54950 7 1 2 106593 54949
0 54951 5 1 1 54950
0 54952 7 1 2 54948 54951
0 54953 5 1 1 54952
0 54954 7 1 2 76101 54953
0 54955 5 1 1 54954
0 54956 7 1 2 88337 106464
0 54957 5 1 1 54956
0 54958 7 1 2 93723 94529
0 54959 5 1 1 54958
0 54960 7 1 2 54957 54959
0 54961 5 1 1 54960
0 54962 7 1 2 69654 54961
0 54963 5 1 1 54962
0 54964 7 1 2 98328 84581
0 54965 7 1 2 87589 54964
0 54966 5 1 1 54965
0 54967 7 1 2 54963 54966
0 54968 5 1 1 54967
0 54969 7 1 2 93024 54968
0 54970 5 1 1 54969
0 54971 7 1 2 85338 95845
0 54972 5 1 1 54971
0 54973 7 1 2 87342 95744
0 54974 7 1 2 78336 54973
0 54975 5 1 1 54974
0 54976 7 1 2 54972 54975
0 54977 5 1 1 54976
0 54978 7 1 2 70554 54977
0 54979 5 1 1 54978
0 54980 7 1 2 91867 89932
0 54981 7 1 2 92405 75650
0 54982 7 1 2 54980 54981
0 54983 5 1 1 54982
0 54984 7 1 2 54979 54983
0 54985 5 1 1 54984
0 54986 7 1 2 71497 54985
0 54987 5 1 1 54986
0 54988 7 1 2 91074 98796
0 54989 7 1 2 105698 54988
0 54990 5 1 1 54989
0 54991 7 1 2 54987 54990
0 54992 5 1 1 54991
0 54993 7 1 2 91489 89132
0 54994 7 1 2 54992 54993
0 54995 5 1 1 54994
0 54996 7 1 2 54970 54995
0 54997 7 1 2 54955 54996
0 54998 7 1 2 54919 54997
0 54999 5 1 1 54998
0 55000 7 1 2 94243 95077
0 55001 7 1 2 54999 55000
0 55002 5 1 1 55001
0 55003 7 1 2 100657 101132
0 55004 7 1 2 90790 55003
0 55005 5 1 1 55004
0 55006 7 1 2 87673 86656
0 55007 7 1 2 106438 55006
0 55008 5 1 1 55007
0 55009 7 1 2 55005 55008
0 55010 5 1 1 55009
0 55011 7 1 2 100069 55010
0 55012 5 1 1 55011
0 55013 7 1 2 75466 94114
0 55014 5 1 1 55013
0 55015 7 1 2 11357 94401
0 55016 5 1 1 55015
0 55017 7 1 2 68192 55016
0 55018 5 1 1 55017
0 55019 7 1 2 91437 93419
0 55020 5 1 1 55019
0 55021 7 1 2 55018 55020
0 55022 5 1 1 55021
0 55023 7 1 2 91602 98871
0 55024 7 1 2 55022 55023
0 55025 5 1 1 55024
0 55026 7 1 2 55014 55025
0 55027 5 1 1 55026
0 55028 7 1 2 71498 55027
0 55029 5 1 1 55028
0 55030 7 1 2 55012 55029
0 55031 5 1 1 55030
0 55032 7 1 2 65512 55031
0 55033 5 1 1 55032
0 55034 7 2 2 66791 100658
0 55035 7 1 2 105166 106594
0 55036 5 1 1 55035
0 55037 7 1 2 71707 105264
0 55038 7 1 2 105534 55037
0 55039 5 1 1 55038
0 55040 7 1 2 55036 55039
0 55041 5 1 1 55040
0 55042 7 1 2 76102 55041
0 55043 5 1 1 55042
0 55044 7 1 2 91606 105435
0 55045 5 1 1 55044
0 55046 7 2 2 90746 93638
0 55047 5 1 1 106596
0 55048 7 1 2 106595 106597
0 55049 5 1 1 55048
0 55050 7 1 2 55045 55049
0 55051 5 1 1 55050
0 55052 7 1 2 78747 55051
0 55053 5 1 1 55052
0 55054 7 1 2 101791 88055
0 55055 7 1 2 104182 105443
0 55056 7 1 2 55054 55055
0 55057 5 1 1 55056
0 55058 7 1 2 55053 55057
0 55059 7 1 2 55043 55058
0 55060 5 1 1 55059
0 55061 7 1 2 85961 55060
0 55062 5 1 1 55061
0 55063 7 1 2 55033 55062
0 55064 5 1 1 55063
0 55065 7 1 2 88619 55064
0 55066 5 1 1 55065
0 55067 7 1 2 91793 106465
0 55068 7 1 2 100684 55067
0 55069 5 1 1 55068
0 55070 7 1 2 55066 55069
0 55071 5 1 1 55070
0 55072 7 1 2 67814 55071
0 55073 5 1 1 55072
0 55074 7 3 2 89144 91246
0 55075 7 1 2 84261 106598
0 55076 5 1 1 55075
0 55077 7 1 2 95891 106320
0 55078 5 1 1 55077
0 55079 7 1 2 55076 55078
0 55080 5 1 1 55079
0 55081 7 1 2 76510 55080
0 55082 5 1 1 55081
0 55083 7 1 2 96039 90985
0 55084 5 1 1 55083
0 55085 7 1 2 55082 55084
0 55086 5 1 1 55085
0 55087 7 1 2 76344 90913
0 55088 7 1 2 55086 55087
0 55089 5 1 1 55088
0 55090 7 1 2 55073 55089
0 55091 5 1 1 55090
0 55092 7 1 2 69655 55091
0 55093 5 1 1 55092
0 55094 7 1 2 87420 91288
0 55095 7 1 2 104976 55094
0 55096 7 1 2 97819 55095
0 55097 7 1 2 95687 55096
0 55098 5 1 1 55097
0 55099 7 1 2 55093 55098
0 55100 7 1 2 55002 55099
0 55101 5 1 1 55100
0 55102 7 1 2 85445 55101
0 55103 5 1 1 55102
0 55104 7 1 2 75467 102022
0 55105 5 1 1 55104
0 55106 7 1 2 75853 83273
0 55107 5 1 1 55106
0 55108 7 1 2 55105 55107
0 55109 5 1 1 55108
0 55110 7 1 2 80766 55109
0 55111 5 1 1 55110
0 55112 7 1 2 91327 96572
0 55113 5 1 1 55112
0 55114 7 1 2 55111 55113
0 55115 5 1 1 55114
0 55116 7 1 2 88620 55115
0 55117 5 1 1 55116
0 55118 7 1 2 74705 101290
0 55119 7 1 2 78915 55118
0 55120 5 1 1 55119
0 55121 7 1 2 98660 105216
0 55122 5 1 1 55121
0 55123 7 1 2 55120 55122
0 55124 5 1 1 55123
0 55125 7 1 2 88260 55124
0 55126 5 1 1 55125
0 55127 7 1 2 55117 55126
0 55128 5 1 1 55127
0 55129 7 1 2 94691 55128
0 55130 5 1 1 55129
0 55131 7 1 2 96573 88261
0 55132 7 1 2 99964 55131
0 55133 5 1 1 55132
0 55134 7 1 2 82877 90553
0 55135 7 1 2 99725 55134
0 55136 5 1 1 55135
0 55137 7 1 2 55133 55136
0 55138 5 1 1 55137
0 55139 7 2 2 67815 55138
0 55140 7 1 2 93439 106601
0 55141 5 1 1 55140
0 55142 7 1 2 55130 55141
0 55143 5 1 1 55142
0 55144 7 1 2 65853 55143
0 55145 5 1 1 55144
0 55146 7 1 2 85339 78131
0 55147 7 1 2 106602 55146
0 55148 5 1 1 55147
0 55149 7 1 2 55145 55148
0 55150 5 1 1 55149
0 55151 7 1 2 71204 89004
0 55152 7 1 2 55150 55151
0 55153 5 1 1 55152
0 55154 7 1 2 55103 55153
0 55155 5 1 1 55154
0 55156 7 1 2 67473 55155
0 55157 5 1 1 55156
0 55158 7 1 2 83948 9927
0 55159 5 1 1 55158
0 55160 7 1 2 105532 55159
0 55161 5 1 1 55160
0 55162 7 4 2 75468 98925
0 55163 7 1 2 97420 91794
0 55164 7 1 2 106603 55163
0 55165 5 1 1 55164
0 55166 7 1 2 55161 55165
0 55167 5 1 1 55166
0 55168 7 1 2 94692 55167
0 55169 5 1 1 55168
0 55170 7 1 2 103916 96574
0 55171 7 1 2 97187 55170
0 55172 5 1 1 55171
0 55173 7 1 2 55169 55172
0 55174 5 1 1 55173
0 55175 7 1 2 69656 55174
0 55176 5 1 1 55175
0 55177 7 2 2 71965 96464
0 55178 7 1 2 95459 90536
0 55179 7 1 2 106607 55178
0 55180 5 1 1 55179
0 55181 7 1 2 63985 74318
0 55182 7 1 2 81288 55181
0 55183 7 1 2 105525 55182
0 55184 5 1 1 55183
0 55185 7 1 2 55180 55184
0 55186 5 1 1 55185
0 55187 7 1 2 70021 55186
0 55188 5 1 1 55187
0 55189 7 1 2 106504 106608
0 55190 5 1 1 55189
0 55191 7 1 2 84178 91833
0 55192 7 1 2 94374 55191
0 55193 5 1 1 55192
0 55194 7 1 2 55190 55193
0 55195 5 1 1 55194
0 55196 7 1 2 71499 55195
0 55197 5 1 1 55196
0 55198 7 1 2 55188 55197
0 55199 5 1 1 55198
0 55200 7 1 2 67816 55199
0 55201 5 1 1 55200
0 55202 7 1 2 71205 86199
0 55203 7 1 2 95753 55202
0 55204 7 1 2 105158 55203
0 55205 5 1 1 55204
0 55206 7 1 2 55201 55205
0 55207 5 1 1 55206
0 55208 7 1 2 94693 55207
0 55209 5 1 1 55208
0 55210 7 1 2 55176 55209
0 55211 5 1 1 55210
0 55212 7 1 2 88262 55211
0 55213 5 1 1 55212
0 55214 7 2 2 76397 90813
0 55215 7 1 2 94002 95765
0 55216 7 1 2 106609 55215
0 55217 5 1 1 55216
0 55218 7 1 2 88330 84685
0 55219 7 1 2 91911 55218
0 55220 5 1 1 55219
0 55221 7 1 2 55217 55220
0 55222 5 1 1 55221
0 55223 7 1 2 71206 55222
0 55224 5 1 1 55223
0 55225 7 1 2 67817 88331
0 55226 7 1 2 94524 55225
0 55227 5 1 1 55226
0 55228 7 1 2 55224 55227
0 55229 5 1 1 55228
0 55230 7 1 2 70555 55229
0 55231 5 1 1 55230
0 55232 7 1 2 87343 90204
0 55233 7 1 2 90791 55232
0 55234 7 1 2 106610 55233
0 55235 5 1 1 55234
0 55236 7 1 2 55231 55235
0 55237 5 1 1 55236
0 55238 7 1 2 106515 55237
0 55239 5 1 1 55238
0 55240 7 1 2 55213 55239
0 55241 5 1 1 55240
0 55242 7 1 2 72485 55241
0 55243 5 1 1 55242
0 55244 7 2 2 72804 96575
0 55245 7 1 2 90214 106611
0 55246 5 1 1 55245
0 55247 7 1 2 92461 106604
0 55248 5 1 1 55247
0 55249 7 1 2 55246 55248
0 55250 5 2 1 55249
0 55251 7 1 2 88263 106613
0 55252 5 1 1 55251
0 55253 7 1 2 84019 90959
0 55254 7 1 2 94601 55253
0 55255 7 1 2 105393 55254
0 55256 7 2 2 106226 55255
0 55257 5 1 1 106615
0 55258 7 1 2 55252 55257
0 55259 5 1 1 55258
0 55260 7 1 2 97421 55259
0 55261 5 1 1 55260
0 55262 7 1 2 80767 100234
0 55263 7 2 2 83336 79529
0 55264 7 1 2 76907 91541
0 55265 7 1 2 106617 55264
0 55266 7 1 2 55262 55265
0 55267 5 1 1 55266
0 55268 7 1 2 69657 55267
0 55269 7 1 2 55261 55268
0 55270 5 1 1 55269
0 55271 7 1 2 84714 75764
0 55272 7 1 2 94060 55271
0 55273 5 1 1 55272
0 55274 7 1 2 94559 55273
0 55275 5 1 1 55274
0 55276 7 1 2 92797 55275
0 55277 5 1 1 55276
0 55278 7 1 2 92310 94438
0 55279 7 1 2 102144 55278
0 55280 7 1 2 105554 55279
0 55281 5 1 1 55280
0 55282 7 1 2 55277 55281
0 55283 5 1 1 55282
0 55284 7 1 2 93353 55283
0 55285 5 1 1 55284
0 55286 7 2 2 66898 84423
0 55287 7 1 2 97422 82766
0 55288 7 1 2 106619 55287
0 55289 7 1 2 96576 96216
0 55290 7 1 2 55288 55289
0 55291 5 1 1 55290
0 55292 7 1 2 64514 55291
0 55293 7 1 2 55285 55292
0 55294 5 1 1 55293
0 55295 7 1 2 55270 55294
0 55296 5 1 1 55295
0 55297 7 1 2 72195 86200
0 55298 7 1 2 93459 55297
0 55299 7 1 2 106527 55298
0 55300 7 1 2 106605 55299
0 55301 5 1 1 55300
0 55302 7 1 2 66090 55301
0 55303 7 1 2 55296 55302
0 55304 5 1 1 55303
0 55305 7 1 2 64515 106614
0 55306 5 1 1 55305
0 55307 7 1 2 80768 104120
0 55308 7 1 2 93553 55307
0 55309 5 1 1 55308
0 55310 7 1 2 55306 55309
0 55311 5 1 1 55310
0 55312 7 1 2 88264 55311
0 55313 5 1 1 55312
0 55314 7 1 2 64516 106616
0 55315 5 1 1 55314
0 55316 7 1 2 55313 55315
0 55317 5 1 1 55316
0 55318 7 1 2 97423 55317
0 55319 5 1 1 55318
0 55320 7 1 2 67818 88343
0 55321 5 1 1 55320
0 55322 7 1 2 23806 55321
0 55323 5 1 1 55322
0 55324 7 1 2 80769 55323
0 55325 5 1 1 55324
0 55326 7 1 2 76511 106612
0 55327 5 1 1 55326
0 55328 7 1 2 55325 55327
0 55329 5 1 1 55328
0 55330 7 1 2 88621 55329
0 55331 5 1 1 55330
0 55332 7 1 2 70022 81289
0 55333 5 1 1 55332
0 55334 7 1 2 81622 55333
0 55335 5 1 1 55334
0 55336 7 1 2 106599 55335
0 55337 5 1 1 55336
0 55338 7 1 2 55331 55337
0 55339 5 1 1 55338
0 55340 7 1 2 76398 92566
0 55341 7 1 2 55339 55340
0 55342 5 1 1 55341
0 55343 7 1 2 71207 55342
0 55344 7 1 2 55319 55343
0 55345 5 1 1 55344
0 55346 7 1 2 55304 55345
0 55347 5 1 1 55346
0 55348 7 1 2 88299 106600
0 55349 5 1 1 55348
0 55350 7 1 2 88642 106606
0 55351 5 1 1 55350
0 55352 7 1 2 55349 55351
0 55353 5 1 1 55352
0 55354 7 1 2 78132 90914
0 55355 7 1 2 55353 55354
0 55356 5 1 1 55355
0 55357 7 1 2 55347 55356
0 55358 5 1 1 55357
0 55359 7 1 2 67474 55358
0 55360 5 1 1 55359
0 55361 7 4 2 72486 84686
0 55362 7 3 2 69304 106621
0 55363 5 1 1 106625
0 55364 7 1 2 41228 55363
0 55365 5 1 1 55364
0 55366 7 2 2 97424 89335
0 55367 7 1 2 55365 106628
0 55368 5 1 1 55367
0 55369 7 1 2 84106 96999
0 55370 5 1 1 55369
0 55371 7 1 2 96978 83942
0 55372 5 1 1 55371
0 55373 7 1 2 55370 55372
0 55374 5 1 1 55373
0 55375 7 1 2 89410 55374
0 55376 5 1 1 55375
0 55377 7 1 2 55368 55376
0 55378 5 1 1 55377
0 55379 7 1 2 71208 55378
0 55380 5 1 1 55379
0 55381 7 1 2 98346 99211
0 55382 7 1 2 106629 55381
0 55383 5 1 1 55382
0 55384 7 1 2 55380 55383
0 55385 5 1 1 55384
0 55386 7 1 2 88086 55385
0 55387 5 1 1 55386
0 55388 7 1 2 99699 79383
0 55389 7 1 2 91917 55388
0 55390 7 1 2 105709 55389
0 55391 5 1 1 55390
0 55392 7 1 2 55387 55391
0 55393 5 1 1 55392
0 55394 7 1 2 82878 55393
0 55395 5 1 1 55394
0 55396 7 1 2 95806 99126
0 55397 5 1 1 55396
0 55398 7 1 2 90916 55397
0 55399 5 1 1 55398
0 55400 7 1 2 69305 93336
0 55401 7 1 2 99279 55400
0 55402 7 1 2 55399 55401
0 55403 5 1 1 55402
0 55404 7 1 2 55395 55403
0 55405 5 1 1 55404
0 55406 7 1 2 84874 55405
0 55407 5 1 1 55406
0 55408 7 1 2 96979 105334
0 55409 5 1 1 55408
0 55410 7 1 2 96938 86602
0 55411 5 1 1 55410
0 55412 7 1 2 55409 55411
0 55413 5 1 1 55412
0 55414 7 1 2 96212 96097
0 55415 5 1 1 55414
0 55416 7 1 2 99117 106346
0 55417 5 1 1 55416
0 55418 7 1 2 55415 55417
0 55419 5 1 1 55418
0 55420 7 1 2 71209 55419
0 55421 5 1 1 55420
0 55422 7 1 2 70732 79481
0 55423 7 1 2 91090 55422
0 55424 7 1 2 99113 55423
0 55425 5 1 1 55424
0 55426 7 1 2 55421 55425
0 55427 5 1 1 55426
0 55428 7 1 2 55413 55427
0 55429 5 1 1 55428
0 55430 7 1 2 55407 55429
0 55431 7 1 2 55360 55430
0 55432 7 1 2 55243 55431
0 55433 5 1 1 55432
0 55434 7 1 2 68193 55433
0 55435 5 1 1 55434
0 55436 7 1 2 69306 100994
0 55437 5 1 1 55436
0 55438 7 1 2 43762 55437
0 55439 5 1 1 55438
0 55440 7 1 2 105717 55439
0 55441 5 1 1 55440
0 55442 7 1 2 87134 99159
0 55443 7 1 2 103878 55442
0 55444 5 1 1 55443
0 55445 7 1 2 55441 55444
0 55446 5 1 1 55445
0 55447 7 1 2 71708 55446
0 55448 5 1 1 55447
0 55449 7 1 2 66607 99834
0 55450 7 1 2 106510 55449
0 55451 5 1 1 55450
0 55452 7 1 2 55448 55451
0 55453 5 1 1 55452
0 55454 7 1 2 85962 55453
0 55455 5 1 1 55454
0 55456 7 1 2 84137 98293
0 55457 5 1 1 55456
0 55458 7 1 2 64517 77978
0 55459 7 1 2 102450 55458
0 55460 5 1 1 55459
0 55461 7 1 2 55457 55460
0 55462 5 1 1 55461
0 55463 7 1 2 69307 55462
0 55464 5 1 1 55463
0 55465 7 1 2 96980 104404
0 55466 5 1 1 55465
0 55467 7 1 2 55464 55466
0 55468 5 1 1 55467
0 55469 7 1 2 85340 76614
0 55470 7 1 2 55468 55469
0 55471 5 1 1 55470
0 55472 7 1 2 55455 55471
0 55473 5 1 1 55472
0 55474 7 1 2 88622 55473
0 55475 5 1 1 55474
0 55476 7 1 2 91872 105087
0 55477 5 1 1 55476
0 55478 7 1 2 66792 98797
0 55479 7 1 2 99700 55478
0 55480 5 1 1 55479
0 55481 7 1 2 55477 55480
0 55482 5 1 1 55481
0 55483 7 1 2 71210 55482
0 55484 5 1 1 55483
0 55485 7 1 2 76966 79482
0 55486 7 1 2 91873 55485
0 55487 5 1 1 55486
0 55488 7 1 2 55484 55487
0 55489 5 1 1 55488
0 55490 7 1 2 70556 55489
0 55491 5 1 1 55490
0 55492 7 1 2 71872 79598
0 55493 7 1 2 98329 55492
0 55494 7 1 2 103917 55493
0 55495 5 1 1 55494
0 55496 7 1 2 55491 55495
0 55497 5 1 1 55496
0 55498 7 1 2 96939 55497
0 55499 5 1 1 55498
0 55500 7 1 2 85341 93489
0 55501 7 1 2 103908 55500
0 55502 7 1 2 99726 55501
0 55503 5 1 1 55502
0 55504 7 1 2 55499 55503
0 55505 5 1 1 55504
0 55506 7 1 2 88265 55505
0 55507 5 1 1 55506
0 55508 7 1 2 55475 55507
0 55509 5 1 1 55508
0 55510 7 1 2 65208 55509
0 55511 5 1 1 55510
0 55512 7 1 2 81290 100391
0 55513 5 1 1 55512
0 55514 7 1 2 96981 79581
0 55515 7 1 2 91826 55514
0 55516 5 1 1 55515
0 55517 7 1 2 55513 55516
0 55518 5 1 1 55517
0 55519 7 1 2 70557 55518
0 55520 5 1 1 55519
0 55521 7 1 2 87349 99301
0 55522 7 1 2 93460 55521
0 55523 5 1 1 55522
0 55524 7 1 2 55520 55523
0 55525 5 1 1 55524
0 55526 7 1 2 88623 55525
0 55527 5 1 1 55526
0 55528 7 1 2 22142 106540
0 55529 5 1 1 55528
0 55530 7 4 2 71500 89190
0 55531 7 1 2 55529 106630
0 55532 5 1 1 55531
0 55533 7 1 2 55527 55532
0 55534 5 1 1 55533
0 55535 7 1 2 70023 55534
0 55536 5 1 1 55535
0 55537 7 1 2 77717 74253
0 55538 7 2 2 103095 55537
0 55539 5 2 1 106634
0 55540 7 1 2 96940 106635
0 55541 5 1 1 55540
0 55542 7 1 2 55536 55541
0 55543 5 1 1 55542
0 55544 7 1 2 81081 55543
0 55545 5 1 1 55544
0 55546 7 1 2 95137 100634
0 55547 5 1 1 55546
0 55548 7 1 2 85342 79918
0 55549 5 1 1 55548
0 55550 7 1 2 55547 55549
0 55551 5 1 1 55550
0 55552 7 1 2 97018 55551
0 55553 5 1 1 55552
0 55554 7 1 2 88344 89191
0 55555 5 1 1 55554
0 55556 7 1 2 55553 55555
0 55557 5 1 1 55556
0 55558 7 1 2 65513 55557
0 55559 5 1 1 55558
0 55560 7 1 2 66793 89885
0 55561 5 1 1 55560
0 55562 7 1 2 84144 88624
0 55563 5 1 1 55562
0 55564 7 1 2 55561 55563
0 55565 5 1 1 55564
0 55566 7 1 2 92104 55565
0 55567 5 1 1 55566
0 55568 7 1 2 55559 55567
0 55569 5 1 1 55568
0 55570 7 1 2 106511 55569
0 55571 5 1 1 55570
0 55572 7 1 2 89157 97482
0 55573 7 1 2 94796 55572
0 55574 7 1 2 104969 104988
0 55575 7 1 2 55573 55574
0 55576 5 1 1 55575
0 55577 7 1 2 67819 55576
0 55578 7 1 2 55571 55577
0 55579 7 1 2 55545 55578
0 55580 7 1 2 55511 55579
0 55581 5 1 1 55580
0 55582 7 1 2 77386 88300
0 55583 5 1 1 55582
0 55584 7 1 2 93345 81082
0 55585 5 1 1 55584
0 55586 7 1 2 55583 55585
0 55587 5 1 1 55586
0 55588 7 1 2 74254 96219
0 55589 7 1 2 55587 55588
0 55590 5 1 1 55589
0 55591 7 1 2 71709 106425
0 55592 5 1 1 55591
0 55593 7 1 2 94448 55592
0 55594 5 1 1 55593
0 55595 7 1 2 100001 104361
0 55596 7 1 2 55594 55595
0 55597 5 1 1 55596
0 55598 7 1 2 55590 55597
0 55599 5 1 1 55598
0 55600 7 1 2 69308 55599
0 55601 5 1 1 55600
0 55602 7 1 2 85343 81291
0 55603 5 1 1 55602
0 55604 7 1 2 99508 99999
0 55605 5 1 1 55604
0 55606 7 1 2 55603 55605
0 55607 5 1 1 55606
0 55608 7 1 2 70558 55607
0 55609 5 1 1 55608
0 55610 7 1 2 93148 84168
0 55611 5 1 1 55610
0 55612 7 1 2 55609 55611
0 55613 5 1 1 55612
0 55614 7 1 2 88625 55613
0 55615 5 1 1 55614
0 55616 7 1 2 96465 106631
0 55617 5 1 1 55616
0 55618 7 1 2 55615 55617
0 55619 5 1 1 55618
0 55620 7 1 2 70024 55619
0 55621 5 1 1 55620
0 55622 7 1 2 106636 55621
0 55623 5 1 1 55622
0 55624 7 1 2 101010 55623
0 55625 5 1 1 55624
0 55626 7 1 2 55601 55625
0 55627 5 1 1 55626
0 55628 7 1 2 67475 55627
0 55629 5 1 1 55628
0 55630 7 1 2 81292 89316
0 55631 5 1 1 55630
0 55632 7 1 2 98577 106632
0 55633 5 1 1 55632
0 55634 7 1 2 55631 55633
0 55635 5 1 1 55634
0 55636 7 1 2 70559 55635
0 55637 5 1 1 55636
0 55638 7 1 2 96555 106633
0 55639 5 1 1 55638
0 55640 7 1 2 55637 55639
0 55641 5 1 1 55640
0 55642 7 1 2 70025 55641
0 55643 5 1 1 55642
0 55644 7 1 2 106637 55643
0 55645 5 1 1 55644
0 55646 7 1 2 104947 55645
0 55647 5 1 1 55646
0 55648 7 1 2 72805 55647
0 55649 7 1 2 55629 55648
0 55650 5 1 1 55649
0 55651 7 1 2 73272 55650
0 55652 7 1 2 55581 55651
0 55653 5 1 1 55652
0 55654 7 1 2 101291 105957
0 55655 5 1 1 55654
0 55656 7 1 2 84138 92828
0 55657 7 1 2 98545 55656
0 55658 5 1 1 55657
0 55659 7 1 2 55655 55658
0 55660 5 1 1 55659
0 55661 7 1 2 67476 55660
0 55662 5 1 1 55661
0 55663 7 1 2 96941 84139
0 55664 7 1 2 80132 90867
0 55665 7 1 2 55663 55664
0 55666 5 1 1 55665
0 55667 7 1 2 55662 55666
0 55668 5 1 1 55667
0 55669 7 1 2 76244 89317
0 55670 7 1 2 55668 55669
0 55671 5 1 1 55670
0 55672 7 1 2 55653 55671
0 55673 5 1 1 55672
0 55674 7 1 2 88087 55673
0 55675 5 1 1 55674
0 55676 7 1 2 98347 105877
0 55677 5 1 1 55676
0 55678 7 1 2 99689 92971
0 55679 5 1 1 55678
0 55680 7 1 2 100105 96771
0 55681 5 2 1 55680
0 55682 7 1 2 55679 106638
0 55683 7 1 2 40450 55682
0 55684 7 1 2 55677 55683
0 55685 5 1 1 55684
0 55686 7 1 2 74578 55685
0 55687 5 1 1 55686
0 55688 7 1 2 81083 105607
0 55689 5 1 1 55688
0 55690 7 1 2 106639 55689
0 55691 5 1 1 55690
0 55692 7 1 2 76345 55691
0 55693 5 1 1 55692
0 55694 7 1 2 69309 99851
0 55695 7 1 2 98390 55694
0 55696 5 1 1 55695
0 55697 7 1 2 55693 55696
0 55698 7 1 2 55687 55697
0 55699 5 1 1 55698
0 55700 7 1 2 70560 55699
0 55701 5 1 1 55700
0 55702 7 1 2 84246 93078
0 55703 7 1 2 106397 55702
0 55704 5 1 1 55703
0 55705 7 1 2 55701 55704
0 55706 5 1 1 55705
0 55707 7 1 2 88266 55706
0 55708 5 1 1 55707
0 55709 7 1 2 71211 106542
0 55710 5 1 1 55709
0 55711 7 1 2 78133 106538
0 55712 5 1 1 55711
0 55713 7 1 2 55710 55712
0 55714 5 1 1 55713
0 55715 7 1 2 101169 90561
0 55716 7 1 2 55714 55715
0 55717 5 1 1 55716
0 55718 7 1 2 55708 55717
0 55719 5 1 1 55718
0 55720 7 1 2 85963 55719
0 55721 5 1 1 55720
0 55722 7 1 2 83764 105088
0 55723 5 1 1 55722
0 55724 7 1 2 76245 78501
0 55725 5 1 1 55724
0 55726 7 1 2 92888 55725
0 55727 7 1 2 55723 55726
0 55728 5 1 1 55727
0 55729 7 2 2 97444 55728
0 55730 7 1 2 96201 106640
0 55731 5 1 1 55730
0 55732 7 1 2 76512 98413
0 55733 5 1 1 55732
0 55734 7 1 2 71212 101969
0 55735 5 1 1 55734
0 55736 7 1 2 55733 55735
0 55737 5 1 1 55736
0 55738 7 1 2 69658 55737
0 55739 5 1 1 55738
0 55740 7 1 2 67477 84730
0 55741 5 1 1 55740
0 55742 7 1 2 55739 55741
0 55743 5 1 1 55742
0 55744 7 1 2 84875 90966
0 55745 7 1 2 55743 55744
0 55746 5 1 1 55745
0 55747 7 1 2 55731 55746
0 55748 5 1 1 55747
0 55749 7 1 2 65209 55748
0 55750 5 1 1 55749
0 55751 7 1 2 83115 93851
0 55752 7 1 2 106641 55751
0 55753 5 1 1 55752
0 55754 7 1 2 55750 55753
0 55755 5 1 1 55754
0 55756 7 1 2 89418 55755
0 55757 5 1 1 55756
0 55758 7 1 2 55721 55757
0 55759 5 1 1 55758
0 55760 7 1 2 89005 55759
0 55761 5 1 1 55760
0 55762 7 1 2 55675 55761
0 55763 7 1 2 55435 55762
0 55764 5 1 1 55763
0 55765 7 1 2 70918 55764
0 55766 5 1 1 55765
0 55767 7 1 2 55157 55766
0 55768 5 1 1 55767
0 55769 7 1 2 68526 55768
0 55770 5 1 1 55769
0 55771 7 1 2 54875 55770
0 55772 7 1 2 53807 55771
0 55773 7 1 2 52545 55772
0 55774 7 1 2 51587 55773
0 55775 5 1 1 55774
0 55776 7 1 2 73786 55775
0 55777 5 1 1 55776
0 55778 7 1 2 51140 55777
0 55779 7 1 2 46321 55778
0 55780 5 1 1 55779
0 55781 7 1 2 72270 55780
0 55782 5 1 1 55781
0 55783 7 1 2 103573 94767
0 55784 5 1 1 55783
0 55785 7 1 2 100329 103158
0 55786 5 1 1 55785
0 55787 7 1 2 84211 83711
0 55788 5 1 1 55787
0 55789 7 1 2 96811 32155
0 55790 5 1 1 55789
0 55791 7 1 2 66389 55790
0 55792 5 1 1 55791
0 55793 7 1 2 32207 55792
0 55794 5 1 1 55793
0 55795 7 1 2 70561 55794
0 55796 5 1 1 55795
0 55797 7 1 2 66390 104395
0 55798 5 1 1 55797
0 55799 7 1 2 68731 91590
0 55800 5 1 1 55799
0 55801 7 1 2 91787 55800
0 55802 5 1 1 55801
0 55803 7 1 2 65514 55802
0 55804 5 1 1 55803
0 55805 7 1 2 55798 55804
0 55806 7 1 2 55796 55805
0 55807 5 1 1 55806
0 55808 7 1 2 68194 55807
0 55809 5 1 1 55808
0 55810 7 1 2 55788 55809
0 55811 5 1 1 55810
0 55812 7 1 2 64898 55811
0 55813 5 1 1 55812
0 55814 7 1 2 55786 55813
0 55815 5 1 1 55814
0 55816 7 1 2 72806 55815
0 55817 5 1 1 55816
0 55818 7 1 2 55784 55817
0 55819 5 1 1 55818
0 55820 7 1 2 65210 55819
0 55821 5 1 1 55820
0 55822 7 1 2 98929 105857
0 55823 5 1 1 55822
0 55824 7 1 2 89259 77051
0 55825 7 1 2 55823 55824
0 55826 5 1 1 55825
0 55827 7 1 2 55821 55826
0 55828 5 1 1 55827
0 55829 7 1 2 102187 104157
0 55830 7 1 2 90397 55829
0 55831 5 1 1 55830
0 55832 7 1 2 103935 77638
0 55833 7 1 2 83205 55832
0 55834 7 1 2 73878 55833
0 55835 5 1 1 55834
0 55836 7 1 2 55831 55835
0 55837 5 1 1 55836
0 55838 7 1 2 55828 55837
0 55839 5 1 1 55838
0 55840 7 28 2 67225 74408
0 55841 5 1 1 106642
0 55842 7 1 2 79741 86315
0 55843 5 1 1 55842
0 55844 7 1 2 68195 103519
0 55845 5 1 1 55844
0 55846 7 1 2 55843 55845
0 55847 5 1 1 55846
0 55848 7 1 2 71501 55847
0 55849 5 1 1 55848
0 55850 7 2 2 79038 77052
0 55851 7 1 2 86901 106670
0 55852 5 1 1 55851
0 55853 7 1 2 55849 55852
0 55854 5 1 1 55853
0 55855 7 1 2 65211 55854
0 55856 5 1 1 55855
0 55857 7 1 2 103022 106034
0 55858 5 1 1 55857
0 55859 7 1 2 55856 55858
0 55860 5 1 1 55859
0 55861 7 1 2 106643 55860
0 55862 5 1 1 55861
0 55863 7 1 2 75299 99642
0 55864 5 1 1 55863
0 55865 7 1 2 74824 106644
0 55866 5 1 1 55865
0 55867 7 1 2 55864 55866
0 55868 5 2 1 55867
0 55869 7 1 2 79210 106672
0 55870 5 1 1 55869
0 55871 7 1 2 72271 100388
0 55872 7 1 2 93128 55871
0 55873 5 1 1 55872
0 55874 7 1 2 55870 55873
0 55875 5 1 1 55874
0 55876 7 1 2 80770 55875
0 55877 5 1 1 55876
0 55878 7 5 2 100140 78296
0 55879 5 2 1 106674
0 55880 7 1 2 106357 106675
0 55881 5 1 1 55880
0 55882 7 1 2 79211 103936
0 55883 7 1 2 101795 55882
0 55884 5 1 1 55883
0 55885 7 2 2 55881 55884
0 55886 5 1 1 106681
0 55887 7 1 2 55877 106682
0 55888 5 1 1 55887
0 55889 7 1 2 76103 55888
0 55890 5 1 1 55889
0 55891 7 1 2 102136 93082
0 55892 5 1 1 55891
0 55893 7 1 2 73606 103970
0 55894 7 1 2 103639 55893
0 55895 5 1 1 55894
0 55896 7 1 2 55892 55895
0 55897 5 1 1 55896
0 55898 7 1 2 74706 55897
0 55899 5 1 1 55898
0 55900 7 1 2 94841 103971
0 55901 7 1 2 93129 55900
0 55902 5 1 1 55901
0 55903 7 1 2 55899 55902
0 55904 5 1 1 55903
0 55905 7 1 2 71502 55904
0 55906 5 1 1 55905
0 55907 7 2 2 82475 101574
0 55908 5 1 1 106683
0 55909 7 1 2 75942 83337
0 55910 7 1 2 106684 55909
0 55911 5 1 1 55910
0 55912 7 1 2 55906 55911
0 55913 5 1 1 55912
0 55914 7 1 2 81791 55913
0 55915 5 1 1 55914
0 55916 7 1 2 100749 101885
0 55917 5 1 1 55916
0 55918 7 1 2 74177 100141
0 55919 7 1 2 55917 55918
0 55920 5 1 1 55919
0 55921 7 1 2 55915 55920
0 55922 5 1 1 55921
0 55923 7 1 2 73787 55922
0 55924 5 1 1 55923
0 55925 7 2 2 81365 103313
0 55926 7 1 2 70026 102838
0 55927 7 1 2 106685 55926
0 55928 5 1 1 55927
0 55929 7 1 2 64899 81650
0 55930 7 1 2 106673 55929
0 55931 5 1 1 55930
0 55932 7 1 2 55928 55931
0 55933 5 1 1 55932
0 55934 7 1 2 80771 55933
0 55935 5 1 1 55934
0 55936 7 1 2 55924 55935
0 55937 7 1 2 55890 55936
0 55938 7 1 2 55862 55937
0 55939 5 2 1 55938
0 55940 7 1 2 74473 106687
0 55941 5 1 1 55940
0 55942 7 1 2 78599 93942
0 55943 5 1 1 55942
0 55944 7 1 2 86740 105559
0 55945 7 1 2 55943 55944
0 55946 5 1 1 55945
0 55947 7 1 2 68196 55946
0 55948 5 1 1 55947
0 55949 7 1 2 65515 55948
0 55950 5 1 1 55949
0 55951 7 1 2 88828 77953
0 55952 5 1 1 55951
0 55953 7 1 2 74891 87116
0 55954 7 1 2 100888 55953
0 55955 5 1 1 55954
0 55956 7 1 2 73273 55955
0 55957 5 1 1 55956
0 55958 7 1 2 86813 81443
0 55959 7 1 2 75658 55958
0 55960 5 1 1 55959
0 55961 7 1 2 55957 55960
0 55962 5 1 1 55961
0 55963 7 1 2 55952 55962
0 55964 5 1 1 55963
0 55965 7 1 2 55950 55964
0 55966 5 1 1 55965
0 55967 7 1 2 30177 55966
0 55968 5 1 1 55967
0 55969 7 1 2 65212 55968
0 55970 5 2 1 55969
0 55971 7 1 2 79431 94407
0 55972 5 1 1 55971
0 55973 7 1 2 82936 87042
0 55974 7 1 2 93299 55973
0 55975 5 1 1 55974
0 55976 7 1 2 55972 55975
0 55977 5 1 1 55976
0 55978 7 1 2 65516 55977
0 55979 5 1 1 55978
0 55980 7 1 2 79432 80143
0 55981 5 1 1 55980
0 55982 7 1 2 64900 95169
0 55983 5 1 1 55982
0 55984 7 1 2 55981 55983
0 55985 5 1 1 55984
0 55986 7 1 2 70562 55985
0 55987 5 1 1 55986
0 55988 7 1 2 55979 55987
0 55989 7 1 2 106689 55988
0 55990 5 1 1 55989
0 55991 7 1 2 106645 55990
0 55992 5 1 1 55991
0 55993 7 1 2 70276 104489
0 55994 5 1 1 55993
0 55995 7 1 2 99012 55994
0 55996 5 1 1 55995
0 55997 7 1 2 99643 55996
0 55998 5 1 1 55997
0 55999 7 1 2 78712 98978
0 56000 5 1 1 55999
0 56001 7 1 2 421 2888
0 56002 5 1 1 56001
0 56003 7 1 2 71710 56002
0 56004 5 1 1 56003
0 56005 7 1 2 75891 99005
0 56006 7 1 2 97765 56005
0 56007 5 1 1 56006
0 56008 7 1 2 86691 56007
0 56009 7 1 2 56004 56008
0 56010 7 1 2 56000 56009
0 56011 5 1 1 56010
0 56012 7 1 2 106646 56011
0 56013 5 1 1 56012
0 56014 7 2 2 55998 56013
0 56015 5 1 1 106691
0 56016 7 1 2 66391 56015
0 56017 5 1 1 56016
0 56018 7 1 2 74409 103244
0 56019 5 1 1 56018
0 56020 7 1 2 55908 56019
0 56021 5 2 1 56020
0 56022 7 1 2 99867 106693
0 56023 5 1 1 56022
0 56024 7 1 2 89803 89660
0 56025 5 1 1 56024
0 56026 7 1 2 68197 56025
0 56027 5 1 1 56026
0 56028 7 1 2 93277 56027
0 56029 5 1 1 56028
0 56030 7 2 2 81792 56029
0 56031 5 1 1 106695
0 56032 7 1 2 99644 106696
0 56033 5 1 1 56032
0 56034 7 1 2 56023 56033
0 56035 7 1 2 56017 56034
0 56036 7 1 2 55992 56035
0 56037 5 1 1 56036
0 56038 7 1 2 82823 56037
0 56039 5 1 1 56038
0 56040 7 1 2 55941 56039
0 56041 5 1 1 56040
0 56042 7 1 2 88626 56041
0 56043 5 1 1 56042
0 56044 7 1 2 99825 85583
0 56045 5 1 1 56044
0 56046 7 1 2 64901 56045
0 56047 5 1 1 56046
0 56048 7 1 2 79201 95962
0 56049 5 1 1 56048
0 56050 7 1 2 56047 56049
0 56051 5 2 1 56050
0 56052 7 1 2 74474 106697
0 56053 5 1 1 56052
0 56054 7 1 2 97425 74475
0 56055 5 1 1 56054
0 56056 7 1 2 86577 56055
0 56057 5 1 1 56056
0 56058 7 1 2 80772 56057
0 56059 5 1 1 56058
0 56060 7 1 2 88308 96609
0 56061 5 1 1 56060
0 56062 7 1 2 3524 56061
0 56063 7 1 2 56059 56062
0 56064 5 1 1 56063
0 56065 7 1 2 73607 56064
0 56066 5 1 1 56065
0 56067 7 1 2 56053 56066
0 56068 5 1 1 56067
0 56069 7 1 2 68198 56068
0 56070 5 1 1 56069
0 56071 7 1 2 98802 100758
0 56072 5 1 1 56071
0 56073 7 1 2 73608 56072
0 56074 5 1 1 56073
0 56075 7 1 2 95090 85584
0 56076 7 1 2 56074 56075
0 56077 5 1 1 56076
0 56078 7 1 2 71503 56077
0 56079 5 1 1 56078
0 56080 7 1 2 100747 56079
0 56081 5 1 1 56080
0 56082 7 1 2 85837 56081
0 56083 5 1 1 56082
0 56084 7 1 2 56070 56083
0 56085 5 1 1 56084
0 56086 7 1 2 74707 56085
0 56087 5 1 1 56086
0 56088 7 1 2 86741 83097
0 56089 5 1 1 56088
0 56090 7 1 2 65517 56089
0 56091 5 1 1 56090
0 56092 7 1 2 83459 102376
0 56093 5 1 1 56092
0 56094 7 1 2 75300 56093
0 56095 5 1 1 56094
0 56096 7 1 2 56091 56095
0 56097 5 1 1 56096
0 56098 7 1 2 64902 56097
0 56099 5 1 1 56098
0 56100 7 1 2 73788 87262
0 56101 5 1 1 56100
0 56102 7 1 2 56099 56101
0 56103 5 1 1 56102
0 56104 7 1 2 68199 56103
0 56105 5 1 1 56104
0 56106 7 2 2 70027 77006
0 56107 7 1 2 102944 106699
0 56108 5 1 1 56107
0 56109 7 1 2 86771 79212
0 56110 5 1 1 56109
0 56111 7 1 2 80773 87392
0 56112 5 1 1 56111
0 56113 7 2 2 56110 56112
0 56114 7 2 2 74883 86162
0 56115 7 1 2 70563 106703
0 56116 5 1 1 56115
0 56117 7 1 2 106701 56116
0 56118 5 2 1 56117
0 56119 7 1 2 76104 106705
0 56120 5 1 1 56119
0 56121 7 1 2 56108 56120
0 56122 7 1 2 56105 56121
0 56123 5 1 1 56122
0 56124 7 1 2 74476 56123
0 56125 5 1 1 56124
0 56126 7 1 2 99503 78757
0 56127 5 1 1 56126
0 56128 7 1 2 85715 82824
0 56129 7 1 2 56127 56128
0 56130 5 1 1 56129
0 56131 7 1 2 56125 56130
0 56132 7 1 2 56087 56131
0 56133 5 1 1 56132
0 56134 7 1 2 106647 56133
0 56135 5 1 1 56134
0 56136 7 1 2 68200 105433
0 56137 5 1 1 56136
0 56138 7 1 2 103212 56137
0 56139 5 1 1 56138
0 56140 7 1 2 82825 56139
0 56141 5 1 1 56140
0 56142 7 1 2 65213 83131
0 56143 5 1 1 56142
0 56144 7 1 2 101814 56143
0 56145 5 1 1 56144
0 56146 7 1 2 70564 56145
0 56147 5 1 1 56146
0 56148 7 1 2 106151 56147
0 56149 5 1 1 56148
0 56150 7 2 2 68201 56149
0 56151 5 1 1 106707
0 56152 7 2 2 83978 86596
0 56153 5 1 1 106709
0 56154 7 1 2 70028 98972
0 56155 7 1 2 104224 56154
0 56156 5 1 1 56155
0 56157 7 1 2 56153 56156
0 56158 5 1 1 56157
0 56159 7 1 2 74708 56158
0 56160 5 1 1 56159
0 56161 7 1 2 56151 56160
0 56162 5 1 1 56161
0 56163 7 1 2 74477 56162
0 56164 5 1 1 56163
0 56165 7 1 2 56141 56164
0 56166 5 1 1 56165
0 56167 7 1 2 66392 56166
0 56168 5 1 1 56167
0 56169 7 1 2 86580 86509
0 56170 5 1 1 56169
0 56171 7 1 2 82836 56170
0 56172 5 1 1 56171
0 56173 7 1 2 65518 56172
0 56174 5 1 1 56173
0 56175 7 1 2 82374 82826
0 56176 5 1 1 56175
0 56177 7 1 2 79773 74478
0 56178 7 1 2 84123 56177
0 56179 5 1 1 56178
0 56180 7 1 2 56176 56179
0 56181 7 1 2 56174 56180
0 56182 5 1 1 56181
0 56183 7 1 2 66608 56182
0 56184 5 1 1 56183
0 56185 7 1 2 85618 82827
0 56186 5 1 1 56185
0 56187 7 1 2 56184 56186
0 56188 5 1 1 56187
0 56189 7 1 2 79433 56188
0 56190 5 1 1 56189
0 56191 7 2 2 88694 74758
0 56192 5 1 1 106711
0 56193 7 1 2 98979 75051
0 56194 5 1 1 56193
0 56195 7 1 2 56192 56194
0 56196 5 1 1 56195
0 56197 7 1 2 64903 56196
0 56198 5 1 1 56197
0 56199 7 1 2 78748 104339
0 56200 5 1 1 56199
0 56201 7 1 2 86288 56200
0 56202 7 1 2 56198 56201
0 56203 5 1 1 56202
0 56204 7 1 2 74479 56203
0 56205 5 1 1 56204
0 56206 7 1 2 64904 86587
0 56207 5 1 1 56206
0 56208 7 1 2 56205 56207
0 56209 5 1 1 56208
0 56210 7 1 2 71504 56209
0 56211 5 1 1 56210
0 56212 7 1 2 56190 56211
0 56213 7 1 2 56168 56212
0 56214 5 1 1 56213
0 56215 7 1 2 99645 56214
0 56216 5 1 1 56215
0 56217 7 1 2 56135 56216
0 56218 5 1 1 56217
0 56219 7 1 2 88267 56218
0 56220 5 1 1 56219
0 56221 7 1 2 56043 56220
0 56222 5 1 1 56221
0 56223 7 1 2 91542 56222
0 56224 5 1 1 56223
0 56225 7 4 2 68527 106648
0 56226 5 2 1 106713
0 56227 7 1 2 88268 106714
0 56228 5 1 1 56227
0 56229 7 2 2 69019 100167
0 56230 7 2 2 96303 106719
0 56231 7 1 2 103051 106721
0 56232 5 1 1 56231
0 56233 7 1 2 56228 56232
0 56234 5 1 1 56233
0 56235 7 1 2 66609 56234
0 56236 5 1 1 56235
0 56237 7 1 2 101575 90960
0 56238 7 1 2 93745 56237
0 56239 5 1 1 56238
0 56240 7 1 2 56236 56239
0 56241 5 1 1 56240
0 56242 7 1 2 76105 56241
0 56243 5 1 1 56242
0 56244 7 1 2 106686 106722
0 56245 5 1 1 56244
0 56246 7 1 2 103947 88269
0 56247 5 2 1 56246
0 56248 7 2 2 74410 104713
0 56249 5 3 1 106725
0 56250 7 1 2 37393 106727
0 56251 5 1 1 56250
0 56252 7 1 2 88627 56251
0 56253 5 1 1 56252
0 56254 7 1 2 106723 56253
0 56255 5 1 1 56254
0 56256 7 1 2 75087 56255
0 56257 5 1 1 56256
0 56258 7 2 2 66610 67226
0 56259 7 1 2 79329 106730
0 56260 7 1 2 102188 56259
0 56261 5 1 1 56260
0 56262 7 1 2 56257 56261
0 56263 5 1 1 56262
0 56264 7 1 2 79414 56263
0 56265 5 1 1 56264
0 56266 7 1 2 56245 56265
0 56267 7 1 2 56243 56266
0 56268 5 1 1 56267
0 56269 7 1 2 65214 56268
0 56270 5 1 1 56269
0 56271 7 3 2 103937 89460
0 56272 5 1 1 106732
0 56273 7 1 2 106724 56272
0 56274 5 1 1 56273
0 56275 7 1 2 97364 78925
0 56276 5 1 1 56275
0 56277 7 1 2 29300 56276
0 56278 5 1 1 56277
0 56279 7 1 2 73609 56278
0 56280 7 1 2 56274 56279
0 56281 5 1 1 56280
0 56282 7 1 2 56270 56281
0 56283 5 2 1 56282
0 56284 7 1 2 80774 106735
0 56285 5 1 1 56284
0 56286 7 1 2 23421 55841
0 56287 5 7 1 56286
0 56288 7 1 2 83451 106737
0 56289 5 1 1 56288
0 56290 7 1 2 100150 79202
0 56291 5 1 1 56290
0 56292 7 1 2 56289 56291
0 56293 5 1 1 56292
0 56294 7 1 2 66611 56293
0 56295 5 1 1 56294
0 56296 7 2 2 99646 79235
0 56297 5 1 1 106744
0 56298 7 2 2 74411 102823
0 56299 5 1 1 106746
0 56300 7 1 2 73992 106747
0 56301 5 1 1 56300
0 56302 7 1 2 56297 56301
0 56303 5 1 1 56302
0 56304 7 1 2 70565 56303
0 56305 5 1 1 56304
0 56306 7 2 2 82476 103247
0 56307 5 2 1 106748
0 56308 7 1 2 106717 106750
0 56309 5 1 1 56308
0 56310 7 1 2 85716 56309
0 56311 5 1 1 56310
0 56312 7 1 2 56305 56311
0 56313 5 1 1 56312
0 56314 7 1 2 73789 56313
0 56315 5 1 1 56314
0 56316 7 1 2 56295 56315
0 56317 5 1 1 56316
0 56318 7 1 2 65215 56317
0 56319 5 1 1 56318
0 56320 7 1 2 73993 106749
0 56321 5 1 1 56320
0 56322 7 1 2 103429 106649
0 56323 5 1 1 56322
0 56324 7 1 2 56321 56323
0 56325 5 1 1 56324
0 56326 7 1 2 81793 56325
0 56327 5 1 1 56326
0 56328 7 1 2 80654 106650
0 56329 5 1 1 56328
0 56330 7 1 2 106751 56329
0 56331 5 1 1 56330
0 56332 7 1 2 78669 56331
0 56333 5 1 1 56332
0 56334 7 1 2 56327 56333
0 56335 5 1 1 56334
0 56336 7 1 2 73790 56335
0 56337 5 1 1 56336
0 56338 7 1 2 56319 56337
0 56339 5 1 1 56338
0 56340 7 1 2 88270 56339
0 56341 5 1 1 56340
0 56342 7 1 2 103945 106679
0 56343 5 3 1 56342
0 56344 7 1 2 93167 106752
0 56345 7 1 2 89051 56344
0 56346 5 1 1 56345
0 56347 7 1 2 56341 56346
0 56348 5 1 1 56347
0 56349 7 1 2 64905 56348
0 56350 5 1 1 56349
0 56351 7 1 2 102960 90268
0 56352 7 1 2 103948 56351
0 56353 5 1 1 56352
0 56354 7 2 2 103927 92077
0 56355 7 1 2 69020 93611
0 56356 7 1 2 106755 56355
0 56357 5 1 1 56356
0 56358 7 1 2 56353 56357
0 56359 5 1 1 56358
0 56360 7 1 2 94355 56359
0 56361 5 1 1 56360
0 56362 7 1 2 56350 56361
0 56363 5 1 1 56362
0 56364 7 1 2 68202 56363
0 56365 5 1 1 56364
0 56366 7 1 2 88628 55886
0 56367 5 1 1 56366
0 56368 7 1 2 64906 106738
0 56369 5 1 1 56368
0 56370 7 1 2 78585 103938
0 56371 5 1 1 56370
0 56372 7 1 2 56369 56371
0 56373 5 1 1 56372
0 56374 7 1 2 80655 56373
0 56375 5 1 1 56374
0 56376 7 1 2 95278 100142
0 56377 5 1 1 56376
0 56378 7 1 2 106718 56377
0 56379 5 1 1 56378
0 56380 7 1 2 95052 56379
0 56381 5 1 1 56380
0 56382 7 1 2 56375 56381
0 56383 5 1 1 56382
0 56384 7 1 2 74709 56383
0 56385 5 1 1 56384
0 56386 7 1 2 106704 106739
0 56387 5 1 1 56386
0 56388 7 1 2 86353 106745
0 56389 5 1 1 56388
0 56390 7 1 2 56387 56389
0 56391 5 1 1 56390
0 56392 7 1 2 70566 56391
0 56393 5 1 1 56392
0 56394 7 1 2 93083 104720
0 56395 5 1 1 56394
0 56396 7 1 2 99647 87394
0 56397 5 1 1 56396
0 56398 7 1 2 56395 56397
0 56399 5 1 1 56398
0 56400 7 1 2 65519 56399
0 56401 5 1 1 56400
0 56402 7 1 2 56393 56401
0 56403 7 1 2 56385 56402
0 56404 5 1 1 56403
0 56405 7 1 2 88271 56404
0 56406 5 1 1 56405
0 56407 7 1 2 56367 56406
0 56408 5 1 1 56407
0 56409 7 1 2 76106 56408
0 56410 5 1 1 56409
0 56411 7 1 2 100642 106733
0 56412 5 1 1 56411
0 56413 7 1 2 79073 90541
0 56414 7 1 2 106740 56413
0 56415 5 1 1 56414
0 56416 7 1 2 56412 56415
0 56417 5 1 1 56416
0 56418 7 1 2 74710 56417
0 56419 5 1 1 56418
0 56420 7 2 2 103939 89424
0 56421 5 1 1 106757
0 56422 7 1 2 103923 106516
0 56423 7 1 2 106353 56422
0 56424 5 1 1 56423
0 56425 7 1 2 56421 56424
0 56426 5 1 1 56425
0 56427 7 1 2 88722 56426
0 56428 5 1 1 56427
0 56429 7 1 2 56419 56428
0 56430 5 1 1 56429
0 56431 7 1 2 70029 56430
0 56432 5 1 1 56431
0 56433 7 1 2 103647 105410
0 56434 7 2 2 67227 74864
0 56435 7 2 2 69021 98335
0 56436 7 1 2 106759 106761
0 56437 7 1 2 56433 56436
0 56438 5 1 1 56437
0 56439 7 1 2 56432 56438
0 56440 5 1 1 56439
0 56441 7 1 2 73274 56440
0 56442 5 1 1 56441
0 56443 7 1 2 56410 56442
0 56444 7 2 2 56365 56443
0 56445 5 1 1 106763
0 56446 7 1 2 56285 106764
0 56447 5 1 1 56446
0 56448 7 1 2 72066 89529
0 56449 7 1 2 56447 56448
0 56450 5 1 1 56449
0 56451 7 1 2 56224 56450
0 56452 5 1 1 56451
0 56453 7 1 2 72807 56452
0 56454 5 1 1 56453
0 56455 7 3 2 103898 98893
0 56456 5 1 1 106765
0 56457 7 1 2 77286 103949
0 56458 7 1 2 90444 56457
0 56459 5 1 1 56458
0 56460 7 1 2 56456 56459
0 56461 5 1 1 56460
0 56462 7 1 2 66794 56461
0 56463 5 1 1 56462
0 56464 7 1 2 90753 106726
0 56465 5 1 1 56464
0 56466 7 1 2 56463 56465
0 56467 5 1 1 56466
0 56468 7 1 2 65520 56467
0 56469 5 1 1 56468
0 56470 7 1 2 88474 106766
0 56471 5 1 1 56470
0 56472 7 1 2 56469 56471
0 56473 5 1 1 56472
0 56474 7 1 2 88272 56473
0 56475 5 1 1 56474
0 56476 7 1 2 74255 103928
0 56477 7 1 2 106388 56476
0 56478 7 1 2 100598 56477
0 56479 5 1 1 56478
0 56480 7 1 2 56475 56479
0 56481 5 1 1 56480
0 56482 7 1 2 65216 56481
0 56483 5 1 1 56482
0 56484 7 1 2 86037 88273
0 56485 5 2 1 56484
0 56486 7 1 2 82937 92619
0 56487 5 1 1 56486
0 56488 7 1 2 106768 56487
0 56489 5 1 1 56488
0 56490 7 1 2 66612 106767
0 56491 7 1 2 56489 56490
0 56492 5 1 1 56491
0 56493 7 1 2 56483 56492
0 56494 5 1 1 56493
0 56495 7 1 2 73610 56494
0 56496 5 1 1 56495
0 56497 7 1 2 67228 86571
0 56498 7 1 2 90054 56497
0 56499 7 1 2 90674 56498
0 56500 7 1 2 98894 56499
0 56501 5 1 1 56500
0 56502 7 1 2 56496 56501
0 56503 5 1 1 56502
0 56504 7 1 2 76246 56503
0 56505 5 1 1 56504
0 56506 7 3 2 76247 90445
0 56507 7 1 2 90484 88629
0 56508 5 1 1 56507
0 56509 7 1 2 94706 56508
0 56510 5 1 1 56509
0 56511 7 1 2 106770 56510
0 56512 5 1 1 56511
0 56513 7 1 2 89471 106771
0 56514 5 1 1 56513
0 56515 7 1 2 95824 90446
0 56516 5 1 1 56515
0 56517 7 1 2 69022 91722
0 56518 7 1 2 95762 56517
0 56519 5 2 1 56518
0 56520 7 1 2 56516 106773
0 56521 5 2 1 56520
0 56522 7 1 2 88309 106775
0 56523 5 1 1 56522
0 56524 7 1 2 88630 106772
0 56525 5 1 1 56524
0 56526 7 1 2 56523 56525
0 56527 5 1 1 56526
0 56528 7 1 2 66795 56527
0 56529 5 1 1 56528
0 56530 7 1 2 56514 56529
0 56531 5 1 1 56530
0 56532 7 1 2 65521 56531
0 56533 5 1 1 56532
0 56534 7 1 2 56512 56533
0 56535 5 1 1 56534
0 56536 7 1 2 78670 56535
0 56537 5 1 1 56536
0 56538 7 1 2 81668 90057
0 56539 7 1 2 90447 56538
0 56540 5 1 1 56539
0 56541 7 1 2 56537 56540
0 56542 5 1 1 56541
0 56543 7 1 2 103950 56542
0 56544 5 1 1 56543
0 56545 7 1 2 77104 106776
0 56546 5 1 1 56545
0 56547 7 1 2 90183 90754
0 56548 5 1 1 56547
0 56549 7 1 2 56546 56548
0 56550 5 1 1 56549
0 56551 7 1 2 76248 56550
0 56552 5 1 1 56551
0 56553 7 1 2 69023 88684
0 56554 5 1 1 56553
0 56555 7 1 2 93871 56554
0 56556 5 1 1 56555
0 56557 7 1 2 106769 56556
0 56558 5 1 1 56557
0 56559 7 1 2 66613 56558
0 56560 5 1 1 56559
0 56561 7 1 2 88372 95825
0 56562 5 1 1 56561
0 56563 7 1 2 56560 56562
0 56564 5 1 1 56563
0 56565 7 1 2 43002 55047
0 56566 5 1 1 56565
0 56567 7 1 2 67010 56566
0 56568 7 1 2 56564 56567
0 56569 5 1 1 56568
0 56570 7 1 2 56552 56569
0 56571 5 1 1 56570
0 56572 7 1 2 73611 56571
0 56573 5 1 1 56572
0 56574 7 1 2 76249 90755
0 56575 7 1 2 94743 56574
0 56576 5 1 1 56575
0 56577 7 1 2 56573 56576
0 56578 5 1 1 56577
0 56579 7 1 2 106651 56578
0 56580 5 1 1 56579
0 56581 7 4 2 93115 102643
0 56582 5 1 1 106777
0 56583 7 1 2 103929 92855
0 56584 5 1 1 56583
0 56585 7 1 2 56582 56584
0 56586 5 1 1 56585
0 56587 7 1 2 90756 56586
0 56588 5 1 1 56587
0 56589 7 1 2 87441 94087
0 56590 5 1 1 56589
0 56591 7 1 2 86510 91543
0 56592 5 1 1 56591
0 56593 7 1 2 56590 56592
0 56594 5 1 1 56593
0 56595 7 1 2 72067 103951
0 56596 7 1 2 89472 56595
0 56597 7 1 2 56594 56596
0 56598 5 1 1 56597
0 56599 7 1 2 56588 56598
0 56600 5 1 1 56599
0 56601 7 1 2 80775 56600
0 56602 5 1 1 56601
0 56603 7 1 2 86354 106778
0 56604 5 1 1 56603
0 56605 7 1 2 90179 89104
0 56606 5 1 1 56605
0 56607 7 1 2 81794 103952
0 56608 7 1 2 56606 56607
0 56609 5 2 1 56608
0 56610 7 1 2 56604 106781
0 56611 5 1 1 56610
0 56612 7 1 2 90448 56611
0 56613 5 1 1 56612
0 56614 7 1 2 56602 56613
0 56615 5 1 1 56614
0 56616 7 1 2 76250 56615
0 56617 5 1 1 56616
0 56618 7 1 2 101356 89858
0 56619 7 1 2 89473 56618
0 56620 7 1 2 98895 56619
0 56621 5 1 1 56620
0 56622 7 1 2 56617 56621
0 56623 5 1 1 56622
0 56624 7 1 2 73994 56623
0 56625 5 1 1 56624
0 56626 7 1 2 101796 88631
0 56627 5 1 1 56626
0 56628 7 1 2 13123 56627
0 56629 5 1 1 56628
0 56630 7 10 2 63986 69310
0 56631 5 1 1 106783
0 56632 7 1 2 99972 100156
0 56633 7 1 2 106784 56632
0 56634 7 1 2 94111 56633
0 56635 7 1 2 56629 56634
0 56636 5 1 1 56635
0 56637 7 1 2 56625 56636
0 56638 7 1 2 56580 56637
0 56639 7 1 2 56544 56638
0 56640 5 1 1 56639
0 56641 7 1 2 73275 56640
0 56642 5 1 1 56641
0 56643 7 1 2 56505 56642
0 56644 5 1 1 56643
0 56645 7 1 2 67820 56644
0 56646 5 1 1 56645
0 56647 7 1 2 94815 78083
0 56648 7 1 2 86149 56647
0 56649 7 2 2 85420 92413
0 56650 7 1 2 95763 106760
0 56651 7 1 2 106793 56650
0 56652 7 1 2 56648 56651
0 56653 5 1 1 56652
0 56654 7 1 2 56646 56653
0 56655 7 1 2 56454 56654
0 56656 5 1 1 56655
0 56657 7 1 2 63812 56656
0 56658 5 1 1 56657
0 56659 7 2 2 103940 74267
0 56660 5 1 1 106795
0 56661 7 1 2 65217 106796
0 56662 5 2 1 56661
0 56663 7 1 2 103953 94843
0 56664 5 1 1 56663
0 56665 7 1 2 56660 56664
0 56666 5 1 1 56665
0 56667 7 1 2 88695 56666
0 56668 5 1 1 56667
0 56669 7 1 2 106797 56668
0 56670 5 1 1 56669
0 56671 7 1 2 73612 56670
0 56672 5 1 1 56671
0 56673 7 1 2 75198 94498
0 56674 5 1 1 56673
0 56675 7 1 2 13348 56674
0 56676 5 1 1 56675
0 56677 7 2 2 103930 56676
0 56678 7 1 2 98336 106799
0 56679 5 1 1 56678
0 56680 7 1 2 56672 56679
0 56681 5 1 1 56680
0 56682 7 1 2 66393 56681
0 56683 5 1 1 56682
0 56684 7 1 2 88711 80105
0 56685 5 1 1 56684
0 56686 7 1 2 68528 90465
0 56687 5 1 1 56686
0 56688 7 1 2 66394 56687
0 56689 5 1 1 56688
0 56690 7 1 2 66796 100058
0 56691 5 1 1 56690
0 56692 7 1 2 56689 56691
0 56693 5 1 1 56692
0 56694 7 1 2 65522 56693
0 56695 5 1 1 56694
0 56696 7 1 2 56685 56695
0 56697 5 1 1 56696
0 56698 7 1 2 76776 56697
0 56699 5 1 1 56698
0 56700 7 1 2 94042 74268
0 56701 5 1 1 56700
0 56702 7 1 2 56699 56701
0 56703 5 1 1 56702
0 56704 7 1 2 103954 56703
0 56705 5 1 1 56704
0 56706 7 1 2 85644 83080
0 56707 5 1 1 56706
0 56708 7 1 2 65218 56707
0 56709 5 1 1 56708
0 56710 7 1 2 105745 56709
0 56711 5 1 1 56710
0 56712 7 1 2 106652 56711
0 56713 5 1 1 56712
0 56714 7 1 2 99570 99973
0 56715 7 1 2 101961 56714
0 56716 5 1 1 56715
0 56717 7 1 2 56713 56716
0 56718 5 1 1 56717
0 56719 7 1 2 75233 56718
0 56720 5 1 1 56719
0 56721 7 2 2 67141 103931
0 56722 7 1 2 83377 90032
0 56723 7 1 2 97112 56722
0 56724 7 1 2 106801 56723
0 56725 5 1 1 56724
0 56726 7 1 2 56720 56725
0 56727 7 1 2 56705 56726
0 56728 5 1 1 56727
0 56729 7 1 2 66614 56728
0 56730 5 1 1 56729
0 56731 7 1 2 56683 56730
0 56732 5 1 1 56731
0 56733 7 1 2 64907 56732
0 56734 5 1 1 56733
0 56735 7 1 2 103955 94847
0 56736 5 1 1 56735
0 56737 7 1 2 106798 56736
0 56738 5 1 1 56737
0 56739 7 1 2 82938 56738
0 56740 5 1 1 56739
0 56741 7 2 2 83378 102189
0 56742 7 1 2 105002 106803
0 56743 5 1 1 56742
0 56744 7 1 2 56740 56743
0 56745 5 1 1 56744
0 56746 7 1 2 65523 56745
0 56747 5 1 1 56746
0 56748 7 3 2 66797 67229
0 56749 7 2 2 74256 106805
0 56750 7 1 2 106804 106808
0 56751 5 1 1 56750
0 56752 7 1 2 56747 56751
0 56753 5 1 1 56752
0 56754 7 1 2 77053 56753
0 56755 5 1 1 56754
0 56756 7 1 2 56734 56755
0 56757 5 1 1 56756
0 56758 7 1 2 73276 56757
0 56759 5 1 1 56758
0 56760 7 2 2 103314 103206
0 56761 7 1 2 106558 106810
0 56762 5 1 1 56761
0 56763 7 1 2 13386 51516
0 56764 5 1 1 56763
0 56765 7 1 2 106653 56764
0 56766 5 1 1 56765
0 56767 7 1 2 56762 56766
0 56768 5 1 1 56767
0 56769 7 1 2 73613 56768
0 56770 5 1 1 56769
0 56771 7 2 2 82477 77836
0 56772 7 1 2 85429 104608
0 56773 7 1 2 106812 56772
0 56774 5 1 1 56773
0 56775 7 1 2 56770 56774
0 56776 5 1 1 56775
0 56777 7 1 2 73791 56776
0 56778 5 1 1 56777
0 56779 7 1 2 92829 75234
0 56780 7 1 2 106811 56779
0 56781 5 1 1 56780
0 56782 7 1 2 56778 56781
0 56783 5 1 1 56782
0 56784 7 1 2 64908 56783
0 56785 5 1 1 56784
0 56786 7 1 2 105003 95536
0 56787 7 1 2 102192 56786
0 56788 5 1 1 56787
0 56789 7 1 2 56785 56788
0 56790 5 1 1 56789
0 56791 7 1 2 87461 56790
0 56792 5 1 1 56791
0 56793 7 2 2 94722 103924
0 56794 5 1 1 106814
0 56795 7 1 2 78558 106815
0 56796 5 1 1 56795
0 56797 7 1 2 64211 106800
0 56798 5 1 1 56797
0 56799 7 1 2 56796 56798
0 56800 5 1 1 56799
0 56801 7 1 2 65219 56800
0 56802 5 1 1 56801
0 56803 7 1 2 75108 102190
0 56804 7 1 2 106809 56803
0 56805 5 1 1 56804
0 56806 7 1 2 56802 56805
0 56807 5 1 1 56806
0 56808 7 1 2 77969 56807
0 56809 5 1 1 56808
0 56810 7 1 2 67821 56809
0 56811 7 1 2 56792 56810
0 56812 7 1 2 56759 56811
0 56813 5 1 1 56812
0 56814 7 1 2 101133 106694
0 56815 5 1 1 56814
0 56816 7 1 2 106692 56815
0 56817 5 1 1 56816
0 56818 7 1 2 75235 56817
0 56819 5 1 1 56818
0 56820 7 1 2 101134 106741
0 56821 5 1 1 56820
0 56822 7 1 2 95170 106654
0 56823 5 1 1 56822
0 56824 7 1 2 56821 56823
0 56825 5 1 1 56824
0 56826 7 1 2 80656 56825
0 56827 5 1 1 56826
0 56828 7 1 2 80776 103956
0 56829 5 1 1 56828
0 56830 7 1 2 106680 56829
0 56831 5 1 1 56830
0 56832 7 1 2 73614 56831
0 56833 5 1 1 56832
0 56834 7 1 2 56794 56833
0 56835 5 1 1 56834
0 56836 7 1 2 70030 56835
0 56837 5 1 1 56836
0 56838 7 1 2 83072 106715
0 56839 5 1 1 56838
0 56840 7 1 2 56837 56839
0 56841 5 1 1 56840
0 56842 7 1 2 68203 56841
0 56843 5 1 1 56842
0 56844 7 1 2 56827 56843
0 56845 5 1 1 56844
0 56846 7 1 2 74711 56845
0 56847 5 1 1 56846
0 56848 7 1 2 99648 106708
0 56849 5 1 1 56848
0 56850 7 1 2 68204 106706
0 56851 5 1 1 56850
0 56852 7 1 2 78749 98799
0 56853 5 1 1 56852
0 56854 7 1 2 56851 56853
0 56855 5 1 1 56854
0 56856 7 1 2 106655 56855
0 56857 5 1 1 56856
0 56858 7 1 2 56849 56857
0 56859 7 1 2 56847 56858
0 56860 5 1 1 56859
0 56861 7 1 2 76777 56860
0 56862 5 1 1 56861
0 56863 7 1 2 56819 56862
0 56864 5 1 1 56863
0 56865 7 1 2 66395 56864
0 56866 5 1 1 56865
0 56867 7 1 2 104148 106656
0 56868 5 1 1 56867
0 56869 7 1 2 83445 83692
0 56870 5 1 1 56869
0 56871 7 1 2 93887 104289
0 56872 7 1 2 56870 56871
0 56873 5 1 1 56872
0 56874 7 1 2 56868 56873
0 56875 5 1 1 56874
0 56876 7 1 2 65220 56875
0 56877 5 1 1 56876
0 56878 7 1 2 104144 106657
0 56879 5 1 1 56878
0 56880 7 1 2 56877 56879
0 56881 5 1 1 56880
0 56882 7 1 2 79434 56881
0 56883 5 1 1 56882
0 56884 7 1 2 68205 97835
0 56885 5 1 1 56884
0 56886 7 1 2 94882 56885
0 56887 5 1 1 56886
0 56888 7 1 2 106658 56887
0 56889 5 1 1 56888
0 56890 7 1 2 99649 106712
0 56891 5 1 1 56890
0 56892 7 1 2 99650 98980
0 56893 5 1 1 56892
0 56894 7 1 2 83481 106659
0 56895 5 1 1 56894
0 56896 7 1 2 56893 56895
0 56897 5 1 1 56896
0 56898 7 1 2 75052 56897
0 56899 5 1 1 56898
0 56900 7 1 2 56891 56899
0 56901 7 1 2 56889 56900
0 56902 5 1 1 56901
0 56903 7 1 2 64909 56902
0 56904 5 1 1 56903
0 56905 7 1 2 101390 96619
0 56906 5 1 1 56905
0 56907 7 1 2 86483 56906
0 56908 5 1 1 56907
0 56909 7 1 2 103957 56908
0 56910 5 1 1 56909
0 56911 7 1 2 81795 106660
0 56912 5 1 1 56911
0 56913 7 1 2 74712 99651
0 56914 5 1 1 56913
0 56915 7 1 2 56912 56914
0 56916 5 1 1 56915
0 56917 7 1 2 106700 56916
0 56918 5 1 1 56917
0 56919 7 1 2 56910 56918
0 56920 5 1 1 56919
0 56921 7 1 2 73615 56920
0 56922 5 1 1 56921
0 56923 7 1 2 100714 101966
0 56924 7 1 2 105303 56923
0 56925 5 1 1 56924
0 56926 7 1 2 56922 56925
0 56927 7 1 2 56904 56926
0 56928 5 1 1 56927
0 56929 7 1 2 71505 56928
0 56930 5 1 1 56929
0 56931 7 1 2 56883 56930
0 56932 5 1 1 56931
0 56933 7 1 2 76778 56932
0 56934 5 1 1 56933
0 56935 7 1 2 71506 101841
0 56936 5 1 1 56935
0 56937 7 1 2 56031 56936
0 56938 5 1 1 56937
0 56939 7 1 2 99652 56938
0 56940 5 1 1 56939
0 56941 7 1 2 100359 83824
0 56942 5 1 1 56941
0 56943 7 1 2 73792 13194
0 56944 5 1 1 56943
0 56945 7 1 2 73277 56944
0 56946 7 1 2 56942 56945
0 56947 5 1 1 56946
0 56948 7 1 2 95174 56947
0 56949 5 1 1 56948
0 56950 7 1 2 71507 56949
0 56951 5 1 1 56950
0 56952 7 1 2 79415 103216
0 56953 5 1 1 56952
0 56954 7 1 2 56951 56953
0 56955 7 1 2 106690 56954
0 56956 5 1 1 56955
0 56957 7 1 2 106661 56956
0 56958 5 1 1 56957
0 56959 7 1 2 56940 56958
0 56960 5 1 1 56959
0 56961 7 1 2 75236 56960
0 56962 5 1 1 56961
0 56963 7 1 2 72808 56962
0 56964 7 1 2 56934 56963
0 56965 7 1 2 56866 56964
0 56966 5 1 1 56965
0 56967 7 1 2 56813 56966
0 56968 5 1 1 56967
0 56969 7 1 2 82478 103052
0 56970 5 1 1 56969
0 56971 7 1 2 106728 56970
0 56972 5 2 1 56971
0 56973 7 1 2 84262 94358
0 56974 5 1 1 56973
0 56975 7 1 2 82204 56974
0 56976 5 1 1 56975
0 56977 7 1 2 81796 93025
0 56978 5 1 1 56977
0 56979 7 1 2 56976 56978
0 56980 5 1 1 56979
0 56981 7 1 2 64910 56980
0 56982 5 1 1 56981
0 56983 7 1 2 100929 79550
0 56984 5 1 1 56983
0 56985 7 1 2 65524 95321
0 56986 7 1 2 56984 56985
0 56987 5 1 1 56986
0 56988 7 1 2 56982 56987
0 56989 5 1 1 56988
0 56990 7 1 2 75237 56989
0 56991 5 1 1 56990
0 56992 7 1 2 69024 89647
0 56993 7 1 2 103411 56992
0 56994 7 1 2 93504 56993
0 56995 5 1 1 56994
0 56996 7 1 2 56991 56995
0 56997 5 1 1 56996
0 56998 7 1 2 106816 56997
0 56999 5 1 1 56998
0 57000 7 1 2 67230 87017
0 57001 7 1 2 102846 57000
0 57002 7 1 2 106794 57001
0 57003 7 1 2 106584 57002
0 57004 5 1 1 57003
0 57005 7 1 2 56999 57004
0 57006 7 1 2 56968 57005
0 57007 5 1 1 57006
0 57008 7 1 2 79645 57007
0 57009 5 1 1 57008
0 57010 7 1 2 72809 106688
0 57011 5 1 1 57010
0 57012 7 2 2 103574 103958
0 57013 7 1 2 99790 106818
0 57014 5 1 1 57013
0 57015 7 1 2 57011 57014
0 57016 5 1 1 57015
0 57017 7 1 2 85990 75884
0 57018 7 1 2 57016 57017
0 57019 5 1 1 57018
0 57020 7 1 2 57009 57019
0 57021 5 1 1 57020
0 57022 7 1 2 73879 57021
0 57023 5 1 1 57022
0 57024 7 2 2 85972 105639
0 57025 7 1 2 95395 106820
0 57026 5 1 1 57025
0 57027 7 1 2 90449 98679
0 57028 5 1 1 57027
0 57029 7 1 2 106774 57028
0 57030 5 1 1 57029
0 57031 7 1 2 65221 57030
0 57032 5 1 1 57031
0 57033 7 1 2 90592 74257
0 57034 7 1 2 87462 57033
0 57035 7 1 2 91357 57034
0 57036 5 1 1 57035
0 57037 7 1 2 57032 57036
0 57038 5 1 1 57037
0 57039 7 1 2 83943 57038
0 57040 5 1 1 57039
0 57041 7 1 2 57026 57040
0 57042 5 1 1 57041
0 57043 7 1 2 73278 57042
0 57044 5 1 1 57043
0 57045 7 1 2 101414 85052
0 57046 5 1 1 57045
0 57047 7 1 2 64911 57046
0 57048 5 1 1 57047
0 57049 7 1 2 92929 85028
0 57050 5 2 1 57049
0 57051 7 1 2 57048 106822
0 57052 5 1 1 57051
0 57053 7 1 2 106821 57052
0 57054 5 1 1 57053
0 57055 7 1 2 57044 57054
0 57056 5 1 1 57055
0 57057 7 1 2 63813 57056
0 57058 5 1 1 57057
0 57059 7 1 2 65694 75943
0 57060 7 1 2 102198 57059
0 57061 7 1 2 91206 84025
0 57062 7 1 2 57060 57061
0 57063 5 1 1 57062
0 57064 7 1 2 57058 57063
0 57065 5 1 1 57064
0 57066 7 1 2 106817 57065
0 57067 5 1 1 57066
0 57068 7 1 2 72810 56445
0 57069 5 1 1 57068
0 57070 7 1 2 95826 106676
0 57071 5 1 1 57070
0 57072 7 1 2 106782 57071
0 57073 5 1 1 57072
0 57074 7 1 2 73995 57073
0 57075 5 1 1 57074
0 57076 7 1 2 78713 87294
0 57077 5 1 1 57076
0 57078 7 1 2 89102 57077
0 57079 5 1 1 57078
0 57080 7 1 2 92695 106571
0 57081 5 1 1 57080
0 57082 7 1 2 57079 57081
0 57083 5 1 1 57082
0 57084 7 1 2 103959 57083
0 57085 5 1 1 57084
0 57086 7 1 2 99427 95827
0 57087 7 1 2 106662 57086
0 57088 5 1 1 57087
0 57089 7 1 2 57085 57088
0 57090 7 1 2 57075 57089
0 57091 5 1 1 57090
0 57092 7 1 2 81159 57091
0 57093 5 1 1 57092
0 57094 7 1 2 66798 81303
0 57095 5 1 1 57094
0 57096 7 1 2 15345 57095
0 57097 5 1 1 57096
0 57098 7 1 2 103960 94007
0 57099 7 1 2 57097 57098
0 57100 5 1 1 57099
0 57101 7 1 2 57093 57100
0 57102 5 1 1 57101
0 57103 7 1 2 67822 57102
0 57104 5 1 1 57103
0 57105 7 1 2 72811 106736
0 57106 5 1 1 57105
0 57107 7 1 2 89889 106819
0 57108 5 1 1 57107
0 57109 7 1 2 57106 57108
0 57110 5 1 1 57109
0 57111 7 1 2 80777 57110
0 57112 5 1 1 57111
0 57113 7 1 2 57104 57112
0 57114 7 1 2 57069 57113
0 57115 5 1 1 57114
0 57116 7 1 2 101988 90323
0 57117 7 1 2 57115 57116
0 57118 5 1 1 57117
0 57119 7 1 2 57067 57118
0 57120 7 1 2 57023 57119
0 57121 7 1 2 56658 57120
0 57122 5 1 1 57121
0 57123 7 1 2 66899 57122
0 57124 5 1 1 57123
0 57125 7 1 2 55839 57124
0 57126 5 1 1 57125
0 57127 7 1 2 67478 57126
0 57128 5 1 1 57127
0 57129 7 1 2 77127 106758
0 57130 5 1 1 57129
0 57131 7 1 2 76691 90176
0 57132 5 1 1 57131
0 57133 7 1 2 74713 90616
0 57134 5 1 1 57133
0 57135 7 1 2 57132 57134
0 57136 5 1 1 57135
0 57137 7 1 2 80657 57136
0 57138 5 1 1 57137
0 57139 7 1 2 93823 92702
0 57140 5 1 1 57139
0 57141 7 1 2 57138 57140
0 57142 5 1 1 57141
0 57143 7 1 2 99653 57142
0 57144 5 1 1 57143
0 57145 7 1 2 57130 57144
0 57146 5 2 1 57145
0 57147 7 2 2 90507 106824
0 57148 7 1 2 89530 106826
0 57149 5 1 1 57148
0 57150 7 1 2 74480 106825
0 57151 5 1 1 57150
0 57152 7 1 2 82828 89297
0 57153 7 1 2 8495 57152
0 57154 7 1 2 103961 57153
0 57155 5 1 1 57154
0 57156 7 1 2 57151 57155
0 57157 5 1 1 57156
0 57158 7 1 2 71508 57157
0 57159 5 1 1 57158
0 57160 7 1 2 68529 90408
0 57161 5 1 1 57160
0 57162 7 1 2 106120 57161
0 57163 5 1 1 57162
0 57164 7 1 2 99654 57163
0 57165 5 1 1 57164
0 57166 7 1 2 92843 84331
0 57167 7 1 2 103097 57166
0 57168 5 1 1 57167
0 57169 7 1 2 57165 57168
0 57170 5 2 1 57169
0 57171 7 1 2 71711 106828
0 57172 5 1 1 57171
0 57173 7 1 2 99655 88274
0 57174 7 1 2 95782 57173
0 57175 5 1 1 57174
0 57176 7 1 2 57172 57175
0 57177 5 1 1 57176
0 57178 7 2 2 67011 57177
0 57179 7 1 2 65614 106830
0 57180 5 1 1 57179
0 57181 7 1 2 57159 57180
0 57182 5 1 1 57181
0 57183 7 1 2 91544 57182
0 57184 5 1 1 57183
0 57185 7 1 2 57149 57184
0 57186 5 1 1 57185
0 57187 7 1 2 70031 57186
0 57188 5 1 1 57187
0 57189 7 1 2 92032 106831
0 57190 5 1 1 57189
0 57191 7 1 2 57188 57190
0 57192 5 1 1 57191
0 57193 7 1 2 63814 57192
0 57194 5 1 1 57193
0 57195 7 1 2 90794 106827
0 57196 5 1 1 57195
0 57197 7 1 2 57194 57196
0 57198 5 1 1 57197
0 57199 7 1 2 66900 57198
0 57200 5 1 1 57199
0 57201 7 1 2 79330 103899
0 57202 7 2 2 83707 57201
0 57203 7 1 2 82879 93612
0 57204 7 1 2 82778 90269
0 57205 7 1 2 57203 57204
0 57206 7 1 2 106832 57205
0 57207 7 1 2 90398 57206
0 57208 5 1 1 57207
0 57209 7 1 2 57200 57208
0 57210 5 1 1 57209
0 57211 7 1 2 68206 57210
0 57212 5 1 1 57211
0 57213 7 1 2 95696 106618
0 57214 7 1 2 106829 57213
0 57215 5 1 1 57214
0 57216 7 1 2 57212 57215
0 57217 5 1 1 57216
0 57218 7 1 2 97062 57217
0 57219 5 1 1 57218
0 57220 7 1 2 96243 104992
0 57221 7 1 2 84239 57220
0 57222 5 1 1 57221
0 57223 7 4 2 67012 102644
0 57224 7 1 2 101874 106834
0 57225 7 1 2 101477 57224
0 57226 5 1 1 57225
0 57227 7 1 2 57222 57226
0 57228 5 1 1 57227
0 57229 7 1 2 66615 57228
0 57230 5 1 1 57229
0 57231 7 1 2 101576 90033
0 57232 7 1 2 103640 57231
0 57233 7 1 2 104315 57232
0 57234 5 1 1 57233
0 57235 7 1 2 57230 57234
0 57236 5 1 1 57235
0 57237 7 1 2 65222 57236
0 57238 5 1 1 57237
0 57239 7 1 2 82175 84269
0 57240 7 1 2 106756 57239
0 57241 5 1 1 57240
0 57242 7 1 2 57238 57241
0 57243 5 1 1 57242
0 57244 7 1 2 68207 57243
0 57245 5 1 1 57244
0 57246 7 1 2 91333 106813
0 57247 7 1 2 106835 57246
0 57248 7 1 2 101306 57247
0 57249 5 1 1 57248
0 57250 7 1 2 57245 57249
0 57251 5 1 1 57250
0 57252 7 1 2 73793 57251
0 57253 5 1 1 57252
0 57254 7 1 2 97426 84560
0 57255 5 1 1 57254
0 57256 7 1 2 84433 57255
0 57257 5 1 1 57256
0 57258 7 1 2 104158 105765
0 57259 7 1 2 57257 57258
0 57260 5 1 1 57259
0 57261 7 1 2 57253 57260
0 57262 5 1 1 57261
0 57263 7 1 2 72812 57262
0 57264 5 1 1 57263
0 57265 7 1 2 70919 89818
0 57266 7 1 2 104999 86432
0 57267 7 2 2 57265 57266
0 57268 7 1 2 105693 106838
0 57269 5 1 1 57268
0 57270 7 1 2 57264 57269
0 57271 5 1 1 57270
0 57272 7 1 2 67479 57271
0 57273 5 1 1 57272
0 57274 7 2 2 98605 78396
0 57275 7 1 2 96805 103765
0 57276 7 2 2 105000 57275
0 57277 7 1 2 69025 106842
0 57278 5 1 1 57277
0 57279 7 1 2 71712 77844
0 57280 5 1 1 57279
0 57281 7 1 2 95239 57280
0 57282 5 1 1 57281
0 57283 7 1 2 106663 57282
0 57284 5 1 1 57283
0 57285 7 1 2 57278 57284
0 57286 5 1 1 57285
0 57287 7 1 2 106840 57286
0 57288 5 1 1 57287
0 57289 7 1 2 57273 57288
0 57290 5 1 1 57289
0 57291 7 1 2 74042 57290
0 57292 5 1 1 57291
0 57293 7 1 2 103941 106266
0 57294 5 1 1 57293
0 57295 7 1 2 101577 95919
0 57296 7 1 2 106559 57295
0 57297 5 1 1 57296
0 57298 7 1 2 57294 57297
0 57299 5 1 1 57298
0 57300 7 1 2 81576 57299
0 57301 5 1 1 57300
0 57302 7 1 2 92466 92067
0 57303 7 1 2 104821 57302
0 57304 7 1 2 94106 57303
0 57305 5 1 1 57304
0 57306 7 1 2 57301 57305
0 57307 5 1 1 57306
0 57308 7 1 2 67480 95423
0 57309 7 1 2 57307 57308
0 57310 5 1 1 57309
0 57311 7 1 2 57292 57310
0 57312 5 1 1 57311
0 57313 7 1 2 73880 57312
0 57314 5 1 1 57313
0 57315 7 1 2 87212 104271
0 57316 5 1 1 57315
0 57317 7 1 2 73794 105731
0 57318 7 1 2 90439 57317
0 57319 7 1 2 57316 57318
0 57320 5 1 1 57319
0 57321 7 1 2 97107 93176
0 57322 7 1 2 95730 57321
0 57323 7 1 2 91664 105468
0 57324 7 1 2 57322 57323
0 57325 5 1 1 57324
0 57326 7 1 2 57320 57325
0 57327 5 1 1 57326
0 57328 7 1 2 68530 57327
0 57329 5 1 1 57328
0 57330 7 1 2 97427 91520
0 57331 5 1 1 57330
0 57332 7 1 2 91581 57331
0 57333 5 1 1 57332
0 57334 7 1 2 86258 57333
0 57335 5 1 1 57334
0 57336 7 1 2 76615 75053
0 57337 7 1 2 91381 57336
0 57338 5 1 1 57337
0 57339 7 1 2 57335 57338
0 57340 5 1 1 57339
0 57341 7 1 2 67481 90851
0 57342 7 1 2 57340 57341
0 57343 5 1 1 57342
0 57344 7 1 2 57329 57343
0 57345 5 1 1 57344
0 57346 7 1 2 68208 57345
0 57347 5 1 1 57346
0 57348 7 1 2 101170 106255
0 57349 5 1 1 57348
0 57350 7 1 2 77287 91256
0 57351 7 1 2 90747 57350
0 57352 5 1 1 57351
0 57353 7 1 2 57349 57352
0 57354 5 1 1 57353
0 57355 7 1 2 65223 57354
0 57356 5 1 1 57355
0 57357 7 1 2 73795 77555
0 57358 7 1 2 89006 57357
0 57359 5 1 1 57358
0 57360 7 1 2 57356 57359
0 57361 5 1 1 57360
0 57362 7 1 2 68531 57361
0 57363 5 1 1 57362
0 57364 7 1 2 100324 84510
0 57365 7 1 2 91931 57364
0 57366 5 1 1 57365
0 57367 7 1 2 57363 57366
0 57368 5 1 1 57367
0 57369 7 1 2 72813 57368
0 57370 5 1 1 57369
0 57371 7 1 2 76692 106384
0 57372 7 1 2 87209 57371
0 57373 5 1 1 57372
0 57374 7 1 2 57370 57373
0 57375 5 1 1 57374
0 57376 7 1 2 88275 57375
0 57377 5 1 1 57376
0 57378 7 1 2 66901 81322
0 57379 7 1 2 95393 57378
0 57380 7 1 2 106479 57379
0 57381 5 1 1 57380
0 57382 7 1 2 57377 57381
0 57383 5 1 1 57382
0 57384 7 1 2 100128 57383
0 57385 5 1 1 57384
0 57386 7 1 2 57347 57385
0 57387 5 1 1 57386
0 57388 7 1 2 106664 57387
0 57389 5 1 1 57388
0 57390 7 1 2 100330 96772
0 57391 5 1 1 57390
0 57392 7 1 2 33966 57391
0 57393 5 1 1 57392
0 57394 7 1 2 65224 57393
0 57395 5 1 1 57394
0 57396 7 1 2 70277 79582
0 57397 7 1 2 98568 57396
0 57398 5 1 1 57397
0 57399 7 1 2 57395 57398
0 57400 5 1 1 57399
0 57401 7 1 2 70032 57400
0 57402 5 1 1 57401
0 57403 7 1 2 72814 101348
0 57404 5 1 1 57403
0 57405 7 1 2 32259 57404
0 57406 5 1 1 57405
0 57407 7 1 2 67482 78326
0 57408 7 1 2 57406 57407
0 57409 5 1 1 57408
0 57410 7 1 2 57402 57409
0 57411 5 1 1 57410
0 57412 7 1 2 73796 91912
0 57413 7 1 2 57411 57412
0 57414 5 1 1 57413
0 57415 7 1 2 90792 106299
0 57416 7 1 2 104661 57415
0 57417 5 1 1 57416
0 57418 7 1 2 57414 57417
0 57419 5 1 1 57418
0 57420 7 1 2 106779 57419
0 57421 5 1 1 57420
0 57422 7 1 2 78906 106734
0 57423 5 1 1 57422
0 57424 7 1 2 81577 106780
0 57425 5 1 1 57424
0 57426 7 1 2 57423 57425
0 57427 5 1 1 57426
0 57428 7 1 2 95936 57427
0 57429 5 1 1 57428
0 57430 7 1 2 101171 106753
0 57431 5 1 1 57430
0 57432 7 1 2 76165 103315
0 57433 7 1 2 103641 57432
0 57434 5 1 1 57433
0 57435 7 1 2 57431 57434
0 57436 5 1 1 57435
0 57437 7 1 2 87752 104316
0 57438 7 1 2 57436 57437
0 57439 5 1 1 57438
0 57440 7 1 2 57429 57439
0 57441 5 1 1 57440
0 57442 7 1 2 65225 57441
0 57443 5 1 1 57442
0 57444 7 1 2 96162 91025
0 57445 7 2 2 67231 76166
0 57446 7 1 2 92856 106844
0 57447 7 1 2 57444 57446
0 57448 5 1 1 57447
0 57449 7 1 2 57443 57448
0 57450 5 1 1 57449
0 57451 7 1 2 68532 57450
0 57452 5 1 1 57451
0 57453 7 1 2 75301 87753
0 57454 7 1 2 94097 57453
0 57455 7 1 2 106754 57454
0 57456 7 1 2 99965 57455
0 57457 5 1 1 57456
0 57458 7 1 2 57452 57457
0 57459 5 1 1 57458
0 57460 7 1 2 72815 57459
0 57461 5 1 1 57460
0 57462 7 1 2 106483 106839
0 57463 5 1 1 57462
0 57464 7 1 2 57461 57463
0 57465 5 1 1 57464
0 57466 7 1 2 67483 57465
0 57467 5 1 1 57466
0 57468 7 1 2 87754 106843
0 57469 5 1 1 57468
0 57470 7 1 2 74223 90625
0 57471 5 1 1 57470
0 57472 7 1 2 68893 92068
0 57473 7 1 2 104317 57472
0 57474 5 1 1 57473
0 57475 7 1 2 57471 57474
0 57476 5 1 1 57475
0 57477 7 1 2 106665 57476
0 57478 5 1 1 57477
0 57479 7 1 2 57469 57478
0 57480 5 1 1 57479
0 57481 7 1 2 57480 106841
0 57482 5 1 1 57481
0 57483 7 1 2 57467 57482
0 57484 5 1 1 57483
0 57485 7 1 2 89588 57484
0 57486 5 1 1 57485
0 57487 7 1 2 57421 57486
0 57488 7 1 2 57389 57487
0 57489 7 1 2 57314 57488
0 57490 5 1 1 57489
0 57491 7 1 2 84876 57490
0 57492 5 1 1 57491
0 57493 7 2 2 72487 106731
0 57494 7 1 2 103434 38338
0 57495 5 1 1 57494
0 57496 7 1 2 76737 57495
0 57497 5 1 1 57496
0 57498 7 1 2 68533 74288
0 57499 7 1 2 91971 57498
0 57500 7 1 2 87602 57499
0 57501 5 1 1 57500
0 57502 7 1 2 57497 57501
0 57503 5 1 1 57502
0 57504 7 1 2 64912 57503
0 57505 5 1 1 57504
0 57506 7 1 2 79094 104243
0 57507 7 1 2 97934 57506
0 57508 5 1 1 57507
0 57509 7 1 2 57505 57508
0 57510 5 1 1 57509
0 57511 7 1 2 68209 57510
0 57512 5 1 1 57511
0 57513 7 1 2 75839 103197
0 57514 7 1 2 104350 57513
0 57515 5 1 1 57514
0 57516 7 1 2 57512 57515
0 57517 5 1 1 57516
0 57518 7 1 2 72816 57517
0 57519 5 1 1 57518
0 57520 7 1 2 96167 105278
0 57521 7 1 2 104351 57520
0 57522 5 1 1 57521
0 57523 7 1 2 57519 57522
0 57524 5 1 1 57523
0 57525 7 1 2 106846 57524
0 57526 5 1 1 57525
0 57527 7 2 2 67142 86572
0 57528 7 2 2 77683 106848
0 57529 7 1 2 95667 106850
0 57530 5 1 1 57529
0 57531 7 1 2 101478 74123
0 57532 5 1 1 57531
0 57533 7 1 2 87622 92376
0 57534 5 1 1 57533
0 57535 7 1 2 57532 57534
0 57536 5 1 1 57535
0 57537 7 1 2 68210 57536
0 57538 5 1 1 57537
0 57539 7 1 2 57530 57538
0 57540 5 1 1 57539
0 57541 7 1 2 66616 57540
0 57542 5 1 1 57541
0 57543 7 1 2 79745 74105
0 57544 7 1 2 93537 57543
0 57545 7 2 2 101924 57544
0 57546 7 1 2 69026 106852
0 57547 5 1 1 57546
0 57548 7 1 2 57542 57547
0 57549 5 1 1 57548
0 57550 7 1 2 72817 57549
0 57551 5 1 1 57550
0 57552 7 1 2 78357 104663
0 57553 7 1 2 106567 57552
0 57554 5 1 1 57553
0 57555 7 1 2 57551 57554
0 57556 5 1 1 57555
0 57557 7 1 2 100429 57556
0 57558 5 1 1 57557
0 57559 7 2 2 102864 104672
0 57560 7 1 2 95379 86017
0 57561 7 1 2 106854 57560
0 57562 5 1 1 57561
0 57563 7 1 2 57558 57562
0 57564 5 1 1 57563
0 57565 7 1 2 84877 57564
0 57566 5 1 1 57565
0 57567 7 1 2 74982 101195
0 57568 5 1 1 57567
0 57569 7 1 2 104279 57568
0 57570 5 1 1 57569
0 57571 7 1 2 70033 57570
0 57572 5 2 1 57571
0 57573 7 1 2 97365 101953
0 57574 5 1 1 57573
0 57575 7 1 2 106856 57574
0 57576 5 1 1 57575
0 57577 7 1 2 86076 57576
0 57578 5 1 1 57577
0 57579 7 2 2 100430 85029
0 57580 7 2 2 66396 87094
0 57581 7 1 2 106858 106860
0 57582 5 1 1 57581
0 57583 7 1 2 57578 57582
0 57584 5 1 1 57583
0 57585 7 1 2 68534 57584
0 57586 5 1 1 57585
0 57587 7 1 2 85717 101520
0 57588 5 1 1 57587
0 57589 7 1 2 99940 57588
0 57590 5 1 1 57589
0 57591 7 1 2 72818 57590
0 57592 5 1 1 57591
0 57593 7 1 2 77684 83944
0 57594 5 1 1 57593
0 57595 7 1 2 57592 57594
0 57596 5 1 1 57595
0 57597 7 1 2 66617 57596
0 57598 5 1 1 57597
0 57599 7 1 2 77601 90814
0 57600 5 1 1 57599
0 57601 7 1 2 85030 101479
0 57602 5 1 1 57601
0 57603 7 1 2 57600 57602
0 57604 5 1 1 57603
0 57605 7 1 2 88408 57604
0 57606 5 1 1 57605
0 57607 7 1 2 57598 57606
0 57608 5 1 1 57607
0 57609 7 1 2 100431 57608
0 57610 5 1 1 57609
0 57611 7 1 2 57586 57610
0 57612 5 2 1 57611
0 57613 7 1 2 76738 106862
0 57614 5 1 1 57613
0 57615 7 1 2 86746 91458
0 57616 5 1 1 57615
0 57617 7 1 2 65525 97271
0 57618 5 1 1 57617
0 57619 7 1 2 57616 57618
0 57620 5 1 1 57619
0 57621 7 1 2 66397 57620
0 57622 5 1 1 57621
0 57623 7 2 2 82126 85031
0 57624 7 1 2 90016 106864
0 57625 5 1 1 57624
0 57626 7 1 2 57622 57625
0 57627 5 1 1 57626
0 57628 7 1 2 64913 57627
0 57629 5 1 1 57628
0 57630 7 1 2 106671 106865
0 57631 5 1 1 57630
0 57632 7 1 2 57629 57631
0 57633 5 1 1 57632
0 57634 7 3 2 100432 57633
0 57635 5 1 1 106866
0 57636 7 1 2 74124 106867
0 57637 5 1 1 57636
0 57638 7 1 2 57614 57637
0 57639 7 1 2 57566 57638
0 57640 5 1 1 57639
0 57641 7 1 2 65226 57640
0 57642 5 1 1 57641
0 57643 7 1 2 57526 57642
0 57644 5 1 1 57643
0 57645 7 1 2 74043 57644
0 57646 5 1 1 57645
0 57647 7 2 2 70034 94900
0 57648 5 1 1 106869
0 57649 7 1 2 79859 74983
0 57650 5 1 1 57649
0 57651 7 1 2 57648 57650
0 57652 5 1 1 57651
0 57653 7 1 2 73616 57652
0 57654 5 1 1 57653
0 57655 7 1 2 73797 78917
0 57656 5 1 1 57655
0 57657 7 1 2 57654 57656
0 57658 5 1 1 57657
0 57659 7 1 2 72819 57658
0 57660 5 1 1 57659
0 57661 7 1 2 91504 103398
0 57662 5 1 1 57661
0 57663 7 1 2 57660 57662
0 57664 5 1 1 57663
0 57665 7 1 2 81797 57664
0 57666 5 1 1 57665
0 57667 7 1 2 68535 81971
0 57668 5 1 1 57667
0 57669 7 1 2 83949 57668
0 57670 5 2 1 57669
0 57671 7 1 2 75302 106871
0 57672 5 1 1 57671
0 57673 7 1 2 87238 90815
0 57674 5 1 1 57673
0 57675 7 1 2 57672 57674
0 57676 5 1 1 57675
0 57677 7 1 2 73279 57676
0 57678 5 1 1 57677
0 57679 7 2 2 75584 79919
0 57680 5 1 1 106873
0 57681 7 1 2 98559 106874
0 57682 5 1 1 57681
0 57683 7 1 2 57678 57682
0 57684 5 1 1 57683
0 57685 7 1 2 80778 57684
0 57686 5 1 1 57685
0 57687 7 1 2 85053 104248
0 57688 5 1 1 57687
0 57689 7 1 2 64914 57688
0 57690 5 2 1 57689
0 57691 7 1 2 106823 106875
0 57692 5 1 1 57691
0 57693 7 1 2 74714 57692
0 57694 5 1 1 57693
0 57695 7 1 2 102093 86722
0 57696 5 1 1 57695
0 57697 7 1 2 57694 57696
0 57698 5 1 1 57697
0 57699 7 1 2 73617 57698
0 57700 5 1 1 57699
0 57701 7 2 2 75610 88723
0 57702 7 1 2 106114 106877
0 57703 5 1 1 57702
0 57704 7 1 2 57700 57703
0 57705 7 1 2 57686 57704
0 57706 7 1 2 57666 57705
0 57707 5 1 1 57706
0 57708 7 1 2 100433 57707
0 57709 5 1 1 57708
0 57710 7 1 2 77546 101196
0 57711 5 1 1 57710
0 57712 7 1 2 101925 102248
0 57713 5 1 1 57712
0 57714 7 1 2 57711 57713
0 57715 5 2 1 57714
0 57716 7 1 2 77128 106879
0 57717 5 1 1 57716
0 57718 7 1 2 99428 76053
0 57719 5 1 1 57718
0 57720 7 1 2 77288 79416
0 57721 5 1 1 57720
0 57722 7 2 2 57719 57721
0 57723 5 1 1 106881
0 57724 7 1 2 65227 57723
0 57725 5 1 1 57724
0 57726 7 1 2 77312 81185
0 57727 5 1 1 57726
0 57728 7 1 2 76107 57727
0 57729 5 1 1 57728
0 57730 7 1 2 4506 57729
0 57731 7 1 2 57725 57730
0 57732 5 1 1 57731
0 57733 7 1 2 101999 57732
0 57734 5 1 1 57733
0 57735 7 1 2 57717 57734
0 57736 5 1 1 57735
0 57737 7 1 2 80658 57736
0 57738 5 1 1 57737
0 57739 7 1 2 57709 57738
0 57740 5 1 1 57739
0 57741 7 1 2 76779 57740
0 57742 5 1 1 57741
0 57743 7 1 2 79882 104978
0 57744 5 1 1 57743
0 57745 7 1 2 66398 87479
0 57746 5 1 1 57745
0 57747 7 1 2 57744 57746
0 57748 5 1 1 57747
0 57749 7 1 2 64915 57748
0 57750 5 1 1 57749
0 57751 7 1 2 95194 87260
0 57752 5 1 1 57751
0 57753 7 1 2 67823 57752
0 57754 7 1 2 57750 57753
0 57755 5 1 1 57754
0 57756 7 1 2 95095 95433
0 57757 5 1 1 57756
0 57758 7 1 2 81798 104961
0 57759 5 1 1 57758
0 57760 7 1 2 72820 57759
0 57761 7 1 2 57757 57760
0 57762 5 1 1 57761
0 57763 7 1 2 73280 57762
0 57764 7 1 2 57755 57763
0 57765 5 1 1 57764
0 57766 7 1 2 92720 105953
0 57767 5 1 1 57766
0 57768 7 1 2 57765 57767
0 57769 5 1 1 57768
0 57770 7 1 2 100434 57769
0 57771 5 1 1 57770
0 57772 7 1 2 82181 105681
0 57773 7 1 2 106138 57772
0 57774 5 1 1 57773
0 57775 7 1 2 66399 57774
0 57776 5 1 1 57775
0 57777 7 1 2 81932 96029
0 57778 5 1 1 57777
0 57779 7 1 2 22566 82182
0 57780 5 1 1 57779
0 57781 7 1 2 85722 57780
0 57782 5 1 1 57781
0 57783 7 1 2 57778 57782
0 57784 7 1 2 57776 57783
0 57785 5 1 1 57784
0 57786 7 1 2 102249 57785
0 57787 5 1 1 57786
0 57788 7 1 2 81799 100435
0 57789 7 1 2 103677 57788
0 57790 5 1 1 57789
0 57791 7 1 2 70035 102166
0 57792 7 1 2 89037 57791
0 57793 5 1 1 57792
0 57794 7 1 2 57790 57793
0 57795 5 1 1 57794
0 57796 7 1 2 71509 57795
0 57797 5 1 1 57796
0 57798 7 1 2 14768 104921
0 57799 5 1 1 57798
0 57800 7 1 2 70278 104926
0 57801 7 1 2 57799 57800
0 57802 5 1 1 57801
0 57803 7 1 2 57797 57802
0 57804 7 1 2 57787 57803
0 57805 5 1 1 57804
0 57806 7 1 2 68211 57805
0 57807 5 1 1 57806
0 57808 7 1 2 101197 106186
0 57809 5 1 1 57808
0 57810 7 3 2 65526 106806
0 57811 7 1 2 82251 105672
0 57812 7 1 2 106883 57811
0 57813 5 1 1 57812
0 57814 7 1 2 57809 57813
0 57815 5 1 1 57814
0 57816 7 1 2 76346 57815
0 57817 5 1 1 57816
0 57818 7 1 2 71510 104051
0 57819 5 1 1 57818
0 57820 7 1 2 92170 57819
0 57821 5 1 1 57820
0 57822 7 1 2 101954 57821
0 57823 5 1 1 57822
0 57824 7 1 2 81619 104280
0 57825 5 1 1 57824
0 57826 7 1 2 70036 104283
0 57827 7 1 2 57825 57826
0 57828 5 1 1 57827
0 57829 7 1 2 57823 57828
0 57830 5 1 1 57829
0 57831 7 1 2 68536 57830
0 57832 5 1 1 57831
0 57833 7 1 2 104281 104922
0 57834 5 1 1 57833
0 57835 7 1 2 103439 57834
0 57836 5 1 1 57835
0 57837 7 1 2 57832 57836
0 57838 7 1 2 57817 57837
0 57839 7 1 2 57807 57838
0 57840 7 1 2 57771 57839
0 57841 5 1 1 57840
0 57842 7 1 2 75238 57841
0 57843 5 1 1 57842
0 57844 7 1 2 57742 57843
0 57845 5 1 1 57844
0 57846 7 1 2 78889 57845
0 57847 5 1 1 57846
0 57848 7 1 2 57646 57847
0 57849 5 1 1 57848
0 57850 7 1 2 73881 57849
0 57851 5 1 1 57850
0 57852 7 1 2 76108 83769
0 57853 5 1 1 57852
0 57854 7 1 2 106882 57853
0 57855 5 1 1 57854
0 57856 7 1 2 102250 57855
0 57857 5 1 1 57856
0 57858 7 1 2 106857 57857
0 57859 5 1 1 57858
0 57860 7 1 2 80659 57859
0 57861 5 1 1 57860
0 57862 7 1 2 99836 93338
0 57863 5 1 1 57862
0 57864 7 1 2 76693 78907
0 57865 5 1 1 57864
0 57866 7 1 2 57863 57865
0 57867 5 1 1 57866
0 57868 7 1 2 72821 57867
0 57869 5 1 1 57868
0 57870 7 1 2 91505 93297
0 57871 5 1 1 57870
0 57872 7 1 2 57869 57871
0 57873 5 1 1 57872
0 57874 7 1 2 81800 57873
0 57875 5 1 1 57874
0 57876 7 1 2 76054 79243
0 57877 5 1 1 57876
0 57878 7 1 2 57877 57680
0 57879 5 1 1 57878
0 57880 7 1 2 72822 57879
0 57881 5 1 1 57880
0 57882 7 1 2 73996 103575
0 57883 5 1 1 57882
0 57884 7 1 2 57881 57883
0 57885 5 1 1 57884
0 57886 7 1 2 80779 57885
0 57887 5 1 1 57886
0 57888 7 1 2 100703 85032
0 57889 5 1 1 57888
0 57890 7 1 2 77602 82205
0 57891 7 1 2 83829 57890
0 57892 5 1 1 57891
0 57893 7 1 2 44624 57892
0 57894 5 1 1 57893
0 57895 7 1 2 64916 57894
0 57896 5 1 1 57895
0 57897 7 1 2 57889 57896
0 57898 7 1 2 57887 57897
0 57899 7 1 2 57875 57898
0 57900 5 1 1 57899
0 57901 7 1 2 100436 57900
0 57902 5 1 1 57901
0 57903 7 1 2 57861 57902
0 57904 5 1 1 57903
0 57905 7 1 2 88276 57904
0 57906 5 1 1 57905
0 57907 7 1 2 88632 106863
0 57908 5 1 1 57907
0 57909 7 1 2 57906 57908
0 57910 5 1 1 57909
0 57911 7 1 2 78278 57910
0 57912 5 1 1 57911
0 57913 7 1 2 91473 106868
0 57914 5 1 1 57913
0 57915 7 1 2 101480 91474
0 57916 5 1 1 57915
0 57917 7 1 2 96246 90628
0 57918 5 1 1 57917
0 57919 7 1 2 57916 57918
0 57920 5 1 1 57919
0 57921 7 1 2 68212 57920
0 57922 5 1 1 57921
0 57923 7 1 2 84493 90871
0 57924 7 1 2 106851 57923
0 57925 5 1 1 57924
0 57926 7 1 2 57922 57925
0 57927 5 1 1 57926
0 57928 7 1 2 66618 57927
0 57929 5 1 1 57928
0 57930 7 1 2 87755 106853
0 57931 5 1 1 57930
0 57932 7 1 2 57929 57931
0 57933 5 1 1 57932
0 57934 7 1 2 72823 57933
0 57935 5 1 1 57934
0 57936 7 1 2 104022 91475
0 57937 5 1 1 57936
0 57938 7 1 2 57935 57937
0 57939 5 1 1 57938
0 57940 7 1 2 100437 57939
0 57941 5 1 1 57940
0 57942 7 1 2 83338 90270
0 57943 7 1 2 90087 57942
0 57944 7 1 2 106855 57943
0 57945 5 1 1 57944
0 57946 7 1 2 57941 57945
0 57947 5 1 1 57946
0 57948 7 1 2 84878 57947
0 57949 5 1 1 57948
0 57950 7 1 2 57914 57949
0 57951 7 1 2 57912 57950
0 57952 5 1 1 57951
0 57953 7 1 2 65228 57952
0 57954 5 1 1 57953
0 57955 7 1 2 77105 106880
0 57956 5 1 1 57955
0 57957 7 1 2 90924 3773
0 57958 5 1 1 57957
0 57959 7 1 2 104924 57958
0 57960 5 1 1 57959
0 57961 7 1 2 57956 57960
0 57962 5 1 1 57961
0 57963 7 1 2 80660 57962
0 57964 5 1 1 57963
0 57965 7 1 2 80780 90816
0 57966 5 1 1 57965
0 57967 7 1 2 89261 57966
0 57968 5 1 1 57967
0 57969 7 1 2 73618 57968
0 57970 5 1 1 57969
0 57971 7 1 2 83073 106872
0 57972 5 1 1 57971
0 57973 7 1 2 57970 57972
0 57974 5 1 1 57973
0 57975 7 1 2 73281 57974
0 57976 5 1 1 57975
0 57977 7 1 2 86297 88310
0 57978 5 1 1 57977
0 57979 7 1 2 27031 57978
0 57980 5 1 1 57979
0 57981 7 1 2 85033 57980
0 57982 5 1 1 57981
0 57983 7 1 2 57976 57982
0 57984 5 1 1 57983
0 57985 7 1 2 66619 57984
0 57986 5 1 1 57985
0 57987 7 1 2 72824 106870
0 57988 5 1 1 57987
0 57989 7 1 2 106876 57988
0 57990 5 1 1 57989
0 57991 7 1 2 85752 57990
0 57992 5 1 1 57991
0 57993 7 1 2 57986 57992
0 57994 5 1 1 57993
0 57995 7 1 2 100438 57994
0 57996 5 1 1 57995
0 57997 7 1 2 57964 57996
0 57998 5 1 1 57997
0 57999 7 1 2 88277 57998
0 58000 5 1 1 57999
0 58001 7 1 2 72825 101462
0 58002 5 1 1 58001
0 58003 7 1 2 103578 58002
0 58004 5 1 1 58003
0 58005 7 1 2 97935 58004
0 58006 5 1 1 58005
0 58007 7 1 2 92760 106861
0 58008 5 1 1 58007
0 58009 7 1 2 58006 58008
0 58010 5 1 1 58009
0 58011 7 1 2 88633 106847
0 58012 7 1 2 58010 58011
0 58013 5 1 1 58012
0 58014 7 1 2 58000 58013
0 58015 5 1 1 58014
0 58016 7 1 2 78279 58015
0 58017 5 1 1 58016
0 58018 7 1 2 87756 93435
0 58019 7 2 2 103900 97483
0 58020 7 1 2 94923 96040
0 58021 7 1 2 106886 58020
0 58022 7 1 2 58018 58021
0 58023 5 1 1 58022
0 58024 7 1 2 58017 58023
0 58025 7 1 2 57954 58024
0 58026 5 1 1 58025
0 58027 7 1 2 89589 58026
0 58028 5 1 1 58027
0 58029 7 1 2 76694 74984
0 58030 7 1 2 100086 83339
0 58031 7 1 2 58029 58030
0 58032 5 1 1 58031
0 58033 7 1 2 102139 58032
0 58034 5 1 1 58033
0 58035 7 1 2 67824 58034
0 58036 5 1 1 58035
0 58037 7 1 2 70037 87297
0 58038 5 1 1 58037
0 58039 7 1 2 97428 77615
0 58040 7 1 2 93339 58039
0 58041 5 1 1 58040
0 58042 7 1 2 83657 58041
0 58043 7 1 2 58038 58042
0 58044 5 1 1 58043
0 58045 7 1 2 102251 58044
0 58046 5 1 1 58045
0 58047 7 1 2 58036 58046
0 58048 5 1 1 58047
0 58049 7 1 2 84879 58048
0 58050 5 1 1 58049
0 58051 7 1 2 57635 58050
0 58052 5 1 1 58051
0 58053 7 1 2 65229 58052
0 58054 5 1 1 58053
0 58055 7 1 2 82014 92601
0 58056 7 1 2 102000 94908
0 58057 7 1 2 58055 58056
0 58058 5 1 1 58057
0 58059 7 1 2 58054 58058
0 58060 5 1 1 58059
0 58061 7 1 2 99115 58060
0 58062 5 1 1 58061
0 58063 7 1 2 80661 79971
0 58064 5 1 1 58063
0 58065 7 1 2 66400 96493
0 58066 5 1 1 58065
0 58067 7 1 2 58064 58066
0 58068 5 1 1 58067
0 58069 7 1 2 68537 58068
0 58070 5 1 1 58069
0 58071 7 1 2 75611 80487
0 58072 5 1 1 58071
0 58073 7 1 2 87658 58072
0 58074 5 1 1 58073
0 58075 7 1 2 66401 58074
0 58076 5 1 1 58075
0 58077 7 1 2 5871 77616
0 58078 5 1 1 58077
0 58079 7 1 2 80781 58078
0 58080 5 1 1 58079
0 58081 7 1 2 71511 629
0 58082 7 1 2 86126 58081
0 58083 7 1 2 58080 58082
0 58084 5 1 1 58083
0 58085 7 1 2 58076 58084
0 58086 5 1 1 58085
0 58087 7 1 2 58070 58086
0 58088 5 1 1 58087
0 58089 7 1 2 85344 58088
0 58090 5 1 1 58089
0 58091 7 1 2 73798 86309
0 58092 5 1 1 58091
0 58093 7 1 2 104146 58092
0 58094 5 1 1 58093
0 58095 7 1 2 76616 58094
0 58096 5 1 1 58095
0 58097 7 1 2 86331 58096
0 58098 5 1 1 58097
0 58099 7 1 2 65230 58098
0 58100 5 1 1 58099
0 58101 7 1 2 95098 103208
0 58102 5 1 1 58101
0 58103 7 1 2 79583 86381
0 58104 5 1 1 58103
0 58105 7 1 2 103465 58104
0 58106 7 1 2 58102 58105
0 58107 5 1 1 58106
0 58108 7 1 2 73619 58107
0 58109 5 1 1 58108
0 58110 7 1 2 66620 106698
0 58111 5 1 1 58110
0 58112 7 1 2 73799 86329
0 58113 5 1 1 58112
0 58114 7 1 2 68213 58113
0 58115 7 1 2 58111 58114
0 58116 7 1 2 58109 58115
0 58117 7 1 2 58100 58116
0 58118 5 1 1 58117
0 58119 7 1 2 97429 77129
0 58120 5 1 1 58119
0 58121 7 1 2 5376 58120
0 58122 5 1 1 58121
0 58123 7 1 2 80662 58122
0 58124 5 1 1 58123
0 58125 7 1 2 80782 79213
0 58126 5 1 1 58125
0 58127 7 1 2 85585 58126
0 58128 5 1 1 58127
0 58129 7 1 2 74715 58128
0 58130 5 1 1 58129
0 58131 7 1 2 106702 58130
0 58132 5 1 1 58131
0 58133 7 1 2 71512 58132
0 58134 5 1 1 58133
0 58135 7 1 2 73282 58134
0 58136 7 1 2 58124 58135
0 58137 5 1 1 58136
0 58138 7 1 2 85964 58137
0 58139 7 1 2 58118 58138
0 58140 5 1 1 58139
0 58141 7 1 2 58090 58140
0 58142 5 1 1 58141
0 58143 7 1 2 88278 58142
0 58144 5 1 1 58143
0 58145 7 1 2 84914 94227
0 58146 5 1 1 58145
0 58147 7 1 2 100063 58146
0 58148 5 1 1 58147
0 58149 7 1 2 96244 58148
0 58150 5 1 1 58149
0 58151 7 1 2 97620 97940
0 58152 5 1 1 58151
0 58153 7 1 2 85965 97430
0 58154 7 1 2 58152 58153
0 58155 5 1 1 58154
0 58156 7 1 2 83225 94653
0 58157 5 1 1 58156
0 58158 7 1 2 58155 58157
0 58159 7 1 2 58150 58158
0 58160 5 1 1 58159
0 58161 7 1 2 65231 58160
0 58162 5 1 1 58161
0 58163 7 1 2 99686 80492
0 58164 5 1 1 58163
0 58165 7 1 2 101335 58164
0 58166 5 1 1 58165
0 58167 7 1 2 65527 58166
0 58168 5 1 1 58167
0 58169 7 1 2 68894 91951
0 58170 7 1 2 100942 58169
0 58171 5 1 1 58170
0 58172 7 1 2 58168 58171
0 58173 5 1 1 58172
0 58174 7 1 2 77966 58173
0 58175 5 1 1 58174
0 58176 7 1 2 75069 103432
0 58177 5 1 1 58176
0 58178 7 1 2 85345 58177
0 58179 5 1 1 58178
0 58180 7 1 2 94606 97936
0 58181 5 1 1 58180
0 58182 7 1 2 58179 58181
0 58183 5 1 1 58182
0 58184 7 1 2 64917 58183
0 58185 5 1 1 58184
0 58186 7 1 2 68214 58185
0 58187 7 1 2 58175 58186
0 58188 7 1 2 58162 58187
0 58189 5 1 1 58188
0 58190 7 2 2 85966 76513
0 58191 7 1 2 93867 106888
0 58192 5 1 1 58191
0 58193 7 1 2 82804 106889
0 58194 5 1 1 58193
0 58195 7 1 2 79546 94057
0 58196 5 1 1 58195
0 58197 7 1 2 58194 58196
0 58198 5 1 1 58197
0 58199 7 1 2 65528 58198
0 58200 5 1 1 58199
0 58201 7 1 2 58192 58200
0 58202 5 1 1 58201
0 58203 7 1 2 73620 58202
0 58204 5 1 1 58203
0 58205 7 1 2 99732 92171
0 58206 5 1 1 58205
0 58207 7 1 2 85346 58206
0 58208 5 1 1 58207
0 58209 7 1 2 24119 58208
0 58210 5 1 1 58209
0 58211 7 1 2 68538 58210
0 58212 5 1 1 58211
0 58213 7 1 2 90723 75527
0 58214 7 1 2 78809 58213
0 58215 7 1 2 89175 58214
0 58216 5 1 1 58215
0 58217 7 1 2 73283 58216
0 58218 7 1 2 58212 58217
0 58219 7 1 2 58204 58218
0 58220 5 1 1 58219
0 58221 7 1 2 88634 58220
0 58222 7 1 2 58189 58221
0 58223 5 1 1 58222
0 58224 7 1 2 72826 58223
0 58225 7 1 2 58144 58224
0 58226 5 1 1 58225
0 58227 7 1 2 81801 92798
0 58228 5 1 1 58227
0 58229 7 1 2 96151 58228
0 58230 5 1 1 58229
0 58231 7 1 2 73621 58230
0 58232 5 1 1 58231
0 58233 7 1 2 89474 106238
0 58234 5 1 1 58233
0 58235 7 1 2 58232 58234
0 58236 5 1 1 58235
0 58237 7 1 2 85967 58236
0 58238 5 1 1 58237
0 58239 7 1 2 98676 106380
0 58240 5 1 1 58239
0 58241 7 1 2 5971 58240
0 58242 5 1 1 58241
0 58243 7 1 2 85718 58242
0 58244 5 1 1 58243
0 58245 7 1 2 58238 58244
0 58246 5 1 1 58245
0 58247 7 1 2 81160 58246
0 58248 5 1 1 58247
0 58249 7 1 2 104377 89859
0 58250 5 1 1 58249
0 58251 7 1 2 81802 81304
0 58252 5 1 1 58251
0 58253 7 1 2 58250 58252
0 58254 5 1 1 58253
0 58255 7 1 2 73622 58254
0 58256 5 1 1 58255
0 58257 7 1 2 85724 89378
0 58258 5 1 1 58257
0 58259 7 1 2 81161 58258
0 58260 5 1 1 58259
0 58261 7 1 2 58256 58260
0 58262 5 1 1 58261
0 58263 7 1 2 89328 58262
0 58264 5 1 1 58263
0 58265 7 1 2 67825 58264
0 58266 7 1 2 58248 58265
0 58267 5 1 1 58266
0 58268 7 1 2 100439 58267
0 58269 7 1 2 58226 58268
0 58270 5 1 1 58269
0 58271 7 1 2 100917 33893
0 58272 5 1 1 58271
0 58273 7 1 2 66402 58272
0 58274 5 1 1 58273
0 58275 7 1 2 75992 87877
0 58276 5 1 1 58275
0 58277 7 1 2 58274 58276
0 58278 5 2 1 58277
0 58279 7 1 2 88635 106890
0 58280 5 1 1 58279
0 58281 7 1 2 79972 89998
0 58282 5 1 1 58281
0 58283 7 1 2 58280 58282
0 58284 5 1 1 58283
0 58285 7 1 2 102252 58284
0 58286 5 1 1 58285
0 58287 7 1 2 101198 88636
0 58288 7 1 2 105757 58287
0 58289 5 1 1 58288
0 58290 7 1 2 58286 58289
0 58291 5 1 1 58290
0 58292 7 1 2 85347 58291
0 58293 5 1 1 58292
0 58294 7 1 2 83912 104919
0 58295 5 1 1 58294
0 58296 7 1 2 77009 102001
0 58297 7 1 2 101926 58296
0 58298 5 1 1 58297
0 58299 7 1 2 58295 58298
0 58300 5 1 1 58299
0 58301 7 1 2 65232 58300
0 58302 5 1 1 58301
0 58303 7 1 2 88324 106859
0 58304 5 1 1 58303
0 58305 7 1 2 58302 58304
0 58306 5 1 1 58305
0 58307 7 1 2 98633 58306
0 58308 5 1 1 58307
0 58309 7 1 2 58293 58308
0 58310 5 1 1 58309
0 58311 7 1 2 81933 58310
0 58312 5 1 1 58311
0 58313 7 1 2 88294 9758
0 58314 5 1 1 58313
0 58315 7 1 2 100616 58314
0 58316 5 1 1 58315
0 58317 7 1 2 85348 90569
0 58318 5 1 1 58317
0 58319 7 1 2 77106 85968
0 58320 7 1 2 89425 58319
0 58321 5 1 1 58320
0 58322 7 1 2 58318 58321
0 58323 7 1 2 58316 58322
0 58324 5 1 1 58323
0 58325 7 1 2 77547 58324
0 58326 5 1 1 58325
0 58327 7 1 2 73930 90409
0 58328 5 1 1 58327
0 58329 7 1 2 94275 92685
0 58330 5 1 1 58329
0 58331 7 1 2 58328 58330
0 58332 5 1 1 58331
0 58333 7 1 2 85349 80181
0 58334 7 1 2 58332 58333
0 58335 5 1 1 58334
0 58336 7 1 2 58326 58335
0 58337 5 1 1 58336
0 58338 7 1 2 101199 58337
0 58339 5 1 1 58338
0 58340 7 1 2 58312 58339
0 58341 7 1 2 58270 58340
0 58342 5 1 1 58341
0 58343 7 1 2 89007 58342
0 58344 5 1 1 58343
0 58345 7 1 2 58062 58344
0 58346 7 1 2 58028 58345
0 58347 7 1 2 57851 58346
0 58348 5 1 1 58347
0 58349 7 1 2 85556 58348
0 58350 5 1 1 58349
0 58351 7 1 2 77313 103657
0 58352 5 1 1 58351
0 58353 7 1 2 97167 58352
0 58354 5 1 1 58353
0 58355 7 1 2 91453 97086
0 58356 5 1 1 58355
0 58357 7 1 2 58354 58356
0 58358 5 1 1 58357
0 58359 7 1 2 78529 103098
0 58360 7 2 2 58358 58359
0 58361 7 1 2 63935 106892
0 58362 5 1 1 58361
0 58363 7 1 2 74579 96400
0 58364 7 1 2 104625 58363
0 58365 7 2 2 98899 58364
0 58366 7 1 2 106720 106894
0 58367 5 1 1 58366
0 58368 7 1 2 58362 58367
0 58369 5 1 1 58368
0 58370 7 1 2 71513 58369
0 58371 5 1 1 58370
0 58372 7 1 2 78331 2414
0 58373 5 1 1 58372
0 58374 7 1 2 75631 96773
0 58375 7 1 2 104244 58374
0 58376 7 1 2 106716 58375
0 58377 7 2 2 58373 58376
0 58378 7 1 2 63936 106896
0 58379 5 1 1 58378
0 58380 7 1 2 58371 58379
0 58381 5 1 1 58380
0 58382 7 1 2 74044 58381
0 58383 5 1 1 58382
0 58384 7 1 2 96774 106891
0 58385 5 1 1 58384
0 58386 7 1 2 97063 105758
0 58387 5 2 1 58386
0 58388 7 1 2 58385 106898
0 58389 5 1 1 58388
0 58390 7 1 2 99656 58389
0 58391 5 1 1 58390
0 58392 7 1 2 66403 100919
0 58393 5 1 1 58392
0 58394 7 1 2 90925 58393
0 58395 5 1 1 58394
0 58396 7 1 2 96775 58395
0 58397 5 1 1 58396
0 58398 7 1 2 106899 58397
0 58399 5 1 1 58398
0 58400 7 1 2 106666 58399
0 58401 5 1 1 58400
0 58402 7 1 2 58391 58401
0 58403 5 1 1 58402
0 58404 7 2 2 72196 58403
0 58405 7 1 2 100882 106900
0 58406 5 1 1 58405
0 58407 7 1 2 58383 58406
0 58408 5 1 1 58407
0 58409 7 1 2 73882 58408
0 58410 5 1 1 58409
0 58411 7 1 2 72827 79973
0 58412 5 1 1 58411
0 58413 7 1 2 100925 6627
0 58414 5 1 1 58413
0 58415 7 1 2 58412 58414
0 58416 5 1 1 58415
0 58417 7 1 2 67484 58416
0 58418 5 1 1 58417
0 58419 7 1 2 102382 58418
0 58420 5 1 1 58419
0 58421 7 1 2 98896 58420
0 58422 5 1 1 58421
0 58423 7 1 2 91300 105528
0 58424 7 1 2 97700 91295
0 58425 7 1 2 58423 58424
0 58426 5 1 1 58425
0 58427 7 1 2 58422 58426
0 58428 5 1 1 58427
0 58429 7 1 2 68539 100414
0 58430 7 1 2 58428 58429
0 58431 5 1 1 58430
0 58432 7 1 2 73800 101986
0 58433 7 1 2 81406 58432
0 58434 7 2 2 100346 90514
0 58435 7 1 2 86119 106445
0 58436 7 1 2 106902 58435
0 58437 7 1 2 58433 58436
0 58438 5 1 1 58437
0 58439 7 1 2 58431 58438
0 58440 5 1 1 58439
0 58441 7 1 2 88279 58440
0 58442 5 1 1 58441
0 58443 7 1 2 91365 106901
0 58444 5 1 1 58443
0 58445 7 1 2 58442 58444
0 58446 5 1 1 58445
0 58447 7 1 2 85350 58446
0 58448 5 1 1 58447
0 58449 7 1 2 79384 106893
0 58450 5 1 1 58449
0 58451 7 1 2 100957 106895
0 58452 5 1 1 58451
0 58453 7 1 2 58450 58452
0 58454 5 1 1 58453
0 58455 7 1 2 71514 58454
0 58456 5 1 1 58455
0 58457 7 1 2 79385 106897
0 58458 5 1 1 58457
0 58459 7 1 2 58456 58458
0 58460 5 1 1 58459
0 58461 7 1 2 89590 58460
0 58462 5 1 1 58461
0 58463 7 1 2 91100 83248
0 58464 5 1 1 58463
0 58465 7 1 2 90926 58464
0 58466 5 1 1 58465
0 58467 7 1 2 96776 58466
0 58468 5 1 1 58467
0 58469 7 1 2 101921 58468
0 58470 5 1 1 58469
0 58471 7 1 2 65233 58470
0 58472 5 1 1 58471
0 58473 7 1 2 100891 97168
0 58474 5 1 1 58473
0 58475 7 1 2 58472 58474
0 58476 5 1 1 58475
0 58477 7 1 2 87421 76399
0 58478 7 1 2 103099 58477
0 58479 7 1 2 98897 58478
0 58480 7 1 2 58476 58479
0 58481 5 1 1 58480
0 58482 7 1 2 58462 58481
0 58483 7 1 2 58448 58482
0 58484 7 1 2 58410 58483
0 58485 5 1 1 58484
0 58486 7 1 2 81934 58485
0 58487 5 1 1 58486
0 58488 7 1 2 93759 74269
0 58489 7 1 2 103962 58488
0 58490 5 1 1 58489
0 58491 7 1 2 74580 106729
0 58492 5 1 1 58491
0 58493 7 1 2 100853 74455
0 58494 7 1 2 106742 58493
0 58495 7 1 2 58492 58494
0 58496 5 1 1 58495
0 58497 7 1 2 58490 58496
0 58498 5 1 1 58497
0 58499 7 1 2 79646 58498
0 58500 5 1 1 58499
0 58501 7 2 2 101571 96304
0 58502 7 1 2 93109 74045
0 58503 7 1 2 106904 58502
0 58504 7 1 2 93837 58503
0 58505 5 1 1 58504
0 58506 7 1 2 58500 58505
0 58507 5 1 1 58506
0 58508 7 1 2 66902 58507
0 58509 5 1 1 58508
0 58510 7 1 2 91885 74046
0 58511 7 1 2 105766 58510
0 58512 7 1 2 106833 58511
0 58513 5 1 1 58512
0 58514 7 1 2 58509 58513
0 58515 5 1 1 58514
0 58516 7 1 2 80154 58515
0 58517 5 1 1 58516
0 58518 7 1 2 68540 78828
0 58519 7 1 2 101189 96231
0 58520 7 1 2 58518 58519
0 58521 7 1 2 103963 58520
0 58522 5 1 1 58521
0 58523 7 1 2 58517 58522
0 58524 5 1 1 58523
0 58525 7 1 2 72488 82070
0 58526 7 1 2 73883 58525
0 58527 7 1 2 58524 58526
0 58528 5 1 1 58527
0 58529 7 1 2 58487 58528
0 58530 7 1 2 58350 58529
0 58531 7 1 2 57492 58530
0 58532 7 1 2 57219 58531
0 58533 7 1 2 57128 58532
0 58534 5 1 1 58533
0 58535 7 1 2 77272 58534
0 58536 5 1 1 58535
0 58537 7 2 2 82531 92414
0 58538 7 1 2 102506 106906
0 58539 5 1 1 58538
0 58540 7 2 2 72272 100736
0 58541 7 1 2 104825 106908
0 58542 5 1 1 58541
0 58543 7 1 2 58539 58542
0 58544 5 1 1 58543
0 58545 7 1 2 64518 58544
0 58546 5 1 1 58545
0 58547 7 1 2 99977 106909
0 58548 5 1 1 58547
0 58549 7 1 2 58546 58548
0 58550 5 1 1 58549
0 58551 7 1 2 100357 58550
0 58552 5 1 1 58551
0 58553 7 1 2 99657 87054
0 58554 5 1 1 58553
0 58555 7 1 2 93242 104714
0 58556 7 1 2 99729 58555
0 58557 5 1 1 58556
0 58558 7 1 2 58554 58557
0 58559 5 1 1 58558
0 58560 7 1 2 64519 58559
0 58561 5 1 1 58560
0 58562 7 1 2 66091 22103
0 58563 5 2 1 58562
0 58564 7 2 2 69659 106910
0 58565 5 1 1 106912
0 58566 7 2 2 85557 103972
0 58567 7 1 2 106913 106914
0 58568 5 1 1 58567
0 58569 7 1 2 58561 58568
0 58570 5 1 1 58569
0 58571 7 1 2 81803 58570
0 58572 5 1 1 58571
0 58573 7 6 2 80382 79774
0 58574 5 4 1 106916
0 58575 7 1 2 76967 106917
0 58576 7 1 2 106915 58575
0 58577 5 1 1 58576
0 58578 7 1 2 71515 58577
0 58579 7 1 2 58572 58578
0 58580 5 1 1 58579
0 58581 7 4 2 68895 104321
0 58582 5 1 1 106926
0 58583 7 1 2 28559 58582
0 58584 5 9 1 58583
0 58585 7 5 2 71966 106930
0 58586 7 1 2 91139 106677
0 58587 5 1 1 58586
0 58588 7 1 2 91676 106667
0 58589 5 1 1 58588
0 58590 7 1 2 58587 58589
0 58591 5 1 1 58590
0 58592 7 1 2 84880 79417
0 58593 7 1 2 58591 58592
0 58594 5 1 1 58593
0 58595 7 1 2 99658 104767
0 58596 5 1 1 58595
0 58597 7 1 2 66404 58596
0 58598 7 1 2 58594 58597
0 58599 5 1 1 58598
0 58600 7 1 2 106939 58599
0 58601 7 1 2 58580 58600
0 58602 5 1 1 58601
0 58603 7 1 2 58552 58602
0 58604 5 1 1 58603
0 58605 7 1 2 72828 58604
0 58606 5 1 1 58605
0 58607 7 1 2 100629 94477
0 58608 5 1 1 58607
0 58609 7 1 2 80447 74319
0 58610 7 1 2 102079 58609
0 58611 5 1 1 58610
0 58612 7 1 2 58608 58611
0 58613 5 1 1 58612
0 58614 7 1 2 69311 58613
0 58615 5 1 1 58614
0 58616 7 1 2 95346 88034
0 58617 7 1 2 105521 58616
0 58618 5 1 1 58617
0 58619 7 1 2 58615 58618
0 58620 5 1 1 58619
0 58621 7 1 2 65529 58620
0 58622 5 1 1 58621
0 58623 7 1 2 93799 94077
0 58624 7 1 2 106124 58623
0 58625 5 1 1 58624
0 58626 7 1 2 58622 58625
0 58627 5 1 1 58626
0 58628 7 1 2 66405 58627
0 58629 5 1 1 58628
0 58630 7 1 2 93562 90271
0 58631 7 1 2 99540 58630
0 58632 7 1 2 100366 58631
0 58633 5 1 1 58632
0 58634 7 1 2 58629 58633
0 58635 5 1 1 58634
0 58636 7 1 2 73284 58635
0 58637 5 1 1 58636
0 58638 7 1 2 93831 87076
0 58639 5 13 1 58638
0 58640 7 11 2 68732 106944
0 58641 7 1 2 76251 106957
0 58642 5 1 1 58641
0 58643 7 1 2 71516 99812
0 58644 5 1 1 58643
0 58645 7 1 2 58642 58644
0 58646 5 1 1 58645
0 58647 7 1 2 68215 103363
0 58648 7 1 2 58646 58647
0 58649 5 1 1 58648
0 58650 7 1 2 58637 58649
0 58651 5 1 1 58650
0 58652 7 1 2 63815 58651
0 58653 5 1 1 58652
0 58654 7 1 2 79418 106958
0 58655 5 1 1 58654
0 58656 7 1 2 104364 58655
0 58657 5 1 1 58656
0 58658 7 1 2 66406 58657
0 58659 5 1 1 58658
0 58660 7 1 2 66092 76425
0 58661 7 1 2 86902 58660
0 58662 5 1 1 58661
0 58663 7 1 2 58659 58662
0 58664 5 1 1 58663
0 58665 7 1 2 71967 85558
0 58666 7 1 2 106927 58665
0 58667 7 1 2 58664 58666
0 58668 5 1 1 58667
0 58669 7 1 2 69660 58668
0 58670 7 1 2 58653 58669
0 58671 5 1 1 58670
0 58672 7 1 2 84915 81143
0 58673 5 1 1 58672
0 58674 7 1 2 97536 58673
0 58675 5 2 1 58674
0 58676 7 1 2 102587 106968
0 58677 5 1 1 58676
0 58678 7 1 2 99574 103976
0 58679 5 1 1 58678
0 58680 7 1 2 58677 58679
0 58681 5 1 1 58680
0 58682 7 1 2 106940 58681
0 58683 5 1 1 58682
0 58684 7 1 2 64520 58683
0 58685 5 1 1 58684
0 58686 7 1 2 101431 58685
0 58687 7 1 2 58671 58686
0 58688 5 1 1 58687
0 58689 7 1 2 58606 58688
0 58690 5 1 1 58689
0 58691 7 1 2 63987 58690
0 58692 5 1 1 58691
0 58693 7 12 2 69068 72273
0 58694 5 2 1 106970
0 58695 7 1 2 80871 102015
0 58696 5 1 1 58695
0 58697 7 1 2 101750 104862
0 58698 5 1 1 58697
0 58699 7 1 2 58696 58698
0 58700 5 1 1 58699
0 58701 7 1 2 71873 58700
0 58702 5 1 1 58701
0 58703 7 1 2 71968 77273
0 58704 7 1 2 102436 58703
0 58705 7 1 2 88468 58704
0 58706 5 1 1 58705
0 58707 7 1 2 58702 58706
0 58708 5 1 1 58707
0 58709 7 1 2 63816 58708
0 58710 5 1 1 58709
0 58711 7 3 2 97725 106928
0 58712 7 1 2 82672 94534
0 58713 5 1 1 58712
0 58714 7 1 2 99797 86531
0 58715 5 1 1 58714
0 58716 7 1 2 58713 58715
0 58717 5 1 1 58716
0 58718 7 1 2 106984 58717
0 58719 5 1 1 58718
0 58720 7 1 2 58710 58719
0 58721 5 1 1 58720
0 58722 7 1 2 70567 58721
0 58723 5 1 1 58722
0 58724 7 1 2 74909 97726
0 58725 7 1 2 101699 58724
0 58726 7 1 2 106931 58725
0 58727 5 1 1 58726
0 58728 7 1 2 58723 58727
0 58729 5 1 1 58728
0 58730 7 1 2 64918 58729
0 58731 5 1 1 58730
0 58732 7 1 2 86409 104763
0 58733 7 2 2 106932 58732
0 58734 7 1 2 65530 106987
0 58735 5 1 1 58734
0 58736 7 1 2 58731 58735
0 58737 5 1 1 58736
0 58738 7 1 2 72829 58737
0 58739 5 1 1 58738
0 58740 7 1 2 91334 96077
0 58741 7 2 2 106933 58740
0 58742 7 1 2 83300 106989
0 58743 5 1 1 58742
0 58744 7 1 2 58739 58743
0 58745 5 1 1 58744
0 58746 7 1 2 66407 58745
0 58747 5 1 1 58746
0 58748 7 4 2 68216 106934
0 58749 7 1 2 83733 85974
0 58750 7 2 2 106991 58749
0 58751 7 1 2 83301 106995
0 58752 5 1 1 58751
0 58753 7 1 2 58747 58752
0 58754 5 1 1 58753
0 58755 7 1 2 64212 58754
0 58756 5 1 1 58755
0 58757 7 1 2 99542 100734
0 58758 5 8 1 58757
0 58759 7 2 2 82252 106997
0 58760 7 1 2 100660 92526
0 58761 7 1 2 107005 58760
0 58762 5 1 1 58761
0 58763 7 1 2 58756 58762
0 58764 5 1 1 58763
0 58765 7 1 2 65854 58764
0 58766 5 1 1 58765
0 58767 7 2 2 80872 101784
0 58768 7 1 2 85846 85421
0 58769 7 1 2 94687 58768
0 58770 7 1 2 94906 58769
0 58771 7 1 2 107007 58770
0 58772 5 1 1 58771
0 58773 7 1 2 58766 58772
0 58774 5 1 1 58773
0 58775 7 1 2 106971 58774
0 58776 5 1 1 58775
0 58777 7 1 2 58692 58776
0 58778 5 1 1 58777
0 58779 7 1 2 65695 58778
0 58780 5 1 1 58779
0 58781 7 2 2 82673 102016
0 58782 5 1 1 107009
0 58783 7 1 2 97727 98877
0 58784 7 1 2 102437 58783
0 58785 5 1 1 58784
0 58786 7 1 2 58782 58785
0 58787 5 1 1 58786
0 58788 7 1 2 63817 58787
0 58789 5 1 1 58788
0 58790 7 1 2 70279 98878
0 58791 7 1 2 106985 58790
0 58792 5 1 1 58791
0 58793 7 1 2 58789 58792
0 58794 5 1 1 58793
0 58795 7 1 2 73801 58794
0 58796 5 1 1 58795
0 58797 7 1 2 84578 107010
0 58798 5 1 1 58797
0 58799 7 1 2 58796 58798
0 58800 5 1 1 58799
0 58801 7 1 2 64521 58800
0 58802 5 1 1 58801
0 58803 7 1 2 87108 93243
0 58804 7 1 2 107008 58803
0 58805 5 1 1 58804
0 58806 7 1 2 58802 58805
0 58807 5 1 1 58806
0 58808 7 1 2 70568 58807
0 58809 5 1 1 58808
0 58810 7 1 2 70280 100973
0 58811 7 1 2 95304 58810
0 58812 7 1 2 106935 58811
0 58813 5 1 1 58812
0 58814 7 1 2 58809 58813
0 58815 5 1 1 58814
0 58816 7 1 2 64919 58815
0 58817 5 1 1 58816
0 58818 7 1 2 93144 106988
0 58819 5 1 1 58818
0 58820 7 1 2 58817 58819
0 58821 5 1 1 58820
0 58822 7 1 2 72830 58821
0 58823 5 1 1 58822
0 58824 7 2 2 65855 83302
0 58825 7 1 2 106990 107011
0 58826 5 1 1 58825
0 58827 7 1 2 58823 58826
0 58828 5 1 1 58827
0 58829 7 1 2 66408 58828
0 58830 5 1 1 58829
0 58831 7 1 2 106996 107012
0 58832 5 1 1 58831
0 58833 7 1 2 58830 58832
0 58834 5 1 1 58833
0 58835 7 2 2 72274 99348
0 58836 7 1 2 64213 107013
0 58837 7 1 2 58834 58836
0 58838 5 1 1 58837
0 58839 7 1 2 67143 58838
0 58840 7 1 2 58780 58839
0 58841 5 1 1 58840
0 58842 7 1 2 103178 105060
0 58843 5 1 1 58842
0 58844 7 1 2 81084 58843
0 58845 5 1 1 58844
0 58846 7 1 2 97888 93026
0 58847 5 1 1 58846
0 58848 7 1 2 58845 58847
0 58849 5 1 1 58848
0 58850 7 3 2 93320 106936
0 58851 7 1 2 58849 107015
0 58852 5 1 1 58851
0 58853 7 1 2 70281 99974
0 58854 7 1 2 86615 58853
0 58855 7 1 2 89643 102181
0 58856 7 1 2 58854 58855
0 58857 5 1 1 58856
0 58858 7 1 2 58852 58857
0 58859 5 1 1 58858
0 58860 7 1 2 66799 58859
0 58861 5 1 1 58860
0 58862 7 3 2 80428 106937
0 58863 7 2 2 71969 107018
0 58864 7 1 2 70920 9426
0 58865 5 1 1 58864
0 58866 7 1 2 74985 98527
0 58867 5 1 1 58866
0 58868 7 1 2 58865 58867
0 58869 5 1 1 58868
0 58870 7 1 2 107021 58869
0 58871 5 1 1 58870
0 58872 7 1 2 117 3177
0 58873 5 1 1 58872
0 58874 7 1 2 100303 90651
0 58875 7 1 2 89783 58874
0 58876 7 1 2 58873 58875
0 58877 5 1 1 58876
0 58878 7 1 2 72831 58877
0 58879 7 1 2 58871 58878
0 58880 5 1 1 58879
0 58881 7 1 2 64522 105314
0 58882 5 1 1 58881
0 58883 7 1 2 93062 84399
0 58884 5 1 1 58883
0 58885 7 1 2 58882 58884
0 58886 5 1 1 58885
0 58887 7 1 2 58886 107022
0 58888 5 1 1 58887
0 58889 7 1 2 91351 101282
0 58890 7 1 2 102364 96580
0 58891 7 1 2 58889 58890
0 58892 5 1 1 58891
0 58893 7 1 2 67826 58892
0 58894 7 1 2 58888 58893
0 58895 5 1 1 58894
0 58896 7 1 2 65531 58895
0 58897 7 1 2 58880 58896
0 58898 5 1 1 58897
0 58899 7 1 2 58861 58898
0 58900 5 1 1 58899
0 58901 7 1 2 69312 58900
0 58902 5 1 1 58901
0 58903 7 1 2 85070 42789
0 58904 5 1 1 58903
0 58905 7 1 2 69661 58904
0 58906 5 1 1 58905
0 58907 7 1 2 85096 58906
0 58908 5 2 1 58907
0 58909 7 1 2 85472 88409
0 58910 7 1 2 106941 58909
0 58911 7 1 2 107023 58910
0 58912 5 1 1 58911
0 58913 7 1 2 58902 58912
0 58914 5 1 1 58913
0 58915 7 1 2 99342 58914
0 58916 5 1 1 58915
0 58917 7 1 2 80429 102177
0 58918 5 1 1 58917
0 58919 7 1 2 82999 102182
0 58920 7 1 2 103370 58919
0 58921 5 1 1 58920
0 58922 7 1 2 58918 58921
0 58923 5 1 1 58922
0 58924 7 1 2 63818 58923
0 58925 5 1 1 58924
0 58926 7 2 2 80430 104322
0 58927 7 2 2 85108 107025
0 58928 7 1 2 106144 107027
0 58929 5 1 1 58928
0 58930 7 1 2 58925 58929
0 58931 5 1 1 58930
0 58932 7 1 2 64523 58931
0 58933 5 1 1 58932
0 58934 7 2 2 80431 106992
0 58935 7 1 2 93063 93571
0 58936 7 1 2 107029 58935
0 58937 5 1 1 58936
0 58938 7 1 2 58933 58937
0 58939 5 1 1 58938
0 58940 7 1 2 71517 58939
0 58941 5 1 1 58940
0 58942 7 1 2 94068 105425
0 58943 7 1 2 107019 58942
0 58944 5 1 1 58943
0 58945 7 1 2 58941 58944
0 58946 5 1 1 58945
0 58947 7 1 2 65532 58946
0 58948 5 1 1 58947
0 58949 7 1 2 93030 44612
0 58950 5 1 1 58949
0 58951 7 1 2 98879 58950
0 58952 7 1 2 107016 58951
0 58953 5 1 1 58952
0 58954 7 1 2 58948 58953
0 58955 5 1 1 58954
0 58956 7 1 2 71213 58955
0 58957 5 1 1 58956
0 58958 7 3 2 104465 106993
0 58959 7 1 2 65856 107031
0 58960 5 1 1 58959
0 58961 7 1 2 93645 93071
0 58962 7 1 2 100968 58961
0 58963 7 1 2 96639 58962
0 58964 5 1 1 58963
0 58965 7 1 2 58960 58964
0 58966 5 1 1 58965
0 58967 7 1 2 92940 58966
0 58968 5 1 1 58967
0 58969 7 1 2 58957 58968
0 58970 5 1 1 58969
0 58971 7 1 2 69313 58970
0 58972 5 1 1 58971
0 58973 7 5 2 70282 83008
0 58974 5 1 1 107034
0 58975 7 1 2 73285 107035
0 58976 5 1 1 58975
0 58977 7 1 2 103123 58976
0 58978 5 1 1 58977
0 58979 7 1 2 103199 58978
0 58980 5 1 1 58979
0 58981 7 1 2 94590 93741
0 58982 7 1 2 99245 58981
0 58983 7 1 2 88410 58982
0 58984 5 1 1 58983
0 58985 7 1 2 58980 58984
0 58986 5 1 1 58985
0 58987 7 1 2 63819 58986
0 58988 5 1 1 58987
0 58989 7 1 2 86027 103270
0 58990 7 1 2 107028 58989
0 58991 5 1 1 58990
0 58992 7 1 2 58988 58991
0 58993 5 1 1 58992
0 58994 7 1 2 71214 58993
0 58995 5 1 1 58994
0 58996 7 1 2 98348 107032
0 58997 5 1 1 58996
0 58998 7 1 2 58995 58997
0 58999 5 1 1 58998
0 59000 7 1 2 64524 58999
0 59001 5 1 1 59000
0 59002 7 1 2 100220 101633
0 59003 5 1 1 59002
0 59004 7 1 2 80432 89133
0 59005 7 1 2 91790 59004
0 59006 5 1 1 59005
0 59007 7 1 2 59003 59006
0 59008 5 1 1 59007
0 59009 7 1 2 63820 59008
0 59010 5 1 1 59009
0 59011 7 1 2 104887 107026
0 59012 5 1 1 59011
0 59013 7 1 2 59010 59012
0 59014 5 1 1 59013
0 59015 7 1 2 103271 59014
0 59016 5 1 1 59015
0 59017 7 1 2 101011 84494
0 59018 7 1 2 107030 59017
0 59019 5 1 1 59018
0 59020 7 1 2 59016 59019
0 59021 5 1 1 59020
0 59022 7 1 2 65533 59021
0 59023 5 1 1 59022
0 59024 7 1 2 101534 3020
0 59025 5 1 1 59024
0 59026 7 1 2 69662 59025
0 59027 7 1 2 107017 59026
0 59028 5 1 1 59027
0 59029 7 1 2 99612 103219
0 59030 7 1 2 100661 59029
0 59031 5 1 1 59030
0 59032 7 1 2 59028 59031
0 59033 5 1 1 59032
0 59034 7 1 2 66800 59033
0 59035 5 1 1 59034
0 59036 7 1 2 59023 59035
0 59037 7 1 2 59001 59036
0 59038 5 1 1 59037
0 59039 7 1 2 72832 59038
0 59040 5 1 1 59039
0 59041 7 2 2 86028 107020
0 59042 7 3 2 89918 104383
0 59043 5 1 1 107041
0 59044 7 1 2 101535 59043
0 59045 5 1 1 59044
0 59046 7 1 2 64525 59045
0 59047 5 1 1 59046
0 59048 7 1 2 78134 84400
0 59049 5 1 1 59048
0 59050 7 1 2 59047 59049
0 59051 5 1 1 59050
0 59052 7 1 2 91707 59051
0 59053 7 1 2 107039 59052
0 59054 5 1 1 59053
0 59055 7 1 2 59040 59054
0 59056 5 1 1 59055
0 59057 7 1 2 70921 59056
0 59058 5 1 1 59057
0 59059 7 1 2 63988 59058
0 59060 7 1 2 58972 59059
0 59061 5 1 1 59060
0 59062 7 1 2 100630 104434
0 59063 5 1 1 59062
0 59064 7 1 2 100221 97860
0 59065 7 1 2 103121 59064
0 59066 5 1 1 59065
0 59067 7 1 2 59063 59066
0 59068 5 1 1 59067
0 59069 7 1 2 63821 59068
0 59070 5 1 1 59069
0 59071 7 1 2 82779 104435
0 59072 7 1 2 106929 59071
0 59073 5 1 1 59072
0 59074 7 1 2 59070 59073
0 59075 5 1 1 59074
0 59076 7 1 2 87887 59075
0 59077 5 1 1 59076
0 59078 7 1 2 87811 96119
0 59079 7 1 2 107040 59078
0 59080 5 1 1 59079
0 59081 7 1 2 59077 59080
0 59082 5 1 1 59081
0 59083 7 1 2 66409 59082
0 59084 5 1 1 59083
0 59085 7 1 2 96169 107033
0 59086 5 1 1 59085
0 59087 7 1 2 59084 59086
0 59088 5 1 1 59087
0 59089 7 1 2 64214 59088
0 59090 5 1 1 59089
0 59091 7 1 2 84794 82015
0 59092 7 1 2 100404 77910
0 59093 7 1 2 59091 59092
0 59094 7 1 2 93498 95956
0 59095 7 1 2 59093 59094
0 59096 5 1 1 59095
0 59097 7 1 2 69069 59096
0 59098 7 1 2 59090 59097
0 59099 5 1 1 59098
0 59100 7 1 2 70733 59099
0 59101 7 1 2 59061 59100
0 59102 5 1 1 59101
0 59103 7 1 2 58916 59102
0 59104 5 1 1 59103
0 59105 7 1 2 67232 59104
0 59106 5 1 1 59105
0 59107 7 1 2 100766 81144
0 59108 5 2 1 59107
0 59109 7 1 2 82510 107044
0 59110 5 1 1 59109
0 59111 7 1 2 93500 59110
0 59112 5 1 1 59111
0 59113 7 1 2 11334 59112
0 59114 5 1 1 59113
0 59115 7 1 2 72833 59114
0 59116 5 1 1 59115
0 59117 7 1 2 105859 59116
0 59118 5 1 1 59117
0 59119 7 1 2 66801 59118
0 59120 5 1 1 59119
0 59121 7 1 2 73802 83507
0 59122 7 1 2 77997 59121
0 59123 7 1 2 99149 59122
0 59124 5 1 1 59123
0 59125 7 1 2 59120 59124
0 59126 5 1 1 59125
0 59127 7 1 2 65534 59126
0 59128 5 1 1 59127
0 59129 7 1 2 84954 98578
0 59130 5 1 1 59129
0 59131 7 1 2 38846 59130
0 59132 5 1 1 59131
0 59133 7 1 2 72834 105894
0 59134 7 1 2 59132 59133
0 59135 5 1 1 59134
0 59136 7 1 2 59128 59135
0 59137 5 1 1 59136
0 59138 7 1 2 71518 59137
0 59139 5 1 1 59138
0 59140 7 1 2 96090 10153
0 59141 5 1 1 59140
0 59142 7 1 2 103272 59141
0 59143 7 1 2 106959 59142
0 59144 5 1 1 59143
0 59145 7 1 2 73286 59144
0 59146 7 1 2 59139 59145
0 59147 5 1 1 59146
0 59148 7 1 2 96085 101490
0 59149 5 1 1 59148
0 59150 7 1 2 105860 59149
0 59151 5 1 1 59150
0 59152 7 1 2 95495 59151
0 59153 5 1 1 59152
0 59154 7 1 2 68217 59153
0 59155 5 1 1 59154
0 59156 7 4 2 72275 89519
0 59157 7 1 2 100662 107046
0 59158 7 1 2 59155 59157
0 59159 7 1 2 59147 59158
0 59160 5 1 1 59159
0 59161 7 1 2 72197 59160
0 59162 7 1 2 59106 59161
0 59163 5 1 1 59162
0 59164 7 1 2 67485 59163
0 59165 7 1 2 58841 59164
0 59166 5 1 1 59165
0 59167 7 3 2 72276 99343
0 59168 5 1 1 107050
0 59169 7 1 2 102386 97837
0 59170 5 1 1 59169
0 59171 7 1 2 66802 84301
0 59172 7 1 2 102582 59171
0 59173 5 1 1 59172
0 59174 7 1 2 59170 59173
0 59175 5 1 1 59174
0 59176 7 1 2 81085 59175
0 59177 5 1 1 59176
0 59178 7 1 2 66803 102020
0 59179 5 1 1 59178
0 59180 7 1 2 59177 59179
0 59181 5 1 1 59180
0 59182 7 1 2 65535 59181
0 59183 5 1 1 59182
0 59184 7 1 2 82939 95477
0 59185 7 1 2 105917 59184
0 59186 5 1 1 59185
0 59187 7 1 2 59183 59186
0 59188 5 1 1 59187
0 59189 7 1 2 107051 59188
0 59190 5 1 1 59189
0 59191 7 5 2 65696 67233
0 59192 5 2 1 107053
0 59193 7 3 2 70734 72277
0 59194 5 1 1 107060
0 59195 7 2 2 107058 59194
0 59196 5 4 1 107063
0 59197 7 1 2 98546 107065
0 59198 5 2 1 59197
0 59199 7 2 2 90458 107054
0 59200 5 1 1 107071
0 59201 7 1 2 77274 107072
0 59202 5 1 1 59201
0 59203 7 2 2 72278 91603
0 59204 5 1 1 107073
0 59205 7 2 2 64526 107074
0 59206 5 1 1 107075
0 59207 7 1 2 59202 59206
0 59208 5 1 1 59207
0 59209 7 1 2 67827 59208
0 59210 5 1 1 59209
0 59211 7 1 2 107069 59210
0 59212 5 1 1 59211
0 59213 7 1 2 75944 59212
0 59214 5 1 1 59213
0 59215 7 1 2 85046 107076
0 59216 5 2 1 59215
0 59217 7 1 2 59214 107077
0 59218 5 1 1 59217
0 59219 7 1 2 69314 59218
0 59220 5 1 1 59219
0 59221 7 5 2 64215 70735
0 59222 5 1 1 107079
0 59223 7 2 2 72279 107024
0 59224 7 1 2 107080 107084
0 59225 5 1 1 59224
0 59226 7 1 2 59220 59225
0 59227 5 1 1 59226
0 59228 7 1 2 66804 59227
0 59229 5 1 1 59228
0 59230 7 2 2 73803 104764
0 59231 7 1 2 107061 107086
0 59232 5 1 1 59231
0 59233 7 3 2 83140 107055
0 59234 7 1 2 82675 107088
0 59235 5 1 1 59234
0 59236 7 1 2 59232 59235
0 59237 5 1 1 59236
0 59238 7 1 2 66410 93354
0 59239 7 1 2 59237 59238
0 59240 5 1 1 59239
0 59241 7 1 2 59229 59240
0 59242 5 1 1 59241
0 59243 7 1 2 65536 59242
0 59244 5 1 1 59243
0 59245 7 2 2 103341 107087
0 59246 7 2 2 106376 107091
0 59247 7 1 2 69315 107093
0 59248 5 1 1 59247
0 59249 7 1 2 84107 94478
0 59250 5 2 1 59249
0 59251 7 1 2 80036 101405
0 59252 5 1 1 59251
0 59253 7 1 2 107095 59252
0 59254 5 1 1 59253
0 59255 7 1 2 80212 107089
0 59256 7 1 2 59254 59255
0 59257 5 1 1 59256
0 59258 7 1 2 65857 59257
0 59259 7 1 2 59248 59258
0 59260 7 1 2 59244 59259
0 59261 5 1 1 59260
0 59262 7 1 2 59200 59204
0 59263 5 1 1 59262
0 59264 7 1 2 81539 59263
0 59265 5 1 1 59264
0 59266 7 1 2 107070 59265
0 59267 5 1 1 59266
0 59268 7 1 2 75945 59267
0 59269 5 1 1 59268
0 59270 7 1 2 107078 59269
0 59271 5 1 1 59270
0 59272 7 1 2 64216 59271
0 59273 5 1 1 59272
0 59274 7 3 2 69316 65697
0 59275 7 1 2 107085 107097
0 59276 5 1 1 59275
0 59277 7 1 2 59273 59276
0 59278 5 1 1 59277
0 59279 7 1 2 66805 59278
0 59280 5 1 1 59279
0 59281 7 2 2 66411 107081
0 59282 7 1 2 107092 107100
0 59283 5 1 1 59282
0 59284 7 1 2 59280 59283
0 59285 5 1 1 59284
0 59286 7 1 2 65537 59285
0 59287 5 1 1 59286
0 59288 7 1 2 64217 107094
0 59289 5 1 1 59288
0 59290 7 1 2 70922 59289
0 59291 7 1 2 59287 59290
0 59292 5 1 1 59291
0 59293 7 1 2 63989 59292
0 59294 7 1 2 59261 59293
0 59295 5 1 1 59294
0 59296 7 1 2 59190 59295
0 59297 5 1 1 59296
0 59298 7 1 2 106942 59297
0 59299 5 1 1 59298
0 59300 7 8 2 71874 80873
0 59301 7 2 2 93622 77529
0 59302 7 1 2 107102 107110
0 59303 5 1 1 59302
0 59304 7 1 2 96444 84365
0 59305 5 1 1 59304
0 59306 7 1 2 59303 59305
0 59307 5 1 1 59306
0 59308 7 2 2 63990 107066
0 59309 5 1 1 107112
0 59310 7 1 2 59168 59309
0 59311 5 2 1 59310
0 59312 7 2 2 76921 96058
0 59313 7 1 2 102183 107116
0 59314 7 1 2 107114 59313
0 59315 7 1 2 59307 59314
0 59316 5 1 1 59315
0 59317 7 1 2 59299 59316
0 59318 5 1 1 59317
0 59319 7 1 2 67144 59318
0 59320 5 1 1 59319
0 59321 7 3 2 72280 85034
0 59322 7 1 2 95725 104592
0 59323 7 2 2 107118 59322
0 59324 7 1 2 93651 107121
0 59325 5 1 1 59324
0 59326 7 1 2 71215 100960
0 59327 7 1 2 77036 59326
0 59328 7 8 2 63991 67234
0 59329 5 1 1 107123
0 59330 7 1 2 106982 59329
0 59331 5 1 1 59330
0 59332 7 1 2 99225 59331
0 59333 7 1 2 59327 59332
0 59334 5 1 1 59333
0 59335 7 1 2 59325 59334
0 59336 5 1 1 59335
0 59337 7 1 2 70736 59336
0 59338 5 1 1 59337
0 59339 7 3 2 65698 92451
0 59340 7 1 2 107122 107131
0 59341 5 1 1 59340
0 59342 7 1 2 59338 59341
0 59343 5 1 1 59342
0 59344 7 1 2 76514 59343
0 59345 5 1 1 59344
0 59346 7 2 2 99359 84302
0 59347 7 1 2 87934 103044
0 59348 7 1 2 107134 59347
0 59349 5 1 1 59348
0 59350 7 1 2 59345 59349
0 59351 5 1 1 59350
0 59352 7 1 2 69663 59351
0 59353 5 1 1 59352
0 59354 7 5 2 67235 67828
0 59355 7 1 2 100809 96703
0 59356 7 1 2 107136 59355
0 59357 7 2 2 73287 77779
0 59358 7 1 2 97869 107141
0 59359 7 1 2 59356 59358
0 59360 5 1 1 59359
0 59361 7 1 2 71970 96551
0 59362 7 1 2 73810 59361
0 59363 7 1 2 97712 107119
0 59364 7 1 2 59362 59363
0 59365 5 1 1 59364
0 59366 7 1 2 59360 59365
0 59367 5 1 1 59366
0 59368 7 1 2 76515 59367
0 59369 5 1 1 59368
0 59370 7 1 2 96401 102645
0 59371 7 1 2 91398 59370
0 59372 7 1 2 88035 84303
0 59373 7 1 2 82059 59372
0 59374 7 1 2 59371 59373
0 59375 5 1 1 59374
0 59376 7 1 2 63992 59375
0 59377 7 1 2 59369 59376
0 59378 5 1 1 59377
0 59379 7 1 2 97870 78397
0 59380 7 1 2 107067 59379
0 59381 5 1 1 59380
0 59382 7 2 2 70737 67236
0 59383 5 1 1 107143
0 59384 7 1 2 87888 107144
0 59385 7 1 2 93207 59384
0 59386 5 1 1 59385
0 59387 7 1 2 59381 59386
0 59388 5 1 1 59387
0 59389 7 1 2 91311 107142
0 59390 7 1 2 59388 59389
0 59391 5 1 1 59390
0 59392 7 1 2 96413 104615
0 59393 7 2 2 85035 92443
0 59394 7 1 2 92520 107145
0 59395 7 1 2 59392 59394
0 59396 5 1 1 59395
0 59397 7 1 2 69070 59396
0 59398 7 1 2 59391 59397
0 59399 5 1 1 59398
0 59400 7 1 2 69317 59399
0 59401 7 1 2 59378 59400
0 59402 5 1 1 59401
0 59403 7 1 2 59353 59402
0 59404 5 1 1 59403
0 59405 7 1 2 63822 59404
0 59406 5 1 1 59405
0 59407 7 1 2 74441 88933
0 59408 5 1 1 59407
0 59409 7 1 2 99354 82511
0 59410 5 1 1 59409
0 59411 7 1 2 59408 59410
0 59412 7 1 2 92727 59411
0 59413 5 1 1 59412
0 59414 7 1 2 99344 98349
0 59415 7 1 2 95324 59414
0 59416 5 1 1 59415
0 59417 7 1 2 59413 59416
0 59418 5 1 1 59417
0 59419 7 1 2 102646 106986
0 59420 7 1 2 59418 59419
0 59421 5 1 1 59420
0 59422 7 1 2 59406 59421
0 59423 5 1 1 59422
0 59424 7 1 2 106945 59423
0 59425 5 1 1 59424
0 59426 7 2 2 78135 90817
0 59427 5 1 1 107147
0 59428 7 1 2 104914 59427
0 59429 5 1 1 59428
0 59430 7 1 2 74910 59429
0 59431 5 1 1 59430
0 59432 7 1 2 64527 104647
0 59433 5 1 1 59432
0 59434 7 1 2 104915 59433
0 59435 5 1 1 59434
0 59436 7 1 2 96563 59435
0 59437 5 1 1 59436
0 59438 7 1 2 59431 59437
0 59439 5 1 1 59438
0 59440 7 1 2 65858 59439
0 59441 5 1 1 59440
0 59442 7 1 2 72835 99975
0 59443 7 1 2 96564 59442
0 59444 7 1 2 105307 59443
0 59445 5 1 1 59444
0 59446 7 1 2 59441 59445
0 59447 5 1 1 59446
0 59448 7 1 2 68218 96844
0 59449 7 1 2 107056 59448
0 59450 7 1 2 106943 59449
0 59451 7 1 2 59447 59450
0 59452 5 1 1 59451
0 59453 7 1 2 59425 59452
0 59454 5 1 1 59453
0 59455 7 1 2 68733 59454
0 59456 5 1 1 59455
0 59457 7 1 2 100631 88927
0 59458 7 1 2 99128 59457
0 59459 5 1 1 59458
0 59460 7 1 2 100810 91712
0 59461 7 1 2 96704 59460
0 59462 7 2 2 87812 74224
0 59463 7 1 2 74161 107149
0 59464 7 1 2 59461 59463
0 59465 5 1 1 59464
0 59466 7 1 2 59459 59465
0 59467 5 1 1 59466
0 59468 7 1 2 69664 59467
0 59469 5 1 1 59468
0 59470 7 1 2 83412 90272
0 59471 7 1 2 73833 59470
0 59472 7 1 2 91549 59471
0 59473 7 1 2 92294 59472
0 59474 5 1 1 59473
0 59475 7 1 2 59469 59474
0 59476 5 1 1 59475
0 59477 7 1 2 64218 59476
0 59478 5 1 1 59477
0 59479 7 2 2 99093 73827
0 59480 5 1 1 107151
0 59481 7 3 2 77911 89871
0 59482 7 1 2 63993 107150
0 59483 7 1 2 107153 59482
0 59484 7 1 2 107152 59483
0 59485 5 1 1 59484
0 59486 7 1 2 59478 59485
0 59487 5 1 1 59486
0 59488 7 1 2 67237 59487
0 59489 5 1 1 59488
0 59490 7 1 2 76922 100961
0 59491 7 1 2 101432 89520
0 59492 7 1 2 59490 59491
0 59493 7 2 2 85847 74225
0 59494 7 1 2 78007 107156
0 59495 7 1 2 59492 59494
0 59496 5 1 1 59495
0 59497 7 1 2 59489 59496
0 59498 5 1 1 59497
0 59499 7 1 2 70283 59498
0 59500 5 1 1 59499
0 59501 7 1 2 84366 107062
0 59502 5 1 1 59501
0 59503 7 1 2 76516 103932
0 59504 7 1 2 92592 59503
0 59505 5 1 1 59504
0 59506 7 1 2 59502 59505
0 59507 5 1 1 59506
0 59508 7 1 2 63994 59507
0 59509 5 1 1 59508
0 59510 7 2 2 101283 106972
0 59511 7 1 2 107098 107158
0 59512 5 1 1 59511
0 59513 7 1 2 59509 59512
0 59514 5 1 1 59513
0 59515 7 1 2 84943 102971
0 59516 7 1 2 96640 59515
0 59517 7 1 2 59514 59516
0 59518 5 1 1 59517
0 59519 7 1 2 59500 59518
0 59520 5 1 1 59519
0 59521 7 1 2 63823 59520
0 59522 5 1 1 59521
0 59523 7 1 2 104593 94000
0 59524 7 1 2 107090 59523
0 59525 7 1 2 104323 59524
0 59526 7 1 2 107148 59525
0 59527 5 1 1 59526
0 59528 7 1 2 59522 59527
0 59529 5 1 1 59528
0 59530 7 1 2 84881 59529
0 59531 5 1 1 59530
0 59532 7 1 2 82479 107068
0 59533 5 1 1 59532
0 59534 7 1 2 70738 103942
0 59535 5 1 1 59534
0 59536 7 1 2 59533 59535
0 59537 5 1 1 59536
0 59538 7 1 2 69071 59537
0 59539 5 1 1 59538
0 59540 7 4 2 93473 106785
0 59541 5 1 1 107160
0 59542 7 1 2 67238 107161
0 59543 5 1 1 59542
0 59544 7 1 2 59539 59543
0 59545 5 1 1 59544
0 59546 7 1 2 93663 59545
0 59547 5 1 1 59546
0 59548 7 2 2 69072 100581
0 59549 7 1 2 70739 107164
0 59550 7 1 2 103452 59549
0 59551 5 1 1 59550
0 59552 7 1 2 59547 59551
0 59553 5 1 1 59552
0 59554 7 1 2 76109 97305
0 59555 7 1 2 98066 59554
0 59556 7 1 2 59553 59555
0 59557 5 1 1 59556
0 59558 7 1 2 59531 59557
0 59559 7 1 2 59456 59558
0 59560 7 1 2 59320 59559
0 59561 5 1 1 59560
0 59562 7 1 2 72489 59561
0 59563 5 1 1 59562
0 59564 7 1 2 87193 90818
0 59565 5 1 1 59564
0 59566 7 1 2 83979 101406
0 59567 5 1 1 59566
0 59568 7 1 2 59565 59567
0 59569 5 1 1 59568
0 59570 7 1 2 69665 59569
0 59571 5 1 1 59570
0 59572 7 2 2 76517 95322
0 59573 5 1 1 107166
0 59574 7 1 2 77530 107167
0 59575 5 1 1 59574
0 59576 7 1 2 59571 59575
0 59577 5 1 1 59576
0 59578 7 1 2 70284 59577
0 59579 5 1 1 59578
0 59580 7 1 2 92873 106918
0 59581 5 1 1 59580
0 59582 7 1 2 59579 59581
0 59583 5 1 1 59582
0 59584 7 1 2 99360 59583
0 59585 5 1 1 59584
0 59586 7 1 2 106922 58974
0 59587 5 2 1 59586
0 59588 7 1 2 99349 90831
0 59589 7 1 2 107168 59588
0 59590 5 1 1 59589
0 59591 7 1 2 59585 59590
0 59592 5 1 1 59591
0 59593 7 1 2 67239 59592
0 59594 5 1 1 59593
0 59595 7 1 2 90834 92729
0 59596 5 2 1 59595
0 59597 7 1 2 107170 106960
0 59598 5 1 1 59597
0 59599 7 1 2 84687 105208
0 59600 5 1 1 59599
0 59601 7 1 2 59598 59600
0 59602 5 1 1 59601
0 59603 7 1 2 107047 59602
0 59604 5 1 1 59603
0 59605 7 1 2 59594 59604
0 59606 5 1 1 59605
0 59607 7 1 2 70923 59606
0 59608 5 1 1 59607
0 59609 7 1 2 79775 84001
0 59610 7 1 2 103933 89521
0 59611 7 1 2 59609 59610
0 59612 7 1 2 93539 59611
0 59613 5 1 1 59612
0 59614 7 1 2 59608 59613
0 59615 5 1 1 59614
0 59616 7 1 2 85367 59615
0 59617 5 1 1 59616
0 59618 7 1 2 101433 97534
0 59619 7 1 2 99064 59618
0 59620 5 1 1 59619
0 59621 7 1 2 88928 106884
0 59622 5 1 1 59621
0 59623 7 2 2 72281 99361
0 59624 5 1 1 107172
0 59625 7 1 2 88411 107173
0 59626 5 1 1 59625
0 59627 7 1 2 59622 59626
0 59628 5 1 1 59627
0 59629 7 1 2 65859 98849
0 59630 7 1 2 59628 59629
0 59631 5 1 1 59630
0 59632 7 1 2 59620 59631
0 59633 5 1 1 59632
0 59634 7 2 2 77912 92078
0 59635 7 1 2 59633 107174
0 59636 5 1 1 59635
0 59637 7 1 2 69318 59636
0 59638 7 1 2 59617 59637
0 59639 5 1 1 59638
0 59640 7 1 2 64528 107096
0 59641 5 1 1 59640
0 59642 7 1 2 80433 92721
0 59643 5 1 1 59642
0 59644 7 1 2 59573 59643
0 59645 5 1 1 59644
0 59646 7 1 2 92844 59645
0 59647 7 1 2 59641 59646
0 59648 5 1 1 59647
0 59649 7 1 2 103179 41368
0 59650 5 1 1 59649
0 59651 7 1 2 65234 104909
0 59652 7 1 2 59650 59651
0 59653 5 1 1 59652
0 59654 7 1 2 59648 59653
0 59655 5 1 1 59654
0 59656 7 1 2 70569 59655
0 59657 5 1 1 59656
0 59658 7 1 2 93064 90819
0 59659 7 1 2 107036 59658
0 59660 5 1 1 59659
0 59661 7 1 2 59657 59660
0 59662 5 1 1 59661
0 59663 7 1 2 102607 89522
0 59664 7 1 2 59662 59663
0 59665 5 1 1 59664
0 59666 7 2 2 70924 98850
0 59667 5 1 1 107176
0 59668 7 1 2 98817 59667
0 59669 5 1 1 59668
0 59670 7 1 2 107115 59669
0 59671 5 1 1 59670
0 59672 7 1 2 90599 92444
0 59673 7 1 2 107137 59672
0 59674 5 1 1 59673
0 59675 7 1 2 59671 59674
0 59676 5 1 1 59675
0 59677 7 1 2 81804 59676
0 59678 5 1 1 59677
0 59679 7 2 2 99798 103342
0 59680 7 1 2 63995 80783
0 59681 7 1 2 93474 59680
0 59682 7 1 2 107178 59681
0 59683 5 1 1 59682
0 59684 7 1 2 88373 107052
0 59685 7 1 2 107177 59684
0 59686 5 1 1 59685
0 59687 7 1 2 59683 59686
0 59688 7 1 2 59678 59687
0 59689 5 1 1 59688
0 59690 7 1 2 107175 59689
0 59691 5 1 1 59690
0 59692 7 1 2 64219 59691
0 59693 7 1 2 59665 59692
0 59694 5 1 1 59693
0 59695 7 1 2 59639 59694
0 59696 5 1 1 59695
0 59697 7 1 2 68219 59696
0 59698 5 1 1 59697
0 59699 7 1 2 99743 101434
0 59700 5 1 1 59699
0 59701 7 1 2 35268 59700
0 59702 5 1 1 59701
0 59703 7 1 2 106961 59702
0 59704 5 1 1 59703
0 59705 7 1 2 84715 101435
0 59706 7 1 2 106591 59705
0 59707 5 1 1 59706
0 59708 7 1 2 59704 59707
0 59709 5 1 1 59708
0 59710 7 1 2 69319 59709
0 59711 5 1 1 59710
0 59712 7 1 2 64220 93421
0 59713 5 1 1 59712
0 59714 7 1 2 10938 59713
0 59715 5 1 1 59714
0 59716 7 1 2 67829 59715
0 59717 5 1 1 59716
0 59718 7 1 2 84532 90832
0 59719 5 1 1 59718
0 59720 7 1 2 59717 59719
0 59721 5 1 1 59720
0 59722 7 1 2 84916 59721
0 59723 5 1 1 59722
0 59724 7 1 2 68734 102232
0 59725 7 1 2 84721 59724
0 59726 5 1 1 59725
0 59727 7 1 2 59723 59726
0 59728 5 1 1 59727
0 59729 7 1 2 70285 59728
0 59730 5 1 1 59729
0 59731 7 1 2 81805 93664
0 59732 7 1 2 102583 59731
0 59733 5 1 1 59732
0 59734 7 1 2 59730 59733
0 59735 5 1 1 59734
0 59736 7 1 2 67240 59735
0 59737 5 1 1 59736
0 59738 7 1 2 59711 59737
0 59739 5 1 1 59738
0 59740 7 1 2 65699 59739
0 59741 5 1 1 59740
0 59742 7 1 2 85088 102395
0 59743 7 2 2 106969 59742
0 59744 7 1 2 107082 107180
0 59745 5 1 1 59744
0 59746 7 1 2 59741 59745
0 59747 5 1 1 59746
0 59748 7 1 2 63996 59747
0 59749 5 1 1 59748
0 59750 7 1 2 107132 107181
0 59751 5 1 1 59750
0 59752 7 1 2 59749 59751
0 59753 5 1 1 59752
0 59754 7 1 2 98011 59753
0 59755 5 1 1 59754
0 59756 7 1 2 102580 92027
0 59757 5 2 1 59756
0 59758 7 2 2 87931 102551
0 59759 7 1 2 70646 93627
0 59760 7 1 2 107184 59759
0 59761 5 1 1 59760
0 59762 7 1 2 107182 59761
0 59763 5 1 1 59762
0 59764 7 1 2 64529 59763
0 59765 5 1 1 59764
0 59766 7 1 2 69666 90515
0 59767 7 1 2 107185 59766
0 59768 5 1 1 59767
0 59769 7 1 2 107183 59768
0 59770 5 1 1 59769
0 59771 7 1 2 66093 59770
0 59772 5 1 1 59771
0 59773 7 1 2 59765 59772
0 59774 5 1 1 59773
0 59775 7 1 2 72836 59774
0 59776 5 1 1 59775
0 59777 7 2 2 92137 90516
0 59778 7 1 2 67241 81540
0 59779 7 1 2 99765 59778
0 59780 7 1 2 107186 59779
0 59781 5 1 1 59780
0 59782 7 1 2 59776 59781
0 59783 5 1 1 59782
0 59784 7 1 2 69073 59783
0 59785 5 1 1 59784
0 59786 7 1 2 77275 81972
0 59787 7 1 2 98012 59786
0 59788 7 1 2 107113 59787
0 59789 5 1 1 59788
0 59790 7 1 2 59785 59789
0 59791 5 1 1 59790
0 59792 7 1 2 81806 59791
0 59793 5 1 1 59792
0 59794 7 1 2 80784 86201
0 59795 7 1 2 75675 59794
0 59796 7 1 2 99362 59795
0 59797 7 1 2 107179 59796
0 59798 5 1 1 59797
0 59799 7 1 2 59793 59798
0 59800 5 1 1 59799
0 59801 7 1 2 85559 59800
0 59802 5 1 1 59801
0 59803 7 1 2 83413 85089
0 59804 7 1 2 84511 94479
0 59805 7 1 2 59803 59804
0 59806 7 2 2 76893 102552
0 59807 7 1 2 107162 107188
0 59808 7 1 2 59805 59807
0 59809 5 1 1 59808
0 59810 7 1 2 73288 59809
0 59811 7 1 2 59802 59810
0 59812 7 1 2 59755 59811
0 59813 5 1 1 59812
0 59814 7 1 2 59698 59813
0 59815 5 1 1 59814
0 59816 7 1 2 72490 59815
0 59817 5 1 1 59816
0 59818 7 2 2 96709 97642
0 59819 5 1 1 107190
0 59820 7 3 2 90517 91343
0 59821 7 1 2 70286 75537
0 59822 7 1 2 105108 59821
0 59823 7 1 2 107192 59822
0 59824 5 1 1 59823
0 59825 7 1 2 59819 59824
0 59826 5 1 1 59825
0 59827 7 1 2 66412 59826
0 59828 5 1 1 59827
0 59829 7 2 2 92138 90378
0 59830 7 1 2 81094 107195
0 59831 5 1 1 59830
0 59832 7 1 2 59828 59831
0 59833 5 1 1 59832
0 59834 7 1 2 67830 59833
0 59835 5 1 1 59834
0 59836 7 1 2 81973 92139
0 59837 7 1 2 107193 59836
0 59838 7 1 2 106911 59837
0 59839 5 1 1 59838
0 59840 7 1 2 59835 59839
0 59841 5 1 1 59840
0 59842 7 1 2 66806 59841
0 59843 5 1 1 59842
0 59844 7 1 2 91140 74289
0 59845 7 1 2 89523 59844
0 59846 7 1 2 67831 87870
0 59847 7 1 2 91976 59846
0 59848 7 1 2 59845 59847
0 59849 5 1 1 59848
0 59850 7 1 2 59843 59849
0 59851 5 1 1 59850
0 59852 7 1 2 65538 59851
0 59853 5 1 1 59852
0 59854 7 1 2 94535 103702
0 59855 7 1 2 90820 59854
0 59856 5 1 1 59855
0 59857 7 1 2 84716 91506
0 59858 7 1 2 105019 59857
0 59859 5 1 1 59858
0 59860 7 1 2 59856 59859
0 59861 5 1 1 59860
0 59862 7 1 2 98073 107187
0 59863 7 1 2 59861 59862
0 59864 5 1 1 59863
0 59865 7 1 2 59853 59864
0 59866 5 1 1 59865
0 59867 7 1 2 68220 59866
0 59868 5 1 1 59867
0 59869 7 1 2 71519 107191
0 59870 5 1 1 59869
0 59871 7 1 2 76876 92140
0 59872 7 1 2 107194 59871
0 59873 5 1 1 59872
0 59874 7 1 2 59870 59873
0 59875 5 1 1 59874
0 59876 7 1 2 106192 59875
0 59877 5 1 1 59876
0 59878 7 1 2 59868 59877
0 59879 5 1 1 59878
0 59880 7 1 2 72282 59879
0 59881 5 1 1 59880
0 59882 7 1 2 76518 80548
0 59883 7 1 2 100582 94237
0 59884 7 1 2 59882 59883
0 59885 7 2 2 83913 92141
0 59886 7 1 2 99363 107197
0 59887 7 1 2 59884 59886
0 59888 5 1 1 59887
0 59889 7 1 2 59881 59888
0 59890 5 1 1 59889
0 59891 7 1 2 85560 59890
0 59892 5 1 1 59891
0 59893 7 1 2 97345 96109
0 59894 5 1 1 59893
0 59895 7 1 2 75109 83122
0 59896 7 1 2 98005 59895
0 59897 5 1 1 59896
0 59898 7 1 2 59894 59897
0 59899 5 1 1 59898
0 59900 7 1 2 91914 59899
0 59901 5 1 1 59900
0 59902 7 2 2 70647 93475
0 59903 7 1 2 99556 79522
0 59904 7 1 2 83921 59903
0 59905 7 1 2 107199 59904
0 59906 5 1 1 59905
0 59907 7 1 2 59901 59906
0 59908 5 1 1 59907
0 59909 7 1 2 76252 59908
0 59910 5 1 1 59909
0 59911 7 1 2 78810 97433
0 59912 7 2 2 84344 90518
0 59913 7 1 2 106382 107201
0 59914 7 1 2 59911 59913
0 59915 5 1 1 59914
0 59916 7 1 2 59910 59915
0 59917 5 1 1 59916
0 59918 7 1 2 66807 59917
0 59919 5 1 1 59918
0 59920 7 1 2 75612 93639
0 59921 7 2 2 98013 59920
0 59922 7 1 2 96110 107037
0 59923 5 1 1 59922
0 59924 7 1 2 97861 80213
0 59925 7 1 2 105235 59924
0 59926 5 1 1 59925
0 59927 7 1 2 59923 59926
0 59928 5 1 1 59927
0 59929 7 1 2 107203 59928
0 59930 5 1 1 59929
0 59931 7 1 2 103320 93205
0 59932 7 1 2 107198 107200
0 59933 7 1 2 59931 59932
0 59934 5 1 1 59933
0 59935 7 1 2 59930 59934
0 59936 7 1 2 59919 59935
0 59937 5 1 1 59936
0 59938 7 1 2 63997 59937
0 59939 5 1 1 59938
0 59940 7 2 2 99615 102032
0 59941 5 1 1 107205
0 59942 7 1 2 75787 83671
0 59943 7 1 2 102109 59942
0 59944 5 1 1 59943
0 59945 7 1 2 59941 59944
0 59946 5 1 1 59945
0 59947 7 1 2 69320 99061
0 59948 5 1 1 59947
0 59949 7 1 2 64221 10695
0 59950 5 1 1 59949
0 59951 7 4 2 59948 59950
0 59952 7 1 2 94805 95658
0 59953 7 1 2 107207 59952
0 59954 7 1 2 59946 59953
0 59955 5 1 1 59954
0 59956 7 1 2 59939 59955
0 59957 5 1 1 59956
0 59958 7 1 2 100583 59957
0 59959 5 1 1 59958
0 59960 7 1 2 80841 75594
0 59961 7 2 2 99050 59960
0 59962 7 1 2 93476 107211
0 59963 5 1 1 59962
0 59964 7 1 2 92343 93640
0 59965 7 1 2 91550 59964
0 59966 5 1 1 59965
0 59967 7 1 2 59963 59966
0 59968 5 1 1 59967
0 59969 7 1 2 69074 59968
0 59970 5 1 1 59969
0 59971 7 1 2 99350 81162
0 59972 7 1 2 95654 59971
0 59973 5 1 1 59972
0 59974 7 1 2 59970 59973
0 59975 5 1 1 59974
0 59976 7 1 2 64222 59975
0 59977 5 1 1 59976
0 59978 7 1 2 76034 87966
0 59979 7 1 2 105470 59978
0 59980 7 1 2 103642 59979
0 59981 5 1 1 59980
0 59982 7 1 2 59977 59981
0 59983 5 1 1 59982
0 59984 7 1 2 84917 59983
0 59985 5 1 1 59984
0 59986 7 1 2 106786 107204
0 59987 5 1 1 59986
0 59988 7 1 2 70740 92452
0 59989 7 1 2 107212 59988
0 59990 5 1 1 59989
0 59991 7 1 2 59987 59990
0 59992 5 1 1 59991
0 59993 7 1 2 100120 59992
0 59994 5 1 1 59993
0 59995 7 1 2 59985 59994
0 59996 5 1 1 59995
0 59997 7 1 2 70287 59996
0 59998 5 1 1 59997
0 59999 7 1 2 94661 107042
0 60000 5 1 1 59999
0 60001 7 1 2 83914 98579
0 60002 7 1 2 107111 60001
0 60003 5 1 1 60002
0 60004 7 1 2 60000 60003
0 60005 5 1 1 60004
0 60006 7 1 2 107196 60005
0 60007 5 1 1 60006
0 60008 7 1 2 76110 99813
0 60009 5 1 1 60008
0 60010 7 1 2 81163 106919
0 60011 5 1 1 60010
0 60012 7 1 2 60009 60011
0 60013 5 1 1 60012
0 60014 7 1 2 91915 106787
0 60015 7 1 2 60013 60014
0 60016 5 1 1 60015
0 60017 7 1 2 60007 60016
0 60018 5 1 1 60017
0 60019 7 1 2 70925 60018
0 60020 5 1 1 60019
0 60021 7 1 2 74320 84602
0 60022 7 1 2 99364 60021
0 60023 7 1 2 76111 98060
0 60024 7 1 2 60022 60023
0 60025 5 1 1 60024
0 60026 7 1 2 72837 60025
0 60027 7 1 2 60020 60026
0 60028 7 1 2 59998 60027
0 60029 5 1 1 60028
0 60030 7 1 2 66903 94075
0 60031 7 1 2 89678 60030
0 60032 7 1 2 105621 60031
0 60033 7 1 2 106946 60032
0 60034 5 1 1 60033
0 60035 7 1 2 96133 96514
0 60036 7 1 2 107202 60035
0 60037 5 1 1 60036
0 60038 7 1 2 60034 60037
0 60039 5 1 1 60038
0 60040 7 1 2 107043 60039
0 60041 5 1 1 60040
0 60042 7 1 2 67832 60041
0 60043 5 1 1 60042
0 60044 7 1 2 72283 60043
0 60045 7 1 2 60029 60044
0 60046 5 1 1 60045
0 60047 7 1 2 67486 60046
0 60048 7 1 2 59959 60047
0 60049 7 1 2 59892 60048
0 60050 5 1 1 60049
0 60051 7 1 2 63824 60050
0 60052 7 1 2 59817 60051
0 60053 5 1 1 60052
0 60054 7 1 2 103046 91512
0 60055 7 1 2 84401 60054
0 60056 5 1 1 60055
0 60057 7 1 2 64223 76112
0 60058 5 1 1 60057
0 60059 7 1 2 80858 99785
0 60060 5 1 1 60059
0 60061 7 1 2 60058 60060
0 60062 5 1 1 60061
0 60063 7 1 2 79647 106167
0 60064 7 1 2 60062 60063
0 60065 5 1 1 60064
0 60066 7 1 2 60056 60065
0 60067 5 1 1 60066
0 60068 7 1 2 69075 60067
0 60069 5 1 1 60068
0 60070 7 1 2 76113 107208
0 60071 5 1 1 60070
0 60072 7 2 2 70288 79742
0 60073 5 1 1 107213
0 60074 7 1 2 65700 104826
0 60075 7 1 2 107214 60074
0 60076 5 1 1 60075
0 60077 7 1 2 60071 60076
0 60078 5 1 1 60077
0 60079 7 1 2 92281 98014
0 60080 7 1 2 60078 60079
0 60081 5 1 1 60080
0 60082 7 1 2 60069 60081
0 60083 5 1 1 60082
0 60084 7 1 2 66808 60083
0 60085 5 1 1 60084
0 60086 7 1 2 73289 56631
0 60087 7 1 2 99365 60086
0 60088 7 1 2 99777 94973
0 60089 7 1 2 60087 60088
0 60090 7 1 2 99331 60089
0 60091 5 1 1 60090
0 60092 7 1 2 60085 60091
0 60093 5 1 1 60092
0 60094 7 1 2 65539 60093
0 60095 5 1 1 60094
0 60096 7 1 2 91454 107099
0 60097 7 1 2 82421 60096
0 60098 5 1 1 60097
0 60099 7 1 2 82016 97632
0 60100 7 1 2 107101 60099
0 60101 5 1 1 60100
0 60102 7 1 2 60098 60101
0 60103 5 1 1 60102
0 60104 7 1 2 63998 60103
0 60105 5 1 1 60104
0 60106 7 1 2 99778 86532
0 60107 5 1 1 60106
0 60108 7 1 2 65860 105236
0 60109 5 1 1 60108
0 60110 7 1 2 60107 60109
0 60111 5 1 1 60110
0 60112 7 1 2 99345 101284
0 60113 7 1 2 60111 60112
0 60114 5 1 1 60113
0 60115 7 1 2 60105 60114
0 60116 5 1 1 60115
0 60117 7 2 2 78187 84382
0 60118 7 1 2 86616 107215
0 60119 7 1 2 60116 60118
0 60120 5 1 1 60119
0 60121 7 1 2 60095 60120
0 60122 5 1 1 60121
0 60123 7 1 2 72284 60122
0 60124 5 1 1 60123
0 60125 7 1 2 95652 94816
0 60126 7 1 2 107057 60125
0 60127 7 1 2 87135 87442
0 60128 7 1 2 95117 60127
0 60129 7 1 2 87112 60128
0 60130 7 1 2 60126 60129
0 60131 5 1 1 60130
0 60132 7 1 2 60124 60131
0 60133 5 1 1 60132
0 60134 7 1 2 99212 60133
0 60135 5 1 1 60134
0 60136 7 2 2 63999 99744
0 60137 7 1 2 71216 86800
0 60138 5 1 1 60137
0 60139 7 1 2 104752 60138
0 60140 5 1 1 60139
0 60141 7 1 2 107217 60140
0 60142 5 1 1 60141
0 60143 7 1 2 73290 92415
0 60144 7 1 2 91713 60143
0 60145 7 1 2 95181 60144
0 60146 5 1 1 60145
0 60147 7 1 2 60142 60146
0 60148 5 1 1 60147
0 60149 7 1 2 65235 60148
0 60150 5 1 1 60149
0 60151 7 2 2 66413 88698
0 60152 7 1 2 99599 105529
0 60153 7 1 2 107219 60152
0 60154 5 1 1 60153
0 60155 7 1 2 60150 60154
0 60156 5 1 1 60155
0 60157 7 1 2 69321 60156
0 60158 5 1 1 60157
0 60159 7 1 2 99425 106878
0 60160 5 1 1 60159
0 60161 7 1 2 100824 92389
0 60162 5 1 1 60161
0 60163 7 1 2 60160 60162
0 60164 5 1 1 60163
0 60165 7 1 2 87988 60164
0 60166 5 1 1 60165
0 60167 7 1 2 92845 80037
0 60168 7 1 2 107220 60167
0 60169 5 1 1 60168
0 60170 7 1 2 60166 60169
0 60171 5 1 1 60170
0 60172 7 1 2 92453 60171
0 60173 5 1 1 60172
0 60174 7 1 2 60158 60173
0 60175 5 1 1 60174
0 60176 7 1 2 97064 60175
0 60177 5 1 1 60176
0 60178 7 2 2 69076 99268
0 60179 7 1 2 65236 106710
0 60180 5 1 1 60179
0 60181 7 1 2 104365 60180
0 60182 5 1 1 60181
0 60183 7 1 2 64530 60182
0 60184 5 1 1 60183
0 60185 7 1 2 77979 96605
0 60186 5 1 1 60185
0 60187 7 1 2 60184 60186
0 60188 5 1 1 60187
0 60189 7 1 2 107221 60188
0 60190 5 1 1 60189
0 60191 7 3 2 67487 90600
0 60192 7 1 2 85594 80155
0 60193 7 1 2 107223 60192
0 60194 5 1 1 60193
0 60195 7 1 2 60190 60194
0 60196 5 1 1 60195
0 60197 7 1 2 85561 60196
0 60198 5 1 1 60197
0 60199 7 1 2 96942 107169
0 60200 5 1 1 60199
0 60201 7 2 2 71875 96982
0 60202 7 1 2 79706 107226
0 60203 5 1 1 60202
0 60204 7 1 2 60200 60203
0 60205 5 1 1 60204
0 60206 7 1 2 98945 107218
0 60207 7 1 2 60205 60206
0 60208 5 1 1 60207
0 60209 7 2 2 75110 87018
0 60210 7 1 2 98598 107228
0 60211 5 1 1 60210
0 60212 7 1 2 80303 101165
0 60213 5 1 1 60212
0 60214 7 1 2 60211 60213
0 60215 5 1 1 60214
0 60216 7 1 2 76519 60215
0 60217 5 1 1 60216
0 60218 7 1 2 67488 107206
0 60219 5 1 1 60218
0 60220 7 1 2 60217 60219
0 60221 5 1 1 60220
0 60222 7 1 2 66809 60221
0 60223 5 1 1 60222
0 60224 7 1 2 93969 98477
0 60225 7 1 2 103057 60224
0 60226 5 1 1 60225
0 60227 7 1 2 60223 60226
0 60228 5 1 1 60227
0 60229 7 1 2 11222 11302
0 60230 7 1 2 85479 60229
0 60231 7 1 2 60228 60230
0 60232 5 1 1 60231
0 60233 7 1 2 60208 60232
0 60234 7 1 2 60198 60233
0 60235 5 1 1 60234
0 60236 7 1 2 72838 60235
0 60237 5 1 1 60236
0 60238 7 1 2 60177 60237
0 60239 5 1 1 60238
0 60240 7 1 2 70741 60239
0 60241 5 1 1 60240
0 60242 7 1 2 83074 97147
0 60243 5 1 1 60242
0 60244 7 1 2 101089 60243
0 60245 5 1 1 60244
0 60246 7 1 2 87989 60245
0 60247 5 1 1 60246
0 60248 7 1 2 43130 45510
0 60249 5 1 1 60248
0 60250 7 1 2 83141 98699
0 60251 7 1 2 60249 60250
0 60252 5 1 1 60251
0 60253 7 1 2 60247 60252
0 60254 5 1 1 60253
0 60255 7 1 2 76520 60254
0 60256 5 1 1 60255
0 60257 7 1 2 89197 97230
0 60258 5 1 1 60257
0 60259 7 3 2 70289 86869
0 60260 5 1 1 107230
0 60261 7 1 2 97076 107231
0 60262 5 1 1 60261
0 60263 7 1 2 60258 60262
0 60264 5 1 1 60263
0 60265 7 1 2 80047 60264
0 60266 5 1 1 60265
0 60267 7 1 2 60256 60266
0 60268 5 1 1 60267
0 60269 7 1 2 70926 60268
0 60270 5 1 1 60269
0 60271 7 1 2 99527 76968
0 60272 7 1 2 105223 60271
0 60273 5 1 1 60272
0 60274 7 1 2 60270 60273
0 60275 5 1 1 60274
0 60276 7 1 2 69322 60275
0 60277 5 1 1 60276
0 60278 7 1 2 80555 85036
0 60279 7 1 2 105946 60278
0 60280 5 1 1 60279
0 60281 7 1 2 60277 60280
0 60282 5 1 1 60281
0 60283 7 1 2 99346 60282
0 60284 5 1 1 60283
0 60285 7 1 2 60241 60284
0 60286 5 1 1 60285
0 60287 7 1 2 76011 60286
0 60288 5 1 1 60287
0 60289 7 1 2 83734 80038
0 60290 5 1 1 60289
0 60291 7 1 2 64531 84309
0 60292 7 1 2 9719 60291
0 60293 7 1 2 83765 60292
0 60294 5 1 1 60293
0 60295 7 1 2 60290 60294
0 60296 5 1 1 60295
0 60297 7 1 2 66414 60296
0 60298 5 1 1 60297
0 60299 7 1 2 84944 99234
0 60300 5 1 1 60299
0 60301 7 1 2 60298 60300
0 60302 5 1 1 60301
0 60303 7 1 2 96983 89554
0 60304 7 1 2 92445 60303
0 60305 7 1 2 94502 60304
0 60306 7 1 2 60302 60305
0 60307 5 1 1 60306
0 60308 7 1 2 60288 60307
0 60309 5 1 1 60308
0 60310 7 1 2 67242 60309
0 60311 5 1 1 60310
0 60312 7 1 2 78498 104967
0 60313 5 1 1 60312
0 60314 7 1 2 7631 60313
0 60315 5 1 1 60314
0 60316 7 1 2 69667 60315
0 60317 5 1 1 60316
0 60318 7 1 2 42864 60317
0 60319 5 1 1 60318
0 60320 7 1 2 85562 60319
0 60321 5 1 1 60320
0 60322 7 1 2 93613 84002
0 60323 7 1 2 95519 60322
0 60324 5 1 1 60323
0 60325 7 1 2 60321 60324
0 60326 5 1 1 60325
0 60327 7 1 2 67489 60326
0 60328 5 1 1 60327
0 60329 7 1 2 58565 107045
0 60330 5 1 1 60329
0 60331 7 1 2 72839 60330
0 60332 5 1 1 60331
0 60333 7 1 2 78503 60332
0 60334 5 1 1 60333
0 60335 7 1 2 71520 60334
0 60336 5 1 1 60335
0 60337 7 2 2 69668 84188
0 60338 7 1 2 95138 107233
0 60339 5 1 1 60338
0 60340 7 1 2 60336 60339
0 60341 5 1 1 60340
0 60342 7 1 2 99398 60341
0 60343 5 1 1 60342
0 60344 7 1 2 60328 60343
0 60345 5 1 1 60344
0 60346 7 1 2 68221 60345
0 60347 5 1 1 60346
0 60348 7 1 2 69669 98823
0 60349 5 1 1 60348
0 60350 7 1 2 105799 60349
0 60351 5 1 1 60350
0 60352 7 1 2 69323 60351
0 60353 5 1 1 60352
0 60354 7 1 2 101050 60353
0 60355 5 1 1 60354
0 60356 7 1 2 102483 60355
0 60357 5 1 1 60356
0 60358 7 1 2 60347 60357
0 60359 5 1 1 60358
0 60360 7 1 2 66810 60359
0 60361 5 1 1 60360
0 60362 7 2 2 85473 78420
0 60363 5 1 1 107235
0 60364 7 1 2 29266 60363
0 60365 5 1 1 60364
0 60366 7 1 2 76521 60365
0 60367 5 1 1 60366
0 60368 7 1 2 96086 104385
0 60369 5 1 1 60368
0 60370 7 1 2 60367 60369
0 60371 5 1 1 60370
0 60372 7 1 2 70290 97956
0 60373 7 1 2 83606 60372
0 60374 7 1 2 60371 60373
0 60375 5 1 1 60374
0 60376 7 1 2 60361 60375
0 60377 5 1 1 60376
0 60378 7 1 2 65540 60377
0 60379 5 1 1 60378
0 60380 7 1 2 98580 105050
0 60381 5 1 1 60380
0 60382 7 1 2 70291 104191
0 60383 5 1 1 60382
0 60384 7 1 2 60381 60383
0 60385 5 1 1 60384
0 60386 7 1 2 85563 60385
0 60387 5 1 1 60386
0 60388 7 1 2 93981 105239
0 60389 5 3 1 60388
0 60390 7 1 2 107236 107237
0 60391 5 1 1 60390
0 60392 7 1 2 60387 60391
0 60393 5 1 1 60392
0 60394 7 1 2 76522 60393
0 60395 5 1 1 60394
0 60396 7 1 2 103627 95300
0 60397 5 1 1 60396
0 60398 7 1 2 69670 98842
0 60399 7 1 2 105583 60398
0 60400 5 1 1 60399
0 60401 7 1 2 60397 60400
0 60402 5 1 1 60401
0 60403 7 1 2 69324 60402
0 60404 5 1 1 60403
0 60405 7 1 2 102356 84189
0 60406 7 1 2 106518 60405
0 60407 5 1 1 60406
0 60408 7 1 2 60404 60407
0 60409 5 1 1 60408
0 60410 7 1 2 76253 60409
0 60411 5 1 1 60410
0 60412 7 1 2 60395 60411
0 60413 5 1 1 60412
0 60414 7 1 2 67490 60413
0 60415 5 1 1 60414
0 60416 7 1 2 98380 92830
0 60417 7 1 2 102357 60416
0 60418 7 1 2 107171 60417
0 60419 5 1 1 60418
0 60420 7 1 2 60415 60419
0 60421 5 1 1 60420
0 60422 7 1 2 81444 60421
0 60423 5 1 1 60422
0 60424 7 1 2 60379 60423
0 60425 5 1 1 60424
0 60426 7 1 2 76012 107048
0 60427 7 1 2 60425 60426
0 60428 5 1 1 60427
0 60429 7 1 2 60311 60428
0 60430 5 1 1 60429
0 60431 7 1 2 85109 60430
0 60432 5 1 1 60431
0 60433 7 1 2 60135 60432
0 60434 7 1 2 60053 60433
0 60435 5 1 1 60434
0 60436 7 1 2 102268 60435
0 60437 5 1 1 60436
0 60438 7 1 2 59563 60437
0 60439 7 1 2 59166 60438
0 60440 5 1 1 60439
0 60441 7 1 2 67013 60440
0 60442 5 1 1 60441
0 60443 7 1 2 87194 83351
0 60444 5 1 1 60443
0 60445 7 1 2 103124 60444
0 60446 5 1 1 60445
0 60447 7 2 2 64532 102253
0 60448 5 1 1 107240
0 60449 7 1 2 69671 101200
0 60450 5 1 1 60449
0 60451 7 1 2 60448 60450
0 60452 5 2 1 60451
0 60453 7 1 2 60446 107242
0 60454 5 1 1 60453
0 60455 7 1 2 91141 102730
0 60456 7 1 2 104285 60455
0 60457 5 1 1 60456
0 60458 7 1 2 60454 60457
0 60459 5 1 1 60458
0 60460 7 1 2 70742 60459
0 60461 5 1 1 60460
0 60462 7 5 2 67833 103296
0 60463 7 1 2 73291 105618
0 60464 7 1 2 107244 60463
0 60465 7 1 2 106998 60464
0 60466 5 1 1 60465
0 60467 7 1 2 60461 60466
0 60468 5 1 1 60467
0 60469 7 1 2 72198 60468
0 60470 5 1 1 60469
0 60471 7 1 2 103359 97171
0 60472 7 1 2 107006 60471
0 60473 5 1 1 60472
0 60474 7 1 2 60470 60473
0 60475 5 1 1 60474
0 60476 7 1 2 69077 60475
0 60477 5 1 1 60476
0 60478 7 1 2 64533 104770
0 60479 5 1 1 60478
0 60480 7 1 2 90868 104513
0 60481 5 1 1 60480
0 60482 7 1 2 60479 60481
0 60483 5 1 1 60482
0 60484 7 1 2 70743 60483
0 60485 7 1 2 106999 60484
0 60486 5 1 1 60485
0 60487 7 2 2 98776 102647
0 60488 7 1 2 105619 107249
0 60489 7 1 2 86077 60488
0 60490 5 1 1 60489
0 60491 7 1 2 60486 60490
0 60492 5 1 1 60491
0 60493 7 1 2 94817 60492
0 60494 5 1 1 60493
0 60495 7 1 2 60477 60494
0 60496 5 1 1 60495
0 60497 7 1 2 70692 60496
0 60498 5 1 1 60497
0 60499 7 1 2 70744 99674
0 60500 5 2 1 60499
0 60501 7 1 2 99355 107251
0 60502 5 1 1 60501
0 60503 7 2 2 59624 60502
0 60504 7 1 2 81935 107253
0 60505 5 1 1 60504
0 60506 7 2 2 80663 107049
0 60507 5 1 1 107255
0 60508 7 1 2 60505 60507
0 60509 5 1 1 60508
0 60510 7 2 2 73292 60509
0 60511 7 2 2 103759 107257
0 60512 7 1 2 96583 107259
0 60513 5 1 1 60512
0 60514 7 1 2 60498 60513
0 60515 5 1 1 60514
0 60516 7 1 2 69027 60515
0 60517 5 1 1 60516
0 60518 7 1 2 69672 106277
0 60519 7 1 2 107260 60518
0 60520 5 1 1 60519
0 60521 7 1 2 60517 60520
0 60522 5 1 1 60521
0 60523 7 1 2 76813 60522
0 60524 5 1 1 60523
0 60525 7 3 2 99366 81936
0 60526 7 2 2 67243 107261
0 60527 5 1 1 107264
0 60528 7 1 2 100811 107265
0 60529 5 2 1 60528
0 60530 7 1 2 72285 86078
0 60531 7 1 2 96374 60530
0 60532 5 1 1 60531
0 60533 7 1 2 107266 60532
0 60534 5 1 1 60533
0 60535 7 1 2 99088 98015
0 60536 7 1 2 60534 60535
0 60537 5 1 1 60536
0 60538 7 1 2 60524 60537
0 60539 5 1 1 60538
0 60540 7 1 2 68896 60539
0 60541 5 1 1 60540
0 60542 7 1 2 104324 107254
0 60543 5 1 1 60542
0 60544 7 2 2 65701 72286
0 60545 5 1 1 107268
0 60546 7 2 2 68735 107269
0 60547 5 1 1 107270
0 60548 7 1 2 102269 89555
0 60549 7 1 2 107271 60548
0 60550 5 1 1 60549
0 60551 7 1 2 60543 60550
0 60552 5 1 1 60551
0 60553 7 1 2 81937 60552
0 60554 5 1 1 60553
0 60555 7 4 2 72287 80664
0 60556 7 1 2 96387 107272
0 60557 5 1 1 60556
0 60558 7 1 2 60554 60557
0 60559 5 1 1 60558
0 60560 7 1 2 98777 103150
0 60561 7 1 2 91853 60560
0 60562 7 1 2 60559 60561
0 60563 5 1 1 60562
0 60564 7 1 2 60541 60563
0 60565 5 1 1 60564
0 60566 7 1 2 72068 60565
0 60567 5 1 1 60566
0 60568 7 1 2 96445 98309
0 60569 5 1 1 60568
0 60570 7 1 2 106923 60569
0 60571 5 4 1 60570
0 60572 7 1 2 99089 102648
0 60573 7 1 2 107276 60572
0 60574 7 1 2 97193 60573
0 60575 5 1 1 60574
0 60576 7 1 2 60567 60575
0 60577 5 1 1 60576
0 60578 7 1 2 85564 60577
0 60579 5 1 1 60578
0 60580 7 1 2 166 93832
0 60581 5 5 1 60580
0 60582 7 2 2 97466 92142
0 60583 7 1 2 74412 91561
0 60584 7 1 2 91647 60583
0 60585 7 1 2 107285 60584
0 60586 5 1 1 60585
0 60587 7 2 2 84304 97484
0 60588 7 1 2 100975 107287
0 60589 5 1 1 60588
0 60590 7 1 2 99096 98570
0 60591 5 1 1 60590
0 60592 7 1 2 60589 60591
0 60593 5 1 1 60592
0 60594 7 1 2 63937 60593
0 60595 5 1 1 60594
0 60596 7 1 2 103304 107286
0 60597 5 1 1 60596
0 60598 7 1 2 60595 60597
0 60599 5 1 1 60598
0 60600 7 1 2 70927 99367
0 60601 7 1 2 60599 60600
0 60602 5 1 1 60601
0 60603 7 1 2 60586 60602
0 60604 5 1 1 60603
0 60605 7 1 2 107280 60604
0 60606 5 1 1 60605
0 60607 7 2 2 91399 106622
0 60608 7 1 2 98880 107289
0 60609 5 1 1 60608
0 60610 7 1 2 70745 96777
0 60611 7 1 2 106440 60610
0 60612 5 1 1 60611
0 60613 7 1 2 60609 60612
0 60614 5 1 1 60613
0 60615 7 1 2 70292 60614
0 60616 5 1 1 60615
0 60617 7 2 2 74442 91156
0 60618 7 1 2 98778 105452
0 60619 7 1 2 107291 60618
0 60620 5 1 1 60619
0 60621 7 1 2 65541 60620
0 60622 7 1 2 60616 60621
0 60623 5 1 1 60622
0 60624 7 1 2 65861 98581
0 60625 7 1 2 107290 60624
0 60626 5 1 1 60625
0 60627 7 1 2 102451 93477
0 60628 7 1 2 97355 60627
0 60629 5 1 1 60628
0 60630 7 1 2 70570 60629
0 60631 7 1 2 60626 60630
0 60632 5 1 1 60631
0 60633 7 1 2 64000 60632
0 60634 7 1 2 60623 60633
0 60635 5 1 1 60634
0 60636 7 1 2 77998 105919
0 60637 5 1 1 60636
0 60638 7 1 2 69325 90454
0 60639 5 1 1 60638
0 60640 7 1 2 43255 60639
0 60641 5 1 1 60640
0 60642 7 1 2 65542 74443
0 60643 7 1 2 60641 60642
0 60644 5 1 1 60643
0 60645 7 1 2 60637 60644
0 60646 5 1 1 60645
0 60647 7 1 2 91562 105802
0 60648 7 1 2 60646 60647
0 60649 5 1 1 60648
0 60650 7 1 2 60635 60649
0 60651 5 1 1 60650
0 60652 7 1 2 72199 60651
0 60653 5 1 1 60652
0 60654 7 1 2 91249 92446
0 60655 7 1 2 100997 60654
0 60656 5 1 1 60655
0 60657 7 1 2 60653 60656
0 60658 5 1 1 60657
0 60659 7 1 2 100304 60658
0 60660 5 1 1 60659
0 60661 7 1 2 60606 60660
0 60662 5 1 1 60661
0 60663 7 1 2 63825 60662
0 60664 5 1 1 60663
0 60665 7 6 2 99368 102270
0 60666 7 1 2 82480 107293
0 60667 5 1 1 60666
0 60668 7 1 2 64224 91563
0 60669 7 1 2 105784 60668
0 60670 5 1 1 60669
0 60671 7 1 2 60667 60670
0 60672 5 1 1 60671
0 60673 7 1 2 65615 60672
0 60674 5 1 1 60673
0 60675 7 2 2 93310 92607
0 60676 5 1 1 107299
0 60677 7 1 2 90292 107300
0 60678 5 1 1 60677
0 60679 7 1 2 60674 60678
0 60680 5 1 1 60679
0 60681 7 1 2 85110 107288
0 60682 7 1 2 107281 60681
0 60683 7 1 2 60680 60682
0 60684 5 1 1 60683
0 60685 7 1 2 60664 60684
0 60686 5 1 1 60685
0 60687 7 1 2 67014 60686
0 60688 5 1 1 60687
0 60689 7 1 2 69078 107209
0 60690 5 1 1 60689
0 60691 7 1 2 59541 60690
0 60692 5 1 1 60691
0 60693 7 2 2 73293 104536
0 60694 7 2 2 94591 78999
0 60695 7 2 2 98140 90886
0 60696 7 1 2 107303 107305
0 60697 7 1 2 107301 60696
0 60698 7 1 2 107282 60697
0 60699 7 1 2 60692 60698
0 60700 5 1 1 60699
0 60701 7 1 2 67244 60700
0 60702 7 1 2 60688 60701
0 60703 5 1 1 60702
0 60704 7 1 2 84688 92473
0 60705 5 1 1 60704
0 60706 7 1 2 96497 60705
0 60707 5 1 1 60706
0 60708 7 1 2 67491 60707
0 60709 5 1 1 60708
0 60710 7 1 2 89092 102119
0 60711 7 2 2 70746 96402
0 60712 7 1 2 88044 107307
0 60713 7 1 2 60710 60712
0 60714 5 1 1 60713
0 60715 7 1 2 60709 60714
0 60716 5 1 1 60715
0 60717 7 1 2 69326 60716
0 60718 5 1 1 60717
0 60719 7 1 2 101096 105622
0 60720 5 1 1 60719
0 60721 7 1 2 99356 99457
0 60722 5 1 1 60721
0 60723 7 1 2 19238 88934
0 60724 5 1 1 60723
0 60725 7 1 2 81541 60724
0 60726 7 1 2 60722 60725
0 60727 5 1 1 60726
0 60728 7 1 2 60720 60727
0 60729 5 1 1 60728
0 60730 7 1 2 85351 88906
0 60731 7 1 2 60729 60730
0 60732 5 1 1 60731
0 60733 7 1 2 60718 60732
0 60734 5 1 1 60733
0 60735 7 1 2 84383 60734
0 60736 5 1 1 60735
0 60737 7 1 2 94592 104789
0 60738 7 1 2 83206 60737
0 60739 7 1 2 107135 60738
0 60740 5 1 1 60739
0 60741 7 1 2 60736 60740
0 60742 5 1 1 60741
0 60743 7 1 2 69028 60742
0 60744 5 1 1 60743
0 60745 7 3 2 65862 99369
0 60746 7 2 2 95588 107216
0 60747 7 1 2 70693 107312
0 60748 5 1 1 60747
0 60749 7 1 2 96316 106420
0 60750 7 1 2 99057 60749
0 60751 5 2 1 60750
0 60752 7 1 2 60748 107314
0 60753 5 1 1 60752
0 60754 7 1 2 107309 60753
0 60755 5 1 1 60754
0 60756 7 1 2 82481 96226
0 60757 7 1 2 90399 60756
0 60758 5 1 1 60757
0 60759 7 1 2 60755 60758
0 60760 5 1 1 60759
0 60761 7 1 2 75199 97065
0 60762 7 1 2 60760 60761
0 60763 5 1 1 60762
0 60764 7 1 2 60744 60763
0 60765 5 1 1 60764
0 60766 7 1 2 106947 60765
0 60767 5 1 1 60766
0 60768 7 1 2 87828 90276
0 60769 5 1 1 60768
0 60770 7 1 2 92864 90887
0 60771 7 1 2 83085 60770
0 60772 5 1 1 60771
0 60773 7 1 2 60769 60772
0 60774 5 1 1 60773
0 60775 7 1 2 107310 60774
0 60776 5 1 1 60775
0 60777 7 1 2 84076 84305
0 60778 7 1 2 95623 102796
0 60779 7 1 2 88929 60778
0 60780 7 1 2 60777 60779
0 60781 5 1 1 60780
0 60782 7 1 2 60776 60781
0 60783 5 1 1 60782
0 60784 7 1 2 72491 60783
0 60785 5 1 1 60784
0 60786 7 2 2 67145 94818
0 60787 7 1 2 100371 90607
0 60788 7 1 2 107316 60787
0 60789 7 1 2 105206 60788
0 60790 5 1 1 60789
0 60791 7 1 2 60785 60790
0 60792 5 1 1 60791
0 60793 7 1 2 65658 60792
0 60794 5 1 1 60793
0 60795 7 2 2 70747 93577
0 60796 7 1 2 70928 78084
0 60797 7 1 2 107318 60796
0 60798 5 1 1 60797
0 60799 7 1 2 64225 75168
0 60800 7 1 2 107311 60799
0 60801 5 1 1 60800
0 60802 7 1 2 60798 60801
0 60803 5 1 1 60802
0 60804 7 2 2 97066 89398
0 60805 7 1 2 96500 107320
0 60806 7 1 2 60803 60805
0 60807 5 1 1 60806
0 60808 7 1 2 60794 60807
0 60809 5 1 1 60808
0 60810 7 1 2 63826 60809
0 60811 5 1 1 60810
0 60812 7 1 2 74413 107294
0 60813 5 1 1 60812
0 60814 7 2 2 70929 89550
0 60815 7 2 2 69029 106788
0 60816 7 1 2 107322 107324
0 60817 5 1 1 60816
0 60818 7 1 2 60813 60817
0 60819 5 1 1 60818
0 60820 7 1 2 101989 107321
0 60821 7 1 2 60819 60820
0 60822 5 1 1 60821
0 60823 7 1 2 60811 60822
0 60824 5 1 1 60823
0 60825 7 1 2 106582 60824
0 60826 5 1 1 60825
0 60827 7 1 2 84882 104139
0 60828 5 1 1 60827
0 60829 7 1 2 81938 96790
0 60830 5 1 1 60829
0 60831 7 1 2 60828 60830
0 60832 5 1 1 60831
0 60833 7 1 2 82482 96668
0 60834 5 1 1 60833
0 60835 7 1 2 99370 84444
0 60836 5 1 1 60835
0 60837 7 1 2 60834 60836
0 60838 5 1 1 60837
0 60839 7 1 2 87495 107304
0 60840 7 1 2 60838 60839
0 60841 7 1 2 60832 60840
0 60842 5 1 1 60841
0 60843 7 1 2 72288 60842
0 60844 7 1 2 60826 60843
0 60845 7 1 2 60767 60844
0 60846 5 1 1 60845
0 60847 7 1 2 68736 60846
0 60848 7 1 2 60703 60847
0 60849 5 1 1 60848
0 60850 7 1 2 94663 93368
0 60851 5 1 1 60850
0 60852 7 1 2 99779 90610
0 60853 7 1 2 92468 60852
0 60854 5 1 1 60853
0 60855 7 1 2 60851 60854
0 60856 5 1 1 60855
0 60857 7 1 2 67245 60856
0 60858 5 1 1 60857
0 60859 7 1 2 101436 95624
0 60860 7 1 2 93321 91179
0 60861 7 1 2 60859 60860
0 60862 7 1 2 97181 60861
0 60863 5 1 1 60862
0 60864 7 1 2 60858 60863
0 60865 5 1 1 60864
0 60866 7 1 2 69673 60865
0 60867 5 1 1 60866
0 60868 7 1 2 81542 90608
0 60869 7 2 2 103351 60868
0 60870 7 1 2 99780 107124
0 60871 7 1 2 107326 60870
0 60872 5 1 1 60871
0 60873 7 1 2 60867 60872
0 60874 5 1 1 60873
0 60875 7 1 2 90130 60874
0 60876 5 1 1 60875
0 60877 7 1 2 102553 93311
0 60878 7 1 2 95731 60877
0 60879 7 1 2 106145 106492
0 60880 7 1 2 60878 60879
0 60881 5 1 1 60880
0 60882 7 1 2 60876 60881
0 60883 5 1 1 60882
0 60884 7 1 2 84883 60883
0 60885 5 1 1 60884
0 60886 7 1 2 80785 99659
0 60887 7 1 2 91383 60886
0 60888 5 1 1 60887
0 60889 7 1 2 70748 93244
0 60890 7 1 2 103145 74226
0 60891 7 1 2 60889 60890
0 60892 7 1 2 106433 60891
0 60893 5 1 1 60892
0 60894 7 1 2 60888 60893
0 60895 5 1 1 60894
0 60896 7 1 2 85969 60895
0 60897 5 1 1 60896
0 60898 7 1 2 76167 80214
0 60899 7 1 2 104159 60898
0 60900 7 1 2 95732 93363
0 60901 7 1 2 60899 60900
0 60902 5 1 1 60901
0 60903 7 1 2 60897 60902
0 60904 5 1 1 60903
0 60905 7 1 2 67834 60904
0 60906 5 1 1 60905
0 60907 7 2 2 72840 96620
0 60908 7 1 2 102554 93485
0 60909 7 1 2 101607 60908
0 60910 7 1 2 107328 60909
0 60911 5 1 1 60910
0 60912 7 1 2 60906 60911
0 60913 7 1 2 60885 60912
0 60914 5 1 1 60913
0 60915 7 1 2 70293 60914
0 60916 5 1 1 60915
0 60917 7 1 2 94664 106973
0 60918 7 1 2 106403 107308
0 60919 7 1 2 60917 60918
0 60920 5 1 1 60919
0 60921 7 2 2 103901 88930
0 60922 7 1 2 103352 105506
0 60923 7 1 2 107330 60922
0 60924 5 1 1 60923
0 60925 7 1 2 60920 60924
0 60926 5 1 1 60925
0 60927 7 1 2 81242 88280
0 60928 7 1 2 60926 60927
0 60929 5 1 1 60928
0 60930 7 1 2 84306 90427
0 60931 7 1 2 103893 60930
0 60932 7 1 2 103318 107323
0 60933 7 1 2 60931 60932
0 60934 5 1 1 60933
0 60935 7 1 2 60929 60934
0 60936 5 1 1 60935
0 60937 7 1 2 107103 60936
0 60938 5 1 1 60937
0 60939 7 2 2 93387 107138
0 60940 7 1 2 91384 107332
0 60941 5 1 1 60940
0 60942 7 1 2 60938 60941
0 60943 5 1 1 60942
0 60944 7 1 2 70571 60943
0 60945 5 1 1 60944
0 60946 7 1 2 101824 94088
0 60947 7 1 2 105518 60946
0 60948 5 1 1 60947
0 60949 7 1 2 8450 60948
0 60950 5 1 1 60949
0 60951 7 1 2 90554 60950
0 60952 5 1 1 60951
0 60953 7 1 2 103703 91620
0 60954 7 1 2 91574 60953
0 60955 5 1 1 60954
0 60956 7 1 2 60952 60955
0 60957 5 1 1 60956
0 60958 7 1 2 107333 60957
0 60959 5 1 1 60958
0 60960 7 1 2 60945 60959
0 60961 7 1 2 60916 60960
0 60962 5 1 1 60961
0 60963 7 1 2 72492 60962
0 60964 5 1 1 60963
0 60965 7 1 2 67835 94176
0 60966 7 1 2 103287 60965
0 60967 5 1 1 60966
0 60968 7 3 2 74444 96778
0 60969 7 1 2 91718 89872
0 60970 7 1 2 102824 60969
0 60971 7 1 2 107334 60970
0 60972 5 1 1 60971
0 60973 7 1 2 60967 60972
0 60974 5 1 1 60973
0 60975 7 1 2 86588 60974
0 60976 5 1 1 60975
0 60977 7 1 2 78543 104680
0 60978 7 1 2 83086 60977
0 60979 7 1 2 102522 60978
0 60980 5 1 1 60979
0 60981 7 1 2 60976 60980
0 60982 5 1 1 60981
0 60983 7 1 2 70294 60982
0 60984 5 1 1 60983
0 60985 7 1 2 69674 75513
0 60986 7 1 2 100965 60985
0 60987 7 1 2 101357 104899
0 60988 7 1 2 60986 60987
0 60989 5 1 1 60988
0 60990 7 2 2 102396 107104
0 60991 7 1 2 70572 103039
0 60992 7 1 2 107337 60991
0 60993 5 1 1 60992
0 60994 7 1 2 30678 60993
0 60995 5 1 1 60994
0 60996 7 1 2 70648 81939
0 60997 7 1 2 102120 60996
0 60998 7 1 2 60995 60997
0 60999 5 1 1 60998
0 61000 7 1 2 60989 60999
0 61001 5 1 1 61000
0 61002 7 1 2 63938 61001
0 61003 5 1 1 61002
0 61004 7 1 2 103284 105296
0 61005 5 1 1 61004
0 61006 7 1 2 96317 80215
0 61007 7 1 2 107338 61006
0 61008 5 1 1 61007
0 61009 7 1 2 61005 61008
0 61010 5 1 1 61009
0 61011 7 1 2 81940 107306
0 61012 7 1 2 61010 61011
0 61013 5 1 1 61012
0 61014 7 1 2 61003 61013
0 61015 5 1 1 61014
0 61016 7 1 2 68222 61015
0 61017 5 1 1 61016
0 61018 7 1 2 60984 61017
0 61019 5 1 1 61018
0 61020 7 1 2 63827 61019
0 61021 5 1 1 61020
0 61022 7 1 2 81941 102491
0 61023 5 1 1 61022
0 61024 7 1 2 99543 96452
0 61025 5 8 1 61024
0 61026 7 1 2 103250 107339
0 61027 5 1 1 61026
0 61028 7 1 2 61023 61027
0 61029 5 1 1 61028
0 61030 7 1 2 63939 61029
0 61031 5 1 1 61030
0 61032 7 3 2 72289 107340
0 61033 7 1 2 65659 84445
0 61034 7 1 2 107347 61033
0 61035 5 1 1 61034
0 61036 7 1 2 61031 61035
0 61037 5 1 1 61036
0 61038 7 1 2 101990 97467
0 61039 7 1 2 61037 61038
0 61040 5 1 1 61039
0 61041 7 1 2 61021 61040
0 61042 5 1 1 61041
0 61043 7 1 2 72200 61042
0 61044 5 1 1 61043
0 61045 7 1 2 80786 92846
0 61046 5 1 1 61045
0 61047 7 1 2 22158 61046
0 61048 5 1 1 61047
0 61049 7 2 2 98967 106836
0 61050 7 1 2 90899 93590
0 61051 7 1 2 107350 61050
0 61052 7 1 2 61048 61051
0 61053 5 1 1 61052
0 61054 7 1 2 66904 61053
0 61055 7 1 2 61044 61054
0 61056 5 1 1 61055
0 61057 7 1 2 81942 74481
0 61058 7 1 2 99213 61057
0 61059 5 1 1 61058
0 61060 7 1 2 97957 78367
0 61061 7 1 2 87675 61060
0 61062 5 1 1 61061
0 61063 7 1 2 61059 61062
0 61064 5 1 1 61063
0 61065 7 1 2 73294 61064
0 61066 5 2 1 61065
0 61067 7 1 2 68223 97108
0 61068 7 1 2 103367 61067
0 61069 7 1 2 86687 103329
0 61070 7 1 2 61068 61069
0 61071 5 1 1 61070
0 61072 7 1 2 107352 61071
0 61073 5 1 1 61072
0 61074 7 1 2 103073 61073
0 61075 5 1 1 61074
0 61076 7 1 2 98560 98905
0 61077 5 1 1 61076
0 61078 7 1 2 102297 61077
0 61079 5 1 1 61078
0 61080 7 1 2 65543 61079
0 61081 5 1 1 61080
0 61082 7 1 2 80304 97067
0 61083 7 1 2 103505 61082
0 61084 5 1 1 61083
0 61085 7 1 2 61081 61084
0 61086 5 1 1 61085
0 61087 7 1 2 102271 83107
0 61088 7 1 2 61086 61087
0 61089 5 1 1 61088
0 61090 7 1 2 61075 61089
0 61091 5 1 1 61090
0 61092 7 1 2 67146 61091
0 61093 5 1 1 61092
0 61094 7 1 2 82940 83123
0 61095 5 3 1 61094
0 61096 7 1 2 102304 107354
0 61097 5 1 1 61096
0 61098 7 1 2 65544 61097
0 61099 5 1 1 61098
0 61100 7 1 2 80305 90099
0 61101 5 1 1 61100
0 61102 7 1 2 61099 61101
0 61103 5 1 1 61102
0 61104 7 1 2 83885 104140
0 61105 7 1 2 98124 61104
0 61106 7 1 2 61103 61105
0 61107 5 1 1 61106
0 61108 7 1 2 61093 61107
0 61109 5 1 1 61108
0 61110 7 1 2 103018 61109
0 61111 5 1 1 61110
0 61112 7 2 2 67836 107341
0 61113 7 1 2 98619 107357
0 61114 5 1 1 61113
0 61115 7 1 2 34524 61114
0 61116 5 1 1 61115
0 61117 7 1 2 72069 102028
0 61118 7 1 2 104609 61117
0 61119 7 1 2 106579 61118
0 61120 7 1 2 61116 61119
0 61121 5 1 1 61120
0 61122 7 1 2 71971 61121
0 61123 7 1 2 61111 61122
0 61124 5 1 1 61123
0 61125 7 1 2 99371 61124
0 61126 7 1 2 61056 61125
0 61127 5 1 1 61126
0 61128 7 1 2 102137 95527
0 61129 7 1 2 75683 61128
0 61130 5 1 1 61129
0 61131 7 1 2 70930 93742
0 61132 7 1 2 103973 61131
0 61133 7 1 2 85368 61132
0 61134 5 1 1 61133
0 61135 7 1 2 61130 61134
0 61136 5 1 1 61135
0 61137 7 1 2 106948 61136
0 61138 5 1 1 61137
0 61139 7 1 2 102949 104822
0 61140 7 1 2 77761 61139
0 61141 7 1 2 107283 61140
0 61142 5 1 1 61141
0 61143 7 1 2 61138 61142
0 61144 5 1 1 61143
0 61145 7 1 2 72493 61144
0 61146 5 1 1 61145
0 61147 7 1 2 77913 102756
0 61148 7 1 2 103066 61147
0 61149 7 1 2 107292 61148
0 61150 7 1 2 106949 61149
0 61151 5 1 1 61150
0 61152 7 1 2 61146 61151
0 61153 5 1 1 61152
0 61154 7 1 2 67837 61153
0 61155 5 1 1 61154
0 61156 7 1 2 74445 100087
0 61157 5 1 1 61156
0 61158 7 1 2 104841 61157
0 61159 5 1 1 61158
0 61160 7 1 2 72201 106950
0 61161 7 4 2 61159 61160
0 61162 7 1 2 82253 107154
0 61163 7 1 2 107359 61162
0 61164 5 1 1 61163
0 61165 7 1 2 61155 61164
0 61166 5 1 1 61165
0 61167 7 1 2 68737 61166
0 61168 5 1 1 61167
0 61169 7 1 2 102555 97087
0 61170 7 1 2 102993 61169
0 61171 5 1 1 61170
0 61172 7 2 2 82512 100440
0 61173 5 1 1 107363
0 61174 7 1 2 84689 107364
0 61175 5 1 1 61174
0 61176 7 2 2 69675 72290
0 61177 7 1 2 101097 107365
0 61178 5 1 1 61177
0 61179 7 1 2 61175 61178
0 61180 5 1 1 61179
0 61181 7 1 2 76923 107157
0 61182 7 1 2 61180 61181
0 61183 5 1 1 61182
0 61184 7 1 2 61171 61183
0 61185 5 1 1 61184
0 61186 7 1 2 84884 61185
0 61187 5 1 1 61186
0 61188 7 1 2 102731 97485
0 61189 7 1 2 85383 61188
0 61190 7 1 2 102994 61189
0 61191 5 1 1 61190
0 61192 7 1 2 61187 61191
0 61193 5 1 1 61192
0 61194 7 1 2 70295 61193
0 61195 5 1 1 61194
0 61196 7 1 2 98883 106762
0 61197 7 2 2 97135 95295
0 61198 7 1 2 107189 107367
0 61199 7 1 2 61196 61198
0 61200 5 1 1 61199
0 61201 7 1 2 61195 61200
0 61202 7 1 2 61168 61201
0 61203 5 1 1 61202
0 61204 7 1 2 67015 61203
0 61205 5 1 1 61204
0 61206 7 2 2 74414 102507
0 61207 5 3 1 107369
0 61208 7 1 2 99660 107000
0 61209 5 1 1 61208
0 61210 7 1 2 107371 61209
0 61211 5 1 1 61210
0 61212 7 1 2 102121 77785
0 61213 7 2 2 61211 61212
0 61214 7 1 2 75169 107374
0 61215 5 1 1 61214
0 61216 7 1 2 63828 61215
0 61217 7 1 2 61205 61216
0 61218 5 1 1 61217
0 61219 7 4 2 72070 94238
0 61220 7 1 2 83278 107376
0 61221 5 1 1 61220
0 61222 7 1 2 82829 104863
0 61223 5 1 1 61222
0 61224 7 1 2 61221 61223
0 61225 5 1 1 61224
0 61226 7 1 2 71876 61225
0 61227 5 1 1 61226
0 61228 7 1 2 85603 107377
0 61229 5 1 1 61228
0 61230 7 1 2 61227 61229
0 61231 5 1 1 61230
0 61232 7 1 2 70573 61231
0 61233 5 1 1 61232
0 61234 7 1 2 96621 107378
0 61235 5 1 1 61234
0 61236 7 1 2 94487 83022
0 61237 5 1 1 61236
0 61238 7 1 2 61235 61237
0 61239 5 1 1 61238
0 61240 7 1 2 70296 61239
0 61241 5 1 1 61240
0 61242 7 1 2 72071 102365
0 61243 7 1 2 105519 61242
0 61244 5 1 1 61243
0 61245 7 1 2 61241 61244
0 61246 7 1 2 61233 61245
0 61247 5 1 1 61246
0 61248 7 1 2 97068 61247
0 61249 5 1 1 61248
0 61250 7 1 2 84945 85838
0 61251 7 1 2 100988 61250
0 61252 5 1 1 61251
0 61253 7 1 2 61249 61252
0 61254 5 1 1 61253
0 61255 7 1 2 99661 61254
0 61256 5 1 1 61255
0 61257 7 1 2 106924 60260
0 61258 5 1 1 61257
0 61259 7 1 2 82830 97088
0 61260 7 1 2 61258 61259
0 61261 5 1 1 61260
0 61262 7 1 2 107353 61261
0 61263 5 1 1 61262
0 61264 7 1 2 106668 61263
0 61265 5 1 1 61264
0 61266 7 1 2 61256 61265
0 61267 5 1 1 61266
0 61268 7 1 2 77639 61267
0 61269 5 1 1 61268
0 61270 7 1 2 76924 107375
0 61271 5 1 1 61270
0 61272 7 1 2 68897 61271
0 61273 7 1 2 61269 61272
0 61274 5 1 1 61273
0 61275 7 1 2 73884 61274
0 61276 7 1 2 61218 61275
0 61277 5 1 1 61276
0 61278 7 1 2 94737 106669
0 61279 7 1 2 107368 61278
0 61280 7 1 2 95947 61279
0 61281 5 1 1 61280
0 61282 7 1 2 101437 81445
0 61283 7 1 2 102349 61282
0 61284 7 1 2 95579 61283
0 61285 5 1 1 61284
0 61286 7 1 2 61281 61285
0 61287 5 1 1 61286
0 61288 7 1 2 65237 61287
0 61289 5 1 1 61288
0 61290 7 1 2 88696 91476
0 61291 7 1 2 107370 61290
0 61292 5 1 1 61291
0 61293 7 1 2 95577 101867
0 61294 7 1 2 106905 61293
0 61295 5 1 1 61294
0 61296 7 1 2 61292 61295
0 61297 5 1 1 61296
0 61298 7 1 2 70297 61297
0 61299 5 1 1 61298
0 61300 7 1 2 80665 106678
0 61301 5 1 1 61300
0 61302 7 1 2 107372 61301
0 61303 5 1 1 61302
0 61304 7 1 2 90629 61303
0 61305 5 1 1 61304
0 61306 7 1 2 61299 61305
0 61307 5 1 1 61306
0 61308 7 1 2 97089 61307
0 61309 5 1 1 61308
0 61310 7 1 2 61289 61309
0 61311 5 1 1 61310
0 61312 7 1 2 89591 61311
0 61313 5 1 1 61312
0 61314 7 1 2 80666 99662
0 61315 5 2 1 61314
0 61316 7 1 2 107373 107380
0 61317 5 1 1 61316
0 61318 7 1 2 92485 61317
0 61319 5 1 1 61318
0 61320 7 1 2 70931 99541
0 61321 5 1 1 61320
0 61322 7 1 2 80787 99946
0 61323 5 1 1 61322
0 61324 7 1 2 61321 61323
0 61325 5 3 1 61324
0 61326 7 1 2 89008 107366
0 61327 7 1 2 107382 61326
0 61328 5 1 1 61327
0 61329 7 1 2 67246 86355
0 61330 7 1 2 82780 61329
0 61331 7 2 2 81807 107083
0 61332 7 1 2 88045 107385
0 61333 7 1 2 61330 61332
0 61334 5 1 1 61333
0 61335 7 1 2 61328 61334
0 61336 5 1 1 61335
0 61337 7 1 2 85352 61336
0 61338 5 1 1 61337
0 61339 7 1 2 61319 61338
0 61340 5 1 1 61339
0 61341 7 1 2 72841 61340
0 61342 5 1 1 61341
0 61343 7 7 2 64001 72291
0 61344 5 1 1 107387
0 61345 7 1 2 107327 107388
0 61346 7 1 2 107383 61345
0 61347 5 1 1 61346
0 61348 7 1 2 61342 61347
0 61349 5 1 1 61348
0 61350 7 1 2 88281 61349
0 61351 5 1 1 61350
0 61352 7 1 2 95564 95697
0 61353 5 1 1 61352
0 61354 7 1 2 69327 96520
0 61355 7 1 2 105147 61354
0 61356 5 1 1 61355
0 61357 7 1 2 61353 61356
0 61358 5 1 1 61357
0 61359 7 1 2 99135 103343
0 61360 7 1 2 88637 61359
0 61361 7 1 2 84918 61360
0 61362 7 1 2 61358 61361
0 61363 5 1 1 61362
0 61364 7 1 2 61351 61363
0 61365 5 1 1 61364
0 61366 7 1 2 97136 61365
0 61367 5 1 1 61366
0 61368 7 1 2 61313 61367
0 61369 7 1 2 61277 61368
0 61370 7 1 2 61127 61369
0 61371 7 1 2 60964 61370
0 61372 7 1 2 60849 61371
0 61373 7 1 2 60579 61372
0 61374 5 1 1 61373
0 61375 7 1 2 96260 61374
0 61376 5 1 1 61375
0 61377 7 1 2 102829 107342
0 61378 5 1 1 61377
0 61379 7 1 2 100291 81243
0 61380 7 1 2 106962 61379
0 61381 5 1 1 61380
0 61382 7 1 2 61378 61381
0 61383 5 1 1 61382
0 61384 7 1 2 72842 61383
0 61385 5 1 1 61384
0 61386 7 1 2 84512 104890
0 61387 7 1 2 101810 61386
0 61388 5 1 1 61387
0 61389 7 1 2 61385 61388
0 61390 5 1 1 61389
0 61391 7 1 2 97000 61390
0 61392 5 1 1 61391
0 61393 7 1 2 60073 107355
0 61394 5 1 1 61393
0 61395 7 1 2 96984 61394
0 61396 5 1 1 61395
0 61397 7 1 2 69328 86533
0 61398 7 1 2 104631 61397
0 61399 5 1 1 61398
0 61400 7 1 2 61396 61399
0 61401 5 1 1 61400
0 61402 7 2 2 97238 103335
0 61403 7 1 2 65545 107394
0 61404 7 1 2 61401 61403
0 61405 5 1 1 61404
0 61406 7 1 2 61392 61405
0 61407 5 1 1 61406
0 61408 7 1 2 68898 61407
0 61409 5 1 1 61408
0 61410 7 2 2 68224 107343
0 61411 7 1 2 95542 97001
0 61412 7 1 2 104325 61411
0 61413 7 1 2 107396 61412
0 61414 5 1 1 61413
0 61415 7 1 2 61409 61414
0 61416 5 1 1 61415
0 61417 7 1 2 106974 61416
0 61418 5 1 1 61417
0 61419 7 2 2 73295 107344
0 61420 7 1 2 107398 107395
0 61421 5 1 1 61420
0 61422 7 1 2 102830 105069
0 61423 5 1 1 61422
0 61424 7 1 2 61421 61423
0 61425 5 1 1 61424
0 61426 7 1 2 96985 61425
0 61427 5 1 1 61426
0 61428 7 2 2 70298 83712
0 61429 5 1 1 107400
0 61430 7 1 2 103125 61429
0 61431 5 1 1 61430
0 61432 7 1 2 100292 106626
0 61433 7 1 2 61431 61432
0 61434 5 1 1 61433
0 61435 7 1 2 61427 61434
0 61436 5 1 1 61435
0 61437 7 1 2 68899 61436
0 61438 5 1 1 61437
0 61439 7 2 2 81943 104326
0 61440 7 1 2 96986 104676
0 61441 7 1 2 107402 61440
0 61442 5 1 1 61441
0 61443 7 1 2 61438 61442
0 61444 5 1 1 61443
0 61445 7 1 2 107125 61444
0 61446 5 1 1 61445
0 61447 7 1 2 61418 61446
0 61448 5 1 1 61447
0 61449 7 1 2 71217 61448
0 61450 5 1 1 61449
0 61451 7 4 2 64534 107105
0 61452 5 1 1 107404
0 61453 7 1 2 70574 105608
0 61454 7 1 2 107405 61453
0 61455 5 1 1 61454
0 61456 7 1 2 96446 81489
0 61457 7 1 2 97002 61456
0 61458 5 1 1 61457
0 61459 7 1 2 61455 61458
0 61460 5 1 1 61459
0 61461 7 1 2 68225 103883
0 61462 7 2 2 61460 61461
0 61463 7 1 2 63829 104327
0 61464 5 1 1 61463
0 61465 7 1 2 25507 61464
0 61466 5 4 1 61465
0 61467 7 1 2 69079 107410
0 61468 7 1 2 107408 61467
0 61469 5 1 1 61468
0 61470 7 1 2 61450 61469
0 61471 5 1 1 61470
0 61472 7 1 2 70749 61471
0 61473 5 1 1 61472
0 61474 7 1 2 103135 88931
0 61475 7 1 2 107409 61474
0 61476 5 1 1 61475
0 61477 7 1 2 61473 61476
0 61478 5 1 1 61477
0 61479 7 1 2 76523 61478
0 61480 5 1 1 61479
0 61481 7 4 2 66905 107411
0 61482 7 2 2 88646 107414
0 61483 5 1 1 107418
0 61484 7 1 2 94593 88652
0 61485 7 1 2 97708 61484
0 61486 5 1 1 61485
0 61487 7 1 2 61483 61486
0 61488 5 1 1 61487
0 61489 7 1 2 96943 61488
0 61490 5 1 1 61489
0 61491 7 1 2 84947 102432
0 61492 7 1 2 102473 61491
0 61493 7 1 2 104904 106580
0 61494 7 1 2 61492 61493
0 61495 5 1 1 61494
0 61496 7 1 2 61490 61495
0 61497 5 1 1 61496
0 61498 7 1 2 71218 61497
0 61499 5 1 1 61498
0 61500 7 1 2 103616 107419
0 61501 5 1 1 61500
0 61502 7 1 2 61499 61501
0 61503 5 1 1 61502
0 61504 7 1 2 76524 61503
0 61505 5 1 1 61504
0 61506 7 1 2 34545 18987
0 61507 5 1 1 61506
0 61508 7 1 2 83915 103273
0 61509 7 1 2 61507 61508
0 61510 7 1 2 107415 61509
0 61511 5 1 1 61510
0 61512 7 1 2 61505 61511
0 61513 5 1 1 61512
0 61514 7 1 2 89524 61513
0 61515 5 1 1 61514
0 61516 7 1 2 98620 90821
0 61517 5 1 1 61516
0 61518 7 1 2 76254 97756
0 61519 5 1 1 61518
0 61520 7 1 2 61517 61519
0 61521 5 1 1 61520
0 61522 7 1 2 83916 91257
0 61523 7 1 2 106789 61522
0 61524 7 1 2 103136 61523
0 61525 7 1 2 61521 61524
0 61526 5 1 1 61525
0 61527 7 1 2 61515 61526
0 61528 5 1 1 61527
0 61529 7 1 2 72292 61528
0 61530 5 1 1 61529
0 61531 7 1 2 99696 106623
0 61532 5 1 1 61531
0 61533 7 1 2 84533 104787
0 61534 5 1 1 61533
0 61535 7 1 2 61532 61534
0 61536 5 1 1 61535
0 61537 7 1 2 78750 74090
0 61538 7 1 2 103252 107126
0 61539 7 1 2 61537 61538
0 61540 7 1 2 93632 61539
0 61541 7 1 2 61536 61540
0 61542 5 1 1 61541
0 61543 7 1 2 61530 61542
0 61544 5 1 1 61543
0 61545 7 1 2 84885 61544
0 61546 5 1 1 61545
0 61547 7 1 2 80874 103712
0 61548 5 1 1 61547
0 61549 7 2 2 96447 90869
0 61550 7 1 2 72494 107420
0 61551 5 1 1 61550
0 61552 7 1 2 61548 61551
0 61553 5 2 1 61552
0 61554 7 1 2 69329 107422
0 61555 7 1 2 105358 61554
0 61556 5 1 1 61555
0 61557 7 1 2 98700 80216
0 61558 7 1 2 74047 61557
0 61559 7 1 2 107295 61558
0 61560 7 1 2 107406 61559
0 61561 5 1 1 61560
0 61562 7 1 2 61556 61561
0 61563 5 1 1 61562
0 61564 7 1 2 80048 103884
0 61565 7 1 2 61563 61564
0 61566 5 1 1 61565
0 61567 7 1 2 61546 61566
0 61568 7 1 2 61480 61567
0 61569 5 1 1 61568
0 61570 7 1 2 70932 61569
0 61571 5 1 1 61570
0 61572 7 2 2 64002 102508
0 61573 5 1 1 107424
0 61574 7 1 2 106975 107001
0 61575 5 1 1 61574
0 61576 7 1 2 61573 61575
0 61577 5 1 1 61576
0 61578 7 1 2 66094 61577
0 61579 5 1 1 61578
0 61580 7 1 2 80875 96515
0 61581 7 1 2 107273 61580
0 61582 5 1 1 61581
0 61583 7 1 2 61579 61582
0 61584 5 1 1 61583
0 61585 7 1 2 96779 61584
0 61586 5 1 1 61585
0 61587 7 1 2 104141 106976
0 61588 7 1 2 100737 61587
0 61589 5 1 1 61588
0 61590 7 1 2 61586 61589
0 61591 5 1 1 61590
0 61592 7 1 2 65702 61591
0 61593 5 1 1 61592
0 61594 7 1 2 100099 61452
0 61595 5 1 1 61594
0 61596 7 1 2 96780 61595
0 61597 5 1 1 61596
0 61598 7 1 2 84746 97077
0 61599 5 1 1 61598
0 61600 7 1 2 61597 61599
0 61601 5 1 1 61600
0 61602 7 1 2 70575 61601
0 61603 5 1 1 61602
0 61604 7 2 2 85599 96453
0 61605 5 5 1 107426
0 61606 7 1 2 80556 98391
0 61607 5 1 1 61606
0 61608 7 1 2 97079 61607
0 61609 5 1 1 61608
0 61610 7 1 2 107428 61609
0 61611 5 1 1 61610
0 61612 7 1 2 61603 61611
0 61613 5 1 1 61612
0 61614 7 1 2 107014 61613
0 61615 5 1 1 61614
0 61616 7 1 2 61593 61615
0 61617 5 1 1 61616
0 61618 7 1 2 76255 61617
0 61619 5 1 1 61618
0 61620 7 1 2 81490 107429
0 61621 5 1 1 61620
0 61622 7 1 2 84003 88881
0 61623 5 1 1 61622
0 61624 7 1 2 80876 105190
0 61625 5 1 1 61624
0 61626 7 1 2 61623 61625
0 61627 5 1 1 61626
0 61628 7 1 2 70576 61627
0 61629 5 1 1 61628
0 61630 7 1 2 61621 61629
0 61631 5 1 1 61630
0 61632 7 1 2 99277 103248
0 61633 7 1 2 99372 61632
0 61634 7 1 2 61631 61633
0 61635 5 1 1 61634
0 61636 7 1 2 61619 61635
0 61637 5 1 1 61636
0 61638 7 1 2 64226 61637
0 61639 5 1 1 61638
0 61640 7 3 2 72843 100143
0 61641 7 1 2 76525 107224
0 61642 5 1 1 61641
0 61643 7 1 2 82532 107222
0 61644 5 1 1 61643
0 61645 7 1 2 61642 61644
0 61646 5 1 1 61645
0 61647 7 1 2 96448 61646
0 61648 5 1 1 61647
0 61649 7 1 2 77276 107106
0 61650 5 1 1 61649
0 61651 7 1 2 100100 61650
0 61652 5 1 1 61651
0 61653 7 1 2 70577 61652
0 61654 5 1 1 61653
0 61655 7 1 2 66095 80557
0 61656 5 1 1 61655
0 61657 7 1 2 61654 61656
0 61658 5 1 1 61657
0 61659 7 1 2 99269 91714
0 61660 7 1 2 61658 61659
0 61661 5 1 1 61660
0 61662 7 1 2 61648 61661
0 61663 5 1 1 61662
0 61664 7 1 2 65703 61663
0 61665 5 1 1 61664
0 61666 7 1 2 99351 99270
0 61667 7 1 2 103654 61666
0 61668 7 1 2 94209 61667
0 61669 5 1 1 61668
0 61670 7 1 2 61665 61669
0 61671 5 1 1 61670
0 61672 7 1 2 107433 61671
0 61673 5 1 1 61672
0 61674 7 1 2 61639 61673
0 61675 5 1 1 61674
0 61676 7 1 2 103137 61675
0 61677 5 1 1 61676
0 61678 7 1 2 70750 91344
0 61679 7 1 2 77815 61678
0 61680 7 1 2 106475 107434
0 61681 7 1 2 61679 61680
0 61682 7 1 2 107412 61681
0 61683 5 1 1 61682
0 61684 7 1 2 61677 61683
0 61685 5 1 1 61684
0 61686 7 1 2 68226 84229
0 61687 7 1 2 61685 61686
0 61688 5 1 1 61687
0 61689 7 1 2 72202 61688
0 61690 7 1 2 61571 61689
0 61691 5 1 1 61690
0 61692 7 1 2 91352 107146
0 61693 7 1 2 107159 61692
0 61694 5 1 1 61693
0 61695 7 1 2 87813 103146
0 61696 7 1 2 103985 61695
0 61697 7 1 2 91699 93491
0 61698 7 1 2 61696 61697
0 61699 5 1 1 61698
0 61700 7 1 2 61694 61699
0 61701 5 1 1 61700
0 61702 7 1 2 96944 61701
0 61703 5 1 1 61702
0 61704 7 1 2 69080 22402
0 61705 5 1 1 61704
0 61706 7 1 2 84690 61344
0 61707 7 2 2 61705 61706
0 61708 7 1 2 70751 93564
0 61709 7 1 2 102475 61708
0 61710 7 1 2 107436 61709
0 61711 5 1 1 61710
0 61712 7 1 2 61703 61711
0 61713 5 1 1 61712
0 61714 7 1 2 63940 61713
0 61715 5 1 1 61714
0 61716 7 1 2 96987 107437
0 61717 5 1 1 61716
0 61718 7 1 2 64535 106790
0 61719 7 1 2 104934 61718
0 61720 5 1 1 61719
0 61721 7 1 2 61717 61720
0 61722 5 1 1 61721
0 61723 7 1 2 73811 106907
0 61724 5 1 1 61723
0 61725 7 2 2 59480 61724
0 61726 5 2 1 107438
0 61727 7 1 2 101647 107440
0 61728 7 1 2 61722 61727
0 61729 5 1 1 61728
0 61730 7 1 2 61715 61729
0 61731 5 1 1 61730
0 61732 7 1 2 81944 61731
0 61733 5 1 1 61732
0 61734 7 1 2 96945 107002
0 61735 5 2 1 61734
0 61736 7 1 2 67492 85379
0 61737 5 1 1 61736
0 61738 7 1 2 107442 61737
0 61739 5 1 1 61738
0 61740 7 1 2 69030 107439
0 61741 5 1 1 61740
0 61742 7 2 2 99745 91624
0 61743 5 1 1 107444
0 61744 7 1 2 63941 61743
0 61745 5 1 1 61744
0 61746 7 1 2 75865 106977
0 61747 7 1 2 106245 61746
0 61748 7 1 2 61745 61747
0 61749 7 1 2 61741 61748
0 61750 7 1 2 61739 61749
0 61751 5 1 1 61750
0 61752 7 1 2 61733 61751
0 61753 5 1 1 61752
0 61754 7 1 2 68900 61753
0 61755 5 1 1 61754
0 61756 7 1 2 101285 105793
0 61757 5 1 1 61756
0 61758 7 1 2 65616 107445
0 61759 5 1 1 61758
0 61760 7 1 2 61757 61759
0 61761 5 1 1 61760
0 61762 7 1 2 63942 61761
0 61763 5 1 1 61762
0 61764 7 1 2 78085 107441
0 61765 5 1 1 61764
0 61766 7 1 2 61763 61765
0 61767 5 1 1 61766
0 61768 7 1 2 103344 95852
0 61769 7 1 2 106446 61768
0 61770 7 1 2 61767 61769
0 61771 5 1 1 61770
0 61772 7 1 2 67147 61771
0 61773 7 1 2 61755 61772
0 61774 5 1 1 61773
0 61775 7 1 2 72072 61774
0 61776 7 1 2 61691 61775
0 61777 5 1 1 61776
0 61778 7 2 2 69330 97445
0 61779 7 1 2 102509 89551
0 61780 7 2 2 107446 61779
0 61781 5 1 1 107448
0 61782 7 3 2 64227 100441
0 61783 5 3 1 107450
0 61784 7 1 2 23349 107453
0 61785 5 3 1 61784
0 61786 7 1 2 70299 87195
0 61787 5 1 1 61786
0 61788 7 1 2 106925 61787
0 61789 5 1 1 61788
0 61790 7 1 2 107456 61789
0 61791 5 1 1 61790
0 61792 7 1 2 104387 107451
0 61793 5 1 1 61792
0 61794 7 1 2 61791 61793
0 61795 5 1 1 61794
0 61796 7 1 2 96437 61795
0 61797 5 1 1 61796
0 61798 7 2 2 100144 97211
0 61799 5 1 1 107459
0 61800 7 1 2 107454 61799
0 61801 5 1 1 61800
0 61802 7 1 2 81945 61801
0 61803 5 1 1 61802
0 61804 7 1 2 100145 101062
0 61805 5 1 1 61804
0 61806 7 1 2 61803 61805
0 61807 5 1 1 61806
0 61808 7 1 2 96282 61807
0 61809 5 1 1 61808
0 61810 7 1 2 61797 61809
0 61811 5 1 1 61810
0 61812 7 1 2 70752 61811
0 61813 5 1 1 61812
0 61814 7 1 2 61781 61813
0 61815 5 1 1 61814
0 61816 7 1 2 73296 61815
0 61817 5 1 1 61816
0 61818 7 1 2 82941 89399
0 61819 7 1 2 105780 61818
0 61820 7 1 2 107457 61819
0 61821 5 1 1 61820
0 61822 7 1 2 61817 61821
0 61823 5 1 1 61822
0 61824 7 1 2 69081 61823
0 61825 5 1 1 61824
0 61826 7 1 2 96266 73812
0 61827 7 1 2 102510 61826
0 61828 5 1 1 61827
0 61829 7 1 2 73813 107274
0 61830 5 1 1 61829
0 61831 7 1 2 70694 60547
0 61832 5 1 1 61831
0 61833 7 1 2 65660 59383
0 61834 5 1 1 61833
0 61835 7 1 2 81946 61834
0 61836 7 1 2 61832 61835
0 61837 5 1 1 61836
0 61838 7 1 2 61830 61837
0 61839 5 2 1 61838
0 61840 7 1 2 102323 107461
0 61841 5 1 1 61840
0 61842 7 1 2 61828 61841
0 61843 5 1 1 61842
0 61844 7 1 2 107317 61843
0 61845 5 1 1 61844
0 61846 7 1 2 61825 61845
0 61847 5 1 1 61846
0 61848 7 1 2 69031 61847
0 61849 5 1 1 61848
0 61850 7 1 2 107059 107252
0 61851 5 1 1 61850
0 61852 7 1 2 102324 61851
0 61853 5 1 1 61852
0 61854 7 1 2 70753 107452
0 61855 5 1 1 61854
0 61856 7 1 2 61853 61855
0 61857 5 1 1 61856
0 61858 7 1 2 69082 61857
0 61859 5 1 1 61858
0 61860 7 2 2 69331 99352
0 61861 7 1 2 103297 107463
0 61862 5 1 1 61861
0 61863 7 1 2 61859 61862
0 61864 5 1 1 61863
0 61865 7 1 2 81947 61864
0 61866 5 1 1 61865
0 61867 7 1 2 102325 107256
0 61868 5 1 1 61867
0 61869 7 1 2 61866 61868
0 61870 5 1 1 61869
0 61871 7 1 2 78727 106278
0 61872 7 1 2 61870 61871
0 61873 5 1 1 61872
0 61874 7 1 2 61849 61873
0 61875 5 1 1 61874
0 61876 7 1 2 96521 61875
0 61877 5 1 1 61876
0 61878 7 1 2 93852 89552
0 61879 7 1 2 93652 61878
0 61880 7 1 2 106887 107229
0 61881 7 1 2 61879 61880
0 61882 5 1 1 61881
0 61883 7 1 2 67838 61882
0 61884 7 1 2 61877 61883
0 61885 5 1 1 61884
0 61886 7 1 2 102487 102865
0 61887 7 1 2 89221 61886
0 61888 5 1 1 61887
0 61889 7 1 2 96593 107458
0 61890 5 1 1 61889
0 61891 7 4 2 72495 104823
0 61892 7 1 2 86907 107465
0 61893 5 1 1 61892
0 61894 7 1 2 61890 61893
0 61895 5 1 1 61894
0 61896 7 1 2 65238 96438
0 61897 7 1 2 61895 61896
0 61898 5 1 1 61897
0 61899 7 1 2 61888 61898
0 61900 5 1 1 61899
0 61901 7 1 2 70754 61900
0 61902 5 1 1 61901
0 61903 7 1 2 73297 107449
0 61904 5 1 1 61903
0 61905 7 1 2 61902 61904
0 61906 5 1 1 61905
0 61907 7 1 2 69083 61906
0 61908 5 1 1 61907
0 61909 7 1 2 67493 78728
0 61910 7 1 2 106791 61909
0 61911 7 1 2 107462 61910
0 61912 5 1 1 61911
0 61913 7 1 2 61908 61912
0 61914 5 1 1 61913
0 61915 7 1 2 69032 61914
0 61916 5 1 1 61915
0 61917 7 1 2 106279 107447
0 61918 7 1 2 107258 61917
0 61919 5 1 1 61918
0 61920 7 1 2 61916 61919
0 61921 5 1 1 61920
0 61922 7 1 2 69676 72073
0 61923 7 1 2 61921 61922
0 61924 5 1 1 61923
0 61925 7 1 2 101084 105813
0 61926 7 1 2 106392 106837
0 61927 7 1 2 61925 61926
0 61928 5 1 1 61927
0 61929 7 1 2 97958 100146
0 61930 5 1 1 61929
0 61931 7 1 2 107455 61930
0 61932 5 1 1 61931
0 61933 7 1 2 84886 61932
0 61934 5 1 1 61933
0 61935 7 1 2 83708 107466
0 61936 5 1 1 61935
0 61937 7 1 2 81808 107460
0 61938 5 1 1 61937
0 61939 7 1 2 61936 61938
0 61940 7 1 2 61934 61939
0 61941 5 1 1 61940
0 61942 7 1 2 91180 74300
0 61943 7 1 2 107302 61942
0 61944 7 1 2 61941 61943
0 61945 5 1 1 61944
0 61946 7 1 2 61928 61945
0 61947 5 1 1 61946
0 61948 7 1 2 69084 61947
0 61949 5 1 1 61948
0 61950 7 1 2 84779 100093
0 61951 5 1 1 61950
0 61952 7 1 2 84758 107467
0 61953 5 1 1 61952
0 61954 7 1 2 96267 102825
0 61955 5 1 1 61954
0 61956 7 1 2 61953 61955
0 61957 5 1 1 61956
0 61958 7 1 2 65546 61957
0 61959 5 1 1 61958
0 61960 7 1 2 61951 61959
0 61961 5 1 1 61960
0 61962 7 1 2 65704 61961
0 61963 5 1 1 61962
0 61964 7 1 2 102813 107386
0 61965 5 1 1 61964
0 61966 7 1 2 61963 61965
0 61967 5 1 1 61966
0 61968 7 2 2 100812 99016
0 61969 7 1 2 64003 107469
0 61970 7 1 2 61967 61969
0 61971 5 1 1 61970
0 61972 7 1 2 61949 61971
0 61973 5 1 1 61972
0 61974 7 1 2 70300 61973
0 61975 5 1 1 61974
0 61976 7 1 2 99635 107133
0 61977 5 1 1 61976
0 61978 7 1 2 102328 107064
0 61979 5 1 1 61978
0 61980 7 1 2 16808 60545
0 61981 5 1 1 61980
0 61982 7 1 2 64004 61981
0 61983 7 1 2 61979 61982
0 61984 5 1 1 61983
0 61985 7 1 2 61977 61984
0 61986 5 1 1 61985
0 61987 7 1 2 106920 107470
0 61988 7 1 2 61986 61987
0 61989 5 1 1 61988
0 61990 7 1 2 72844 61989
0 61991 7 1 2 61975 61990
0 61992 7 1 2 61924 61991
0 61993 5 1 1 61992
0 61994 7 1 2 68901 61993
0 61995 7 1 2 61885 61994
0 61996 5 1 1 61995
0 61997 7 1 2 74014 61996
0 61998 5 1 1 61997
0 61999 7 1 2 65239 88661
0 62000 5 2 1 61999
0 62001 7 1 2 85037 107038
0 62002 5 1 1 62001
0 62003 7 1 2 107471 62002
0 62004 5 1 1 62003
0 62005 7 1 2 107468 62004
0 62006 5 1 1 62005
0 62007 7 1 2 99081 107435
0 62008 7 1 2 107277 62007
0 62009 5 1 1 62008
0 62010 7 1 2 62006 62009
0 62011 5 1 1 62010
0 62012 7 1 2 96331 62011
0 62013 5 1 1 62012
0 62014 7 2 2 103298 102488
0 62015 5 1 1 107473
0 62016 7 1 2 80549 107474
0 62017 5 1 1 62016
0 62018 7 2 2 72496 103237
0 62019 7 1 2 70695 107475
0 62020 7 1 2 106951 62019
0 62021 5 1 1 62020
0 62022 7 1 2 62017 62021
0 62023 5 1 1 62022
0 62024 7 1 2 69033 62023
0 62025 5 1 1 62024
0 62026 7 1 2 63943 99571
0 62027 7 1 2 101755 103299
0 62028 7 1 2 62026 62027
0 62029 5 1 1 62028
0 62030 7 1 2 62025 62029
0 62031 5 1 1 62030
0 62032 7 1 2 99373 104882
0 62033 7 1 2 62031 62032
0 62034 5 1 1 62033
0 62035 7 1 2 62013 62034
0 62036 5 1 1 62035
0 62037 7 1 2 74106 62036
0 62038 5 1 1 62037
0 62039 7 1 2 79006 62038
0 62040 5 1 1 62039
0 62041 7 1 2 71972 62040
0 62042 7 1 2 61998 62041
0 62043 5 1 1 62042
0 62044 7 1 2 103138 77786
0 62045 5 1 1 62044
0 62046 7 1 2 94594 78729
0 62047 7 1 2 97259 62046
0 62048 5 1 1 62047
0 62049 7 1 2 62045 62048
0 62050 5 1 1 62049
0 62051 7 1 2 72845 62050
0 62052 5 1 1 62051
0 62053 7 1 2 78730 103336
0 62054 7 1 2 94977 62053
0 62055 5 1 1 62054
0 62056 7 1 2 62052 62055
0 62057 5 1 1 62056
0 62058 7 1 2 107476 62057
0 62059 5 1 1 62058
0 62060 7 1 2 101079 92149
0 62061 7 2 2 71973 102699
0 62062 7 1 2 105284 107477
0 62063 7 1 2 62060 62062
0 62064 5 1 1 62063
0 62065 7 1 2 62059 62064
0 62066 5 1 1 62065
0 62067 7 1 2 72074 62066
0 62068 5 1 1 62067
0 62069 7 3 2 88901 107117
0 62070 7 1 2 107351 107479
0 62071 5 1 1 62070
0 62072 7 1 2 62068 62071
0 62073 5 1 1 62072
0 62074 7 1 2 99374 62073
0 62075 5 1 1 62074
0 62076 7 1 2 102194 95470
0 62077 7 2 2 66906 74107
0 62078 7 1 2 91545 107482
0 62079 7 1 2 62076 62078
0 62080 5 1 1 62079
0 62081 7 1 2 62075 62080
0 62082 5 1 1 62081
0 62083 7 1 2 107003 62082
0 62084 5 1 1 62083
0 62085 7 1 2 106952 107243
0 62086 7 1 2 96375 62085
0 62087 5 1 1 62086
0 62088 7 1 2 65661 89873
0 62089 7 1 2 99375 62088
0 62090 7 1 2 84887 107245
0 62091 7 1 2 62089 62090
0 62092 5 1 1 62091
0 62093 7 1 2 62087 62092
0 62094 5 1 1 62093
0 62095 7 1 2 68738 62094
0 62096 5 1 1 62095
0 62097 7 2 2 84888 96376
0 62098 7 1 2 84037 107241
0 62099 7 1 2 107484 62098
0 62100 5 1 1 62099
0 62101 7 1 2 62096 62100
0 62102 5 1 1 62101
0 62103 7 1 2 91075 62102
0 62104 5 1 1 62103
0 62105 7 1 2 89525 107348
0 62106 5 1 1 62105
0 62107 7 1 2 60527 62106
0 62108 5 1 1 62107
0 62109 7 1 2 93743 96501
0 62110 7 1 2 103731 62109
0 62111 7 1 2 62108 62110
0 62112 5 1 1 62111
0 62113 7 1 2 62104 62112
0 62114 5 1 1 62113
0 62115 7 1 2 79648 62114
0 62116 5 1 1 62115
0 62117 7 1 2 96377 107349
0 62118 5 1 1 62117
0 62119 7 1 2 107267 62118
0 62120 5 1 1 62119
0 62121 7 1 2 72846 95745
0 62122 7 1 2 102326 62121
0 62123 7 1 2 74048 62122
0 62124 7 1 2 62120 62123
0 62125 5 1 1 62124
0 62126 7 1 2 62116 62125
0 62127 5 1 1 62126
0 62128 7 1 2 72203 62127
0 62129 5 1 1 62128
0 62130 7 1 2 72075 103974
0 62131 7 3 2 107262 62130
0 62132 7 1 2 93312 107486
0 62133 5 1 1 62132
0 62134 7 1 2 95589 107331
0 62135 7 1 2 107399 62134
0 62136 5 1 1 62135
0 62137 7 1 2 62133 62136
0 62138 5 1 1 62137
0 62139 7 1 2 100813 62138
0 62140 5 1 1 62139
0 62141 7 1 2 84332 89497
0 62142 7 1 2 107487 62141
0 62143 5 1 1 62142
0 62144 7 1 2 62140 62143
0 62145 5 1 1 62144
0 62146 7 1 2 63830 62145
0 62147 5 1 1 62146
0 62148 7 1 2 100814 92560
0 62149 7 1 2 107488 62148
0 62150 5 1 1 62149
0 62151 7 1 2 62147 62150
0 62152 5 1 1 62151
0 62153 7 1 2 99196 62152
0 62154 5 1 1 62153
0 62155 7 1 2 62129 62154
0 62156 5 1 1 62155
0 62157 7 1 2 66907 62156
0 62158 5 1 1 62157
0 62159 7 1 2 62084 62158
0 62160 7 1 2 62043 62159
0 62161 5 1 1 62160
0 62162 7 1 2 92334 62161
0 62163 5 1 1 62162
0 62164 7 9 2 69085 67247
0 62165 7 1 2 84384 107416
0 62166 5 1 1 62165
0 62167 7 2 2 68227 102272
0 62168 7 1 2 79117 85369
0 62169 7 1 2 107498 62168
0 62170 5 1 1 62169
0 62171 7 1 2 62166 62170
0 62172 5 1 1 62171
0 62173 7 1 2 97748 62172
0 62174 5 1 1 62173
0 62175 7 1 2 76814 97486
0 62176 7 1 2 104442 62175
0 62177 7 1 2 107499 62176
0 62178 5 1 1 62177
0 62179 7 1 2 62174 62178
0 62180 5 1 1 62179
0 62181 7 1 2 72847 62180
0 62182 5 1 1 62181
0 62183 7 2 2 104471 107417
0 62184 5 1 1 107500
0 62185 7 1 2 72204 107501
0 62186 5 1 1 62185
0 62187 7 1 2 62182 62186
0 62188 5 1 1 62187
0 62189 7 1 2 107489 62188
0 62190 5 1 1 62189
0 62191 7 1 2 99675 92480
0 62192 7 2 2 70696 90428
0 62193 7 1 2 97757 99051
0 62194 7 1 2 107502 62193
0 62195 7 1 2 62191 62194
0 62196 5 1 1 62195
0 62197 7 1 2 62190 62196
0 62198 5 1 1 62197
0 62199 7 1 2 81948 62198
0 62200 5 1 1 62199
0 62201 7 3 2 103885 90748
0 62202 7 1 2 98927 107504
0 62203 5 1 1 62202
0 62204 7 2 2 96414 104538
0 62205 7 1 2 90801 98074
0 62206 7 1 2 107507 62205
0 62207 5 1 1 62206
0 62208 7 1 2 62203 62207
0 62209 5 1 1 62208
0 62210 7 1 2 70301 62209
0 62211 5 1 1 62210
0 62212 7 1 2 91267 88656
0 62213 7 1 2 107508 62212
0 62214 5 1 1 62213
0 62215 7 1 2 62211 62214
0 62216 5 1 1 62215
0 62217 7 1 2 98621 62216
0 62218 5 1 1 62217
0 62219 7 2 2 96781 83279
0 62220 7 1 2 94210 107505
0 62221 7 1 2 107509 62220
0 62222 5 1 1 62221
0 62223 7 1 2 62218 62222
0 62224 5 1 1 62223
0 62225 7 1 2 69034 62224
0 62226 5 1 1 62225
0 62227 7 2 2 72293 107423
0 62228 7 1 2 75671 89498
0 62229 7 1 2 94819 62228
0 62230 7 1 2 107511 62229
0 62231 5 1 1 62230
0 62232 7 1 2 62226 62231
0 62233 5 1 1 62232
0 62234 7 1 2 68902 62233
0 62235 5 1 1 62234
0 62236 7 2 2 78188 89556
0 62237 7 1 2 73298 102273
0 62238 7 1 2 107513 62237
0 62239 7 1 2 107512 62238
0 62240 5 1 1 62239
0 62241 7 1 2 62235 62240
0 62242 5 1 1 62241
0 62243 7 1 2 72205 62242
0 62244 5 1 1 62243
0 62245 7 2 2 73299 98414
0 62246 7 1 2 102523 107514
0 62247 7 2 2 107515 62246
0 62248 5 1 1 107517
0 62249 7 2 2 102274 107516
0 62250 7 3 2 77914 107389
0 62251 7 1 2 107519 107521
0 62252 5 1 1 62251
0 62253 7 1 2 85038 103147
0 62254 7 1 2 91319 62253
0 62255 7 1 2 100772 62254
0 62256 5 1 1 62255
0 62257 7 1 2 62252 62256
0 62258 5 1 1 62257
0 62259 7 1 2 68903 62258
0 62260 5 1 1 62259
0 62261 7 1 2 62248 62260
0 62262 5 1 1 62261
0 62263 7 1 2 72206 62262
0 62264 5 1 1 62263
0 62265 7 1 2 72497 90430
0 62266 7 1 2 91641 97248
0 62267 7 1 2 107120 62266
0 62268 7 1 2 62265 62267
0 62269 5 1 1 62268
0 62270 7 1 2 62264 62269
0 62271 5 1 1 62270
0 62272 7 1 2 107284 62271
0 62273 5 1 1 62272
0 62274 7 1 2 98803 3860
0 62275 5 2 1 62274
0 62276 7 2 2 97200 96050
0 62277 7 1 2 101826 107526
0 62278 5 1 1 62277
0 62279 7 1 2 98016 107520
0 62280 5 1 1 62279
0 62281 7 1 2 62278 62280
0 62282 5 1 1 62281
0 62283 7 1 2 107390 62282
0 62284 5 1 1 62283
0 62285 7 1 2 91274 79678
0 62286 7 1 2 96516 62285
0 62287 7 1 2 103732 107478
0 62288 7 1 2 62286 62287
0 62289 5 1 1 62288
0 62290 7 1 2 62284 62289
0 62291 5 1 1 62290
0 62292 7 1 2 68904 62291
0 62293 5 1 1 62292
0 62294 7 1 2 72207 107518
0 62295 5 1 1 62294
0 62296 7 1 2 62293 62295
0 62297 5 1 1 62296
0 62298 7 1 2 107524 62297
0 62299 5 1 1 62298
0 62300 7 1 2 86097 99022
0 62301 7 1 2 92150 97454
0 62302 7 1 2 62300 62301
0 62303 5 1 1 62302
0 62304 7 1 2 62184 62303
0 62305 5 1 1 62304
0 62306 7 1 2 89421 107391
0 62307 7 1 2 62305 62306
0 62308 5 1 1 62307
0 62309 7 1 2 62299 62308
0 62310 7 1 2 62273 62309
0 62311 7 1 2 62244 62310
0 62312 7 1 2 62200 62311
0 62313 5 1 1 62312
0 62314 7 1 2 72076 62313
0 62315 5 1 1 62314
0 62316 7 2 2 64005 102649
0 62317 7 1 2 100769 107528
0 62318 5 1 1 62317
0 62319 7 2 2 91677 98599
0 62320 5 1 1 107530
0 62321 7 1 2 72498 101540
0 62322 5 1 1 62321
0 62323 7 1 2 62320 62322
0 62324 5 2 1 62323
0 62325 7 1 2 69086 102700
0 62326 7 1 2 107532 62325
0 62327 5 1 1 62326
0 62328 7 1 2 62318 62327
0 62329 5 1 1 62328
0 62330 7 1 2 83087 62329
0 62331 5 1 1 62330
0 62332 7 1 2 99799 91845
0 62333 7 1 2 102866 86589
0 62334 7 1 2 62332 62333
0 62335 5 1 1 62334
0 62336 7 1 2 62331 62335
0 62337 5 1 1 62336
0 62338 7 1 2 72848 62337
0 62339 5 1 1 62338
0 62340 7 1 2 82831 91846
0 62341 7 1 2 104716 62340
0 62342 7 1 2 88653 62341
0 62343 5 1 1 62342
0 62344 7 1 2 70697 62343
0 62345 7 1 2 62339 62344
0 62346 5 1 1 62345
0 62347 7 1 2 103368 107490
0 62348 7 1 2 104627 62347
0 62349 7 1 2 101143 62348
0 62350 5 1 1 62349
0 62351 7 1 2 65662 62350
0 62352 5 1 1 62351
0 62353 7 1 2 69035 62352
0 62354 7 1 2 62346 62353
0 62355 5 1 1 62354
0 62356 7 2 2 89499 107491
0 62357 5 1 1 107534
0 62358 7 2 2 72294 73804
0 62359 7 1 2 65663 89557
0 62360 7 2 2 107536 62359
0 62361 5 1 1 107538
0 62362 7 1 2 62357 62361
0 62363 5 1 1 62362
0 62364 7 1 2 98415 62363
0 62365 5 1 1 62364
0 62366 7 1 2 104142 107535
0 62367 5 1 1 62366
0 62368 7 1 2 96791 107539
0 62369 5 1 1 62368
0 62370 7 1 2 62367 62369
0 62371 7 1 2 62365 62370
0 62372 5 1 1 62371
0 62373 7 1 2 75810 104628
0 62374 7 1 2 62372 62373
0 62375 5 1 1 62374
0 62376 7 1 2 62355 62375
0 62377 5 1 1 62376
0 62378 7 1 2 68905 62377
0 62379 5 1 1 62378
0 62380 7 1 2 102275 107492
0 62381 7 1 2 101144 62380
0 62382 5 1 1 62381
0 62383 7 1 2 107537 107503
0 62384 7 1 2 104127 62383
0 62385 5 1 1 62384
0 62386 7 1 2 62382 62385
0 62387 5 1 1 62386
0 62388 7 2 2 74009 104629
0 62389 7 1 2 70302 107540
0 62390 7 1 2 62387 62389
0 62391 5 1 1 62390
0 62392 7 1 2 62379 62391
0 62393 5 1 1 62392
0 62394 7 1 2 71974 62393
0 62395 5 1 1 62394
0 62396 7 1 2 79743 107392
0 62397 7 2 2 101145 62396
0 62398 7 1 2 75840 103139
0 62399 7 1 2 107542 62398
0 62400 5 1 1 62399
0 62401 7 1 2 62395 62400
0 62402 5 1 1 62401
0 62403 7 1 2 84889 62402
0 62404 5 1 1 62403
0 62405 7 1 2 104128 103122
0 62406 5 2 1 62405
0 62407 7 1 2 101146 107401
0 62408 5 1 1 62407
0 62409 7 1 2 107544 62408
0 62410 5 1 1 62409
0 62411 7 1 2 103140 107493
0 62412 7 1 2 62410 62411
0 62413 5 1 1 62412
0 62414 7 1 2 106938 106953
0 62415 7 1 2 107543 62414
0 62416 5 1 1 62415
0 62417 7 1 2 62413 62416
0 62418 5 1 1 62417
0 62419 7 1 2 75775 62418
0 62420 5 1 1 62419
0 62421 7 1 2 62404 62420
0 62422 7 1 2 62315 62421
0 62423 5 1 1 62422
0 62424 7 1 2 107210 62423
0 62425 5 1 1 62424
0 62426 7 1 2 70303 101705
0 62427 5 1 1 62426
0 62428 7 1 2 91678 93828
0 62429 5 1 1 62428
0 62430 7 1 2 62427 62429
0 62431 5 1 1 62430
0 62432 7 1 2 98701 98046
0 62433 7 1 2 62431 62432
0 62434 5 1 1 62433
0 62435 7 1 2 98779 95565
0 62436 7 1 2 107296 62435
0 62437 7 1 2 100738 62436
0 62438 5 1 1 62437
0 62439 7 1 2 62434 62438
0 62440 5 1 1 62439
0 62441 7 1 2 91076 62440
0 62442 5 1 1 62441
0 62443 7 1 2 8266 47675
0 62444 5 1 1 62443
0 62445 7 1 2 81000 20269
0 62446 7 2 2 62444 62445
0 62447 7 1 2 69087 107546
0 62448 5 1 1 62447
0 62449 7 1 2 93628 107225
0 62450 5 1 1 62449
0 62451 7 1 2 62448 62450
0 62452 5 1 1 62451
0 62453 7 1 2 102276 62452
0 62454 5 1 1 62453
0 62455 7 1 2 98464 73814
0 62456 7 1 2 105795 62455
0 62457 5 1 1 62456
0 62458 7 1 2 62454 62457
0 62459 5 1 1 62458
0 62460 7 1 2 83088 105070
0 62461 7 1 2 62459 62460
0 62462 5 1 1 62461
0 62463 7 1 2 62442 62462
0 62464 5 1 1 62463
0 62465 7 1 2 67148 62464
0 62466 5 1 1 62465
0 62467 7 1 2 97285 88699
0 62468 5 1 1 62467
0 62469 7 1 2 107472 62468
0 62470 5 1 1 62469
0 62471 7 1 2 97239 90254
0 62472 7 1 2 98142 62471
0 62473 7 1 2 62470 62472
0 62474 5 1 1 62473
0 62475 7 1 2 62466 62474
0 62476 5 1 1 62475
0 62477 7 1 2 67248 62476
0 62478 5 1 1 62477
0 62479 7 1 2 91077 98052
0 62480 5 1 1 62479
0 62481 7 1 2 74482 103690
0 62482 7 1 2 98130 62481
0 62483 5 1 1 62482
0 62484 7 1 2 62480 62483
0 62485 5 1 1 62484
0 62486 7 1 2 107278 62485
0 62487 5 1 1 62486
0 62488 7 1 2 96537 107379
0 62489 7 1 2 86079 62488
0 62490 7 1 2 96332 62489
0 62491 5 1 1 62490
0 62492 7 1 2 62487 62491
0 62493 5 1 1 62492
0 62494 7 1 2 71219 62493
0 62495 5 1 1 62494
0 62496 7 1 2 91291 97308
0 62497 7 1 2 106963 62496
0 62498 7 1 2 98047 62497
0 62499 5 1 1 62498
0 62500 7 1 2 62495 62499
0 62501 5 1 1 62500
0 62502 7 1 2 100088 62501
0 62503 5 1 1 62502
0 62504 7 1 2 62478 62503
0 62505 5 1 1 62504
0 62506 7 1 2 68906 62505
0 62507 5 1 1 62506
0 62508 7 2 2 103300 107297
0 62509 7 1 2 107234 107548
0 62510 5 1 1 62509
0 62511 7 1 2 101438 103909
0 62512 5 2 1 62511
0 62513 7 1 2 100442 98851
0 62514 5 1 1 62513
0 62515 7 1 2 107550 62514
0 62516 5 1 1 62515
0 62517 7 1 2 84038 62516
0 62518 7 1 2 96333 62517
0 62519 5 1 1 62518
0 62520 7 1 2 62510 62519
0 62521 5 1 1 62520
0 62522 7 1 2 84890 62521
0 62523 5 1 1 62522
0 62524 7 1 2 107549 107421
0 62525 5 1 1 62524
0 62526 7 1 2 100584 98465
0 62527 5 2 1 62526
0 62528 7 1 2 77492 101201
0 62529 5 1 1 62528
0 62530 7 1 2 107552 62529
0 62531 5 1 1 62530
0 62532 7 1 2 106964 62531
0 62533 7 1 2 96334 62532
0 62534 5 1 1 62533
0 62535 7 1 2 62525 62534
0 62536 7 1 2 62523 62535
0 62537 5 1 1 62536
0 62538 7 1 2 107541 62537
0 62539 5 1 1 62538
0 62540 7 1 2 62507 62539
0 62541 5 1 1 62540
0 62542 7 1 2 71975 62541
0 62543 5 1 1 62542
0 62544 7 1 2 83735 102862
0 62545 5 1 1 62544
0 62546 7 1 2 104620 107246
0 62547 5 1 1 62546
0 62548 7 1 2 62545 62547
0 62549 5 1 1 62548
0 62550 7 1 2 107413 62549
0 62551 5 1 1 62550
0 62552 7 2 2 103345 98631
0 62553 7 1 2 70578 107554
0 62554 7 1 2 103141 62553
0 62555 7 1 2 107407 62554
0 62556 5 1 1 62555
0 62557 7 1 2 62551 62556
0 62558 5 1 1 62557
0 62559 7 1 2 107263 62558
0 62560 5 1 1 62559
0 62561 7 1 2 107551 107553
0 62562 5 1 1 62561
0 62563 7 1 2 93899 62562
0 62564 7 1 2 98084 62563
0 62565 5 1 1 62564
0 62566 7 1 2 62560 62565
0 62567 5 1 1 62566
0 62568 7 1 2 95445 62567
0 62569 5 1 1 62568
0 62570 7 1 2 104160 99069
0 62571 5 1 1 62570
0 62572 7 1 2 86859 107555
0 62573 5 1 1 62572
0 62574 7 1 2 62571 62573
0 62575 5 1 1 62574
0 62576 7 1 2 73300 103142
0 62577 7 1 2 62575 62576
0 62578 5 1 1 62577
0 62579 7 1 2 39669 104830
0 62580 5 1 1 62579
0 62581 7 1 2 70698 101191
0 62582 7 1 2 96540 62581
0 62583 7 1 2 62580 62582
0 62584 5 1 1 62583
0 62585 7 1 2 62578 62584
0 62586 5 1 1 62585
0 62587 7 1 2 99376 107004
0 62588 7 1 2 62586 62587
0 62589 5 1 1 62588
0 62590 7 1 2 62569 62589
0 62591 7 1 2 62543 62590
0 62592 5 1 1 62591
0 62593 7 1 2 85565 62592
0 62594 5 1 1 62593
0 62595 7 1 2 99340 102776
0 62596 7 1 2 102057 62595
0 62597 5 2 1 62596
0 62598 7 1 2 82513 104771
0 62599 7 1 2 101608 62598
0 62600 5 1 1 62599
0 62601 7 1 2 107556 62600
0 62602 5 1 1 62601
0 62603 7 1 2 73805 62602
0 62604 5 1 1 62603
0 62605 7 2 2 103774 107483
0 62606 7 1 2 101785 107558
0 62607 5 1 1 62606
0 62608 7 1 2 100351 75827
0 62609 7 1 2 87430 107247
0 62610 7 1 2 62608 62609
0 62611 5 1 1 62610
0 62612 7 1 2 62607 62611
0 62613 5 1 1 62612
0 62614 7 1 2 64228 62613
0 62615 5 1 1 62614
0 62616 7 1 2 102711 97212
0 62617 5 1 1 62616
0 62618 7 1 2 102743 62617
0 62619 5 1 1 62618
0 62620 7 1 2 100663 78368
0 62621 7 1 2 62619 62620
0 62622 5 1 1 62621
0 62623 7 1 2 100976 107139
0 62624 7 1 2 89336 62623
0 62625 7 1 2 98388 62624
0 62626 5 1 1 62625
0 62627 7 1 2 62622 62626
0 62628 7 1 2 62615 62627
0 62629 5 1 1 62628
0 62630 7 1 2 65240 62629
0 62631 5 1 1 62630
0 62632 7 1 2 62604 62631
0 62633 5 1 1 62632
0 62634 7 1 2 71877 62633
0 62635 5 1 1 62634
0 62636 7 1 2 96504 93716
0 62637 7 1 2 107248 62636
0 62638 5 1 1 62637
0 62639 7 1 2 100157 79649
0 62640 7 1 2 101615 62639
0 62641 7 1 2 105735 62640
0 62642 5 1 1 62641
0 62643 7 1 2 62638 62642
0 62644 5 1 1 62643
0 62645 7 1 2 63944 62644
0 62646 5 1 1 62645
0 62647 7 1 2 103040 102814
0 62648 5 1 1 62647
0 62649 7 1 2 62015 62648
0 62650 5 1 1 62649
0 62651 7 1 2 89385 105099
0 62652 7 1 2 62650 62651
0 62653 5 1 1 62652
0 62654 7 1 2 62646 62653
0 62655 5 1 1 62654
0 62656 7 1 2 65863 62655
0 62657 5 1 1 62656
0 62658 7 2 2 102277 97003
0 62659 7 1 2 96403 84020
0 62660 7 1 2 103993 62659
0 62661 7 1 2 107560 62660
0 62662 5 1 1 62661
0 62663 7 1 2 62657 62662
0 62664 5 1 1 62663
0 62665 7 1 2 67149 62664
0 62666 5 1 1 62665
0 62667 7 1 2 101609 107335
0 62668 5 1 1 62667
0 62669 7 1 2 74483 97141
0 62670 7 2 2 105317 62669
0 62671 7 1 2 70699 107562
0 62672 5 1 1 62671
0 62673 7 1 2 62668 62672
0 62674 5 2 1 62673
0 62675 7 1 2 88431 107564
0 62676 5 1 1 62675
0 62677 7 1 2 88036 87422
0 62678 7 2 2 90199 62677
0 62679 7 1 2 99417 79057
0 62680 7 1 2 107566 62679
0 62681 5 1 1 62680
0 62682 7 1 2 62676 62681
0 62683 5 1 1 62682
0 62684 7 1 2 102701 62683
0 62685 5 1 1 62684
0 62686 7 1 2 62666 62685
0 62687 7 1 2 62635 62686
0 62688 5 1 1 62687
0 62689 7 1 2 70579 62688
0 62690 5 1 1 62689
0 62691 7 1 2 76136 92161
0 62692 7 1 2 106155 107336
0 62693 7 1 2 62691 62692
0 62694 5 1 1 62693
0 62695 7 1 2 79000 100347
0 62696 7 1 2 76865 62695
0 62697 7 1 2 105609 62696
0 62698 5 1 1 62697
0 62699 7 1 2 62694 62698
0 62700 5 1 1 62699
0 62701 7 1 2 63945 62700
0 62702 5 1 1 62701
0 62703 7 1 2 13061 17969
0 62704 7 1 2 105689 62703
0 62705 7 1 2 107563 62704
0 62706 5 1 1 62705
0 62707 7 1 2 62702 62706
0 62708 5 1 1 62707
0 62709 7 1 2 67249 62708
0 62710 5 1 1 62709
0 62711 7 1 2 75135 79001
0 62712 7 1 2 91708 62711
0 62713 7 1 2 102030 104674
0 62714 7 1 2 62712 62713
0 62715 5 1 1 62714
0 62716 7 1 2 62710 62715
0 62717 5 1 1 62716
0 62718 7 1 2 71878 62717
0 62719 5 1 1 62718
0 62720 7 1 2 102964 107559
0 62721 5 1 1 62720
0 62722 7 1 2 107557 62721
0 62723 5 1 1 62722
0 62724 7 1 2 107430 62723
0 62725 5 1 1 62724
0 62726 7 1 2 74911 103063
0 62727 7 1 2 107565 62726
0 62728 5 1 1 62727
0 62729 7 1 2 62725 62728
0 62730 7 1 2 62719 62729
0 62731 7 1 2 62690 62730
0 62732 5 1 1 62731
0 62733 7 1 2 68228 62732
0 62734 5 1 1 62733
0 62735 7 1 2 73301 86559
0 62736 7 1 2 78297 62735
0 62737 7 1 2 97692 104963
0 62738 7 1 2 106169 62737
0 62739 7 1 2 62736 62738
0 62740 5 1 1 62739
0 62741 7 1 2 62734 62740
0 62742 5 1 1 62741
0 62743 7 1 2 99377 62742
0 62744 5 1 1 62743
0 62745 7 1 2 104286 106885
0 62746 5 1 1 62745
0 62747 7 1 2 70580 84307
0 62748 7 1 2 99680 62747
0 62749 5 1 1 62748
0 62750 7 1 2 62746 62749
0 62751 5 1 1 62750
0 62752 7 1 2 65241 62751
0 62753 5 1 1 62752
0 62754 7 1 2 83142 102167
0 62755 7 1 2 95205 62754
0 62756 5 1 1 62755
0 62757 7 1 2 62753 62756
0 62758 5 1 1 62757
0 62759 7 1 2 96439 62758
0 62760 5 1 1 62759
0 62761 7 3 2 89181 107250
0 62762 7 1 2 65664 107568
0 62763 5 1 1 62762
0 62764 7 1 2 62760 62763
0 62765 5 1 1 62764
0 62766 7 1 2 89526 62765
0 62767 5 1 1 62766
0 62768 7 1 2 73822 107569
0 62769 5 1 1 62768
0 62770 7 1 2 62767 62769
0 62771 5 1 1 62770
0 62772 7 1 2 69036 62771
0 62773 5 1 1 62772
0 62774 7 1 2 91575 107570
0 62775 5 1 1 62774
0 62776 7 1 2 62773 62775
0 62777 5 1 1 62776
0 62778 7 1 2 85566 62777
0 62779 5 1 1 62778
0 62780 7 1 2 99663 107238
0 62781 5 1 1 62780
0 62782 7 1 2 103943 102723
0 62783 5 1 1 62782
0 62784 7 1 2 62781 62783
0 62785 5 1 1 62784
0 62786 7 1 2 70581 62785
0 62787 5 1 1 62786
0 62788 7 1 2 84759 103964
0 62789 5 1 1 62788
0 62790 7 1 2 56299 62789
0 62791 5 1 1 62790
0 62792 7 1 2 74912 62791
0 62793 5 1 1 62792
0 62794 7 1 2 62787 62793
0 62795 5 1 1 62794
0 62796 7 1 2 98125 62795
0 62797 5 1 1 62796
0 62798 7 1 2 81949 106743
0 62799 5 1 1 62798
0 62800 7 1 2 107381 62799
0 62801 5 2 1 62800
0 62802 7 1 2 102894 107571
0 62803 5 1 1 62802
0 62804 7 1 2 62797 62803
0 62805 5 1 1 62804
0 62806 7 1 2 89527 62805
0 62807 5 1 1 62806
0 62808 7 1 2 73823 74456
0 62809 7 1 2 107572 62808
0 62810 5 1 1 62809
0 62811 7 1 2 62807 62810
0 62812 5 1 1 62811
0 62813 7 1 2 97090 62812
0 62814 5 1 1 62813
0 62815 7 1 2 62779 62814
0 62816 5 1 1 62815
0 62817 7 1 2 98132 62816
0 62818 5 1 1 62817
0 62819 7 1 2 70700 107360
0 62820 5 1 1 62819
0 62821 7 1 2 65665 99772
0 62822 7 1 2 106802 62821
0 62823 5 1 1 62822
0 62824 7 1 2 62820 62823
0 62825 5 1 1 62824
0 62826 7 1 2 88932 62825
0 62827 5 1 1 62826
0 62828 7 1 2 73834 107361
0 62829 5 1 1 62828
0 62830 7 1 2 62827 62829
0 62831 5 1 1 62830
0 62832 7 1 2 63946 62831
0 62833 5 1 1 62832
0 62834 7 1 2 96357 107362
0 62835 5 1 1 62834
0 62836 7 1 2 62833 62835
0 62837 5 1 1 62836
0 62838 7 1 2 68739 62837
0 62839 5 1 1 62838
0 62840 7 1 2 104846 61173
0 62841 5 1 1 62840
0 62842 7 1 2 70304 74227
0 62843 7 1 2 62841 62842
0 62844 7 1 2 96378 62843
0 62845 5 1 1 62844
0 62846 7 1 2 84955 102867
0 62847 7 1 2 96489 62846
0 62848 5 1 1 62847
0 62849 7 1 2 62845 62848
0 62850 5 1 1 62849
0 62851 7 1 2 84891 62850
0 62852 5 1 1 62851
0 62853 7 1 2 100089 107384
0 62854 5 1 1 62853
0 62855 7 1 2 80667 104838
0 62856 5 1 1 62855
0 62857 7 1 2 62854 62856
0 62858 5 1 1 62857
0 62859 7 1 2 105648 62858
0 62860 5 1 1 62859
0 62861 7 1 2 62852 62860
0 62862 7 1 2 62839 62861
0 62863 5 1 1 62862
0 62864 7 1 2 85039 79650
0 62865 7 1 2 92512 62864
0 62866 7 1 2 62863 62865
0 62867 5 1 1 62866
0 62868 7 1 2 62818 62867
0 62869 7 1 2 62744 62868
0 62870 5 1 1 62869
0 62871 7 1 2 81086 62870
0 62872 5 1 1 62871
0 62873 7 1 2 97332 93480
0 62874 5 1 1 62873
0 62875 7 1 2 60676 62874
0 62876 5 4 1 62875
0 62877 7 1 2 90630 107107
0 62878 5 1 1 62877
0 62879 7 1 2 86534 74290
0 62880 7 1 2 99014 62879
0 62881 5 1 1 62880
0 62882 7 1 2 62878 62881
0 62883 5 1 1 62882
0 62884 7 1 2 70582 62883
0 62885 5 1 1 62884
0 62886 7 1 2 86102 92682
0 62887 7 1 2 106849 62886
0 62888 5 1 1 62887
0 62889 7 1 2 62885 62888
0 62890 5 1 1 62889
0 62891 7 1 2 107573 62890
0 62892 5 1 1 62891
0 62893 7 1 2 87423 101974
0 62894 7 1 2 103132 98068
0 62895 7 1 2 62893 62894
0 62896 5 1 1 62895
0 62897 7 1 2 74360 75170
0 62898 7 2 2 93481 62897
0 62899 5 1 1 107577
0 62900 7 1 2 70305 106563
0 62901 7 1 2 107578 62900
0 62902 5 1 1 62901
0 62903 7 1 2 62896 62902
0 62904 5 1 1 62903
0 62905 7 1 2 73806 62904
0 62906 5 1 1 62905
0 62907 7 1 2 100235 103173
0 62908 7 1 2 92608 99291
0 62909 7 1 2 62907 62908
0 62910 5 1 1 62909
0 62911 7 1 2 62906 62910
0 62912 7 1 2 62892 62911
0 62913 5 1 1 62912
0 62914 7 1 2 106978 62913
0 62915 5 1 1 62914
0 62916 7 2 2 89411 107163
0 62917 7 2 2 79776 103245
0 62918 7 1 2 94595 85192
0 62919 7 1 2 107581 62918
0 62920 7 1 2 107579 62919
0 62921 5 1 1 62920
0 62922 7 1 2 87583 99122
0 62923 7 1 2 107582 62922
0 62924 7 1 2 107574 62923
0 62925 5 1 1 62924
0 62926 7 1 2 62921 62925
0 62927 7 1 2 62915 62926
0 62928 5 1 1 62927
0 62929 7 1 2 104129 62928
0 62930 5 1 1 62929
0 62931 7 1 2 106979 106954
0 62932 5 1 1 62931
0 62933 7 1 2 74913 107127
0 62934 5 1 1 62933
0 62935 7 1 2 62932 62934
0 62936 5 1 1 62935
0 62937 7 1 2 68740 62936
0 62938 5 1 1 62937
0 62939 7 1 2 86688 91847
0 62940 7 1 2 102511 62939
0 62941 5 1 1 62940
0 62942 7 1 2 62938 62941
0 62943 5 1 1 62942
0 62944 7 2 2 87757 107575
0 62945 5 1 1 107583
0 62946 7 1 2 62899 62945
0 62947 5 1 1 62946
0 62948 7 1 2 77842 62947
0 62949 7 1 2 62943 62948
0 62950 5 1 1 62949
0 62951 7 1 2 98889 105394
0 62952 5 1 1 62951
0 62953 7 2 2 63831 107576
0 62954 5 1 1 107585
0 62955 7 1 2 96701 107586
0 62956 5 1 1 62955
0 62957 7 1 2 62952 62956
0 62958 5 1 1 62957
0 62959 7 1 2 100739 103894
0 62960 7 1 2 62958 62959
0 62961 5 1 1 62960
0 62962 7 1 2 62950 62961
0 62963 5 1 1 62962
0 62964 7 1 2 101147 62963
0 62965 5 1 1 62964
0 62966 7 1 2 86356 102099
0 62967 7 1 2 107464 62966
0 62968 7 1 2 104605 62967
0 62969 7 1 2 107567 62968
0 62970 5 1 1 62969
0 62971 7 1 2 102650 91564
0 62972 7 1 2 105940 62971
0 62973 5 1 1 62972
0 62974 7 1 2 98416 88638
0 62975 7 1 2 107425 62974
0 62976 5 1 1 62975
0 62977 7 1 2 62973 62976
0 62978 5 1 1 62977
0 62979 7 1 2 92561 92609
0 62980 5 1 1 62979
0 62981 7 1 2 62954 62980
0 62982 5 1 1 62981
0 62983 7 1 2 66908 62982
0 62984 7 1 2 62978 62983
0 62985 5 1 1 62984
0 62986 7 1 2 62970 62985
0 62987 5 1 1 62986
0 62988 7 1 2 72077 62987
0 62989 5 1 1 62988
0 62990 7 1 2 73302 62989
0 62991 7 1 2 62965 62990
0 62992 7 1 2 62930 62991
0 62993 5 1 1 62992
0 62994 7 1 2 74321 96256
0 62995 7 1 2 107140 62994
0 62996 7 1 2 63832 97109
0 62997 7 1 2 98890 62996
0 62998 7 1 2 62995 62997
0 62999 5 1 1 62998
0 63000 7 1 2 98261 107128
0 63001 5 1 1 63000
0 63002 7 1 2 106980 107531
0 63003 5 1 1 63002
0 63004 7 1 2 63001 63003
0 63005 5 1 1 63004
0 63006 7 2 2 93717 96344
0 63007 7 1 2 106903 107587
0 63008 7 1 2 63005 63007
0 63009 5 1 1 63008
0 63010 7 1 2 62999 63009
0 63011 5 1 1 63010
0 63012 7 1 2 81950 63011
0 63013 5 1 1 63012
0 63014 7 2 2 95353 91700
0 63015 7 1 2 107588 107589
0 63016 5 1 1 63015
0 63017 7 2 2 91353 92182
0 63018 7 1 2 65705 98001
0 63019 7 1 2 107591 63018
0 63020 5 1 1 63019
0 63021 7 1 2 63016 63020
0 63022 5 1 1 63021
0 63023 7 1 2 69088 63022
0 63024 5 1 1 63023
0 63025 7 1 2 77387 93328
0 63026 5 2 1 63025
0 63027 7 1 2 65706 105662
0 63028 5 1 1 63027
0 63029 7 1 2 107593 63028
0 63030 5 1 1 63029
0 63031 7 1 2 84424 92469
0 63032 7 1 2 63030 63031
0 63033 5 1 1 63032
0 63034 7 1 2 63024 63033
0 63035 5 1 1 63034
0 63036 7 1 2 72499 63035
0 63037 5 1 1 63036
0 63038 7 1 2 98530 106513
0 63039 5 1 1 63038
0 63040 7 1 2 63037 63039
0 63041 5 1 1 63040
0 63042 7 1 2 100740 63041
0 63043 5 1 1 63042
0 63044 7 1 2 70933 98262
0 63045 5 1 1 63044
0 63046 7 1 2 77196 106178
0 63047 5 1 1 63046
0 63048 7 1 2 63045 63047
0 63049 5 1 1 63048
0 63050 7 1 2 64006 63049
0 63051 5 1 1 63050
0 63052 7 1 2 99357 63051
0 63053 5 1 1 63052
0 63054 7 1 2 72500 98006
0 63055 5 1 1 63054
0 63056 7 1 2 88935 63055
0 63057 5 1 1 63056
0 63058 7 1 2 107592 63057
0 63059 7 1 2 63053 63058
0 63060 5 1 1 63059
0 63061 7 1 2 96541 106449
0 63062 7 1 2 107590 63061
0 63063 5 1 1 63062
0 63064 7 1 2 63060 63063
0 63065 5 1 1 63064
0 63066 7 1 2 80877 63065
0 63067 5 1 1 63066
0 63068 7 1 2 96505 98715
0 63069 7 1 2 98751 107319
0 63070 7 1 2 63068 63069
0 63071 5 1 1 63070
0 63072 7 1 2 63067 63071
0 63073 5 1 1 63072
0 63074 7 1 2 80668 63073
0 63075 5 1 1 63074
0 63076 7 1 2 63043 63075
0 63077 5 1 1 63076
0 63078 7 1 2 72295 63077
0 63079 5 1 1 63078
0 63080 7 1 2 63013 63079
0 63081 5 1 1 63080
0 63082 7 1 2 88282 63081
0 63083 5 1 1 63082
0 63084 7 3 2 84590 85982
0 63085 7 1 2 98002 73815
0 63086 5 1 1 63085
0 63087 7 1 2 70755 95285
0 63088 7 1 2 96584 63087
0 63089 5 1 1 63088
0 63090 7 1 2 63086 63089
0 63091 5 1 1 63090
0 63092 7 1 2 64007 63091
0 63093 5 1 1 63092
0 63094 7 1 2 95646 92593
0 63095 5 1 1 63094
0 63096 7 1 2 107594 63095
0 63097 5 1 1 63096
0 63098 7 1 2 69089 65666
0 63099 7 1 2 63097 63098
0 63100 5 1 1 63099
0 63101 7 1 2 63093 63100
0 63102 5 1 1 63101
0 63103 7 1 2 63947 63102
0 63104 5 1 1 63103
0 63105 7 1 2 65667 105797
0 63106 5 1 1 63105
0 63107 7 1 2 63104 63106
0 63108 5 1 1 63107
0 63109 7 1 2 106965 63108
0 63110 5 1 1 63109
0 63111 7 1 2 84039 98007
0 63112 7 1 2 107485 63111
0 63113 5 1 1 63112
0 63114 7 1 2 63110 63113
0 63115 5 1 1 63114
0 63116 7 1 2 72501 63115
0 63117 5 1 1 63116
0 63118 7 1 2 82514 107108
0 63119 5 1 1 63118
0 63120 7 1 2 65864 84747
0 63121 5 1 1 63120
0 63122 7 1 2 63119 63121
0 63123 5 1 1 63122
0 63124 7 1 2 70583 63123
0 63125 5 1 1 63124
0 63126 7 1 2 65865 107431
0 63127 5 1 1 63126
0 63128 7 1 2 63125 63127
0 63129 5 1 1 63128
0 63130 7 1 2 77197 63129
0 63131 5 1 1 63130
0 63132 7 1 2 100741 101321
0 63133 5 1 1 63132
0 63134 7 1 2 63131 63133
0 63135 5 1 1 63134
0 63136 7 1 2 99378 102513
0 63137 7 1 2 63135 63136
0 63138 5 1 1 63137
0 63139 7 1 2 63117 63138
0 63140 5 1 1 63139
0 63141 7 1 2 107595 63140
0 63142 5 1 1 63141
0 63143 7 1 2 99379 101786
0 63144 7 2 2 106620 63143
0 63145 5 1 1 107598
0 63146 7 1 2 87073 27048
0 63147 5 1 1 63146
0 63148 7 1 2 69332 96565
0 63149 5 1 1 63148
0 63150 7 1 2 63147 63149
0 63151 5 1 1 63150
0 63152 7 1 2 68741 63151
0 63153 5 1 1 63152
0 63154 7 1 2 84919 101541
0 63155 5 1 1 63154
0 63156 7 1 2 63153 63155
0 63157 5 1 1 63156
0 63158 7 1 2 72502 63157
0 63159 5 1 1 63158
0 63160 7 1 2 94945 107427
0 63161 5 1 1 63160
0 63162 7 1 2 98225 63161
0 63163 5 1 1 63162
0 63164 7 1 2 63159 63163
0 63165 5 1 1 63164
0 63166 7 1 2 107599 63165
0 63167 5 1 1 63166
0 63168 7 2 2 79002 97184
0 63169 7 2 2 107325 107600
0 63170 5 1 1 107602
0 63171 7 1 2 63170 63145
0 63172 5 1 1 63171
0 63173 7 1 2 96566 63172
0 63174 5 1 1 63173
0 63175 7 1 2 70649 102715
0 63176 7 1 2 90431 63175
0 63177 7 1 2 97185 63176
0 63178 5 1 1 63177
0 63179 7 1 2 63174 63178
0 63180 5 1 1 63179
0 63181 7 1 2 100773 63180
0 63182 5 1 1 63181
0 63183 7 1 2 84892 107533
0 63184 5 1 1 63183
0 63185 7 1 2 98282 107525
0 63186 5 1 1 63185
0 63187 7 1 2 70584 83193
0 63188 7 1 2 100783 63187
0 63189 5 1 1 63188
0 63190 7 1 2 63186 63189
0 63191 7 1 2 63184 63190
0 63192 5 1 1 63191
0 63193 7 1 2 107603 63192
0 63194 5 1 1 63193
0 63195 7 1 2 63182 63194
0 63196 7 1 2 63167 63195
0 63197 5 1 1 63196
0 63198 7 1 2 70934 63197
0 63199 5 1 1 63198
0 63200 7 1 2 67250 63199
0 63201 7 1 2 63142 63200
0 63202 5 1 1 63201
0 63203 7 1 2 96379 46665
0 63204 5 1 1 63203
0 63205 7 2 2 72503 107298
0 63206 7 1 2 96111 107604
0 63207 5 1 1 63206
0 63208 7 1 2 63204 63207
0 63209 5 1 1 63208
0 63210 7 1 2 106966 63209
0 63211 5 1 1 63210
0 63212 7 1 2 64008 107547
0 63213 5 1 1 63212
0 63214 7 1 2 69090 98466
0 63215 7 1 2 97172 63214
0 63216 5 1 1 63215
0 63217 7 1 2 63213 63216
0 63218 5 1 1 63217
0 63219 7 1 2 102278 63218
0 63220 5 1 1 63219
0 63221 7 1 2 103910 73828
0 63222 7 1 2 91652 63221
0 63223 5 1 1 63222
0 63224 7 1 2 63220 63223
0 63225 5 1 1 63224
0 63226 7 1 2 82515 63225
0 63227 5 1 1 63226
0 63228 7 1 2 74415 107605
0 63229 5 1 1 63228
0 63230 7 1 2 63227 63229
0 63231 5 1 1 63230
0 63232 7 1 2 84893 84040
0 63233 7 1 2 63231 63232
0 63234 5 1 1 63233
0 63235 7 1 2 63211 63234
0 63236 5 1 1 63235
0 63237 7 1 2 63236 107596
0 63238 5 1 1 63237
0 63239 7 1 2 84425 102346
0 63240 7 1 2 106967 63239
0 63241 7 1 2 96380 63240
0 63242 5 1 1 63241
0 63243 7 1 2 98869 107601
0 63244 5 1 1 63243
0 63245 7 1 2 96381 107597
0 63246 5 1 1 63245
0 63247 7 1 2 63244 63246
0 63248 5 1 1 63247
0 63249 7 1 2 70935 107279
0 63250 7 1 2 63248 63249
0 63251 5 1 1 63250
0 63252 7 1 2 63242 63251
0 63253 5 1 1 63252
0 63254 7 1 2 98263 63253
0 63255 5 1 1 63254
0 63256 7 1 2 72296 63255
0 63257 7 1 2 63238 63256
0 63258 5 1 1 63257
0 63259 7 1 2 72208 63258
0 63260 7 1 2 63202 63259
0 63261 5 1 1 63260
0 63262 7 1 2 68229 63261
0 63263 7 1 2 63083 63262
0 63264 5 1 1 63263
0 63265 7 1 2 62993 63264
0 63266 5 1 1 63265
0 63267 7 1 2 86410 102173
0 63268 7 1 2 106845 63267
0 63269 7 1 2 107580 63268
0 63270 5 1 1 63269
0 63271 7 1 2 71976 107129
0 63272 7 1 2 82279 63271
0 63273 7 1 2 96852 63272
0 63274 7 1 2 107584 63273
0 63275 5 1 1 63274
0 63276 7 1 2 63270 63275
0 63277 5 1 1 63276
0 63278 7 1 2 104130 63277
0 63279 5 1 1 63278
0 63280 7 1 2 104131 107109
0 63281 5 1 1 63280
0 63282 7 1 2 84748 101148
0 63283 5 1 1 63282
0 63284 7 1 2 63281 63283
0 63285 5 1 1 63284
0 63286 7 1 2 81350 63285
0 63287 5 1 1 63286
0 63288 7 1 2 97069 98207
0 63289 7 1 2 99289 63288
0 63290 5 1 1 63289
0 63291 7 1 2 63287 63290
0 63292 5 1 1 63291
0 63293 7 1 2 85848 63292
0 63294 5 1 1 63293
0 63295 7 1 2 99577 98250
0 63296 5 1 1 63295
0 63297 7 1 2 98231 63296
0 63298 5 1 1 63297
0 63299 7 1 2 69037 91247
0 63300 7 1 2 93970 63299
0 63301 7 1 2 79157 63300
0 63302 7 1 2 63298 63301
0 63303 5 1 1 63302
0 63304 7 1 2 63294 63303
0 63305 5 1 1 63304
0 63306 7 1 2 70585 63305
0 63307 5 1 1 63306
0 63308 7 1 2 97578 107527
0 63309 5 1 1 63308
0 63310 7 2 2 73303 101149
0 63311 7 1 2 97706 107606
0 63312 5 1 1 63311
0 63313 7 1 2 63309 63312
0 63314 5 1 1 63313
0 63315 7 1 2 107432 63314
0 63316 5 1 1 63315
0 63317 7 1 2 72849 89193
0 63318 7 1 2 97450 63317
0 63319 5 1 1 63318
0 63320 7 1 2 63316 63319
0 63321 7 1 2 63307 63320
0 63322 5 1 1 63321
0 63323 7 1 2 72078 63322
0 63324 5 1 1 63323
0 63325 7 1 2 84920 104132
0 63326 5 1 1 63325
0 63327 7 1 2 95026 101150
0 63328 5 1 1 63327
0 63329 7 1 2 63326 63328
0 63330 5 1 1 63329
0 63331 7 1 2 70306 63330
0 63332 5 1 1 63331
0 63333 7 1 2 101151 106921
0 63334 5 1 1 63333
0 63335 7 1 2 63332 63334
0 63336 5 1 1 63335
0 63337 7 1 2 95235 87269
0 63338 7 1 2 63336 63337
0 63339 5 1 1 63338
0 63340 7 1 2 63324 63339
0 63341 5 1 1 63340
0 63342 7 1 2 106981 63341
0 63343 5 1 1 63342
0 63344 7 1 2 107232 107607
0 63345 5 1 1 63344
0 63346 7 1 2 107545 63345
0 63347 5 1 1 63346
0 63348 7 1 2 83207 63347
0 63349 5 1 1 63348
0 63350 7 1 2 83886 85040
0 63351 7 1 2 102214 63350
0 63352 5 1 1 63351
0 63353 7 1 2 63349 63352
0 63354 5 1 1 63353
0 63355 7 1 2 77640 63354
0 63356 5 1 1 63355
0 63357 7 1 2 81951 95446
0 63358 7 1 2 98417 63357
0 63359 7 1 2 81351 63358
0 63360 5 1 1 63359
0 63361 7 1 2 63356 63360
0 63362 5 1 1 63361
0 63363 7 1 2 107130 63362
0 63364 5 1 1 63363
0 63365 7 1 2 63343 63364
0 63366 5 1 1 63365
0 63367 7 1 2 23671 31925
0 63368 7 1 2 99062 59222
0 63369 7 1 2 63367 63368
0 63370 7 1 2 63366 63369
0 63371 5 1 1 63370
0 63372 7 1 2 63279 63371
0 63373 7 1 2 63266 63372
0 63374 7 1 2 62872 63373
0 63375 7 1 2 62594 63374
0 63376 7 1 2 62425 63375
0 63377 5 1 1 63376
0 63378 7 1 2 97431 63377
0 63379 5 1 1 63378
0 63380 7 1 2 65707 99094
0 63381 5 1 1 63380
0 63382 7 1 2 82539 93329
0 63383 5 1 1 63382
0 63384 7 1 2 63381 63383
0 63385 5 1 1 63384
0 63386 7 1 2 91427 90451
0 63387 7 2 2 98355 63386
0 63388 5 1 1 107608
0 63389 7 1 2 106955 107609
0 63390 5 1 1 63389
0 63391 7 1 2 103042 96227
0 63392 5 1 1 63391
0 63393 7 1 2 90593 77780
0 63394 7 1 2 95258 63393
0 63395 5 1 1 63394
0 63396 7 1 2 63392 63395
0 63397 5 1 1 63396
0 63398 7 1 2 63833 63397
0 63399 5 1 1 63398
0 63400 7 1 2 94596 77758
0 63401 7 1 2 92562 63400
0 63402 5 1 1 63401
0 63403 7 1 2 69038 63402
0 63404 7 1 2 63399 63403
0 63405 5 1 1 63404
0 63406 7 1 2 63948 107315
0 63407 5 1 1 63406
0 63408 7 1 2 67494 63407
0 63409 7 1 2 63405 63408
0 63410 5 1 1 63409
0 63411 7 1 2 65668 76815
0 63412 7 1 2 87758 63411
0 63413 7 1 2 106522 63412
0 63414 5 1 1 63413
0 63415 7 1 2 63410 63414
0 63416 5 1 1 63415
0 63417 7 1 2 106956 63416
0 63418 5 1 1 63417
0 63419 7 1 2 98041 96134
0 63420 7 1 2 100410 63419
0 63421 5 1 1 63420
0 63422 7 1 2 84603 102433
0 63423 5 1 1 63422
0 63424 7 1 2 17809 63423
0 63425 5 1 1 63424
0 63426 7 1 2 97137 106525
0 63427 7 1 2 63425 63426
0 63428 5 1 1 63427
0 63429 7 1 2 63421 63428
0 63430 5 1 1 63429
0 63431 7 1 2 63834 63430
0 63432 5 1 1 63431
0 63433 7 1 2 70307 87424
0 63434 7 1 2 86411 89500
0 63435 7 1 2 63433 63434
0 63436 7 1 2 106523 63435
0 63437 5 1 1 63436
0 63438 7 1 2 63432 63437
0 63439 5 1 1 63438
0 63440 7 1 2 65547 63439
0 63441 5 1 1 63440
0 63442 7 1 2 78731 98600
0 63443 7 1 2 101616 63442
0 63444 7 1 2 101739 63443
0 63445 5 1 1 63444
0 63446 7 1 2 63441 63445
0 63447 7 1 2 63418 63446
0 63448 5 1 1 63447
0 63449 7 1 2 72850 63448
0 63450 5 1 1 63449
0 63451 7 1 2 63390 63450
0 63452 5 1 1 63451
0 63453 7 1 2 68742 63452
0 63454 5 1 1 63453
0 63455 7 1 2 102279 107313
0 63456 5 1 1 63455
0 63457 7 1 2 67150 106421
0 63458 7 1 2 106994 63457
0 63459 5 1 1 63458
0 63460 7 1 2 63456 63459
0 63461 5 1 1 63460
0 63462 7 1 2 96782 63461
0 63463 5 1 1 63462
0 63464 7 1 2 63463 63388
0 63465 5 1 1 63464
0 63466 7 1 2 84921 63465
0 63467 5 1 1 63466
0 63468 7 1 2 97446 107329
0 63469 7 1 2 107480 63468
0 63470 5 1 1 63469
0 63471 7 1 2 63467 63470
0 63472 5 1 1 63471
0 63473 7 1 2 70308 63472
0 63474 5 1 1 63473
0 63475 7 1 2 88357 101787
0 63476 7 1 2 106232 63475
0 63477 7 1 2 107510 63476
0 63478 5 1 1 63477
0 63479 7 1 2 63474 63478
0 63480 7 1 2 63454 63479
0 63481 5 1 1 63480
0 63482 7 1 2 107393 63481
0 63483 5 1 1 63482
0 63484 7 1 2 90466 85041
0 63485 5 1 1 63484
0 63486 7 1 2 86549 88654
0 63487 5 1 1 63486
0 63488 7 1 2 63485 63487
0 63489 5 1 1 63488
0 63490 7 1 2 96946 63489
0 63491 5 1 1 63490
0 63492 7 1 2 104883 107227
0 63493 5 1 1 63492
0 63494 7 1 2 63491 63493
0 63495 5 1 1 63494
0 63496 7 1 2 102913 63495
0 63497 5 1 1 63496
0 63498 7 2 2 63949 72851
0 63499 7 1 2 96947 97094
0 63500 7 1 2 107610 63499
0 63501 7 1 2 97804 63500
0 63502 5 1 1 63501
0 63503 7 1 2 63497 63502
0 63504 5 1 1 63503
0 63505 7 1 2 103020 63504
0 63506 5 1 1 63505
0 63507 7 1 2 27524 107356
0 63508 5 1 1 63507
0 63509 7 1 2 96783 78116
0 63510 7 1 2 107481 63509
0 63511 7 1 2 63508 63510
0 63512 5 1 1 63511
0 63513 7 1 2 63506 63512
0 63514 5 1 1 63513
0 63515 7 1 2 107494 63514
0 63516 5 1 1 63515
0 63517 7 1 2 99226 107155
0 63518 7 1 2 107239 63517
0 63519 5 1 1 63518
0 63520 7 1 2 92831 89695
0 63521 7 1 2 104884 63520
0 63522 7 1 2 85370 63521
0 63523 5 1 1 63522
0 63524 7 1 2 63519 63523
0 63525 5 1 1 63524
0 63526 7 1 2 63835 63525
0 63527 5 1 1 63526
0 63528 7 1 2 98582 92143
0 63529 7 1 2 88647 63528
0 63530 7 1 2 106520 63529
0 63531 5 1 1 63530
0 63532 7 1 2 63527 63531
0 63533 5 1 1 63532
0 63534 7 1 2 70586 63533
0 63535 5 1 1 63534
0 63536 7 1 2 83352 95471
0 63537 7 1 2 84636 63536
0 63538 7 1 2 84763 63537
0 63539 5 1 1 63538
0 63540 7 1 2 63535 63539
0 63541 5 1 1 63540
0 63542 7 1 2 72504 63541
0 63543 5 1 1 63542
0 63544 7 1 2 96784 77781
0 63545 7 1 2 103174 63544
0 63546 7 1 2 102366 95957
0 63547 7 1 2 63545 63546
0 63548 5 1 1 63547
0 63549 7 1 2 63543 63548
0 63550 5 1 1 63549
0 63551 7 1 2 32689 7068
0 63552 7 1 2 106983 63551
0 63553 7 1 2 63550 63552
0 63554 5 1 1 63553
0 63555 7 1 2 63516 63554
0 63556 7 1 2 63483 63555
0 63557 5 1 1 63556
0 63558 7 1 2 67016 63557
0 63559 5 1 1 63558
0 63560 7 1 2 104514 92454
0 63561 5 1 1 63560
0 63562 7 1 2 96948 107529
0 63563 5 1 1 63562
0 63564 7 1 2 63561 63563
0 63565 5 1 1 63564
0 63566 7 1 2 107403 63565
0 63567 5 1 1 63566
0 63568 7 1 2 96988 107345
0 63569 5 1 1 63568
0 63570 7 1 2 107443 63569
0 63571 5 1 1 63570
0 63572 7 1 2 64009 102280
0 63573 7 1 2 102570 63572
0 63574 7 1 2 63571 63573
0 63575 5 1 1 63574
0 63576 7 1 2 63567 63575
0 63577 5 1 1 63576
0 63578 7 1 2 104677 63577
0 63579 5 1 1 63578
0 63580 7 1 2 102702 91183
0 63581 5 1 1 63580
0 63582 7 1 2 99676 96845
0 63583 5 1 1 63582
0 63584 7 1 2 63581 63583
0 63585 5 1 1 63584
0 63586 7 1 2 73304 88037
0 63587 7 1 2 106246 63586
0 63588 7 1 2 63585 63587
0 63589 5 1 1 63588
0 63590 7 1 2 72209 104885
0 63591 7 1 2 107506 63590
0 63592 5 1 1 63591
0 63593 7 1 2 63589 63592
0 63594 5 1 1 63593
0 63595 7 1 2 96949 63594
0 63596 5 1 1 63595
0 63597 7 1 2 102777 79011
0 63598 7 1 2 104891 93316
0 63599 7 1 2 63597 63598
0 63600 5 1 1 63599
0 63601 7 1 2 63596 63600
0 63602 5 1 1 63601
0 63603 7 1 2 84894 63602
0 63604 5 1 1 63603
0 63605 7 2 2 84691 98070
0 63606 7 1 2 99677 107612
0 63607 5 1 1 63606
0 63608 7 1 2 96585 107165
0 63609 5 1 1 63608
0 63610 7 1 2 63607 63609
0 63611 5 1 1 63610
0 63612 7 1 2 81952 63611
0 63613 5 1 1 63612
0 63614 7 1 2 107275 107613
0 63615 5 1 1 63614
0 63616 7 1 2 63613 63615
0 63617 5 1 1 63616
0 63618 7 1 2 96989 63617
0 63619 5 1 1 63618
0 63620 7 1 2 100147 98071
0 63621 7 1 2 106624 63620
0 63622 7 1 2 107346 63621
0 63623 5 1 1 63622
0 63624 7 1 2 63619 63623
0 63625 5 1 1 63624
0 63626 7 1 2 67151 63625
0 63627 5 1 1 63626
0 63628 7 1 2 104828 107358
0 63629 5 1 1 63628
0 63630 7 1 2 83693 98584
0 63631 5 1 1 63630
0 63632 7 1 2 93800 63631
0 63633 7 1 2 106627 63632
0 63634 5 1 1 63633
0 63635 7 1 2 63629 63634
0 63636 5 1 1 63635
0 63637 7 1 2 96440 107495
0 63638 7 1 2 63636 63637
0 63639 5 1 1 63638
0 63640 7 1 2 63627 63639
0 63641 5 1 1 63640
0 63642 7 1 2 73305 63641
0 63643 5 1 1 63642
0 63644 7 1 2 91778 87613
0 63645 7 1 2 106807 63644
0 63646 7 1 2 106447 63645
0 63647 7 1 2 96294 63646
0 63648 5 1 1 63647
0 63649 7 1 2 63643 63648
0 63650 5 1 1 63649
0 63651 7 1 2 76816 63650
0 63652 5 1 1 63651
0 63653 7 1 2 63604 63652
0 63654 5 1 1 63653
0 63655 7 1 2 69039 63654
0 63656 5 1 1 63655
0 63657 7 1 2 91490 107522
0 63658 7 1 2 107397 63657
0 63659 5 1 1 63658
0 63660 7 1 2 96533 107496
0 63661 7 1 2 87217 63660
0 63662 7 1 2 105100 63661
0 63663 5 1 1 63662
0 63664 7 1 2 63659 63663
0 63665 5 1 1 63664
0 63666 7 1 2 107561 63665
0 63667 5 1 1 63666
0 63668 7 1 2 68230 106792
0 63669 7 1 2 103130 63668
0 63670 7 1 2 97491 63669
0 63671 5 1 1 63670
0 63672 7 1 2 73306 92144
0 63673 7 1 2 97249 63672
0 63674 5 1 1 63673
0 63675 7 1 2 90594 91423
0 63676 5 1 1 63675
0 63677 7 1 2 63674 63676
0 63678 5 1 1 63677
0 63679 7 1 2 96990 107497
0 63680 7 1 2 63678 63679
0 63681 5 1 1 63680
0 63682 7 1 2 63671 63681
0 63683 5 1 1 63682
0 63684 7 1 2 81953 63683
0 63685 5 1 1 63684
0 63686 7 1 2 96950 96441
0 63687 7 1 2 107523 63686
0 63688 7 1 2 87543 63687
0 63689 5 1 1 63688
0 63690 7 1 2 63685 63689
0 63691 5 1 1 63690
0 63692 7 1 2 107611 63691
0 63693 5 1 1 63692
0 63694 7 1 2 63667 63693
0 63695 7 1 2 63656 63694
0 63696 5 1 1 63695
0 63697 7 1 2 68907 63696
0 63698 5 1 1 63697
0 63699 7 1 2 63579 63698
0 63700 5 1 1 63699
0 63701 7 1 2 72079 63700
0 63702 5 1 1 63701
0 63703 7 1 2 63559 63702
0 63704 5 1 1 63703
0 63705 7 1 2 63385 63704
0 63706 5 1 1 63705
0 63707 7 1 2 63379 63706
0 63708 7 1 2 62163 63707
0 63709 7 1 2 61777 63708
0 63710 7 1 2 61376 63709
0 63711 7 1 2 60442 63710
0 63712 5 1 1 63711
0 63713 7 1 2 103629 63712
0 63714 5 1 1 63713
0 63715 7 1 2 58536 63714
0 63716 7 1 2 55782 63715
0 63717 7 1 2 42233 63716
0 63718 7 1 2 22010 63717
3 129999 5 0 1 63718
