1 0 0 8 0
2 32 1 0
2 1959 1 0
2 1960 1 0
2 1961 1 0
2 1962 1 0
2 1963 1 0
2 1964 1 0
2 1965 1 0
1 1 0 10 0
2 1966 1 1
2 1967 1 1
2 1968 1 1
2 1969 1 1
2 1970 1 1
2 1971 1 1
2 1972 1 1
2 1973 1 1
2 1974 1 1
2 1975 1 1
1 2 0 10 0
2 1976 1 2
2 1977 1 2
2 1978 1 2
2 1979 1 2
2 1980 1 2
2 1981 1 2
2 1982 1 2
2 1983 1 2
2 1984 1 2
2 1985 1 2
1 3 0 11 0
2 1986 1 3
2 1987 1 3
2 1988 1 3
2 1989 1 3
2 1990 1 3
2 1991 1 3
2 1992 1 3
2 1993 1 3
2 1994 1 3
2 1995 1 3
2 1996 1 3
1 4 0 10 0
2 1997 1 4
2 1998 1 4
2 1999 1 4
2 2000 1 4
2 2001 1 4
2 2002 1 4
2 2003 1 4
2 2004 1 4
2 2005 1 4
2 2006 1 4
1 5 0 11 0
2 2007 1 5
2 2008 1 5
2 2009 1 5
2 2010 1 5
2 2011 1 5
2 2012 1 5
2 2013 1 5
2 2014 1 5
2 2015 1 5
2 2016 1 5
2 2017 1 5
1 6 0 10 0
2 2018 1 6
2 2019 1 6
2 2020 1 6
2 2021 1 6
2 2022 1 6
2 2023 1 6
2 2024 1 6
2 2025 1 6
2 2026 1 6
2 2027 1 6
1 7 0 10 0
2 2028 1 7
2 2029 1 7
2 2030 1 7
2 2031 1 7
2 2032 1 7
2 2033 1 7
2 2034 1 7
2 2035 1 7
2 2036 1 7
2 2037 1 7
1 8 0 10 0
2 2038 1 8
2 2039 1 8
2 2040 1 8
2 2041 1 8
2 2042 1 8
2 2043 1 8
2 2044 1 8
2 2045 1 8
2 2046 1 8
2 2047 1 8
1 9 0 10 0
2 2048 1 9
2 2049 1 9
2 2050 1 9
2 2051 1 9
2 2052 1 9
2 2053 1 9
2 2054 1 9
2 2055 1 9
2 2056 1 9
2 2057 1 9
1 10 0 11 0
2 2058 1 10
2 2059 1 10
2 2060 1 10
2 2061 1 10
2 2062 1 10
2 2063 1 10
2 2064 1 10
2 2065 1 10
2 2066 1 10
2 2067 1 10
2 2068 1 10
1 11 0 10 0
2 2069 1 11
2 2070 1 11
2 2071 1 11
2 2072 1 11
2 2073 1 11
2 2074 1 11
2 2075 1 11
2 2076 1 11
2 2077 1 11
2 2078 1 11
1 12 0 10 0
2 2079 1 12
2 2080 1 12
2 2081 1 12
2 2082 1 12
2 2083 1 12
2 2084 1 12
2 2085 1 12
2 2086 1 12
2 2087 1 12
2 2088 1 12
1 13 0 10 0
2 2089 1 13
2 2090 1 13
2 2091 1 13
2 2092 1 13
2 2093 1 13
2 2094 1 13
2 2095 1 13
2 2096 1 13
2 2097 1 13
2 2098 1 13
1 14 0 10 0
2 2099 1 14
2 2100 1 14
2 2101 1 14
2 2102 1 14
2 2103 1 14
2 2104 1 14
2 2105 1 14
2 2106 1 14
2 2107 1 14
2 2108 1 14
1 15 0 10 0
2 2109 1 15
2 2110 1 15
2 2111 1 15
2 2112 1 15
2 2113 1 15
2 2114 1 15
2 2115 1 15
2 2116 1 15
2 2117 1 15
2 2118 1 15
1 16 0 3 0
2 2119 1 16
2 2120 1 16
2 2121 1 16
1 17 0 3 0
2 2122 1 17
2 2123 1 17
2 2124 1 17
1 18 0 3 0
2 2125 1 18
2 2126 1 18
2 2127 1 18
1 19 0 3 0
2 2128 1 19
2 2129 1 19
2 2130 1 19
1 20 0 3 0
2 2131 1 20
2 2132 1 20
2 2133 1 20
1 21 0 3 0
2 2134 1 21
2 2135 1 21
2 2136 1 21
1 22 0 3 0
2 2137 1 22
2 2138 1 22
2 2139 1 22
1 23 0 3 0
2 2140 1 23
2 2141 1 23
2 2142 1 23
1 24 0 3 0
2 2143 1 24
2 2144 1 24
2 2145 1 24
1 25 0 3 0
2 2146 1 25
2 2147 1 25
2 2148 1 25
1 26 0 3 0
2 2149 1 26
2 2150 1 26
2 2151 1 26
1 27 0 3 0
2 2152 1 27
2 2153 1 27
2 2154 1 27
1 28 0 4 0
2 2155 1 28
2 2156 1 28
2 2157 1 28
2 2158 1 28
1 29 0 3 0
2 2159 1 29
2 2160 1 29
2 2161 1 29
1 30 0 4 0
2 2162 1 30
2 2163 1 30
2 2164 1 30
2 2165 1 30
1 31 0 4 0
2 2166 1 31
2 2167 1 31
2 2168 1 31
2 2169 1 31
2 2170 1 33
2 2171 1 33
2 2172 1 34
2 2173 1 34
2 2174 1 35
2 2175 1 35
2 2176 1 36
2 2177 1 36
2 2178 1 37
2 2179 1 37
2 2180 1 38
2 2181 1 38
2 2182 1 39
2 2183 1 39
2 2184 1 40
2 2185 1 40
2 2186 1 41
2 2187 1 41
2 2188 1 42
2 2189 1 42
2 2190 1 43
2 2191 1 43
2 2192 1 44
2 2193 1 44
2 2194 1 45
2 2195 1 45
2 2196 1 46
2 2197 1 46
2 2198 1 47
2 2199 1 47
2 2200 1 48
2 2201 1 48
2 2202 1 48
2 2203 1 49
2 2204 1 49
2 2205 1 49
2 2206 1 50
2 2207 1 50
2 2208 1 50
2 2209 1 51
2 2210 1 51
2 2211 1 51
2 2212 1 52
2 2213 1 52
2 2214 1 52
2 2215 1 53
2 2216 1 53
2 2217 1 53
2 2218 1 54
2 2219 1 54
2 2220 1 54
2 2221 1 55
2 2222 1 55
2 2223 1 55
2 2224 1 56
2 2225 1 56
2 2226 1 56
2 2227 1 57
2 2228 1 57
2 2229 1 57
2 2230 1 58
2 2231 1 58
2 2232 1 58
2 2233 1 59
2 2234 1 59
2 2235 1 59
2 2236 1 60
2 2237 1 60
2 2238 1 60
2 2239 1 60
2 2240 1 61
2 2241 1 61
2 2242 1 61
2 2243 1 62
2 2244 1 62
2 2245 1 63
2 2246 1 63
2 2247 1 64
2 2248 1 64
2 2249 1 66
2 2250 1 66
2 2251 1 66
2 2252 1 68
2 2253 1 68
2 2254 1 74
2 2255 1 74
2 2256 1 76
2 2257 1 76
2 2258 1 81
2 2259 1 81
2 2260 1 84
2 2261 1 84
2 2262 1 87
2 2263 1 87
2 2264 1 89
2 2265 1 89
2 2266 1 90
2 2267 1 90
2 2268 1 95
2 2269 1 95
2 2270 1 98
2 2271 1 98
2 2272 1 103
2 2273 1 103
2 2274 1 104
2 2275 1 104
2 2276 1 105
2 2277 1 105
2 2278 1 108
2 2279 1 108
2 2280 1 111
2 2281 1 111
2 2282 1 113
2 2283 1 113
2 2284 1 114
2 2285 1 114
2 2286 1 119
2 2287 1 119
2 2288 1 122
2 2289 1 122
2 2290 1 127
2 2291 1 127
2 2292 1 127
2 2293 1 129
2 2294 1 129
2 2295 1 132
2 2296 1 132
2 2297 1 135
2 2298 1 135
2 2299 1 137
2 2300 1 137
2 2301 1 138
2 2302 1 138
2 2303 1 143
2 2304 1 143
2 2305 1 146
2 2306 1 146
2 2307 1 151
2 2308 1 151
2 2309 1 151
2 2310 1 153
2 2311 1 153
2 2312 1 156
2 2313 1 156
2 2314 1 159
2 2315 1 159
2 2316 1 161
2 2317 1 161
2 2318 1 162
2 2319 1 162
2 2320 1 167
2 2321 1 167
2 2322 1 170
2 2323 1 170
2 2324 1 175
2 2325 1 175
2 2326 1 175
2 2327 1 177
2 2328 1 177
2 2329 1 180
2 2330 1 180
2 2331 1 183
2 2332 1 183
2 2333 1 185
2 2334 1 185
2 2335 1 186
2 2336 1 186
2 2337 1 191
2 2338 1 191
2 2339 1 194
2 2340 1 194
2 2341 1 199
2 2342 1 199
2 2343 1 199
2 2344 1 201
2 2345 1 201
2 2346 1 204
2 2347 1 204
2 2348 1 207
2 2349 1 207
2 2350 1 209
2 2351 1 209
2 2352 1 210
2 2353 1 210
2 2354 1 215
2 2355 1 215
2 2356 1 218
2 2357 1 218
2 2358 1 223
2 2359 1 223
2 2360 1 223
2 2361 1 225
2 2362 1 225
2 2363 1 228
2 2364 1 228
2 2365 1 231
2 2366 1 231
2 2367 1 233
2 2368 1 233
2 2369 1 234
2 2370 1 234
2 2371 1 239
2 2372 1 239
2 2373 1 242
2 2374 1 242
2 2375 1 247
2 2376 1 247
2 2377 1 247
2 2378 1 249
2 2379 1 249
2 2380 1 252
2 2381 1 252
2 2382 1 255
2 2383 1 255
2 2384 1 257
2 2385 1 257
2 2386 1 258
2 2387 1 258
2 2388 1 263
2 2389 1 263
2 2390 1 266
2 2391 1 266
2 2392 1 271
2 2393 1 271
2 2394 1 271
2 2395 1 273
2 2396 1 273
2 2397 1 276
2 2398 1 276
2 2399 1 279
2 2400 1 279
2 2401 1 281
2 2402 1 281
2 2403 1 282
2 2404 1 282
2 2405 1 287
2 2406 1 287
2 2407 1 290
2 2408 1 290
2 2409 1 295
2 2410 1 295
2 2411 1 295
2 2412 1 297
2 2413 1 297
2 2414 1 300
2 2415 1 300
2 2416 1 303
2 2417 1 303
2 2418 1 305
2 2419 1 305
2 2420 1 306
2 2421 1 306
2 2422 1 311
2 2423 1 311
2 2424 1 314
2 2425 1 314
2 2426 1 319
2 2427 1 319
2 2428 1 319
2 2429 1 321
2 2430 1 321
2 2431 1 324
2 2432 1 324
2 2433 1 327
2 2434 1 327
2 2435 1 329
2 2436 1 329
2 2437 1 330
2 2438 1 330
2 2439 1 335
2 2440 1 335
2 2441 1 338
2 2442 1 338
2 2443 1 343
2 2444 1 343
2 2445 1 343
2 2446 1 345
2 2447 1 345
2 2448 1 348
2 2449 1 348
2 2450 1 351
2 2451 1 351
2 2452 1 353
2 2453 1 353
2 2454 1 354
2 2455 1 354
2 2456 1 359
2 2457 1 359
2 2458 1 362
2 2459 1 362
2 2460 1 367
2 2461 1 367
2 2462 1 367
2 2463 1 369
2 2464 1 369
2 2465 1 372
2 2466 1 372
2 2467 1 375
2 2468 1 375
2 2469 1 377
2 2470 1 377
2 2471 1 378
2 2472 1 378
2 2473 1 383
2 2474 1 383
2 2475 1 386
2 2476 1 386
2 2477 1 391
2 2478 1 391
2 2479 1 391
2 2480 1 393
2 2481 1 393
2 2482 1 396
2 2483 1 396
2 2484 1 399
2 2485 1 399
2 2486 1 401
2 2487 1 401
2 2488 1 402
2 2489 1 402
2 2490 1 407
2 2491 1 407
2 2492 1 410
2 2493 1 410
2 2494 1 415
2 2495 1 415
2 2496 1 415
2 2497 1 417
2 2498 1 417
2 2499 1 420
2 2500 1 420
2 2501 1 423
2 2502 1 423
2 2503 1 425
2 2504 1 425
2 2505 1 426
2 2506 1 426
2 2507 1 431
2 2508 1 431
2 2509 1 434
2 2510 1 434
2 2511 1 439
2 2512 1 439
2 2513 1 439
2 2514 1 441
2 2515 1 441
2 2516 1 444
2 2517 1 444
2 2518 1 447
2 2519 1 447
2 2520 1 449
2 2521 1 449
2 2522 1 450
2 2523 1 450
2 2524 1 455
2 2525 1 455
2 2526 1 458
2 2527 1 458
2 2528 1 463
2 2529 1 463
2 2530 1 463
2 2531 1 465
2 2532 1 465
2 2533 1 468
2 2534 1 468
2 2535 1 471
2 2536 1 471
2 2537 1 473
2 2538 1 473
2 2539 1 474
2 2540 1 474
2 2541 1 479
2 2542 1 479
2 2543 1 482
2 2544 1 482
2 2545 1 487
2 2546 1 487
2 2547 1 487
2 2548 1 489
2 2549 1 489
2 2550 1 492
2 2551 1 492
2 2552 1 495
2 2553 1 495
2 2554 1 497
2 2555 1 497
2 2556 1 498
2 2557 1 498
2 2558 1 503
2 2559 1 503
2 2560 1 506
2 2561 1 506
2 2562 1 511
2 2563 1 511
2 2564 1 511
2 2565 1 513
2 2566 1 513
2 2567 1 516
2 2568 1 516
2 2569 1 519
2 2570 1 519
2 2571 1 521
2 2572 1 521
2 2573 1 522
2 2574 1 522
2 2575 1 527
2 2576 1 527
2 2577 1 530
2 2578 1 530
2 2579 1 535
2 2580 1 535
2 2581 1 535
2 2582 1 537
2 2583 1 537
2 2584 1 540
2 2585 1 540
2 2586 1 543
2 2587 1 543
2 2588 1 545
2 2589 1 545
2 2590 1 546
2 2591 1 546
2 2592 1 551
2 2593 1 551
2 2594 1 554
2 2595 1 554
2 2596 1 559
2 2597 1 559
2 2598 1 559
2 2599 1 561
2 2600 1 561
2 2601 1 564
2 2602 1 564
2 2603 1 567
2 2604 1 567
2 2605 1 569
2 2606 1 569
2 2607 1 570
2 2608 1 570
2 2609 1 575
2 2610 1 575
2 2611 1 578
2 2612 1 578
2 2613 1 583
2 2614 1 583
2 2615 1 583
2 2616 1 585
2 2617 1 585
2 2618 1 588
2 2619 1 588
2 2620 1 591
2 2621 1 591
2 2622 1 593
2 2623 1 593
2 2624 1 594
2 2625 1 594
2 2626 1 599
2 2627 1 599
2 2628 1 602
2 2629 1 602
2 2630 1 607
2 2631 1 607
2 2632 1 607
2 2633 1 609
2 2634 1 609
2 2635 1 612
2 2636 1 612
2 2637 1 615
2 2638 1 615
2 2639 1 617
2 2640 1 617
2 2641 1 618
2 2642 1 618
2 2643 1 623
2 2644 1 623
2 2645 1 626
2 2646 1 626
2 2647 1 631
2 2648 1 631
2 2649 1 631
2 2650 1 633
2 2651 1 633
2 2652 1 636
2 2653 1 636
2 2654 1 639
2 2655 1 639
2 2656 1 641
2 2657 1 641
2 2658 1 642
2 2659 1 642
2 2660 1 647
2 2661 1 647
2 2662 1 650
2 2663 1 650
2 2664 1 655
2 2665 1 655
2 2666 1 655
2 2667 1 657
2 2668 1 657
2 2669 1 660
2 2670 1 660
2 2671 1 663
2 2672 1 663
2 2673 1 665
2 2674 1 665
2 2675 1 666
2 2676 1 666
2 2677 1 671
2 2678 1 671
2 2679 1 674
2 2680 1 674
2 2681 1 679
2 2682 1 679
2 2683 1 679
2 2684 1 681
2 2685 1 681
2 2686 1 686
2 2687 1 686
2 2688 1 687
2 2689 1 687
2 2690 1 687
2 2691 1 688
2 2692 1 688
2 2693 1 689
2 2694 1 689
2 2695 1 690
2 2696 1 690
2 2697 1 695
2 2698 1 695
2 2699 1 698
2 2700 1 698
2 2701 1 703
2 2702 1 703
2 2703 1 703
2 2704 1 711
2 2705 1 711
2 2706 1 714
2 2707 1 714
2 2708 1 717
2 2709 1 717
2 2710 1 728
2 2711 1 728
2 2712 1 739
2 2713 1 739
2 2714 1 741
2 2715 1 741
2 2716 1 743
2 2717 1 743
2 2718 1 744
2 2719 1 744
2 2720 1 745
2 2721 1 745
2 2722 1 747
2 2723 1 747
2 2724 1 750
2 2725 1 750
2 2726 1 753
2 2727 1 753
2 2728 1 756
2 2729 1 756
2 2730 1 757
2 2731 1 757
2 2732 1 759
2 2733 1 759
2 2734 1 761
2 2735 1 761
2 2736 1 767
2 2737 1 767
2 2738 1 770
2 2739 1 770
2 2740 1 770
2 2741 1 774
2 2742 1 774
2 2743 1 775
2 2744 1 775
2 2745 1 777
2 2746 1 777
2 2747 1 780
2 2748 1 780
2 2749 1 781
2 2750 1 781
2 2751 1 785
2 2752 1 785
2 2753 1 788
2 2754 1 788
2 2755 1 789
2 2756 1 789
2 2757 1 793
2 2758 1 793
2 2759 1 796
2 2760 1 796
2 2761 1 797
2 2762 1 797
2 2763 1 801
2 2764 1 801
2 2765 1 804
2 2766 1 804
2 2767 1 805
2 2768 1 805
2 2769 1 807
2 2770 1 807
2 2771 1 810
2 2772 1 810
2 2773 1 811
2 2774 1 811
2 2775 1 815
2 2776 1 815
2 2777 1 818
2 2778 1 818
2 2779 1 819
2 2780 1 819
2 2781 1 823
2 2782 1 823
2 2783 1 826
2 2784 1 826
2 2785 1 827
2 2786 1 827
2 2787 1 831
2 2788 1 831
2 2789 1 834
2 2790 1 834
2 2791 1 835
2 2792 1 835
2 2793 1 839
2 2794 1 839
2 2795 1 842
2 2796 1 842
2 2797 1 843
2 2798 1 843
2 2799 1 847
2 2800 1 847
2 2801 1 850
2 2802 1 850
2 2803 1 851
2 2804 1 851
2 2805 1 855
2 2806 1 855
2 2807 1 858
2 2808 1 858
2 2809 1 859
2 2810 1 859
2 2811 1 863
2 2812 1 863
2 2813 1 866
2 2814 1 866
2 2815 1 867
2 2816 1 867
2 2817 1 869
2 2818 1 869
2 2819 1 871
2 2820 1 871
2 2821 1 872
2 2822 1 872
2 2823 1 873
2 2824 1 873
2 2825 1 874
2 2826 1 874
2 2827 1 875
2 2828 1 875
2 2829 1 878
2 2830 1 878
2 2831 1 879
2 2832 1 879
2 2833 1 883
2 2834 1 883
2 2835 1 886
2 2836 1 886
2 2837 1 887
2 2838 1 887
2 2839 1 891
2 2840 1 891
2 2841 1 894
2 2842 1 894
2 2843 1 895
2 2844 1 895
2 2845 1 899
2 2846 1 899
2 2847 1 902
2 2848 1 902
2 2849 1 903
2 2850 1 903
2 2851 1 907
2 2852 1 907
2 2853 1 910
2 2854 1 910
2 2855 1 911
2 2856 1 911
2 2857 1 915
2 2858 1 915
2 2859 1 918
2 2860 1 918
2 2861 1 919
2 2862 1 919
2 2863 1 923
2 2864 1 923
2 2865 1 926
2 2866 1 926
2 2867 1 927
2 2868 1 927
2 2869 1 931
2 2870 1 931
2 2871 1 934
2 2872 1 934
2 2873 1 935
2 2874 1 935
2 2875 1 937
2 2876 1 937
2 2877 1 940
2 2878 1 940
2 2879 1 943
2 2880 1 943
2 2881 1 947
2 2882 1 947
2 2883 1 950
2 2884 1 950
2 2885 1 951
2 2886 1 951
2 2887 1 955
2 2888 1 955
2 2889 1 958
2 2890 1 958
2 2891 1 959
2 2892 1 959
2 2893 1 961
2 2894 1 961
2 2895 1 964
2 2896 1 964
2 2897 1 965
2 2898 1 965
2 2899 1 967
2 2900 1 967
2 2901 1 973
2 2902 1 973
2 2903 1 976
2 2904 1 976
2 2905 1 979
2 2906 1 979
2 2907 1 982
2 2908 1 982
2 2909 1 985
2 2910 1 985
2 2911 1 989
2 2912 1 989
2 2913 1 992
2 2914 1 992
2 2915 1 993
2 2916 1 993
2 2917 1 997
2 2918 1 997
2 2919 1 1000
2 2920 1 1000
2 2921 1 1001
2 2922 1 1001
2 2923 1 1003
2 2924 1 1003
2 2925 1 1006
2 2926 1 1006
2 2927 1 1009
2 2928 1 1009
2 2929 1 1013
2 2930 1 1013
2 2931 1 1016
2 2932 1 1016
2 2933 1 1017
2 2934 1 1017
2 2935 1 1021
2 2936 1 1021
2 2937 1 1024
2 2938 1 1024
2 2939 1 1025
2 2940 1 1025
2 2941 1 1029
2 2942 1 1029
2 2943 1 1032
2 2944 1 1032
2 2945 1 1033
2 2946 1 1033
2 2947 1 1037
2 2948 1 1037
2 2949 1 1040
2 2950 1 1040
2 2951 1 1041
2 2952 1 1041
2 2953 1 1045
2 2954 1 1045
2 2955 1 1048
2 2956 1 1048
2 2957 1 1049
2 2958 1 1049
2 2959 1 1051
2 2960 1 1051
2 2961 1 1054
2 2962 1 1054
2 2963 1 1055
2 2964 1 1055
2 2965 1 1059
2 2966 1 1059
2 2967 1 1062
2 2968 1 1062
2 2969 1 1063
2 2970 1 1063
2 2971 1 1065
2 2972 1 1065
2 2973 1 1067
2 2974 1 1067
2 2975 1 1070
2 2976 1 1070
2 2977 1 1071
2 2978 1 1071
2 2979 1 1073
2 2980 1 1073
2 2981 1 1075
2 2982 1 1075
2 2983 1 1077
2 2984 1 1077
2 2985 1 1079
2 2986 1 1079
2 2987 1 1080
2 2988 1 1080
2 2989 1 1081
2 2990 1 1081
2 2991 1 1082
2 2992 1 1082
2 2993 1 1083
2 2994 1 1083
2 2995 1 1084
2 2996 1 1084
2 2997 1 1085
2 2998 1 1085
2 2999 1 1086
2 3000 1 1086
2 3001 1 1088
2 3002 1 1088
2 3003 1 1091
2 3004 1 1091
2 3005 1 1095
2 3006 1 1095
2 3007 1 1098
2 3008 1 1098
2 3009 1 1101
2 3010 1 1101
2 3011 1 1105
2 3012 1 1105
2 3013 1 1108
2 3014 1 1108
2 3015 1 1109
2 3016 1 1109
2 3017 1 1112
2 3018 1 1112
2 3019 1 1113
2 3020 1 1113
2 3021 1 1117
2 3022 1 1117
2 3023 1 1120
2 3024 1 1120
2 3025 1 1121
2 3026 1 1121
2 3027 1 1125
2 3028 1 1125
2 3029 1 1128
2 3030 1 1128
2 3031 1 1129
2 3032 1 1129
2 3033 1 1133
2 3034 1 1133
2 3035 1 1136
2 3036 1 1136
2 3037 1 1139
2 3038 1 1139
2 3039 1 1143
2 3040 1 1143
2 3041 1 1146
2 3042 1 1146
2 3043 1 1149
2 3044 1 1149
2 3045 1 1153
2 3046 1 1153
2 3047 1 1156
2 3048 1 1156
2 3049 1 1157
2 3050 1 1157
2 3051 1 1159
2 3052 1 1159
2 3053 1 1162
2 3054 1 1162
2 3055 1 1163
2 3056 1 1163
2 3057 1 1167
2 3058 1 1167
2 3059 1 1170
2 3060 1 1170
2 3061 1 1171
2 3062 1 1171
2 3063 1 1175
2 3064 1 1175
2 3065 1 1178
2 3066 1 1178
2 3067 1 1179
2 3068 1 1179
2 3069 1 1183
2 3070 1 1183
2 3071 1 1186
2 3072 1 1186
2 3073 1 1187
2 3074 1 1187
2 3075 1 1191
2 3076 1 1191
2 3077 1 1194
2 3078 1 1194
2 3079 1 1195
2 3080 1 1195
2 3081 1 1199
2 3082 1 1199
2 3083 1 1202
2 3084 1 1202
2 3085 1 1203
2 3086 1 1203
2 3087 1 1205
2 3088 1 1205
2 3089 1 1211
2 3090 1 1211
2 3091 1 1214
2 3092 1 1214
2 3093 1 1217
2 3094 1 1217
2 3095 1 1220
2 3096 1 1220
2 3097 1 1223
2 3098 1 1223
2 3099 1 1227
2 3100 1 1227
2 3101 1 1230
2 3102 1 1230
2 3103 1 1231
2 3104 1 1231
2 3105 1 1235
2 3106 1 1235
2 3107 1 1238
2 3108 1 1238
2 3109 1 1239
2 3110 1 1239
2 3111 1 1243
2 3112 1 1243
2 3113 1 1246
2 3114 1 1246
2 3115 1 1247
2 3116 1 1247
2 3117 1 1251
2 3118 1 1251
2 3119 1 1254
2 3120 1 1254
2 3121 1 1255
2 3122 1 1255
2 3123 1 1259
2 3124 1 1259
2 3125 1 1262
2 3126 1 1262
2 3127 1 1263
2 3128 1 1263
2 3129 1 1267
2 3130 1 1267
2 3131 1 1270
2 3132 1 1270
2 3133 1 1271
2 3134 1 1271
2 3135 1 1275
2 3136 1 1275
2 3137 1 1278
2 3138 1 1278
2 3139 1 1279
2 3140 1 1279
2 3141 1 1281
2 3142 1 1281
2 3143 1 1284
2 3144 1 1284
2 3145 1 1287
2 3146 1 1287
2 3147 1 1291
2 3148 1 1291
2 3149 1 1294
2 3150 1 1294
2 3151 1 1295
2 3152 1 1295
2 3153 1 1299
2 3154 1 1299
2 3155 1 1302
2 3156 1 1302
2 3157 1 1303
2 3158 1 1303
2 3159 1 1307
2 3160 1 1307
2 3161 1 1310
2 3162 1 1310
2 3163 1 1311
2 3164 1 1311
2 3165 1 1315
2 3166 1 1315
2 3167 1 1318
2 3168 1 1318
2 3169 1 1319
2 3170 1 1319
2 3171 1 1325
2 3172 1 1325
2 3173 1 1328
2 3174 1 1328
2 3175 1 1329
2 3176 1 1329
2 3177 1 1333
2 3178 1 1333
2 3179 1 1336
2 3180 1 1336
2 3181 1 1337
2 3182 1 1337
2 3183 1 1341
2 3184 1 1341
2 3185 1 1344
2 3186 1 1344
2 3187 1 1345
2 3188 1 1345
2 3189 1 1349
2 3190 1 1349
2 3191 1 1352
2 3192 1 1352
2 3193 1 1353
2 3194 1 1353
2 3195 1 1355
2 3196 1 1355
2 3197 1 1358
2 3198 1 1358
2 3199 1 1361
2 3200 1 1361
2 3201 1 1365
2 3202 1 1365
2 3203 1 1368
2 3204 1 1368
2 3205 1 1369
2 3206 1 1369
2 3207 1 1373
2 3208 1 1373
2 3209 1 1376
2 3210 1 1376
2 3211 1 1379
2 3212 1 1379
2 3213 1 1381
2 3214 1 1381
2 3215 1 1383
2 3216 1 1383
2 3217 1 1385
2 3218 1 1385
2 3219 1 1387
2 3220 1 1387
2 3221 1 1389
2 3222 1 1389
2 3223 1 1391
2 3224 1 1391
2 3225 1 1392
2 3226 1 1392
2 3227 1 1393
2 3228 1 1393
2 3229 1 1393
2 3230 1 1396
2 3231 1 1396
2 3232 1 1399
2 3233 1 1399
2 3234 1 1407
2 3235 1 1407
2 3236 1 1410
2 3237 1 1410
2 3238 1 1411
2 3239 1 1411
2 3240 1 1415
2 3241 1 1415
2 3242 1 1418
2 3243 1 1418
2 3244 1 1421
2 3245 1 1421
2 3246 1 1423
2 3247 1 1423
2 3248 1 1425
2 3249 1 1425
2 3250 1 1427
2 3251 1 1427
2 3252 1 1428
2 3253 1 1428
2 3254 1 1430
2 3255 1 1430
2 3256 1 1431
2 3257 1 1431
2 3258 1 1435
2 3259 1 1435
2 3260 1 1438
2 3261 1 1438
2 3262 1 1439
2 3263 1 1439
2 3264 1 1443
2 3265 1 1443
2 3266 1 1446
2 3267 1 1446
2 3268 1 1447
2 3269 1 1447
2 3270 1 1451
2 3271 1 1451
2 3272 1 1454
2 3273 1 1454
2 3274 1 1455
2 3275 1 1455
2 3276 1 1459
2 3277 1 1459
2 3278 1 1462
2 3279 1 1462
2 3280 1 1463
2 3281 1 1463
2 3282 1 1467
2 3283 1 1467
2 3284 1 1470
2 3285 1 1470
2 3286 1 1471
2 3287 1 1471
2 3288 1 1475
2 3289 1 1475
2 3290 1 1478
2 3291 1 1478
2 3292 1 1479
2 3293 1 1479
2 3294 1 1483
2 3295 1 1483
2 3296 1 1486
2 3297 1 1486
2 3298 1 1487
2 3299 1 1487
2 3300 1 1491
2 3301 1 1491
2 3302 1 1494
2 3303 1 1494
2 3304 1 1495
2 3305 1 1495
2 3306 1 1499
2 3307 1 1499
2 3308 1 1502
2 3309 1 1502
2 3310 1 1503
2 3311 1 1503
2 3312 1 1507
2 3313 1 1507
2 3314 1 1510
2 3315 1 1510
2 3316 1 1511
2 3317 1 1511
2 3318 1 1515
2 3319 1 1515
2 3320 1 1518
2 3321 1 1518
2 3322 1 1519
2 3323 1 1519
2 3324 1 1523
2 3325 1 1523
2 3326 1 1526
2 3327 1 1526
2 3328 1 1527
2 3329 1 1527
2 3330 1 1529
2 3331 1 1529
2 3332 1 1530
2 3333 1 1530
2 3334 1 1530
2 3335 1 1533
2 3336 1 1533
2 3337 1 1536
2 3338 1 1536
2 3339 1 1536
2 3340 1 1537
2 3341 1 1537
2 3342 1 1539
2 3343 1 1539
2 3344 1 1542
2 3345 1 1542
2 3346 1 1545
2 3347 1 1545
2 3348 1 1548
2 3349 1 1548
2 3350 1 1548
2 3351 1 1551
2 3352 1 1551
2 3353 1 1554
2 3354 1 1554
2 3355 1 1554
2 3356 1 1554
2 3357 1 1554
2 3358 1 1554
2 3359 1 1557
2 3360 1 1557
2 3361 1 1560
2 3362 1 1560
2 3363 1 1560
2 3364 1 1560
2 3365 1 1563
2 3366 1 1563
2 3367 1 1566
2 3368 1 1566
2 3369 1 1566
2 3370 1 1566
2 3371 1 1568
2 3372 1 1568
2 3373 1 1568
2 3374 1 1568
2 3375 1 1571
2 3376 1 1571
2 3377 1 1574
2 3378 1 1574
2 3379 1 1574
2 3380 1 1576
2 3381 1 1576
2 3382 1 1576
2 3383 1 1576
2 3384 1 1579
2 3385 1 1579
2 3386 1 1582
2 3387 1 1582
2 3388 1 1582
2 3389 1 1582
2 3390 1 1582
2 3391 1 1584
2 3392 1 1584
2 3393 1 1584
2 3394 1 1584
2 3395 1 1587
2 3396 1 1587
2 3397 1 1590
2 3398 1 1590
2 3399 1 1590
2 3400 1 1590
2 3401 1 1592
2 3402 1 1592
2 3403 1 1592
2 3404 1 1592
2 3405 1 1595
2 3406 1 1595
2 3407 1 1598
2 3408 1 1598
2 3409 1 1598
2 3410 1 1598
2 3411 1 1600
2 3412 1 1600
2 3413 1 1600
2 3414 1 1600
2 3415 1 1603
2 3416 1 1603
2 3417 1 1606
2 3418 1 1606
2 3419 1 1606
2 3420 1 1606
2 3421 1 1608
2 3422 1 1608
2 3423 1 1608
2 3424 1 1608
2 3425 1 1611
2 3426 1 1611
2 3427 1 1614
2 3428 1 1614
2 3429 1 1614
2 3430 1 1616
2 3431 1 1616
2 3432 1 1616
2 3433 1 1616
2 3434 1 1619
2 3435 1 1619
2 3436 1 1622
2 3437 1 1622
2 3438 1 1622
2 3439 1 1624
2 3440 1 1624
2 3441 1 1624
2 3442 1 1624
2 3443 1 1627
2 3444 1 1627
2 3445 1 1630
2 3446 1 1630
2 3447 1 1630
2 3448 1 1632
2 3449 1 1632
2 3450 1 1632
2 3451 1 1635
2 3452 1 1635
2 3453 1 1638
2 3454 1 1638
2 3455 1 1639
2 3456 1 1639
2 3457 1 1641
2 3458 1 1641
2 3459 1 1645
2 3460 1 1645
2 3461 1 1650
2 3462 1 1650
2 3463 1 1651
2 3464 1 1651
2 3465 1 1654
2 3466 1 1654
2 3467 1 1655
2 3468 1 1655
2 3469 1 1658
2 3470 1 1658
2 3471 1 1659
2 3472 1 1659
2 3473 1 1662
2 3474 1 1662
2 3475 1 1663
2 3476 1 1663
2 3477 1 1666
2 3478 1 1666
2 3479 1 1667
2 3480 1 1667
2 3481 1 1670
2 3482 1 1670
2 3483 1 1672
2 3484 1 1672
2 3485 1 1674
2 3486 1 1674
2 3487 1 1675
2 3488 1 1675
2 3489 1 1678
2 3490 1 1678
2 3491 1 1680
2 3492 1 1680
2 3493 1 1682
2 3494 1 1682
2 3495 1 1686
2 3496 1 1686
2 3497 1 1688
2 3498 1 1688
2 3499 1 1688
2 3500 1 1688
2 3501 1 1688
2 3502 1 1689
2 3503 1 1689
2 3504 1 1689
2 3505 1 1690
2 3506 1 1690
2 3507 1 1692
2 3508 1 1692
2 3509 1 1693
2 3510 1 1693
2 3511 1 1695
2 3512 1 1695
2 3513 1 1695
2 3514 1 1695
2 3515 1 1698
2 3516 1 1698
2 3517 1 1701
2 3518 1 1701
2 3519 1 1701
2 3520 1 1701
2 3521 1 1705
2 3522 1 1705
2 3523 1 1705
2 3524 1 1709
2 3525 1 1709
2 3526 1 1717
2 3527 1 1717
2 3528 1 1719
2 3529 1 1719
2 3530 1 1719
2 3531 1 1720
2 3532 1 1720
2 3533 1 1730
2 3534 1 1730
2 3535 1 1735
2 3536 1 1735
2 3537 1 1736
2 3538 1 1736
2 3539 1 1741
2 3540 1 1741
2 3541 1 1741
2 3542 1 1747
2 3543 1 1747
2 3544 1 1748
2 3545 1 1748
2 3546 1 1754
2 3547 1 1754
2 3548 1 1754
2 3549 1 1758
2 3550 1 1758
2 3551 1 1759
2 3552 1 1759
2 3553 1 1759
2 3554 1 1760
2 3555 1 1760
2 3556 1 1769
2 3557 1 1769
2 3558 1 1769
2 3559 1 1770
2 3560 1 1770
2 3561 1 1792
2 3562 1 1792
2 3563 1 1793
2 3564 1 1793
2 3565 1 1801
2 3566 1 1801
2 3567 1 1801
2 3568 1 1802
2 3569 1 1802
2 3570 1 1811
2 3571 1 1811
2 3572 1 1821
2 3573 1 1821
2 3574 1 1822
2 3575 1 1822
2 3576 1 1825
2 3577 1 1825
2 3578 1 1826
2 3579 1 1826
2 3580 1 1829
2 3581 1 1829
2 3582 1 1832
2 3583 1 1832
2 3584 1 1844
2 3585 1 1844
2 3586 1 1847
2 3587 1 1847
2 3588 1 1848
2 3589 1 1848
2 3590 1 1851
2 3591 1 1851
2 3592 1 1852
2 3593 1 1852
2 3594 1 1853
2 3595 1 1853
2 3596 1 1855
2 3597 1 1855
2 3598 1 1858
2 3599 1 1858
2 3600 1 1861
2 3601 1 1861
0 33 5 2 1 1966
0 34 5 2 1 1976
0 35 5 2 1 1986
0 36 5 2 1 1997
0 37 5 2 1 2007
0 38 5 2 1 2018
0 39 5 2 1 2028
0 40 5 2 1 2038
0 41 5 2 1 2048
0 42 5 2 1 2058
0 43 5 2 1 2069
0 44 5 2 1 2079
0 45 5 2 1 2089
0 46 5 2 1 2099
0 47 5 2 1 2109
0 48 5 3 1 2119
0 49 5 3 1 2122
0 50 5 3 1 2125
0 51 5 3 1 2128
0 52 5 3 1 2131
0 53 5 3 1 2134
0 54 5 3 1 2137
0 55 5 3 1 2140
0 56 5 3 1 2143
0 57 5 3 1 2146
0 58 5 3 1 2149
0 59 5 3 1 2152
0 60 5 4 1 2155
0 61 5 3 1 2159
0 62 5 2 1 2162
0 63 5 2 1 2166
0 64 7 2 2 2240 2243
0 65 5 1 1 2247
0 66 7 3 2 2167 2248
0 67 5 1 1 2249
0 68 7 2 2 2241 2168
0 69 5 1 1 2252
0 70 7 1 2 65 2253
0 71 5 1 1 70
0 72 7 1 2 2160 2245
0 73 5 1 1 72
0 74 7 2 2 71 73
0 75 5 1 1 2254
0 76 7 2 2 2236 2255
0 77 5 1 1 2256
0 78 7 1 2 2163 69
0 79 7 1 2 77 78
0 80 5 1 1 79
0 81 7 2 2 67 80
0 82 5 1 1 2258
0 83 7 1 2 2237 82
0 84 5 2 1 83
0 85 7 1 2 2156 2259
0 86 5 1 1 85
0 87 7 2 2 2260 86
0 88 5 1 1 2262
0 89 7 2 2 2233 2263
0 90 5 2 1 2264
0 91 7 1 2 75 2261
0 92 5 1 1 91
0 93 7 1 2 2238 2250
0 94 5 1 1 93
0 95 7 2 2 92 94
0 96 5 1 1 2268
0 97 7 1 2 2266 96
0 98 5 2 1 97
0 99 7 1 2 2164 2257
0 100 5 1 1 99
0 101 7 1 2 2157 2251
0 102 5 1 1 101
0 103 7 2 2 100 102
0 104 5 2 1 2272
0 105 7 2 2 2270 2273
0 106 5 1 1 2276
0 107 7 1 2 2234 106
0 108 5 2 1 107
0 109 7 1 2 2153 2277
0 110 5 1 1 109
0 111 7 2 2 2278 110
0 112 5 1 1 2280
0 113 7 2 2 2230 2281
0 114 5 2 1 2282
0 115 7 1 2 88 2279
0 116 5 1 1 115
0 117 7 1 2 2265 2274
0 118 5 1 1 117
0 119 7 2 2 116 118
0 120 5 1 1 2286
0 121 7 1 2 2284 120
0 122 5 2 1 121
0 123 7 1 2 2267 2275
0 124 5 1 1 123
0 125 7 1 2 2269 124
0 126 5 1 1 125
0 127 7 3 2 2271 126
0 128 5 1 1 2290
0 129 7 2 2 2288 128
0 130 5 1 1 2293
0 131 7 1 2 2231 130
0 132 5 2 1 131
0 133 7 1 2 2150 2294
0 134 5 1 1 133
0 135 7 2 2 2295 134
0 136 5 1 1 2297
0 137 7 2 2 2227 2298
0 138 5 2 1 2299
0 139 7 1 2 112 2296
0 140 5 1 1 139
0 141 7 1 2 2283 2291
0 142 5 1 1 141
0 143 7 2 2 140 142
0 144 5 1 1 2303
0 145 7 1 2 2301 144
0 146 5 2 1 145
0 147 7 1 2 2285 2292
0 148 5 1 1 147
0 149 7 1 2 2287 148
0 150 5 1 1 149
0 151 7 3 2 2289 150
0 152 5 1 1 2307
0 153 7 2 2 2305 152
0 154 5 1 1 2310
0 155 7 1 2 2228 154
0 156 5 2 1 155
0 157 7 1 2 2147 2311
0 158 5 1 1 157
0 159 7 2 2 2312 158
0 160 5 1 1 2314
0 161 7 2 2 2224 2315
0 162 5 2 1 2316
0 163 7 1 2 136 2313
0 164 5 1 1 163
0 165 7 1 2 2300 2308
0 166 5 1 1 165
0 167 7 2 2 164 166
0 168 5 1 1 2320
0 169 7 1 2 2318 168
0 170 5 2 1 169
0 171 7 1 2 2302 2309
0 172 5 1 1 171
0 173 7 1 2 2304 172
0 174 5 1 1 173
0 175 7 3 2 2306 174
0 176 5 1 1 2324
0 177 7 2 2 2322 176
0 178 5 1 1 2327
0 179 7 1 2 2225 178
0 180 5 2 1 179
0 181 7 1 2 2144 2328
0 182 5 1 1 181
0 183 7 2 2 2329 182
0 184 5 1 1 2331
0 185 7 2 2 2221 2332
0 186 5 2 1 2333
0 187 7 1 2 160 2330
0 188 5 1 1 187
0 189 7 1 2 2317 2325
0 190 5 1 1 189
0 191 7 2 2 188 190
0 192 5 1 1 2337
0 193 7 1 2 2335 192
0 194 5 2 1 193
0 195 7 1 2 2319 2326
0 196 5 1 1 195
0 197 7 1 2 2321 196
0 198 5 1 1 197
0 199 7 3 2 2323 198
0 200 5 1 1 2341
0 201 7 2 2 2339 200
0 202 5 1 1 2344
0 203 7 1 2 2222 202
0 204 5 2 1 203
0 205 7 1 2 2141 2345
0 206 5 1 1 205
0 207 7 2 2 2346 206
0 208 5 1 1 2348
0 209 7 2 2 2218 2349
0 210 5 2 1 2350
0 211 7 1 2 184 2347
0 212 5 1 1 211
0 213 7 1 2 2334 2342
0 214 5 1 1 213
0 215 7 2 2 212 214
0 216 5 1 1 2354
0 217 7 1 2 2352 216
0 218 5 2 1 217
0 219 7 1 2 2336 2343
0 220 5 1 1 219
0 221 7 1 2 2338 220
0 222 5 1 1 221
0 223 7 3 2 2340 222
0 224 5 1 1 2358
0 225 7 2 2 2356 224
0 226 5 1 1 2361
0 227 7 1 2 2219 226
0 228 5 2 1 227
0 229 7 1 2 2138 2362
0 230 5 1 1 229
0 231 7 2 2 2363 230
0 232 5 1 1 2365
0 233 7 2 2 2215 2366
0 234 5 2 1 2367
0 235 7 1 2 208 2364
0 236 5 1 1 235
0 237 7 1 2 2351 2359
0 238 5 1 1 237
0 239 7 2 2 236 238
0 240 5 1 1 2371
0 241 7 1 2 2369 240
0 242 5 2 1 241
0 243 7 1 2 2353 2360
0 244 5 1 1 243
0 245 7 1 2 2355 244
0 246 5 1 1 245
0 247 7 3 2 2357 246
0 248 5 1 1 2375
0 249 7 2 2 2373 248
0 250 5 1 1 2378
0 251 7 1 2 2216 250
0 252 5 2 1 251
0 253 7 1 2 2135 2379
0 254 5 1 1 253
0 255 7 2 2 2380 254
0 256 5 1 1 2382
0 257 7 2 2 2212 2383
0 258 5 2 1 2384
0 259 7 1 2 232 2381
0 260 5 1 1 259
0 261 7 1 2 2368 2376
0 262 5 1 1 261
0 263 7 2 2 260 262
0 264 5 1 1 2388
0 265 7 1 2 2386 264
0 266 5 2 1 265
0 267 7 1 2 2370 2377
0 268 5 1 1 267
0 269 7 1 2 2372 268
0 270 5 1 1 269
0 271 7 3 2 2374 270
0 272 5 1 1 2392
0 273 7 2 2 2390 272
0 274 5 1 1 2395
0 275 7 1 2 2213 274
0 276 5 2 1 275
0 277 7 1 2 2132 2396
0 278 5 1 1 277
0 279 7 2 2 2397 278
0 280 5 1 1 2399
0 281 7 2 2 2209 2400
0 282 5 2 1 2401
0 283 7 1 2 256 2398
0 284 5 1 1 283
0 285 7 1 2 2385 2393
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 2405
0 289 7 1 2 2403 288
0 290 5 2 1 289
0 291 7 1 2 2387 2394
0 292 5 1 1 291
0 293 7 1 2 2389 292
0 294 5 1 1 293
0 295 7 3 2 2391 294
0 296 5 1 1 2409
0 297 7 2 2 2407 296
0 298 5 1 1 2412
0 299 7 1 2 2210 298
0 300 5 2 1 299
0 301 7 1 2 2129 2413
0 302 5 1 1 301
0 303 7 2 2 2414 302
0 304 5 1 1 2416
0 305 7 2 2 2206 2417
0 306 5 2 1 2418
0 307 7 1 2 280 2415
0 308 5 1 1 307
0 309 7 1 2 2402 2410
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 2422
0 313 7 1 2 2420 312
0 314 5 2 1 313
0 315 7 1 2 2404 2411
0 316 5 1 1 315
0 317 7 1 2 2406 316
0 318 5 1 1 317
0 319 7 3 2 2408 318
0 320 5 1 1 2426
0 321 7 2 2 2424 320
0 322 5 1 1 2429
0 323 7 1 2 2207 322
0 324 5 2 1 323
0 325 7 1 2 2126 2430
0 326 5 1 1 325
0 327 7 2 2 2431 326
0 328 5 1 1 2433
0 329 7 2 2 2203 2434
0 330 5 2 1 2435
0 331 7 1 2 304 2432
0 332 5 1 1 331
0 333 7 1 2 2419 2427
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 2439
0 337 7 1 2 2437 336
0 338 5 2 1 337
0 339 7 1 2 2421 2428
0 340 5 1 1 339
0 341 7 1 2 2423 340
0 342 5 1 1 341
0 343 7 3 2 2425 342
0 344 5 1 1 2443
0 345 7 2 2 2441 344
0 346 5 1 1 2446
0 347 7 1 2 2204 346
0 348 5 2 1 347
0 349 7 1 2 2123 2447
0 350 5 1 1 349
0 351 7 2 2 2448 350
0 352 5 1 1 2450
0 353 7 2 2 2200 2451
0 354 5 2 1 2452
0 355 7 1 2 328 2449
0 356 5 1 1 355
0 357 7 1 2 2436 2444
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 2456
0 361 7 1 2 2454 360
0 362 5 2 1 361
0 363 7 1 2 2438 2445
0 364 5 1 1 363
0 365 7 1 2 2440 364
0 366 5 1 1 365
0 367 7 3 2 2442 366
0 368 5 1 1 2460
0 369 7 2 2 2458 368
0 370 5 1 1 2463
0 371 7 1 2 2201 370
0 372 5 2 1 371
0 373 7 1 2 2120 2464
0 374 5 1 1 373
0 375 7 2 2 2465 374
0 376 5 1 1 2467
0 377 7 2 2 2198 2468
0 378 5 2 1 2469
0 379 7 1 2 352 2466
0 380 5 1 1 379
0 381 7 1 2 2453 2461
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 2473
0 385 7 1 2 2471 384
0 386 5 2 1 385
0 387 7 1 2 2455 2462
0 388 5 1 1 387
0 389 7 1 2 2457 388
0 390 5 1 1 389
0 391 7 3 2 2459 390
0 392 5 1 1 2477
0 393 7 2 2 2475 392
0 394 5 1 1 2480
0 395 7 1 2 2199 394
0 396 5 2 1 395
0 397 7 1 2 2110 2481
0 398 5 1 1 397
0 399 7 2 2 2482 398
0 400 5 1 1 2484
0 401 7 2 2 2196 2485
0 402 5 2 1 2486
0 403 7 1 2 376 2483
0 404 5 1 1 403
0 405 7 1 2 2470 2478
0 406 5 1 1 405
0 407 7 2 2 404 406
0 408 5 1 1 2490
0 409 7 1 2 2488 408
0 410 5 2 1 409
0 411 7 1 2 2472 2479
0 412 5 1 1 411
0 413 7 1 2 2474 412
0 414 5 1 1 413
0 415 7 3 2 2476 414
0 416 5 1 1 2494
0 417 7 2 2 2492 416
0 418 5 1 1 2497
0 419 7 1 2 2197 418
0 420 5 2 1 419
0 421 7 1 2 2100 2498
0 422 5 1 1 421
0 423 7 2 2 2499 422
0 424 5 1 1 2501
0 425 7 2 2 2194 2502
0 426 5 2 1 2503
0 427 7 1 2 400 2500
0 428 5 1 1 427
0 429 7 1 2 2487 2495
0 430 5 1 1 429
0 431 7 2 2 428 430
0 432 5 1 1 2507
0 433 7 1 2 2505 432
0 434 5 2 1 433
0 435 7 1 2 2489 2496
0 436 5 1 1 435
0 437 7 1 2 2491 436
0 438 5 1 1 437
0 439 7 3 2 2493 438
0 440 5 1 1 2511
0 441 7 2 2 2509 440
0 442 5 1 1 2514
0 443 7 1 2 2195 442
0 444 5 2 1 443
0 445 7 1 2 2090 2515
0 446 5 1 1 445
0 447 7 2 2 2516 446
0 448 5 1 1 2518
0 449 7 2 2 2192 2519
0 450 5 2 1 2520
0 451 7 1 2 424 2517
0 452 5 1 1 451
0 453 7 1 2 2504 2512
0 454 5 1 1 453
0 455 7 2 2 452 454
0 456 5 1 1 2524
0 457 7 1 2 2522 456
0 458 5 2 1 457
0 459 7 1 2 2506 2513
0 460 5 1 1 459
0 461 7 1 2 2508 460
0 462 5 1 1 461
0 463 7 3 2 2510 462
0 464 5 1 1 2528
0 465 7 2 2 2526 464
0 466 5 1 1 2531
0 467 7 1 2 2193 466
0 468 5 2 1 467
0 469 7 1 2 2080 2532
0 470 5 1 1 469
0 471 7 2 2 2533 470
0 472 5 1 1 2535
0 473 7 2 2 2190 2536
0 474 5 2 1 2537
0 475 7 1 2 448 2534
0 476 5 1 1 475
0 477 7 1 2 2521 2529
0 478 5 1 1 477
0 479 7 2 2 476 478
0 480 5 1 1 2541
0 481 7 1 2 2539 480
0 482 5 2 1 481
0 483 7 1 2 2523 2530
0 484 5 1 1 483
0 485 7 1 2 2525 484
0 486 5 1 1 485
0 487 7 3 2 2527 486
0 488 5 1 1 2545
0 489 7 2 2 2543 488
0 490 5 1 1 2548
0 491 7 1 2 2191 490
0 492 5 2 1 491
0 493 7 1 2 2070 2549
0 494 5 1 1 493
0 495 7 2 2 2550 494
0 496 5 1 1 2552
0 497 7 2 2 2188 2553
0 498 5 2 1 2554
0 499 7 1 2 472 2551
0 500 5 1 1 499
0 501 7 1 2 2538 2546
0 502 5 1 1 501
0 503 7 2 2 500 502
0 504 5 1 1 2558
0 505 7 1 2 2556 504
0 506 5 2 1 505
0 507 7 1 2 2540 2547
0 508 5 1 1 507
0 509 7 1 2 2542 508
0 510 5 1 1 509
0 511 7 3 2 2544 510
0 512 5 1 1 2562
0 513 7 2 2 2560 512
0 514 5 1 1 2565
0 515 7 1 2 2189 514
0 516 5 2 1 515
0 517 7 1 2 2059 2566
0 518 5 1 1 517
0 519 7 2 2 2567 518
0 520 5 1 1 2569
0 521 7 2 2 2186 2570
0 522 5 2 1 2571
0 523 7 1 2 496 2568
0 524 5 1 1 523
0 525 7 1 2 2555 2563
0 526 5 1 1 525
0 527 7 2 2 524 526
0 528 5 1 1 2575
0 529 7 1 2 2573 528
0 530 5 2 1 529
0 531 7 1 2 2557 2564
0 532 5 1 1 531
0 533 7 1 2 2559 532
0 534 5 1 1 533
0 535 7 3 2 2561 534
0 536 5 1 1 2579
0 537 7 2 2 2577 536
0 538 5 1 1 2582
0 539 7 1 2 2187 538
0 540 5 2 1 539
0 541 7 1 2 2049 2583
0 542 5 1 1 541
0 543 7 2 2 2584 542
0 544 5 1 1 2586
0 545 7 2 2 2184 2587
0 546 5 2 1 2588
0 547 7 1 2 520 2585
0 548 5 1 1 547
0 549 7 1 2 2572 2580
0 550 5 1 1 549
0 551 7 2 2 548 550
0 552 5 1 1 2592
0 553 7 1 2 2590 552
0 554 5 2 1 553
0 555 7 1 2 2574 2581
0 556 5 1 1 555
0 557 7 1 2 2576 556
0 558 5 1 1 557
0 559 7 3 2 2578 558
0 560 5 1 1 2596
0 561 7 2 2 2594 560
0 562 5 1 1 2599
0 563 7 1 2 2185 562
0 564 5 2 1 563
0 565 7 1 2 2039 2600
0 566 5 1 1 565
0 567 7 2 2 2601 566
0 568 5 1 1 2603
0 569 7 2 2 2182 2604
0 570 5 2 1 2605
0 571 7 1 2 544 2602
0 572 5 1 1 571
0 573 7 1 2 2589 2597
0 574 5 1 1 573
0 575 7 2 2 572 574
0 576 5 1 1 2609
0 577 7 1 2 2607 576
0 578 5 2 1 577
0 579 7 1 2 2591 2598
0 580 5 1 1 579
0 581 7 1 2 2593 580
0 582 5 1 1 581
0 583 7 3 2 2595 582
0 584 5 1 1 2613
0 585 7 2 2 2611 584
0 586 5 1 1 2616
0 587 7 1 2 2183 586
0 588 5 2 1 587
0 589 7 1 2 2029 2617
0 590 5 1 1 589
0 591 7 2 2 2618 590
0 592 5 1 1 2620
0 593 7 2 2 2180 2621
0 594 5 2 1 2622
0 595 7 1 2 568 2619
0 596 5 1 1 595
0 597 7 1 2 2606 2614
0 598 5 1 1 597
0 599 7 2 2 596 598
0 600 5 1 1 2626
0 601 7 1 2 2624 600
0 602 5 2 1 601
0 603 7 1 2 2608 2615
0 604 5 1 1 603
0 605 7 1 2 2610 604
0 606 5 1 1 605
0 607 7 3 2 2612 606
0 608 5 1 1 2630
0 609 7 2 2 2628 608
0 610 5 1 1 2633
0 611 7 1 2 2181 610
0 612 5 2 1 611
0 613 7 1 2 2019 2634
0 614 5 1 1 613
0 615 7 2 2 2635 614
0 616 5 1 1 2637
0 617 7 2 2 2178 2638
0 618 5 2 1 2639
0 619 7 1 2 592 2636
0 620 5 1 1 619
0 621 7 1 2 2623 2631
0 622 5 1 1 621
0 623 7 2 2 620 622
0 624 5 1 1 2643
0 625 7 1 2 2641 624
0 626 5 2 1 625
0 627 7 1 2 2625 2632
0 628 5 1 1 627
0 629 7 1 2 2627 628
0 630 5 1 1 629
0 631 7 3 2 2629 630
0 632 5 1 1 2647
0 633 7 2 2 2645 632
0 634 5 1 1 2650
0 635 7 1 2 2179 634
0 636 5 2 1 635
0 637 7 1 2 2008 2651
0 638 5 1 1 637
0 639 7 2 2 2652 638
0 640 5 1 1 2654
0 641 7 2 2 2176 2655
0 642 5 2 1 2656
0 643 7 1 2 616 2653
0 644 5 1 1 643
0 645 7 1 2 2640 2648
0 646 5 1 1 645
0 647 7 2 2 644 646
0 648 5 1 1 2660
0 649 7 1 2 2658 648
0 650 5 2 1 649
0 651 7 1 2 2642 2649
0 652 5 1 1 651
0 653 7 1 2 2644 652
0 654 5 1 1 653
0 655 7 3 2 2646 654
0 656 5 1 1 2664
0 657 7 2 2 2662 656
0 658 5 1 1 2667
0 659 7 1 2 2177 658
0 660 5 2 1 659
0 661 7 1 2 1998 2668
0 662 5 1 1 661
0 663 7 2 2 2669 662
0 664 5 1 1 2671
0 665 7 2 2 2174 2672
0 666 5 2 1 2673
0 667 7 1 2 640 2670
0 668 5 1 1 667
0 669 7 1 2 2657 2665
0 670 5 1 1 669
0 671 7 2 2 668 670
0 672 5 1 1 2677
0 673 7 1 2 2675 672
0 674 5 2 1 673
0 675 7 1 2 2659 2666
0 676 5 1 1 675
0 677 7 1 2 2661 676
0 678 5 1 1 677
0 679 7 3 2 2663 678
0 680 5 1 1 2681
0 681 7 2 2 2679 680
0 682 5 1 1 2684
0 683 7 1 2 1987 2685
0 684 5 1 1 683
0 685 7 1 2 2175 682
0 686 5 2 1 685
0 687 7 3 2 684 2686
0 688 5 2 1 2688
0 689 7 2 2 2172 2689
0 690 5 2 1 2693
0 691 7 1 2 664 2687
0 692 5 1 1 691
0 693 7 1 2 2674 2682
0 694 5 1 1 693
0 695 7 2 2 692 694
0 696 5 1 1 2697
0 697 7 1 2 2695 696
0 698 5 2 1 697
0 699 7 1 2 2676 2683
0 700 5 1 1 699
0 701 7 1 2 2678 700
0 702 5 1 1 701
0 703 7 3 2 2680 702
0 704 5 1 1 2701
0 705 7 1 2 2696 2702
0 706 5 1 1 705
0 707 7 1 2 2698 706
0 708 5 1 1 707
0 709 7 1 2 2699 708
0 710 5 1 1 709
0 711 7 2 2 2700 704
0 712 5 1 1 2704
0 713 7 1 2 2173 712
0 714 5 2 1 713
0 715 7 1 2 1977 2705
0 716 5 1 1 715
0 717 7 2 2 2706 716
0 718 7 1 2 2170 2708
0 719 5 1 1 718
0 720 7 1 2 2691 2707
0 721 5 1 1 720
0 722 7 1 2 2694 2703
0 723 5 1 1 722
0 724 7 1 2 721 723
0 725 5 1 1 724
0 726 7 1 2 719 725
0 727 5 1 1 726
0 728 7 2 2 710 727
0 729 5 1 1 2710
0 730 7 1 2 2171 2690
0 731 5 1 1 730
0 732 7 1 2 2711 731
0 733 5 1 1 732
0 734 7 1 2 1967 2692
0 735 5 1 1 734
0 736 7 1 2 729 735
0 737 5 1 1 736
0 738 7 1 2 2709 737
0 739 7 2 2 733 738
0 740 5 1 1 2712
0 741 7 2 2 2030 2111
0 742 5 1 1 2714
0 743 7 2 2 2020 2101
0 744 5 2 1 2716
0 745 7 2 2 2031 2091
0 746 5 1 1 2720
0 747 7 2 2 2009 2112
0 748 5 1 1 2722
0 749 7 1 2 2721 2723
0 750 5 2 1 749
0 751 7 1 2 746 748
0 752 5 1 1 751
0 753 7 2 2 752 2724
0 754 5 1 1 2726
0 755 7 1 2 2717 2727
0 756 5 2 1 755
0 757 7 2 2 2725 2728
0 758 5 1 1 2730
0 759 7 2 2 2021 2113
0 760 5 1 1 2732
0 761 7 2 2 2032 2102
0 762 5 1 1 2734
0 763 7 1 2 760 2735
0 764 5 1 1 763
0 765 7 1 2 2733 762
0 766 5 1 1 765
0 767 7 2 2 764 766
0 768 5 1 1 2736
0 769 7 1 2 758 768
0 770 5 3 1 769
0 771 7 1 2 2718 2738
0 772 5 1 1 771
0 773 7 1 2 2715 772
0 774 5 2 1 773
0 775 7 2 2 1999 2114
0 776 5 1 1 2743
0 777 7 2 2 2033 2081
0 778 5 1 1 2745
0 779 7 1 2 2744 2746
0 780 5 2 1 779
0 781 7 2 2 2022 2092
0 782 5 1 1 2749
0 783 7 1 2 776 778
0 784 5 1 1 783
0 785 7 2 2 2747 784
0 786 5 1 1 2751
0 787 7 1 2 2750 2752
0 788 5 2 1 787
0 789 7 2 2 2748 2753
0 790 5 1 1 2755
0 791 7 1 2 2719 754
0 792 5 1 1 791
0 793 7 2 2 2729 792
0 794 5 1 1 2757
0 795 7 1 2 790 2758
0 796 5 2 1 795
0 797 7 2 2 2010 2103
0 798 5 1 1 2761
0 799 7 1 2 782 786
0 800 5 1 1 799
0 801 7 2 2 2754 800
0 802 5 1 1 2763
0 803 7 1 2 2762 2764
0 804 5 2 1 803
0 805 7 2 2 1988 2115
0 806 5 1 1 2767
0 807 7 2 2 2034 2071
0 808 5 1 1 2769
0 809 7 1 2 2768 2770
0 810 5 2 1 809
0 811 7 2 2 2023 2082
0 812 5 1 1 2773
0 813 7 1 2 806 808
0 814 5 1 1 813
0 815 7 2 2 2771 814
0 816 5 1 1 2775
0 817 7 1 2 2774 2776
0 818 5 2 1 817
0 819 7 2 2 2772 2777
0 820 5 1 1 2779
0 821 7 1 2 798 802
0 822 5 1 1 821
0 823 7 2 2 2765 822
0 824 5 1 1 2781
0 825 7 1 2 820 2782
0 826 5 2 1 825
0 827 7 2 2 2766 2783
0 828 5 1 1 2785
0 829 7 1 2 2756 794
0 830 5 1 1 829
0 831 7 2 2 2759 830
0 832 5 1 1 2787
0 833 7 1 2 828 2788
0 834 5 2 1 833
0 835 7 2 2 2760 2789
0 836 5 1 1 2791
0 837 7 1 2 2731 2737
0 838 5 1 1 837
0 839 7 2 2 2739 838
0 840 5 1 1 2793
0 841 7 1 2 836 2794
0 842 5 2 1 841
0 843 7 2 2 2000 2104
0 844 5 1 1 2797
0 845 7 1 2 812 816
0 846 5 1 1 845
0 847 7 2 2 2778 846
0 848 5 1 1 2799
0 849 7 1 2 2798 2800
0 850 5 2 1 849
0 851 7 2 2 2011 2093
0 852 5 1 1 2803
0 853 7 1 2 844 848
0 854 5 1 1 853
0 855 7 2 2 2801 854
0 856 5 1 1 2805
0 857 7 1 2 2804 2806
0 858 5 2 1 857
0 859 7 2 2 2802 2807
0 860 5 1 1 2809
0 861 7 1 2 2780 824
0 862 5 1 1 861
0 863 7 2 2 2784 862
0 864 5 1 1 2811
0 865 7 1 2 860 2812
0 866 5 2 1 865
0 867 7 2 2 2035 2040
0 868 5 1 1 2815
0 869 7 2 2 2024 2050
0 870 5 1 1 2817
0 871 7 2 2 2816 2818
0 872 5 2 1 2819
0 873 7 2 2 2060 2820
0 874 5 2 1 2823
0 875 7 2 2 1978 2116
0 876 5 1 1 2827
0 877 7 1 2 2824 2828
0 878 5 2 1 877
0 879 7 2 2 2036 2061
0 880 5 1 1 2831
0 881 7 1 2 2825 876
0 882 5 1 1 881
0 883 7 2 2 2829 882
0 884 5 1 1 2833
0 885 7 1 2 2832 2834
0 886 5 2 1 885
0 887 7 2 2 2830 2835
0 888 5 1 1 2837
0 889 7 1 2 852 856
0 890 5 1 1 889
0 891 7 2 2 2808 890
0 892 5 1 1 2839
0 893 7 1 2 888 2840
0 894 5 2 1 893
0 895 7 2 2 2012 2083
0 896 5 1 1 2843
0 897 7 1 2 880 884
0 898 5 1 1 897
0 899 7 2 2 2836 898
0 900 5 1 1 2845
0 901 7 1 2 2844 2846
0 902 5 2 1 901
0 903 7 2 2 2025 2072
0 904 5 1 1 2849
0 905 7 1 2 896 900
0 906 5 1 1 905
0 907 7 2 2 2847 906
0 908 5 1 1 2851
0 909 7 1 2 2850 2852
0 910 5 2 1 909
0 911 7 2 2 2848 2853
0 912 5 1 1 2855
0 913 7 1 2 2838 892
0 914 5 1 1 913
0 915 7 2 2 2841 914
0 916 5 1 1 2857
0 917 7 1 2 912 2858
0 918 5 2 1 917
0 919 7 2 2 2842 2859
0 920 5 1 1 2861
0 921 7 1 2 2810 864
0 922 5 1 1 921
0 923 7 2 2 2813 922
0 924 5 1 1 2863
0 925 7 1 2 920 2864
0 926 5 2 1 925
0 927 7 2 2 2814 2865
0 928 5 1 1 2867
0 929 7 1 2 2786 832
0 930 5 1 1 929
0 931 7 2 2 2790 930
0 932 5 1 1 2869
0 933 7 1 2 928 2870
0 934 5 2 1 933
0 935 7 2 2 1989 2105
0 936 5 1 1 2873
0 937 7 2 2 2001 2094
0 938 5 1 1 2875
0 939 7 1 2 2874 2876
0 940 5 2 1 939
0 941 7 1 2 904 908
0 942 5 1 1 941
0 943 7 2 2 2854 942
0 944 5 1 1 2879
0 945 7 1 2 936 938
0 946 5 1 1 945
0 947 7 2 2 2877 946
0 948 5 1 1 2881
0 949 7 1 2 2880 2882
0 950 5 2 1 949
0 951 7 2 2 2878 2883
0 952 5 1 1 2885
0 953 7 1 2 2856 916
0 954 5 1 1 953
0 955 7 2 2 2860 954
0 956 5 1 1 2887
0 957 7 1 2 952 2888
0 958 5 2 1 957
0 959 7 2 2 2013 2073
0 960 5 1 1 2891
0 961 7 2 2 1979 2106
0 962 5 1 1 2893
0 963 7 1 2 2892 2894
0 964 5 2 1 963
0 965 7 2 2 1968 2117
0 966 5 1 1 2897
0 967 7 2 2 2002 2084
0 968 5 1 1 2899
0 969 7 1 2 2026 2062
0 970 5 1 1 969
0 971 7 1 2 2821 970
0 972 5 1 1 971
0 973 7 2 2 2826 972
0 974 5 1 1 2901
0 975 7 1 2 2900 2902
0 976 5 2 1 975
0 977 7 1 2 968 974
0 978 5 1 1 977
0 979 7 2 2 2903 978
0 980 5 1 1 2905
0 981 7 1 2 2898 2906
0 982 5 2 1 981
0 983 7 1 2 966 980
0 984 5 1 1 983
0 985 7 2 2 2907 984
0 986 5 1 1 2909
0 987 7 1 2 960 962
0 988 5 1 1 987
0 989 7 2 2 2895 988
0 990 5 1 1 2911
0 991 7 1 2 2910 2912
0 992 5 2 1 991
0 993 7 2 2 2896 2913
0 994 5 1 1 2915
0 995 7 1 2 944 948
0 996 5 1 1 995
0 997 7 2 2 2884 996
0 998 5 1 1 2917
0 999 7 1 2 994 2918
0 1000 5 2 1 999
0 1001 7 2 2 2037 2051
0 1002 5 1 1 2921
0 1003 7 2 2 1990 2095
0 1004 5 1 1 2923
0 1005 7 1 2 2922 2924
0 1006 5 2 1 1005
0 1007 7 1 2 986 990
0 1008 5 1 1 1007
0 1009 7 2 2 2914 1008
0 1010 5 1 1 2927
0 1011 7 1 2 1002 1004
0 1012 5 1 1 1011
0 1013 7 2 2 2925 1012
0 1014 5 1 1 2929
0 1015 7 1 2 2928 2930
0 1016 5 2 1 1015
0 1017 7 2 2 2926 2931
0 1018 5 1 1 2933
0 1019 7 1 2 2916 998
0 1020 5 1 1 1019
0 1021 7 2 2 2919 1020
0 1022 5 1 1 2935
0 1023 7 1 2 1018 2936
0 1024 5 2 1 1023
0 1025 7 2 2 2920 2937
0 1026 5 1 1 2939
0 1027 7 1 2 2886 956
0 1028 5 1 1 1027
0 1029 7 2 2 2889 1028
0 1030 5 1 1 2941
0 1031 7 1 2 1026 2942
0 1032 5 2 1 1031
0 1033 7 2 2 2890 2943
0 1034 5 1 1 2945
0 1035 7 1 2 2862 924
0 1036 5 1 1 1035
0 1037 7 2 2 2866 1036
0 1038 5 1 1 2947
0 1039 7 1 2 1034 2948
0 1040 5 2 1 1039
0 1041 7 2 2 2904 2908
0 1042 5 1 1 2951
0 1043 7 1 2 2934 1022
0 1044 5 1 1 1043
0 1045 7 2 2 2938 1044
0 1046 5 1 1 2953
0 1047 7 1 2 1042 2954
0 1048 5 2 1 1047
0 1049 7 2 2 2014 2063
0 1050 5 1 1 2957
0 1051 7 2 2 2003 2074
0 1052 5 1 1 2959
0 1053 7 1 2 2958 2960
0 1054 5 2 1 1053
0 1055 7 2 2 1969 2107
0 1056 5 1 1 2963
0 1057 7 1 2 1050 1052
0 1058 5 1 1 1057
0 1059 7 2 2 2961 1058
0 1060 5 1 1 2965
0 1061 7 1 2 2964 2966
0 1062 5 2 1 1061
0 1063 7 2 2 2962 2967
0 1064 5 1 1 2969
0 1065 7 2 2 1980 2096
0 1066 5 1 1 2971
0 1067 7 2 2 32 2118
0 1068 5 1 1 2973
0 1069 7 1 2 2972 2974
0 1070 5 2 1 1069
0 1071 7 2 2 1991 2085
0 1072 5 1 1 2977
0 1073 7 2 2 2004 2052
0 1074 5 1 1 2979
0 1075 7 2 2 1959 2075
0 1076 5 1 1 2981
0 1077 7 2 2 1981 2053
0 1078 5 1 1 2983
0 1079 7 2 2 2982 2984
0 1080 5 2 1 2985
0 1081 7 2 2 1992 2986
0 1082 5 2 1 2989
0 1083 7 2 2 2980 2990
0 1084 5 2 1 2993
0 1085 7 2 2 2015 2994
0 1086 5 2 1 2997
0 1087 7 1 2 2978 2998
0 1088 5 2 1 1087
0 1089 7 1 2 1072 2999
0 1090 5 1 1 1089
0 1091 7 2 2 3001 1090
0 1092 5 1 1 3003
0 1093 7 1 2 868 870
0 1094 5 1 1 1093
0 1095 7 2 2 2822 1094
0 1096 5 1 1 3005
0 1097 7 1 2 3004 3006
0 1098 5 2 1 1097
0 1099 7 1 2 1092 1096
0 1100 5 1 1 1099
0 1101 7 2 2 3007 1100
0 1102 5 1 1 3009
0 1103 7 1 2 1066 1068
0 1104 5 1 1 1103
0 1105 7 2 2 2975 1104
0 1106 5 1 1 3011
0 1107 7 1 2 3010 3012
0 1108 5 2 1 1107
0 1109 7 2 2 2976 3013
0 1110 5 1 1 3015
0 1111 7 1 2 1064 1110
0 1112 5 2 1 1111
0 1113 7 2 2 3002 3008
0 1114 5 1 1 3019
0 1115 7 1 2 2970 3016
0 1116 5 1 1 1115
0 1117 7 2 2 3017 1116
0 1118 5 1 1 3021
0 1119 7 1 2 1114 3022
0 1120 5 2 1 1119
0 1121 7 2 2 3018 3023
0 1122 5 1 1 3025
0 1123 7 1 2 2952 1046
0 1124 5 1 1 1123
0 1125 7 2 2 2955 1124
0 1126 5 1 1 3027
0 1127 7 1 2 1122 3028
0 1128 5 2 1 1127
0 1129 7 2 2 2956 3029
0 1130 5 1 1 3031
0 1131 7 1 2 2940 1030
0 1132 5 1 1 1131
0 1133 7 2 2 2944 1132
0 1134 5 1 1 3033
0 1135 7 1 2 1130 3034
0 1136 5 2 1 1135
0 1137 7 1 2 1010 1014
0 1138 5 1 1 1137
0 1139 7 2 2 2932 1138
0 1140 5 1 1 3037
0 1141 7 1 2 3020 1118
0 1142 5 1 1 1141
0 1143 7 2 2 3024 1142
0 1144 5 1 1 3039
0 1145 7 1 2 3038 3040
0 1146 5 2 1 1145
0 1147 7 1 2 1056 1060
0 1148 5 1 1 1147
0 1149 7 2 2 2968 1148
0 1150 5 1 1 3043
0 1151 7 1 2 1102 1106
0 1152 5 1 1 1151
0 1153 7 2 2 3014 1152
0 1154 5 1 1 3045
0 1155 7 1 2 3044 3046
0 1156 5 2 1 1155
0 1157 7 2 2 1993 2076
0 1158 5 1 1 3049
0 1159 7 2 2 1982 2086
0 1160 5 1 1 3051
0 1161 7 1 2 3050 3052
0 1162 5 2 1 1161
0 1163 7 2 2 1970 2097
0 1164 5 1 1 3055
0 1165 7 1 2 1158 1160
0 1166 5 1 1 1165
0 1167 7 2 2 3053 1166
0 1168 5 1 1 3057
0 1169 7 1 2 3056 3058
0 1170 5 2 1 1169
0 1171 7 2 2 3054 3059
0 1172 5 1 1 3061
0 1173 7 1 2 1150 1154
0 1174 5 1 1 1173
0 1175 7 2 2 3047 1174
0 1176 5 1 1 3063
0 1177 7 1 2 1172 3064
0 1178 5 2 1 1177
0 1179 7 2 2 3048 3065
0 1180 5 1 1 3067
0 1181 7 1 2 1140 1144
0 1182 5 1 1 1181
0 1183 7 2 2 3041 1182
0 1184 5 1 1 3069
0 1185 7 1 2 1180 3070
0 1186 5 2 1 1185
0 1187 7 2 2 3042 3071
0 1188 5 1 1 3073
0 1189 7 1 2 3026 1126
0 1190 5 1 1 1189
0 1191 7 2 2 3030 1190
0 1192 5 1 1 3075
0 1193 7 1 2 1188 3076
0 1194 5 2 1 1193
0 1195 7 2 2 1960 2108
0 1196 5 1 1 3079
0 1197 7 1 2 1164 1168
0 1198 5 1 1 1197
0 1199 7 2 2 3060 1198
0 1200 5 1 1 3081
0 1201 7 1 2 3080 3082
0 1202 5 2 1 1201
0 1203 7 2 2 2027 2041
0 1204 5 1 1 3085
0 1205 7 2 2 2005 2064
0 1206 5 1 1 3087
0 1207 7 1 2 2016 2054
0 1208 5 1 1 1207
0 1209 7 1 2 2995 1208
0 1210 5 1 1 1209
0 1211 7 2 2 3000 1210
0 1212 5 1 1 3089
0 1213 7 1 2 3088 3090
0 1214 5 2 1 1213
0 1215 7 1 2 1206 1212
0 1216 5 1 1 1215
0 1217 7 2 2 3091 1216
0 1218 5 1 1 3093
0 1219 7 1 2 3086 3094
0 1220 5 2 1 1219
0 1221 7 1 2 1204 1218
0 1222 5 1 1 1221
0 1223 7 2 2 3095 1222
0 1224 5 1 1 3097
0 1225 7 1 2 1196 1200
0 1226 5 1 1 1225
0 1227 7 2 2 3083 1226
0 1228 5 1 1 3099
0 1229 7 1 2 3098 3100
0 1230 5 2 1 1229
0 1231 7 2 2 3084 3101
0 1232 5 1 1 3103
0 1233 7 1 2 3062 1176
0 1234 5 1 1 1233
0 1235 7 2 2 3066 1234
0 1236 5 1 1 3105
0 1237 7 1 2 1232 3106
0 1238 5 2 1 1237
0 1239 7 2 2 3092 3096
0 1240 5 1 1 3109
0 1241 7 1 2 3104 1236
0 1242 5 1 1 1241
0 1243 7 2 2 3107 1242
0 1244 5 1 1 3111
0 1245 7 1 2 1240 3112
0 1246 5 2 1 1245
0 1247 7 2 2 3108 3113
0 1248 5 1 1 3115
0 1249 7 1 2 3068 1184
0 1250 5 1 1 1249
0 1251 7 2 2 3072 1250
0 1252 5 1 1 3117
0 1253 7 1 2 1248 3118
0 1254 5 2 1 1253
0 1255 7 2 2 1994 2065
0 1256 5 1 1 3121
0 1257 7 1 2 1074 2991
0 1258 5 1 1 1257
0 1259 7 2 2 2996 1258
0 1260 5 1 1 3123
0 1261 7 1 2 3122 3124
0 1262 5 2 1 1261
0 1263 7 2 2 2017 2042
0 1264 5 1 1 3127
0 1265 7 1 2 1256 1260
0 1266 5 1 1 1265
0 1267 7 2 2 3125 1266
0 1268 5 1 1 3129
0 1269 7 1 2 3128 3130
0 1270 5 2 1 1269
0 1271 7 2 2 3126 3131
0 1272 5 1 1 3133
0 1273 7 1 2 1224 1228
0 1274 5 1 1 1273
0 1275 7 2 2 3102 1274
0 1276 5 1 1 3135
0 1277 7 1 2 1272 3136
0 1278 5 2 1 1277
0 1279 7 2 2 1983 2077
0 1280 5 1 1 3139
0 1281 7 2 2 1961 2098
0 1282 5 1 1 3141
0 1283 7 1 2 3140 3142
0 1284 5 2 1 1283
0 1285 7 1 2 1264 1268
0 1286 5 1 1 1285
0 1287 7 2 2 3132 1286
0 1288 5 1 1 3145
0 1289 7 1 2 1280 1282
0 1290 5 1 1 1289
0 1291 7 2 2 3143 1290
0 1292 5 1 1 3147
0 1293 7 1 2 3146 3148
0 1294 5 2 1 1293
0 1295 7 2 2 3144 3149
0 1296 5 1 1 3151
0 1297 7 1 2 3134 1276
0 1298 5 1 1 1297
0 1299 7 2 2 3137 1298
0 1300 5 1 1 3153
0 1301 7 1 2 1296 3154
0 1302 5 2 1 1301
0 1303 7 2 2 3138 3155
0 1304 5 1 1 3157
0 1305 7 1 2 3110 1244
0 1306 5 1 1 1305
0 1307 7 2 2 3114 1306
0 1308 5 1 1 3159
0 1309 7 1 2 1304 3160
0 1310 5 2 1 1309
0 1311 7 2 2 1971 2087
0 1312 5 1 1 3163
0 1313 7 1 2 1288 1292
0 1314 5 1 1 1313
0 1315 7 2 2 3150 1314
0 1316 5 1 1 3165
0 1317 7 1 2 3164 3166
0 1318 5 2 1 1317
0 1319 7 2 2 1984 2066
0 1320 5 1 1 3169
0 1321 7 1 2 1995 2055
0 1322 5 1 1 1321
0 1323 7 1 2 2987 1322
0 1324 5 1 1 1323
0 1325 7 2 2 2992 1324
0 1326 5 1 1 3171
0 1327 7 1 2 3170 3172
0 1328 5 2 1 1327
0 1329 7 2 2 2006 2043
0 1330 5 1 1 3175
0 1331 7 1 2 1320 1326
0 1332 5 1 1 1331
0 1333 7 2 2 3173 1332
0 1334 5 1 1 3177
0 1335 7 1 2 3176 3178
0 1336 5 2 1 1335
0 1337 7 2 2 3174 3179
0 1338 5 1 1 3181
0 1339 7 1 2 1312 1316
0 1340 5 1 1 1339
0 1341 7 2 2 3167 1340
0 1342 5 1 1 3183
0 1343 7 1 2 1338 3184
0 1344 5 2 1 1343
0 1345 7 2 2 3168 3185
0 1346 5 1 1 3187
0 1347 7 1 2 3152 1300
0 1348 5 1 1 1347
0 1349 7 2 2 3156 1348
0 1350 5 1 1 3189
0 1351 7 1 2 1346 3190
0 1352 5 2 1 1351
0 1353 7 2 2 1962 2088
0 1354 5 1 1 3193
0 1355 7 2 2 1972 2078
0 1356 5 1 1 3195
0 1357 7 1 2 3194 3196
0 1358 5 2 1 1357
0 1359 7 1 2 1330 1334
0 1360 5 1 1 1359
0 1361 7 2 2 3180 1360
0 1362 5 1 1 3199
0 1363 7 1 2 1354 1356
0 1364 5 1 1 1363
0 1365 7 2 2 3197 1364
0 1366 5 1 1 3201
0 1367 7 1 2 3200 3202
0 1368 5 2 1 1367
0 1369 7 2 2 3198 3203
0 1370 5 1 1 3205
0 1371 7 1 2 3182 1342
0 1372 5 1 1 1371
0 1373 7 2 2 3186 1372
0 1374 5 1 1 3207
0 1375 7 1 2 1370 3208
0 1376 5 2 1 1375
0 1377 7 1 2 1362 1366
0 1378 5 1 1 1377
0 1379 7 2 2 3204 1378
0 1380 5 1 1 3211
0 1381 7 2 2 1973 2067
0 1382 5 1 1 3213
0 1383 7 2 2 1996 2044
0 1384 5 1 1 3215
0 1385 7 2 2 3214 3216
0 1386 5 1 1 3217
0 1387 7 2 2 1974 2056
0 1388 5 1 1 3219
0 1389 7 2 2 1963 2068
0 1390 5 1 1 3221
0 1391 7 2 2 3220 3222
0 1392 5 2 1 3223
0 1393 7 3 2 1386 3225
0 1394 5 1 1 3227
0 1395 7 1 2 3212 1394
0 1396 5 2 1 1395
0 1397 7 1 2 1076 1078
0 1398 5 1 1 1397
0 1399 7 2 2 2988 1398
0 1400 5 1 1 3232
0 1401 7 1 2 1382 1384
0 1402 5 1 1 1401
0 1403 7 1 2 3228 1402
0 1404 5 1 1 1403
0 1405 7 1 2 3218 3224
0 1406 5 1 1 1405
0 1407 7 2 2 1404 1406
0 1408 5 1 1 3234
0 1409 7 1 2 3233 1408
0 1410 5 2 1 1409
0 1411 7 2 2 1985 2045
0 1412 5 1 1 3238
0 1413 7 1 2 1388 1390
0 1414 5 1 1 1413
0 1415 7 2 2 3226 1414
0 1416 5 1 1 3240
0 1417 7 1 2 3239 3241
0 1418 5 2 1 1417
0 1419 7 1 2 1412 1416
0 1420 5 1 1 1419
0 1421 7 2 2 3242 1420
0 1422 5 1 1 3244
0 1423 7 2 2 1964 2057
0 1424 5 1 1 3246
0 1425 7 2 2 1975 2046
0 1426 5 1 1 3248
0 1427 7 2 2 3247 3249
0 1428 5 2 1 3250
0 1429 7 1 2 3245 3251
0 1430 5 2 1 1429
0 1431 7 2 2 3243 3254
0 1432 5 1 1 3256
0 1433 7 1 2 1400 3235
0 1434 5 1 1 1433
0 1435 7 2 2 3236 1434
0 1436 5 1 1 3258
0 1437 7 1 2 1432 3259
0 1438 5 2 1 1437
0 1439 7 2 2 3237 3260
0 1440 5 1 1 3262
0 1441 7 1 2 1380 3229
0 1442 5 1 1 1441
0 1443 7 2 2 3230 1442
0 1444 5 1 1 3264
0 1445 7 1 2 1440 3265
0 1446 5 2 1 1445
0 1447 7 2 2 3231 3266
0 1448 5 1 1 3268
0 1449 7 1 2 3206 1374
0 1450 5 1 1 1449
0 1451 7 2 2 3209 1450
0 1452 5 1 1 3270
0 1453 7 1 2 1448 3271
0 1454 5 2 1 1453
0 1455 7 2 2 3210 3272
0 1456 5 1 1 3274
0 1457 7 1 2 3188 1350
0 1458 5 1 1 1457
0 1459 7 2 2 3191 1458
0 1460 5 1 1 3276
0 1461 7 1 2 1456 3277
0 1462 5 2 1 1461
0 1463 7 2 2 3192 3278
0 1464 5 1 1 3280
0 1465 7 1 2 3158 1308
0 1466 5 1 1 1465
0 1467 7 2 2 3161 1466
0 1468 5 1 1 3282
0 1469 7 1 2 1464 3283
0 1470 5 2 1 1469
0 1471 7 2 2 3162 3284
0 1472 5 1 1 3286
0 1473 7 1 2 3116 1252
0 1474 5 1 1 1473
0 1475 7 2 2 3119 1474
0 1476 5 1 1 3288
0 1477 7 1 2 1472 3289
0 1478 5 2 1 1477
0 1479 7 2 2 3120 3290
0 1480 5 1 1 3292
0 1481 7 1 2 3074 1192
0 1482 5 1 1 1481
0 1483 7 2 2 3077 1482
0 1484 5 1 1 3294
0 1485 7 1 2 1480 3295
0 1486 5 2 1 1485
0 1487 7 2 2 3078 3296
0 1488 5 1 1 3298
0 1489 7 1 2 3032 1134
0 1490 5 1 1 1489
0 1491 7 2 2 3035 1490
0 1492 5 1 1 3300
0 1493 7 1 2 1488 3301
0 1494 5 2 1 1493
0 1495 7 2 2 3036 3302
0 1496 5 1 1 3304
0 1497 7 1 2 2946 1038
0 1498 5 1 1 1497
0 1499 7 2 2 2949 1498
0 1500 5 1 1 3306
0 1501 7 1 2 1496 3307
0 1502 5 2 1 1501
0 1503 7 2 2 2950 3308
0 1504 5 1 1 3310
0 1505 7 1 2 2868 932
0 1506 5 1 1 1505
0 1507 7 2 2 2871 1506
0 1508 5 1 1 3312
0 1509 7 1 2 1504 3313
0 1510 5 2 1 1509
0 1511 7 2 2 2872 3314
0 1512 5 1 1 3316
0 1513 7 1 2 2792 840
0 1514 5 1 1 1513
0 1515 7 2 2 2795 1514
0 1516 5 1 1 3318
0 1517 7 1 2 1512 3319
0 1518 5 2 1 1517
0 1519 7 2 2 2796 3320
0 1520 5 1 1 3322
0 1521 7 1 2 2740 742
0 1522 5 1 1 1521
0 1523 7 2 2 2741 1522
0 1524 5 1 1 3324
0 1525 7 1 2 1520 3325
0 1526 5 2 1 1525
0 1527 7 2 2 2742 3326
0 1528 5 1 1 3328
0 1529 7 2 2 2246 1528
0 1530 5 3 1 3330
0 1531 7 1 2 3323 1524
0 1532 5 1 1 1531
0 1533 7 2 2 3327 1532
0 1534 5 1 1 3335
0 1535 7 1 2 2165 1534
0 1536 5 3 1 1535
0 1537 7 2 2 2169 3329
0 1538 5 1 1 3340
0 1539 7 2 2 3337 1538
0 1540 5 1 1 3342
0 1541 7 1 2 3332 1540
0 1542 5 2 1 1541
0 1543 7 1 2 3317 1516
0 1544 5 1 1 1543
0 1545 7 2 2 3321 1544
0 1546 5 1 1 3346
0 1547 7 1 2 2161 1546
0 1548 5 3 1 1547
0 1549 7 1 2 3311 1508
0 1550 5 1 1 1549
0 1551 7 2 2 3315 1550
0 1552 5 1 1 3351
0 1553 7 1 2 2158 1552
0 1554 5 6 1 1553
0 1555 7 1 2 3305 1500
0 1556 5 1 1 1555
0 1557 7 2 2 3309 1556
0 1558 5 1 1 3359
0 1559 7 1 2 2154 1558
0 1560 5 4 1 1559
0 1561 7 1 2 3299 1492
0 1562 5 1 1 1561
0 1563 7 2 2 3303 1562
0 1564 5 1 1 3365
0 1565 7 1 2 2151 1564
0 1566 5 4 1 1565
0 1567 7 1 2 2232 3366
0 1568 5 4 1 1567
0 1569 7 1 2 3293 1484
0 1570 5 1 1 1569
0 1571 7 2 2 3297 1570
0 1572 5 1 1 3375
0 1573 7 1 2 2148 1572
0 1574 5 3 1 1573
0 1575 7 1 2 2229 3376
0 1576 5 4 1 1575
0 1577 7 1 2 3287 1476
0 1578 5 1 1 1577
0 1579 7 2 2 3291 1578
0 1580 5 1 1 3384
0 1581 7 1 2 2145 1580
0 1582 5 5 1 1581
0 1583 7 1 2 2226 3385
0 1584 5 4 1 1583
0 1585 7 1 2 3281 1468
0 1586 5 1 1 1585
0 1587 7 2 2 3285 1586
0 1588 5 1 1 3395
0 1589 7 1 2 2142 1588
0 1590 5 4 1 1589
0 1591 7 1 2 2223 3396
0 1592 5 4 1 1591
0 1593 7 1 2 3275 1460
0 1594 5 1 1 1593
0 1595 7 2 2 3279 1594
0 1596 5 1 1 3405
0 1597 7 1 2 2139 1596
0 1598 5 4 1 1597
0 1599 7 1 2 2220 3406
0 1600 5 4 1 1599
0 1601 7 1 2 3269 1452
0 1602 5 1 1 1601
0 1603 7 2 2 3273 1602
0 1604 5 1 1 3415
0 1605 7 1 2 2136 1604
0 1606 5 4 1 1605
0 1607 7 1 2 2217 3416
0 1608 5 4 1 1607
0 1609 7 1 2 3263 1444
0 1610 5 1 1 1609
0 1611 7 2 2 3267 1610
0 1612 5 1 1 3425
0 1613 7 1 2 2133 1612
0 1614 5 3 1 1613
0 1615 7 1 2 2214 3426
0 1616 5 4 1 1615
0 1617 7 1 2 3257 1436
0 1618 5 1 1 1617
0 1619 7 2 2 3261 1618
0 1620 5 1 1 3434
0 1621 7 1 2 2130 1620
0 1622 5 3 1 1621
0 1623 7 1 2 2211 3435
0 1624 5 4 1 1623
0 1625 7 1 2 1422 3252
0 1626 5 1 1 1625
0 1627 7 2 2 3255 1626
0 1628 5 1 1 3443
0 1629 7 1 2 2127 1628
0 1630 5 3 1 1629
0 1631 7 1 2 2208 3444
0 1632 5 3 1 1631
0 1633 7 1 2 1424 1426
0 1634 5 1 1 1633
0 1635 7 2 2 3253 1634
0 1636 5 1 1 3451
0 1637 7 1 2 2205 3452
0 1638 5 2 1 1637
0 1639 7 2 2 2124 1636
0 1640 5 1 1 3455
0 1641 7 2 2 1965 2047
0 1642 5 1 1 3457
0 1643 7 1 2 2121 1642
0 1644 5 1 1 1643
0 1645 7 2 2 1640 1644
0 1646 5 1 1 3459
0 1647 7 1 2 3453 1646
0 1648 7 1 2 3448 1647
0 1649 5 1 1 1648
0 1650 7 2 2 3445 1649
0 1651 5 2 1 3461
0 1652 7 1 2 3439 3463
0 1653 5 1 1 1652
0 1654 7 2 2 3436 1653
0 1655 5 2 1 3465
0 1656 7 1 2 3430 3467
0 1657 5 1 1 1656
0 1658 7 2 2 3427 1657
0 1659 5 2 1 3469
0 1660 7 1 2 3421 3471
0 1661 5 1 1 1660
0 1662 7 2 2 3417 1661
0 1663 5 2 1 3473
0 1664 7 1 2 3411 3475
0 1665 5 1 1 1664
0 1666 7 2 2 3407 1665
0 1667 5 2 1 3477
0 1668 7 1 2 3401 3479
0 1669 5 1 1 1668
0 1670 7 2 2 3397 1669
0 1671 5 1 1 3481
0 1672 7 2 2 3391 1671
0 1673 5 1 1 3483
0 1674 7 2 2 3386 1673
0 1675 5 2 1 3485
0 1676 7 1 2 3380 3487
0 1677 5 1 1 1676
0 1678 7 2 2 3377 1677
0 1679 5 1 1 3489
0 1680 7 2 2 3371 1679
0 1681 5 1 1 3491
0 1682 7 2 2 3367 1681
0 1683 7 1 2 3361 3493
0 1684 5 1 1 1683
0 1685 7 1 2 2239 3352
0 1686 5 2 1 1685
0 1687 7 1 2 2235 3360
0 1688 5 5 1 1687
0 1689 7 3 2 3495 3497
0 1690 7 2 2 1684 3502
0 1691 5 1 1 3505
0 1692 7 2 2 3353 1691
0 1693 5 2 1 3507
0 1694 7 1 2 2242 3347
0 1695 5 4 1 1694
0 1696 7 1 2 3509 3511
0 1697 5 1 1 1696
0 1698 7 2 2 3348 1697
0 1699 5 1 1 3515
0 1700 7 1 2 2244 3336
0 1701 5 4 1 1700
0 1702 7 1 2 3333 3517
0 1703 7 1 2 1699 1702
0 1704 5 1 1 1703
0 1705 7 3 2 3344 1704
0 1706 5 1 1 3521
0 1707 7 1 2 3338 3331
0 1708 5 1 1 1707
0 1709 7 2 2 3354 3496
0 1710 5 1 1 3524
0 1711 7 1 2 3498 3525
0 1712 5 1 1 1711
0 1713 7 1 2 3494 1712
0 1714 5 1 1 1713
0 1715 7 1 2 3355 3506
0 1716 5 1 1 1715
0 1717 7 2 2 3362 1710
0 1718 5 1 1 3526
0 1719 7 3 2 3378 3381
0 1720 5 2 1 3528
0 1721 7 1 2 3486 3531
0 1722 5 1 1 1721
0 1723 7 1 2 3488 3529
0 1724 5 1 1 1723
0 1725 7 1 2 1722 1724
0 1726 5 1 1 1725
0 1727 7 1 2 3387 3484
0 1728 5 1 1 1727
0 1729 7 1 2 3388 3392
0 1730 5 2 1 1729
0 1731 7 1 2 3482 3533
0 1732 5 1 1 1731
0 1733 7 1 2 1728 1732
0 1734 5 1 1 1733
0 1735 7 2 2 3398 3402
0 1736 5 2 1 3535
0 1737 7 1 2 3480 3537
0 1738 5 1 1 1737
0 1739 7 1 2 3478 3536
0 1740 5 1 1 1739
0 1741 7 3 2 3408 3412
0 1742 5 1 1 3539
0 1743 7 1 2 3476 1742
0 1744 5 1 1 1743
0 1745 7 1 2 3474 3540
0 1746 5 1 1 1745
0 1747 7 2 2 3418 3422
0 1748 5 2 1 3542
0 1749 7 1 2 3470 3543
0 1750 5 1 1 1749
0 1751 7 1 2 2202 3458
0 1752 5 1 1 1751
0 1753 7 1 2 3454 1752
0 1754 7 3 2 3449 1753
0 1755 5 1 1 3546
0 1756 7 1 2 3446 3460
0 1757 7 1 2 3547 1756
0 1758 5 2 1 1757
0 1759 7 3 2 3437 3440
0 1760 5 2 1 3551
0 1761 7 1 2 3462 3554
0 1762 5 1 1 1761
0 1763 7 1 2 3464 3552
0 1764 5 1 1 1763
0 1765 7 1 2 1762 1764
0 1766 5 1 1 1765
0 1767 7 1 2 3549 1766
0 1768 5 1 1 1767
0 1769 7 3 2 3428 3431
0 1770 5 2 1 3556
0 1771 7 1 2 3468 3559
0 1772 5 1 1 1771
0 1773 7 1 2 3466 3557
0 1774 5 1 1 1773
0 1775 7 1 2 1772 1774
0 1776 5 1 1 1775
0 1777 7 1 2 1768 1776
0 1778 5 1 1 1777
0 1779 7 1 2 3472 3544
0 1780 5 1 1 1779
0 1781 7 1 2 1778 1780
0 1782 7 1 2 1750 1781
0 1783 7 1 2 1746 1782
0 1784 7 1 2 1744 1783
0 1785 7 1 2 1740 1784
0 1786 7 1 2 1738 1785
0 1787 7 1 2 1734 1786
0 1788 7 1 2 1726 1787
0 1789 5 1 1 1788
0 1790 7 1 2 3368 3492
0 1791 5 1 1 1790
0 1792 7 2 2 3369 3372
0 1793 5 2 1 3561
0 1794 7 1 2 3490 3563
0 1795 5 1 1 1794
0 1796 7 1 2 1791 1795
0 1797 7 1 2 1789 1796
0 1798 7 1 2 1718 1797
0 1799 7 1 2 1716 1798
0 1800 7 1 2 1714 1799
0 1801 7 3 2 3349 3512
0 1802 5 2 1 3565
0 1803 7 1 2 3508 3568
0 1804 5 1 1 1803
0 1805 7 1 2 3510 3566
0 1806 5 1 1 1805
0 1807 7 1 2 1804 1806
0 1808 7 1 2 1800 1807
0 1809 7 1 2 1708 1808
0 1810 7 1 2 3339 3518
0 1811 5 2 1 1810
0 1812 7 1 2 3570 3516
0 1813 5 1 1 1812
0 1814 7 1 2 3345 1813
0 1815 7 1 2 1809 1814
0 1816 7 1 2 3522 1815
0 1817 5 1 1 1816
0 1818 7 1 2 3450 3456
0 1819 5 1 1 1818
0 1820 7 1 2 3447 1755
0 1821 7 2 2 1819 1820
0 1822 5 2 1 3572
0 1823 7 1 2 3441 3574
0 1824 5 1 1 1823
0 1825 7 2 2 3438 1824
0 1826 5 2 1 3576
0 1827 7 1 2 3432 3578
0 1828 5 1 1 1827
0 1829 7 2 2 3429 1828
0 1830 5 1 1 3580
0 1831 7 1 2 3423 1830
0 1832 5 2 1 1831
0 1833 7 1 2 3419 3582
0 1834 7 1 2 3409 1833
0 1835 5 1 1 1834
0 1836 7 1 2 3413 1835
0 1837 7 1 2 3403 1836
0 1838 5 1 1 1837
0 1839 7 1 2 3399 1838
0 1840 5 1 1 1839
0 1841 7 1 2 3393 1840
0 1842 5 1 1 1841
0 1843 7 1 2 3389 1842
0 1844 5 2 1 1843
0 1845 7 1 2 3382 3584
0 1846 5 1 1 1845
0 1847 7 2 2 3379 1846
0 1848 5 2 1 3586
0 1849 7 1 2 3373 3588
0 1850 5 1 1 1849
0 1851 7 2 2 3370 1850
0 1852 5 2 1 3590
0 1853 7 2 2 3363 3591
0 1854 5 1 1 3594
0 1855 7 2 2 3503 1854
0 1856 5 1 1 3596
0 1857 7 1 2 3356 1856
0 1858 5 2 1 1857
0 1859 7 1 2 3513 3598
0 1860 5 1 1 1859
0 1861 7 2 2 3350 1860
0 1862 5 1 1 3600
0 1863 7 1 2 3343 3601
0 1864 5 1 1 1863
0 1865 7 1 2 3341 3519
0 1866 5 1 1 1865
0 1867 7 1 2 3569 3599
0 1868 5 1 1 1867
0 1869 7 1 2 3364 3499
0 1870 5 1 1 1869
0 1871 7 1 2 3592 1870
0 1872 5 1 1 1871
0 1873 7 1 2 3500 3595
0 1874 5 1 1 1873
0 1875 7 1 2 3562 3589
0 1876 5 1 1 1875
0 1877 7 1 2 3564 3587
0 1878 5 1 1 1877
0 1879 7 1 2 1876 1878
0 1880 5 1 1 1879
0 1881 7 1 2 3390 3532
0 1882 5 1 1 1881
0 1883 7 1 2 3530 3585
0 1884 5 1 1 1883
0 1885 7 1 2 3400 3534
0 1886 5 1 1 1885
0 1887 7 1 2 3410 3538
0 1888 5 1 1 1887
0 1889 7 1 2 3541 3583
0 1890 5 1 1 1889
0 1891 7 1 2 3420 1890
0 1892 5 1 1 1891
0 1893 7 1 2 3545 3581
0 1894 5 1 1 1893
0 1895 7 1 2 3558 3577
0 1896 5 1 1 1895
0 1897 7 1 2 3555 3575
0 1898 5 1 1 1897
0 1899 7 1 2 3553 3573
0 1900 5 1 1 1899
0 1901 7 1 2 1898 1900
0 1902 5 1 1 1901
0 1903 7 1 2 3550 1902
0 1904 5 1 1 1903
0 1905 7 1 2 3560 3579
0 1906 5 1 1 1905
0 1907 7 1 2 1904 1906
0 1908 7 1 2 1896 1907
0 1909 5 1 1 1908
0 1910 7 1 2 1894 1909
0 1911 7 1 2 1892 1910
0 1912 7 1 2 1888 1911
0 1913 7 1 2 1886 1912
0 1914 7 1 2 1884 1913
0 1915 7 1 2 1882 1914
0 1916 5 1 1 1915
0 1917 7 1 2 1880 1916
0 1918 7 1 2 1874 1917
0 1919 7 1 2 1872 1918
0 1920 7 1 2 1868 1919
0 1921 7 1 2 1866 1920
0 1922 7 1 2 1864 1921
0 1923 7 1 2 3357 3597
0 1924 5 1 1 1923
0 1925 7 1 2 3358 3567
0 1926 5 1 1 1925
0 1927 7 1 2 3501 3593
0 1928 5 1 1 1927
0 1929 7 1 2 3527 1928
0 1930 7 1 2 1926 1929
0 1931 5 1 1 1930
0 1932 7 1 2 1924 1931
0 1933 5 1 1 1932
0 1934 7 1 2 3571 1862
0 1935 5 1 1 1934
0 1936 7 1 2 1933 1935
0 1937 7 1 2 1922 1936
0 1938 7 1 2 1706 1937
0 1939 5 1 1 1938
0 1940 7 1 2 1817 1939
0 1941 7 1 2 2713 1940
0 1942 5 1 1 1941
0 1943 7 1 2 3442 3548
0 1944 7 1 2 3433 1943
0 1945 7 1 2 3424 1944
0 1946 7 1 2 3414 1945
0 1947 7 1 2 3404 1946
0 1948 7 1 2 3394 1947
0 1949 7 1 2 3383 1948
0 1950 7 1 2 3374 1949
0 1951 7 1 2 3504 1950
0 1952 7 1 2 3514 1951
0 1953 7 1 2 3334 1952
0 1954 7 1 2 3520 1953
0 1955 7 1 2 3523 1954
0 1956 5 1 1 1955
0 1957 7 1 2 740 1956
0 1958 5 1 1 1957
3 4099 7 0 2 1942 1958
