1 0 0 8 0
2 32 1 0
2 1233 1 0
2 1234 1 0
2 1235 1 0
2 1236 1 0
2 1237 1 0
2 1238 1 0
2 1239 1 0
1 1 0 8 0
2 1240 1 1
2 1241 1 1
2 1242 1 1
2 1243 1 1
2 1244 1 1
2 1245 1 1
2 1246 1 1
2 1247 1 1
1 2 0 8 0
2 1248 1 2
2 1249 1 2
2 1250 1 2
2 1251 1 2
2 1252 1 2
2 1253 1 2
2 1254 1 2
2 1255 1 2
1 3 0 9 0
2 1256 1 3
2 1257 1 3
2 1258 1 3
2 1259 1 3
2 1260 1 3
2 1261 1 3
2 1262 1 3
2 1263 1 3
2 1264 1 3
1 4 0 8 0
2 1265 1 4
2 1266 1 4
2 1267 1 4
2 1268 1 4
2 1269 1 4
2 1270 1 4
2 1271 1 4
2 1272 1 4
1 5 0 9 0
2 1273 1 5
2 1274 1 5
2 1275 1 5
2 1276 1 5
2 1277 1 5
2 1278 1 5
2 1279 1 5
2 1280 1 5
2 1281 1 5
1 6 0 8 0
2 1282 1 6
2 1283 1 6
2 1284 1 6
2 1285 1 6
2 1286 1 6
2 1287 1 6
2 1288 1 6
2 1289 1 6
1 7 0 8 0
2 1290 1 7
2 1291 1 7
2 1292 1 7
2 1293 1 7
2 1294 1 7
2 1295 1 7
2 1296 1 7
2 1297 1 7
1 8 0 8 0
2 1298 1 8
2 1299 1 8
2 1300 1 8
2 1301 1 8
2 1302 1 8
2 1303 1 8
2 1304 1 8
2 1305 1 8
1 9 0 8 0
2 1306 1 9
2 1307 1 9
2 1308 1 9
2 1309 1 9
2 1310 1 9
2 1311 1 9
2 1312 1 9
2 1313 1 9
1 10 0 9 0
2 1314 1 10
2 1315 1 10
2 1316 1 10
2 1317 1 10
2 1318 1 10
2 1319 1 10
2 1320 1 10
2 1321 1 10
2 1322 1 10
1 11 0 8 0
2 1323 1 11
2 1324 1 11
2 1325 1 11
2 1326 1 11
2 1327 1 11
2 1328 1 11
2 1329 1 11
2 1330 1 11
1 12 0 8 0
2 1331 1 12
2 1332 1 12
2 1333 1 12
2 1334 1 12
2 1335 1 12
2 1336 1 12
2 1337 1 12
2 1338 1 12
1 13 0 8 0
2 1339 1 13
2 1340 1 13
2 1341 1 13
2 1342 1 13
2 1343 1 13
2 1344 1 13
2 1345 1 13
2 1346 1 13
1 14 0 8 0
2 1347 1 14
2 1348 1 14
2 1349 1 14
2 1350 1 14
2 1351 1 14
2 1352 1 14
2 1353 1 14
2 1354 1 14
1 15 0 8 0
2 1355 1 15
2 1356 1 15
2 1357 1 15
2 1358 1 15
2 1359 1 15
2 1360 1 15
2 1361 1 15
2 1362 1 15
1 16 0 2 0
2 1363 1 16
2 1364 1 16
1 17 0 3 0
2 1365 1 17
2 1366 1 17
2 1367 1 17
1 18 0 3 0
2 1368 1 18
2 1369 1 18
2 1370 1 18
1 19 0 3 0
2 1371 1 19
2 1372 1 19
2 1373 1 19
1 20 0 3 0
2 1374 1 20
2 1375 1 20
2 1376 1 20
1 21 0 3 0
2 1377 1 21
2 1378 1 21
2 1379 1 21
1 22 0 3 0
2 1380 1 22
2 1381 1 22
2 1382 1 22
1 23 0 3 0
2 1383 1 23
2 1384 1 23
2 1385 1 23
1 24 0 3 0
2 1386 1 24
2 1387 1 24
2 1388 1 24
1 25 0 3 0
2 1389 1 25
2 1390 1 25
2 1391 1 25
1 26 0 3 0
2 1392 1 26
2 1393 1 26
2 1394 1 26
1 27 0 3 0
2 1395 1 27
2 1396 1 27
2 1397 1 27
1 28 0 3 0
2 1398 1 28
2 1399 1 28
2 1400 1 28
1 29 0 3 0
2 1401 1 29
2 1402 1 29
2 1403 1 29
1 30 0 3 0
2 1404 1 30
2 1405 1 30
2 1406 1 30
1 31 0 2 0
2 1407 1 31
2 1408 1 31
2 1409 1 35
2 1410 1 35
2 1411 1 36
2 1412 1 36
2 1413 1 37
2 1414 1 37
2 1415 1 38
2 1416 1 38
2 1417 1 39
2 1418 1 39
2 1419 1 40
2 1420 1 40
2 1421 1 41
2 1422 1 41
2 1423 1 42
2 1424 1 42
2 1425 1 43
2 1426 1 43
2 1427 1 44
2 1428 1 44
2 1429 1 45
2 1430 1 45
2 1431 1 46
2 1432 1 46
2 1433 1 47
2 1434 1 47
2 1435 1 48
2 1436 1 48
2 1437 1 48
2 1438 1 49
2 1439 1 49
2 1440 1 51
2 1441 1 51
2 1442 1 54
2 1443 1 54
2 1444 1 55
2 1445 1 55
2 1446 1 59
2 1447 1 59
2 1448 1 62
2 1449 1 62
2 1450 1 63
2 1451 1 63
2 1452 1 65
2 1453 1 65
2 1454 1 66
2 1455 1 66
2 1456 1 67
2 1457 1 67
2 1458 1 69
2 1459 1 69
2 1460 1 74
2 1461 1 74
2 1462 1 75
2 1463 1 75
2 1464 1 78
2 1465 1 78
2 1466 1 81
2 1467 1 81
2 1468 1 84
2 1469 1 84
2 1470 1 85
2 1471 1 85
2 1472 1 89
2 1473 1 89
2 1474 1 92
2 1475 1 92
2 1476 1 93
2 1477 1 93
2 1478 1 95
2 1479 1 95
2 1480 1 98
2 1481 1 98
2 1482 1 99
2 1483 1 99
2 1484 1 103
2 1485 1 103
2 1486 1 106
2 1487 1 106
2 1488 1 107
2 1489 1 107
2 1490 1 111
2 1491 1 111
2 1492 1 114
2 1493 1 114
2 1494 1 115
2 1495 1 115
2 1496 1 119
2 1497 1 119
2 1498 1 122
2 1499 1 122
2 1500 1 123
2 1501 1 123
2 1502 1 125
2 1503 1 125
2 1504 1 127
2 1505 1 127
2 1506 1 129
2 1507 1 129
2 1508 1 135
2 1509 1 135
2 1510 1 138
2 1511 1 138
2 1512 1 138
2 1513 1 141
2 1514 1 141
2 1515 1 144
2 1516 1 144
2 1517 1 145
2 1518 1 145
2 1519 1 149
2 1520 1 149
2 1521 1 152
2 1522 1 152
2 1523 1 153
2 1524 1 153
2 1525 1 157
2 1526 1 157
2 1527 1 160
2 1528 1 160
2 1529 1 161
2 1530 1 161
2 1531 1 165
2 1532 1 165
2 1533 1 168
2 1534 1 168
2 1535 1 169
2 1536 1 169
2 1537 1 171
2 1538 1 171
2 1539 1 173
2 1540 1 173
2 1541 1 175
2 1542 1 175
2 1543 1 176
2 1544 1 176
2 1545 1 177
2 1546 1 177
2 1547 1 178
2 1548 1 178
2 1549 1 180
2 1550 1 180
2 1551 1 181
2 1552 1 181
2 1553 1 185
2 1554 1 185
2 1555 1 188
2 1556 1 188
2 1557 1 189
2 1558 1 189
2 1559 1 193
2 1560 1 193
2 1561 1 196
2 1562 1 196
2 1563 1 197
2 1564 1 197
2 1565 1 201
2 1566 1 201
2 1567 1 204
2 1568 1 204
2 1569 1 205
2 1570 1 205
2 1571 1 209
2 1572 1 209
2 1573 1 212
2 1574 1 212
2 1575 1 213
2 1576 1 213
2 1577 1 217
2 1578 1 217
2 1579 1 220
2 1580 1 220
2 1581 1 221
2 1582 1 221
2 1583 1 225
2 1584 1 225
2 1585 1 228
2 1586 1 228
2 1587 1 229
2 1588 1 229
2 1589 1 233
2 1590 1 233
2 1591 1 236
2 1592 1 236
2 1593 1 237
2 1594 1 237
2 1595 1 239
2 1596 1 239
2 1597 1 242
2 1598 1 242
2 1599 1 245
2 1600 1 245
2 1601 1 249
2 1602 1 249
2 1603 1 252
2 1604 1 252
2 1605 1 253
2 1606 1 253
2 1607 1 257
2 1608 1 257
2 1609 1 260
2 1610 1 260
2 1611 1 261
2 1612 1 261
2 1613 1 263
2 1614 1 263
2 1615 1 266
2 1616 1 266
2 1617 1 267
2 1618 1 267
2 1619 1 269
2 1620 1 269
2 1621 1 275
2 1622 1 275
2 1623 1 278
2 1624 1 278
2 1625 1 281
2 1626 1 281
2 1627 1 284
2 1628 1 284
2 1629 1 287
2 1630 1 287
2 1631 1 291
2 1632 1 291
2 1633 1 294
2 1634 1 294
2 1635 1 295
2 1636 1 295
2 1637 1 299
2 1638 1 299
2 1639 1 302
2 1640 1 302
2 1641 1 303
2 1642 1 303
2 1643 1 305
2 1644 1 305
2 1645 1 308
2 1646 1 308
2 1647 1 311
2 1648 1 311
2 1649 1 315
2 1650 1 315
2 1651 1 318
2 1652 1 318
2 1653 1 319
2 1654 1 319
2 1655 1 323
2 1656 1 323
2 1657 1 326
2 1658 1 326
2 1659 1 327
2 1660 1 327
2 1661 1 331
2 1662 1 331
2 1663 1 334
2 1664 1 334
2 1665 1 335
2 1666 1 335
2 1667 1 339
2 1668 1 339
2 1669 1 342
2 1670 1 342
2 1671 1 343
2 1672 1 343
2 1673 1 347
2 1674 1 347
2 1675 1 350
2 1676 1 350
2 1677 1 351
2 1678 1 351
2 1679 1 353
2 1680 1 353
2 1681 1 356
2 1682 1 356
2 1683 1 357
2 1684 1 357
2 1685 1 361
2 1686 1 361
2 1687 1 364
2 1688 1 364
2 1689 1 365
2 1690 1 365
2 1691 1 367
2 1692 1 367
2 1693 1 369
2 1694 1 369
2 1695 1 372
2 1696 1 372
2 1697 1 373
2 1698 1 373
2 1699 1 375
2 1700 1 375
2 1701 1 377
2 1702 1 377
2 1703 1 379
2 1704 1 379
2 1705 1 381
2 1706 1 381
2 1707 1 382
2 1708 1 382
2 1709 1 383
2 1710 1 383
2 1711 1 384
2 1712 1 384
2 1713 1 385
2 1714 1 385
2 1715 1 386
2 1716 1 386
2 1717 1 387
2 1718 1 387
2 1719 1 388
2 1720 1 388
2 1721 1 390
2 1722 1 390
2 1723 1 393
2 1724 1 393
2 1725 1 397
2 1726 1 397
2 1727 1 400
2 1728 1 400
2 1729 1 403
2 1730 1 403
2 1731 1 407
2 1732 1 407
2 1733 1 410
2 1734 1 410
2 1735 1 411
2 1736 1 411
2 1737 1 414
2 1738 1 414
2 1739 1 415
2 1740 1 415
2 1741 1 419
2 1742 1 419
2 1743 1 422
2 1744 1 422
2 1745 1 423
2 1746 1 423
2 1747 1 427
2 1748 1 427
2 1749 1 430
2 1750 1 430
2 1751 1 431
2 1752 1 431
2 1753 1 435
2 1754 1 435
2 1755 1 438
2 1756 1 438
2 1757 1 441
2 1758 1 441
2 1759 1 445
2 1760 1 445
2 1761 1 448
2 1762 1 448
2 1763 1 451
2 1764 1 451
2 1765 1 455
2 1766 1 455
2 1767 1 458
2 1768 1 458
2 1769 1 459
2 1770 1 459
2 1771 1 461
2 1772 1 461
2 1773 1 464
2 1774 1 464
2 1775 1 465
2 1776 1 465
2 1777 1 469
2 1778 1 469
2 1779 1 472
2 1780 1 472
2 1781 1 473
2 1782 1 473
2 1783 1 477
2 1784 1 477
2 1785 1 480
2 1786 1 480
2 1787 1 481
2 1788 1 481
2 1789 1 485
2 1790 1 485
2 1791 1 488
2 1792 1 488
2 1793 1 489
2 1794 1 489
2 1795 1 493
2 1796 1 493
2 1797 1 496
2 1798 1 496
2 1799 1 497
2 1800 1 497
2 1801 1 501
2 1802 1 501
2 1803 1 504
2 1804 1 504
2 1805 1 505
2 1806 1 505
2 1807 1 507
2 1808 1 507
2 1809 1 513
2 1810 1 513
2 1811 1 516
2 1812 1 516
2 1813 1 519
2 1814 1 519
2 1815 1 522
2 1816 1 522
2 1817 1 525
2 1818 1 525
2 1819 1 529
2 1820 1 529
2 1821 1 532
2 1822 1 532
2 1823 1 533
2 1824 1 533
2 1825 1 537
2 1826 1 537
2 1827 1 540
2 1828 1 540
2 1829 1 541
2 1830 1 541
2 1831 1 545
2 1832 1 545
2 1833 1 548
2 1834 1 548
2 1835 1 549
2 1836 1 549
2 1837 1 553
2 1838 1 553
2 1839 1 556
2 1840 1 556
2 1841 1 557
2 1842 1 557
2 1843 1 561
2 1844 1 561
2 1845 1 564
2 1846 1 564
2 1847 1 565
2 1848 1 565
2 1849 1 569
2 1850 1 569
2 1851 1 572
2 1852 1 572
2 1853 1 573
2 1854 1 573
2 1855 1 577
2 1856 1 577
2 1857 1 580
2 1858 1 580
2 1859 1 581
2 1860 1 581
2 1861 1 583
2 1862 1 583
2 1863 1 586
2 1864 1 586
2 1865 1 589
2 1866 1 589
2 1867 1 593
2 1868 1 593
2 1869 1 596
2 1870 1 596
2 1871 1 597
2 1872 1 597
2 1873 1 601
2 1874 1 601
2 1875 1 604
2 1876 1 604
2 1877 1 605
2 1878 1 605
2 1879 1 609
2 1880 1 609
2 1881 1 612
2 1882 1 612
2 1883 1 613
2 1884 1 613
2 1885 1 617
2 1886 1 617
2 1887 1 620
2 1888 1 620
2 1889 1 621
2 1890 1 621
2 1891 1 627
2 1892 1 627
2 1893 1 630
2 1894 1 630
2 1895 1 631
2 1896 1 631
2 1897 1 635
2 1898 1 635
2 1899 1 638
2 1900 1 638
2 1901 1 639
2 1902 1 639
2 1903 1 643
2 1904 1 643
2 1905 1 646
2 1906 1 646
2 1907 1 647
2 1908 1 647
2 1909 1 651
2 1910 1 651
2 1911 1 654
2 1912 1 654
2 1913 1 655
2 1914 1 655
2 1915 1 657
2 1916 1 657
2 1917 1 660
2 1918 1 660
2 1919 1 663
2 1920 1 663
2 1921 1 667
2 1922 1 667
2 1923 1 670
2 1924 1 670
2 1925 1 671
2 1926 1 671
2 1927 1 675
2 1928 1 675
2 1929 1 678
2 1930 1 678
2 1931 1 681
2 1932 1 681
2 1933 1 683
2 1934 1 683
2 1935 1 685
2 1936 1 685
2 1937 1 687
2 1938 1 687
2 1939 1 689
2 1940 1 689
2 1941 1 691
2 1942 1 691
2 1943 1 693
2 1944 1 693
2 1945 1 694
2 1946 1 694
2 1947 1 695
2 1948 1 695
2 1949 1 695
2 1950 1 698
2 1951 1 698
2 1952 1 701
2 1953 1 701
2 1954 1 709
2 1955 1 709
2 1956 1 712
2 1957 1 712
2 1958 1 713
2 1959 1 713
2 1960 1 717
2 1961 1 717
2 1962 1 720
2 1963 1 720
2 1964 1 723
2 1965 1 723
2 1966 1 725
2 1967 1 725
2 1968 1 727
2 1969 1 727
2 1970 1 729
2 1971 1 729
2 1972 1 730
2 1973 1 730
2 1974 1 732
2 1975 1 732
2 1976 1 733
2 1977 1 733
2 1978 1 737
2 1979 1 737
2 1980 1 740
2 1981 1 740
2 1982 1 741
2 1983 1 741
2 1984 1 745
2 1985 1 745
2 1986 1 748
2 1987 1 748
2 1988 1 749
2 1989 1 749
2 1990 1 753
2 1991 1 753
2 1992 1 756
2 1993 1 756
2 1994 1 757
2 1995 1 757
2 1996 1 761
2 1997 1 761
2 1998 1 764
2 1999 1 764
2 2000 1 765
2 2001 1 765
2 2002 1 769
2 2003 1 769
2 2004 1 772
2 2005 1 772
2 2006 1 773
2 2007 1 773
2 2008 1 777
2 2009 1 777
2 2010 1 780
2 2011 1 780
2 2012 1 781
2 2013 1 781
2 2014 1 785
2 2015 1 785
2 2016 1 788
2 2017 1 788
2 2018 1 789
2 2019 1 789
2 2020 1 793
2 2021 1 793
2 2022 1 796
2 2023 1 796
2 2024 1 797
2 2025 1 797
2 2026 1 801
2 2027 1 801
2 2028 1 804
2 2029 1 804
2 2030 1 805
2 2031 1 805
2 2032 1 809
2 2033 1 809
2 2034 1 812
2 2035 1 812
2 2036 1 813
2 2037 1 813
2 2038 1 817
2 2039 1 817
2 2040 1 820
2 2041 1 820
2 2042 1 821
2 2043 1 821
2 2044 1 823
2 2045 1 823
2 2046 1 828
2 2047 1 828
2 2048 1 831
2 2049 1 831
2 2050 1 834
2 2051 1 834
2 2052 1 834
2 2053 1 836
2 2054 1 836
2 2055 1 837
2 2056 1 837
2 2057 1 838
2 2058 1 838
2 2059 1 841
2 2060 1 841
2 2061 1 842
2 2062 1 842
2 2063 1 844
2 2064 1 844
2 2065 1 846
2 2066 1 846
2 2067 1 849
2 2068 1 849
2 2069 1 850
2 2070 1 850
2 2071 1 852
2 2072 1 852
2 2073 1 854
2 2074 1 854
2 2075 1 857
2 2076 1 857
2 2077 1 858
2 2078 1 858
2 2079 1 860
2 2080 1 860
2 2081 1 862
2 2082 1 862
2 2083 1 865
2 2084 1 865
2 2085 1 865
2 2086 1 868
2 2087 1 868
2 2088 1 870
2 2089 1 870
2 2090 1 873
2 2091 1 873
2 2092 1 874
2 2093 1 874
2 2094 1 876
2 2095 1 876
2 2096 1 878
2 2097 1 878
2 2098 1 881
2 2099 1 881
2 2100 1 881
2 2101 1 884
2 2102 1 884
2 2103 1 886
2 2104 1 886
2 2105 1 889
2 2106 1 889
2 2107 1 890
2 2108 1 890
2 2109 1 892
2 2110 1 892
2 2111 1 894
2 2112 1 894
2 2113 1 897
2 2114 1 897
2 2115 1 897
2 2116 1 900
2 2117 1 900
2 2118 1 902
2 2119 1 902
2 2120 1 905
2 2121 1 905
2 2122 1 906
2 2123 1 906
2 2124 1 908
2 2125 1 908
2 2126 1 910
2 2127 1 910
2 2128 1 913
2 2129 1 913
2 2130 1 913
2 2131 1 916
2 2132 1 916
2 2133 1 918
2 2134 1 918
2 2135 1 919
2 2136 1 919
2 2137 1 921
2 2138 1 921
2 2139 1 921
2 2140 1 924
2 2141 1 924
2 2142 1 926
2 2143 1 926
2 2144 1 927
2 2145 1 927
2 2146 1 929
2 2147 1 929
2 2148 1 930
2 2149 1 930
2 2150 1 933
2 2151 1 933
2 2152 1 934
2 2153 1 934
2 2154 1 937
2 2155 1 937
2 2156 1 938
2 2157 1 938
2 2158 1 941
2 2159 1 941
2 2160 1 942
2 2161 1 942
2 2162 1 945
2 2163 1 945
2 2164 1 948
2 2165 1 948
2 2166 1 950
2 2167 1 950
2 2168 1 953
2 2169 1 953
2 2170 1 953
2 2171 1 954
2 2172 1 954
2 2173 1 957
2 2174 1 957
2 2175 1 960
2 2176 1 960
2 2177 1 962
2 2178 1 962
2 2179 1 965
2 2180 1 965
2 2181 1 965
2 2182 1 969
2 2183 1 969
2 2184 1 969
2 2185 1 973
2 2186 1 973
2 2187 1 974
2 2188 1 974
2 2189 1 977
2 2190 1 977
2 2191 1 978
2 2192 1 978
2 2193 1 981
2 2194 1 981
2 2195 1 982
2 2196 1 982
2 2197 1 985
2 2198 1 985
2 2199 1 986
2 2200 1 986
2 2201 1 989
2 2202 1 989
2 2203 1 990
2 2204 1 990
2 2205 1 993
2 2206 1 993
2 2207 1 994
2 2208 1 994
2 2209 1 997
2 2210 1 997
2 2211 1 997
2 2212 1 997
2 2213 1 1004
2 2214 1 1004
2 2215 1 1016
2 2216 1 1016
2 2217 1 1024
2 2218 1 1024
2 2219 1 1030
2 2220 1 1030
2 2221 1 1036
2 2222 1 1036
2 2223 1 1044
2 2224 1 1044
2 2225 1 1046
2 2226 1 1046
2 2227 1 1048
2 2228 1 1048
2 2229 1 1056
2 2230 1 1056
2 2231 1 1062
2 2232 1 1062
2 2233 1 1070
2 2234 1 1070
2 2235 1 1072
2 2236 1 1072
2 2237 1 1075
2 2238 1 1075
2 2239 1 1076
2 2240 1 1076
2 2241 1 1083
2 2242 1 1083
2 2243 1 1136
2 2244 1 1136
2 2245 1 1148
2 2246 1 1148
2 2247 1 1179
2 2248 1 1179
2 2249 1 1207
2 2250 1 1207
2 2251 1 1216
2 2252 1 1216
0 33 5 1 1 1363
0 34 5 1 1 1365
0 35 5 2 1 1368
0 36 5 2 1 1371
0 37 5 2 1 1374
0 38 5 2 1 1377
0 39 5 2 1 1380
0 40 5 2 1 1383
0 41 5 2 1 1386
0 42 5 2 1 1389
0 43 5 2 1 1392
0 44 5 2 1 1395
0 45 5 2 1 1398
0 46 5 2 1 1401
0 47 5 2 1 1404
0 48 5 3 1 1407
0 49 7 2 2 1265 1355
0 50 5 1 1 1438
0 51 7 2 2 1290 1331
0 52 5 1 1 1440
0 53 7 1 2 1439 1441
0 54 5 2 1 53
0 55 7 2 2 1282 1339
0 56 5 1 1 1444
0 57 7 1 2 50 52
0 58 5 1 1 57
0 59 7 2 2 1442 58
0 60 5 1 1 1446
0 61 7 1 2 1445 1447
0 62 5 2 1 61
0 63 7 2 2 1443 1448
0 64 5 1 1 1450
0 65 7 2 2 1283 1347
0 66 5 2 1 1452
0 67 7 2 2 1273 1356
0 68 5 1 1 1456
0 69 7 2 2 1291 1340
0 70 5 1 1 1458
0 71 7 1 2 68 70
0 72 5 1 1 71
0 73 7 1 2 1457 1459
0 74 5 2 1 73
0 75 7 2 2 72 1460
0 76 5 1 1 1462
0 77 7 1 2 1453 1463
0 78 5 2 1 77
0 79 7 1 2 1454 76
0 80 5 1 1 79
0 81 7 2 2 1464 80
0 82 5 1 1 1466
0 83 7 1 2 64 1467
0 84 5 2 1 83
0 85 7 2 2 1274 1348
0 86 5 1 1 1470
0 87 7 1 2 56 60
0 88 5 1 1 87
0 89 7 2 2 1449 88
0 90 5 1 1 1472
0 91 7 1 2 1471 1473
0 92 5 2 1 91
0 93 7 2 2 1256 1357
0 94 5 1 1 1476
0 95 7 2 2 1292 1323
0 96 5 1 1 1478
0 97 7 1 2 1477 1479
0 98 5 2 1 97
0 99 7 2 2 1284 1332
0 100 5 1 1 1482
0 101 7 1 2 94 96
0 102 5 1 1 101
0 103 7 2 2 1480 102
0 104 5 1 1 1484
0 105 7 1 2 1483 1485
0 106 5 2 1 105
0 107 7 2 2 1481 1486
0 108 5 1 1 1488
0 109 7 1 2 86 90
0 110 5 1 1 109
0 111 7 2 2 1474 110
0 112 5 1 1 1490
0 113 7 1 2 108 1491
0 114 5 2 1 113
0 115 7 2 2 1475 1492
0 116 5 1 1 1494
0 117 7 1 2 1451 82
0 118 5 1 1 117
0 119 7 2 2 1468 118
0 120 5 1 1 1496
0 121 7 1 2 116 1497
0 122 5 2 1 121
0 123 7 2 2 1469 1498
0 124 5 1 1 1500
0 125 7 2 2 1461 1465
0 126 5 1 1 1502
0 127 7 2 2 1285 1358
0 128 5 1 1 1504
0 129 7 2 2 1293 1349
0 130 5 1 1 1506
0 131 7 1 2 128 1507
0 132 5 1 1 131
0 133 7 1 2 1505 130
0 134 5 1 1 133
0 135 7 2 2 132 134
0 136 5 1 1 1508
0 137 7 1 2 126 136
0 138 5 3 1 137
0 139 7 1 2 1503 1509
0 140 5 1 1 139
0 141 7 2 2 1510 140
0 142 5 1 1 1513
0 143 7 1 2 124 1514
0 144 5 2 1 143
0 145 7 2 2 1266 1350
0 146 5 1 1 1517
0 147 7 1 2 100 104
0 148 5 1 1 147
0 149 7 2 2 1487 148
0 150 5 1 1 1519
0 151 7 1 2 1518 1520
0 152 5 2 1 151
0 153 7 2 2 1275 1341
0 154 5 1 1 1523
0 155 7 1 2 146 150
0 156 5 1 1 155
0 157 7 2 2 1521 156
0 158 5 1 1 1525
0 159 7 1 2 1524 1526
0 160 5 2 1 159
0 161 7 2 2 1522 1527
0 162 5 1 1 1529
0 163 7 1 2 1489 112
0 164 5 1 1 163
0 165 7 2 2 1493 164
0 166 5 1 1 1531
0 167 7 1 2 162 1532
0 168 5 2 1 167
0 169 7 2 2 1248 1359
0 170 5 1 1 1535
0 171 7 2 2 1294 1298
0 172 5 1 1 1537
0 173 7 2 2 1286 1306
0 174 5 1 1 1539
0 175 7 2 2 1538 1540
0 176 5 2 1 1541
0 177 7 2 2 1314 1542
0 178 5 2 1 1545
0 179 7 1 2 1536 1546
0 180 5 2 1 179
0 181 7 2 2 1295 1315
0 182 5 1 1 1551
0 183 7 1 2 170 1547
0 184 5 1 1 183
0 185 7 2 2 1549 184
0 186 5 1 1 1553
0 187 7 1 2 1552 1554
0 188 5 2 1 187
0 189 7 2 2 1550 1555
0 190 5 1 1 1557
0 191 7 1 2 154 158
0 192 5 1 1 191
0 193 7 2 2 1528 192
0 194 5 1 1 1559
0 195 7 1 2 190 1560
0 196 5 2 1 195
0 197 7 2 2 1276 1333
0 198 5 1 1 1563
0 199 7 1 2 182 186
0 200 5 1 1 199
0 201 7 2 2 1556 200
0 202 5 1 1 1565
0 203 7 1 2 1564 1566
0 204 5 2 1 203
0 205 7 2 2 1287 1324
0 206 5 1 1 1569
0 207 7 1 2 198 202
0 208 5 1 1 207
0 209 7 2 2 1567 208
0 210 5 1 1 1571
0 211 7 1 2 1570 1572
0 212 5 2 1 211
0 213 7 2 2 1568 1573
0 214 5 1 1 1575
0 215 7 1 2 1558 194
0 216 5 1 1 215
0 217 7 2 2 1561 216
0 218 5 1 1 1577
0 219 7 1 2 214 1578
0 220 5 2 1 219
0 221 7 2 2 1562 1579
0 222 5 1 1 1581
0 223 7 1 2 1530 166
0 224 5 1 1 223
0 225 7 2 2 1533 224
0 226 5 1 1 1583
0 227 7 1 2 222 1584
0 228 5 2 1 227
0 229 7 2 2 1534 1585
0 230 5 1 1 1587
0 231 7 1 2 1495 120
0 232 5 1 1 231
0 233 7 2 2 1499 232
0 234 5 1 1 1589
0 235 7 1 2 230 1590
0 236 5 2 1 235
0 237 7 2 2 1257 1351
0 238 5 1 1 1593
0 239 7 2 2 1267 1342
0 240 5 1 1 1595
0 241 7 1 2 1594 1596
0 242 5 2 1 241
0 243 7 1 2 206 210
0 244 5 1 1 243
0 245 7 2 2 1574 244
0 246 5 1 1 1599
0 247 7 1 2 238 240
0 248 5 1 1 247
0 249 7 2 2 1597 248
0 250 5 1 1 1601
0 251 7 1 2 1600 1602
0 252 5 2 1 251
0 253 7 2 2 1598 1603
0 254 5 1 1 1605
0 255 7 1 2 1576 218
0 256 5 1 1 255
0 257 7 2 2 1580 256
0 258 5 1 1 1607
0 259 7 1 2 254 1608
0 260 5 2 1 259
0 261 7 2 2 1277 1325
0 262 5 1 1 1611
0 263 7 2 2 1249 1352
0 264 5 1 1 1613
0 265 7 1 2 1612 1614
0 266 5 2 1 265
0 267 7 2 2 1240 1360
0 268 5 1 1 1617
0 269 7 2 2 1268 1334
0 270 5 1 1 1619
0 271 7 1 2 1288 1316
0 272 5 1 1 271
0 273 7 1 2 1543 272
0 274 5 1 1 273
0 275 7 2 2 1548 274
0 276 5 1 1 1621
0 277 7 1 2 1620 1622
0 278 5 2 1 277
0 279 7 1 2 270 276
0 280 5 1 1 279
0 281 7 2 2 1623 280
0 282 5 1 1 1625
0 283 7 1 2 1618 1626
0 284 5 2 1 283
0 285 7 1 2 268 282
0 286 5 1 1 285
0 287 7 2 2 1627 286
0 288 5 1 1 1629
0 289 7 1 2 262 264
0 290 5 1 1 289
0 291 7 2 2 1615 290
0 292 5 1 1 1631
0 293 7 1 2 1630 1632
0 294 5 2 1 293
0 295 7 2 2 1616 1633
0 296 5 1 1 1635
0 297 7 1 2 246 250
0 298 5 1 1 297
0 299 7 2 2 1604 298
0 300 5 1 1 1637
0 301 7 1 2 296 1638
0 302 5 2 1 301
0 303 7 2 2 1296 1307
0 304 5 1 1 1641
0 305 7 2 2 1258 1343
0 306 5 1 1 1643
0 307 7 1 2 1642 1644
0 308 5 2 1 307
0 309 7 1 2 288 292
0 310 5 1 1 309
0 311 7 2 2 1634 310
0 312 5 1 1 1647
0 313 7 1 2 304 306
0 314 5 1 1 313
0 315 7 2 2 1645 314
0 316 5 1 1 1649
0 317 7 1 2 1648 1650
0 318 5 2 1 317
0 319 7 2 2 1646 1651
0 320 5 1 1 1653
0 321 7 1 2 1636 300
0 322 5 1 1 321
0 323 7 2 2 1639 322
0 324 5 1 1 1655
0 325 7 1 2 320 1656
0 326 5 2 1 325
0 327 7 2 2 1640 1657
0 328 5 1 1 1659
0 329 7 1 2 1606 258
0 330 5 1 1 329
0 331 7 2 2 1609 330
0 332 5 1 1 1661
0 333 7 1 2 328 1662
0 334 5 2 1 333
0 335 7 2 2 1610 1663
0 336 5 1 1 1665
0 337 7 1 2 1582 226
0 338 5 1 1 337
0 339 7 2 2 1586 338
0 340 5 1 1 1667
0 341 7 1 2 336 1668
0 342 5 2 1 341
0 343 7 2 2 1624 1628
0 344 5 1 1 1671
0 345 7 1 2 1654 324
0 346 5 1 1 345
0 347 7 2 2 1658 346
0 348 5 1 1 1673
0 349 7 1 2 344 1674
0 350 5 2 1 349
0 351 7 2 2 1278 1317
0 352 5 1 1 1677
0 353 7 2 2 1269 1326
0 354 5 1 1 1679
0 355 7 1 2 1678 1680
0 356 5 2 1 355
0 357 7 2 2 1241 1353
0 358 5 1 1 1683
0 359 7 1 2 352 354
0 360 5 1 1 359
0 361 7 2 2 1681 360
0 362 5 1 1 1685
0 363 7 1 2 1684 1686
0 364 5 2 1 363
0 365 7 2 2 1682 1687
0 366 5 1 1 1689
0 367 7 2 2 1250 1344
0 368 5 1 1 1691
0 369 7 2 2 32 1361
0 370 5 1 1 1693
0 371 7 1 2 1692 1694
0 372 5 2 1 371
0 373 7 2 2 1259 1335
0 374 5 1 1 1697
0 375 7 2 2 1270 1308
0 376 5 1 1 1699
0 377 7 2 2 1233 1327
0 378 5 1 1 1701
0 379 7 2 2 1251 1309
0 380 5 1 1 1703
0 381 7 2 2 1702 1704
0 382 5 2 1 1705
0 383 7 2 2 1260 1706
0 384 5 2 1 1709
0 385 7 2 2 1700 1710
0 386 5 2 1 1713
0 387 7 2 2 1279 1714
0 388 5 2 1 1717
0 389 7 1 2 1698 1718
0 390 5 2 1 389
0 391 7 1 2 374 1719
0 392 5 1 1 391
0 393 7 2 2 1721 392
0 394 5 1 1 1723
0 395 7 1 2 172 174
0 396 5 1 1 395
0 397 7 2 2 1544 396
0 398 5 1 1 1725
0 399 7 1 2 1724 1726
0 400 5 2 1 399
0 401 7 1 2 394 398
0 402 5 1 1 401
0 403 7 2 2 1727 402
0 404 5 1 1 1729
0 405 7 1 2 368 370
0 406 5 1 1 405
0 407 7 2 2 1695 406
0 408 5 1 1 1731
0 409 7 1 2 1730 1732
0 410 5 2 1 409
0 411 7 2 2 1696 1733
0 412 5 1 1 1735
0 413 7 1 2 366 412
0 414 5 2 1 413
0 415 7 2 2 1722 1728
0 416 5 1 1 1739
0 417 7 1 2 1690 1736
0 418 5 1 1 417
0 419 7 2 2 1737 418
0 420 5 1 1 1741
0 421 7 1 2 416 1742
0 422 5 2 1 421
0 423 7 2 2 1738 1743
0 424 5 1 1 1745
0 425 7 1 2 1672 348
0 426 5 1 1 425
0 427 7 2 2 1675 426
0 428 5 1 1 1747
0 429 7 1 2 424 1748
0 430 5 2 1 429
0 431 7 2 2 1676 1749
0 432 5 1 1 1751
0 433 7 1 2 1660 332
0 434 5 1 1 433
0 435 7 2 2 1664 434
0 436 5 1 1 1753
0 437 7 1 2 432 1754
0 438 5 2 1 437
0 439 7 1 2 312 316
0 440 5 1 1 439
0 441 7 2 2 1652 440
0 442 5 1 1 1757
0 443 7 1 2 1740 420
0 444 5 1 1 443
0 445 7 2 2 1744 444
0 446 5 1 1 1759
0 447 7 1 2 1758 1760
0 448 5 2 1 447
0 449 7 1 2 358 362
0 450 5 1 1 449
0 451 7 2 2 1688 450
0 452 5 1 1 1763
0 453 7 1 2 404 408
0 454 5 1 1 453
0 455 7 2 2 1734 454
0 456 5 1 1 1765
0 457 7 1 2 1764 1766
0 458 5 2 1 457
0 459 7 2 2 1261 1328
0 460 5 1 1 1769
0 461 7 2 2 1252 1336
0 462 5 1 1 1771
0 463 7 1 2 1770 1772
0 464 5 2 1 463
0 465 7 2 2 1242 1345
0 466 5 1 1 1775
0 467 7 1 2 460 462
0 468 5 1 1 467
0 469 7 2 2 1773 468
0 470 5 1 1 1777
0 471 7 1 2 1776 1778
0 472 5 2 1 471
0 473 7 2 2 1774 1779
0 474 5 1 1 1781
0 475 7 1 2 452 456
0 476 5 1 1 475
0 477 7 2 2 1767 476
0 478 5 1 1 1783
0 479 7 1 2 474 1784
0 480 5 2 1 479
0 481 7 2 2 1768 1785
0 482 5 1 1 1787
0 483 7 1 2 442 446
0 484 5 1 1 483
0 485 7 2 2 1761 484
0 486 5 1 1 1789
0 487 7 1 2 482 1790
0 488 5 2 1 487
0 489 7 2 2 1762 1791
0 490 5 1 1 1793
0 491 7 1 2 1746 428
0 492 5 1 1 491
0 493 7 2 2 1750 492
0 494 5 1 1 1795
0 495 7 1 2 490 1796
0 496 5 2 1 495
0 497 7 2 2 1234 1354
0 498 5 1 1 1799
0 499 7 1 2 466 470
0 500 5 1 1 499
0 501 7 2 2 1780 500
0 502 5 1 1 1801
0 503 7 1 2 1800 1802
0 504 5 2 1 503
0 505 7 2 2 1289 1299
0 506 5 1 1 1805
0 507 7 2 2 1271 1318
0 508 5 1 1 1807
0 509 7 1 2 1280 1310
0 510 5 1 1 509
0 511 7 1 2 1715 510
0 512 5 1 1 511
0 513 7 2 2 1720 512
0 514 5 1 1 1809
0 515 7 1 2 1808 1810
0 516 5 2 1 515
0 517 7 1 2 508 514
0 518 5 1 1 517
0 519 7 2 2 1811 518
0 520 5 1 1 1813
0 521 7 1 2 1806 1814
0 522 5 2 1 521
0 523 7 1 2 506 520
0 524 5 1 1 523
0 525 7 2 2 1815 524
0 526 5 1 1 1817
0 527 7 1 2 498 502
0 528 5 1 1 527
0 529 7 2 2 1803 528
0 530 5 1 1 1819
0 531 7 1 2 1818 1820
0 532 5 2 1 531
0 533 7 2 2 1804 1821
0 534 5 1 1 1823
0 535 7 1 2 1782 478
0 536 5 1 1 535
0 537 7 2 2 1786 536
0 538 5 1 1 1825
0 539 7 1 2 534 1826
0 540 5 2 1 539
0 541 7 2 2 1812 1816
0 542 5 1 1 1829
0 543 7 1 2 1824 538
0 544 5 1 1 543
0 545 7 2 2 1827 544
0 546 5 1 1 1831
0 547 7 1 2 542 1832
0 548 5 2 1 547
0 549 7 2 2 1828 1833
0 550 5 1 1 1835
0 551 7 1 2 1788 486
0 552 5 1 1 551
0 553 7 2 2 1792 552
0 554 5 1 1 1837
0 555 7 1 2 550 1838
0 556 5 2 1 555
0 557 7 2 2 1262 1319
0 558 5 1 1 1841
0 559 7 1 2 376 1711
0 560 5 1 1 559
0 561 7 2 2 1716 560
0 562 5 1 1 1843
0 563 7 1 2 1842 1844
0 564 5 2 1 563
0 565 7 2 2 1281 1300
0 566 5 1 1 1847
0 567 7 1 2 558 562
0 568 5 1 1 567
0 569 7 2 2 1845 568
0 570 5 1 1 1849
0 571 7 1 2 1848 1850
0 572 5 2 1 571
0 573 7 2 2 1846 1851
0 574 5 1 1 1853
0 575 7 1 2 526 530
0 576 5 1 1 575
0 577 7 2 2 1822 576
0 578 5 1 1 1855
0 579 7 1 2 574 1856
0 580 5 2 1 579
0 581 7 2 2 1253 1329
0 582 5 1 1 1859
0 583 7 2 2 1235 1346
0 584 5 1 1 1861
0 585 7 1 2 1860 1862
0 586 5 2 1 585
0 587 7 1 2 566 570
0 588 5 1 1 587
0 589 7 2 2 1852 588
0 590 5 1 1 1865
0 591 7 1 2 582 584
0 592 5 1 1 591
0 593 7 2 2 1863 592
0 594 5 1 1 1867
0 595 7 1 2 1866 1868
0 596 5 2 1 595
0 597 7 2 2 1864 1869
0 598 5 1 1 1871
0 599 7 1 2 1854 578
0 600 5 1 1 599
0 601 7 2 2 1857 600
0 602 5 1 1 1873
0 603 7 1 2 598 1874
0 604 5 2 1 603
0 605 7 2 2 1858 1875
0 606 5 1 1 1877
0 607 7 1 2 1830 546
0 608 5 1 1 607
0 609 7 2 2 1834 608
0 610 5 1 1 1879
0 611 7 1 2 606 1880
0 612 5 2 1 611
0 613 7 2 2 1243 1337
0 614 5 1 1 1883
0 615 7 1 2 590 594
0 616 5 1 1 615
0 617 7 2 2 1870 616
0 618 5 1 1 1885
0 619 7 1 2 1884 1886
0 620 5 2 1 619
0 621 7 2 2 1254 1320
0 622 5 1 1 1889
0 623 7 1 2 1263 1311
0 624 5 1 1 623
0 625 7 1 2 1707 624
0 626 5 1 1 625
0 627 7 2 2 1712 626
0 628 5 1 1 1891
0 629 7 1 2 1890 1892
0 630 5 2 1 629
0 631 7 2 2 1272 1301
0 632 5 1 1 1895
0 633 7 1 2 622 628
0 634 5 1 1 633
0 635 7 2 2 1893 634
0 636 5 1 1 1897
0 637 7 1 2 1896 1898
0 638 5 2 1 637
0 639 7 2 2 1894 1899
0 640 5 1 1 1901
0 641 7 1 2 614 618
0 642 5 1 1 641
0 643 7 2 2 1887 642
0 644 5 1 1 1903
0 645 7 1 2 640 1904
0 646 5 2 1 645
0 647 7 2 2 1888 1905
0 648 5 1 1 1907
0 649 7 1 2 1872 602
0 650 5 1 1 649
0 651 7 2 2 1876 650
0 652 5 1 1 1909
0 653 7 1 2 648 1910
0 654 5 2 1 653
0 655 7 2 2 1236 1338
0 656 5 1 1 1913
0 657 7 2 2 1244 1330
0 658 5 1 1 1915
0 659 7 1 2 1914 1916
0 660 5 2 1 659
0 661 7 1 2 632 636
0 662 5 1 1 661
0 663 7 2 2 1900 662
0 664 5 1 1 1919
0 665 7 1 2 656 658
0 666 5 1 1 665
0 667 7 2 2 1917 666
0 668 5 1 1 1921
0 669 7 1 2 1920 1922
0 670 5 2 1 669
0 671 7 2 2 1918 1923
0 672 5 1 1 1925
0 673 7 1 2 1902 644
0 674 5 1 1 673
0 675 7 2 2 1906 674
0 676 5 1 1 1927
0 677 7 1 2 672 1928
0 678 5 2 1 677
0 679 7 1 2 664 668
0 680 5 1 1 679
0 681 7 2 2 1924 680
0 682 5 1 1 1931
0 683 7 2 2 1245 1321
0 684 5 1 1 1933
0 685 7 2 2 1264 1302
0 686 5 1 1 1935
0 687 7 2 2 1934 1936
0 688 5 1 1 1937
0 689 7 2 2 1246 1312
0 690 5 1 1 1939
0 691 7 2 2 1237 1322
0 692 5 1 1 1941
0 693 7 2 2 1940 1942
0 694 5 2 1 1943
0 695 7 3 2 688 1945
0 696 5 1 1 1947
0 697 7 1 2 1932 696
0 698 5 2 1 697
0 699 7 1 2 378 380
0 700 5 1 1 699
0 701 7 2 2 1708 700
0 702 5 1 1 1952
0 703 7 1 2 684 686
0 704 5 1 1 703
0 705 7 1 2 1948 704
0 706 5 1 1 705
0 707 7 1 2 1938 1944
0 708 5 1 1 707
0 709 7 2 2 706 708
0 710 5 1 1 1954
0 711 7 1 2 1953 710
0 712 5 2 1 711
0 713 7 2 2 1255 1303
0 714 5 1 1 1958
0 715 7 1 2 690 692
0 716 5 1 1 715
0 717 7 2 2 1946 716
0 718 5 1 1 1960
0 719 7 1 2 1959 1961
0 720 5 2 1 719
0 721 7 1 2 714 718
0 722 5 1 1 721
0 723 7 2 2 1962 722
0 724 5 1 1 1964
0 725 7 2 2 1238 1313
0 726 5 1 1 1966
0 727 7 2 2 1247 1304
0 728 5 1 1 1968
0 729 7 2 2 1967 1969
0 730 5 2 1 1970
0 731 7 1 2 1965 1971
0 732 5 2 1 731
0 733 7 2 2 1963 1974
0 734 5 1 1 1976
0 735 7 1 2 702 1955
0 736 5 1 1 735
0 737 7 2 2 1956 736
0 738 5 1 1 1978
0 739 7 1 2 734 1979
0 740 5 2 1 739
0 741 7 2 2 1957 1980
0 742 5 1 1 1982
0 743 7 1 2 682 1949
0 744 5 1 1 743
0 745 7 2 2 1950 744
0 746 5 1 1 1984
0 747 7 1 2 742 1985
0 748 5 2 1 747
0 749 7 2 2 1951 1986
0 750 5 1 1 1988
0 751 7 1 2 1926 676
0 752 5 1 1 751
0 753 7 2 2 1929 752
0 754 5 1 1 1990
0 755 7 1 2 750 1991
0 756 5 2 1 755
0 757 7 2 2 1930 1992
0 758 5 1 1 1994
0 759 7 1 2 1908 652
0 760 5 1 1 759
0 761 7 2 2 1911 760
0 762 5 1 1 1996
0 763 7 1 2 758 1997
0 764 5 2 1 763
0 765 7 2 2 1912 1998
0 766 5 1 1 2000
0 767 7 1 2 1878 610
0 768 5 1 1 767
0 769 7 2 2 1881 768
0 770 5 1 1 2002
0 771 7 1 2 766 2003
0 772 5 2 1 771
0 773 7 2 2 1882 2004
0 774 5 1 1 2006
0 775 7 1 2 1836 554
0 776 5 1 1 775
0 777 7 2 2 1839 776
0 778 5 1 1 2008
0 779 7 1 2 774 2009
0 780 5 2 1 779
0 781 7 2 2 1840 2010
0 782 5 1 1 2012
0 783 7 1 2 1794 494
0 784 5 1 1 783
0 785 7 2 2 1797 784
0 786 5 1 1 2014
0 787 7 1 2 782 2015
0 788 5 2 1 787
0 789 7 2 2 1798 2016
0 790 5 1 1 2018
0 791 7 1 2 1752 436
0 792 5 1 1 791
0 793 7 2 2 1755 792
0 794 5 1 1 2020
0 795 7 1 2 790 2021
0 796 5 2 1 795
0 797 7 2 2 1756 2022
0 798 5 1 1 2024
0 799 7 1 2 1666 340
0 800 5 1 1 799
0 801 7 2 2 1669 800
0 802 5 1 1 2026
0 803 7 1 2 798 2027
0 804 5 2 1 803
0 805 7 2 2 1670 2028
0 806 5 1 1 2030
0 807 7 1 2 1588 234
0 808 5 1 1 807
0 809 7 2 2 1591 808
0 810 5 1 1 2032
0 811 7 1 2 806 2033
0 812 5 2 1 811
0 813 7 2 2 1592 2034
0 814 5 1 1 2036
0 815 7 1 2 1501 142
0 816 5 1 1 815
0 817 7 2 2 1515 816
0 818 5 1 1 2038
0 819 7 1 2 814 2039
0 820 5 2 1 819
0 821 7 2 2 1516 2040
0 822 5 1 1 2042
0 823 7 2 2 1297 1362
0 824 5 1 1 2044
0 825 7 1 2 1455 1511
0 826 5 1 1 825
0 827 7 1 2 2045 826
0 828 5 2 1 827
0 829 7 1 2 1512 824
0 830 5 1 1 829
0 831 7 2 2 2046 830
0 832 5 1 1 2048
0 833 7 1 2 822 2049
0 834 5 3 1 833
0 835 7 1 2 2043 832
0 836 5 2 1 835
0 837 7 2 2 2050 2053
0 838 5 2 1 2055
0 839 7 1 2 2037 818
0 840 5 1 1 839
0 841 7 2 2 2041 840
0 842 5 2 1 2059
0 843 7 1 2 1402 2061
0 844 5 2 1 843
0 845 7 1 2 1431 2060
0 846 5 2 1 845
0 847 7 1 2 2031 810
0 848 5 1 1 847
0 849 7 2 2 2035 848
0 850 5 2 1 2067
0 851 7 1 2 1399 2069
0 852 5 2 1 851
0 853 7 1 2 1429 2068
0 854 5 2 1 853
0 855 7 1 2 2025 802
0 856 5 1 1 855
0 857 7 2 2 2029 856
0 858 5 2 1 2075
0 859 7 1 2 1396 2077
0 860 5 2 1 859
0 861 7 1 2 1427 2076
0 862 5 2 1 861
0 863 7 1 2 2019 794
0 864 5 1 1 863
0 865 7 3 2 2023 864
0 866 5 1 1 2083
0 867 7 1 2 1393 866
0 868 5 2 1 867
0 869 7 1 2 1425 2084
0 870 5 2 1 869
0 871 7 1 2 2013 786
0 872 5 1 1 871
0 873 7 2 2 2017 872
0 874 5 2 1 2090
0 875 7 1 2 1390 2092
0 876 5 2 1 875
0 877 7 1 2 1423 2091
0 878 5 2 1 877
0 879 7 1 2 2007 778
0 880 5 1 1 879
0 881 7 3 2 2011 880
0 882 5 1 1 2098
0 883 7 1 2 1387 882
0 884 5 2 1 883
0 885 7 1 2 1421 2099
0 886 5 2 1 885
0 887 7 1 2 2001 770
0 888 5 1 1 887
0 889 7 2 2 2005 888
0 890 5 2 1 2105
0 891 7 1 2 1384 2107
0 892 5 2 1 891
0 893 7 1 2 1419 2106
0 894 5 2 1 893
0 895 7 1 2 1983 746
0 896 5 1 1 895
0 897 7 3 2 1987 896
0 898 5 1 1 2113
0 899 7 1 2 1375 898
0 900 5 2 1 899
0 901 7 1 2 1413 2114
0 902 5 2 1 901
0 903 7 1 2 1977 738
0 904 5 1 1 903
0 905 7 2 2 1981 904
0 906 5 2 1 2120
0 907 7 1 2 1372 2122
0 908 5 2 1 907
0 909 7 1 2 1411 2121
0 910 5 2 1 909
0 911 7 1 2 724 1972
0 912 5 1 1 911
0 913 7 3 2 1975 912
0 914 5 1 1 2128
0 915 7 1 2 1369 914
0 916 5 2 1 915
0 917 7 1 2 1409 2129
0 918 5 2 1 917
0 919 7 2 2 726 728
0 920 5 1 1 2135
0 921 7 3 2 1973 920
0 922 5 1 1 2137
0 923 7 1 2 1366 922
0 924 5 2 1 923
0 925 7 1 2 34 2138
0 926 5 2 1 925
0 927 7 2 2 1239 1305
0 928 5 1 1 2144
0 929 7 2 2 33 2145
0 930 5 2 1 2146
0 931 7 1 2 2142 2148
0 932 5 1 1 931
0 933 7 2 2 2140 932
0 934 5 2 1 2150
0 935 7 1 2 2133 2152
0 936 5 1 1 935
0 937 7 2 2 2131 936
0 938 5 2 1 2154
0 939 7 1 2 2126 2156
0 940 5 1 1 939
0 941 7 2 2 2124 940
0 942 5 2 1 2158
0 943 7 1 2 2118 2160
0 944 5 1 1 943
0 945 7 2 2 2116 944
0 946 5 1 1 2162
0 947 7 1 2 1415 2163
0 948 5 2 1 947
0 949 7 1 2 1378 946
0 950 5 2 1 949
0 951 7 1 2 1989 754
0 952 5 1 1 951
0 953 7 3 2 1993 952
0 954 5 2 1 2168
0 955 7 1 2 2166 2169
0 956 5 1 1 955
0 957 7 2 2 2164 956
0 958 5 1 1 2173
0 959 7 1 2 1417 958
0 960 5 2 1 959
0 961 7 1 2 1381 2174
0 962 5 2 1 961
0 963 7 1 2 1995 762
0 964 5 1 1 963
0 965 7 3 2 1999 964
0 966 5 1 1 2179
0 967 7 1 2 2177 2180
0 968 5 1 1 967
0 969 7 3 2 2175 968
0 970 5 1 1 2182
0 971 7 1 2 2111 2183
0 972 5 1 1 971
0 973 7 2 2 2109 972
0 974 5 2 1 2185
0 975 7 1 2 2103 2187
0 976 5 1 1 975
0 977 7 2 2 2101 976
0 978 5 2 1 2189
0 979 7 1 2 2096 2191
0 980 5 1 1 979
0 981 7 2 2 2094 980
0 982 5 2 1 2193
0 983 7 1 2 2088 2195
0 984 5 1 1 983
0 985 7 2 2 2086 984
0 986 5 2 1 2197
0 987 7 1 2 2081 2199
0 988 5 1 1 987
0 989 7 2 2 2079 988
0 990 5 2 1 2201
0 991 7 1 2 2073 2203
0 992 5 1 1 991
0 993 7 2 2 2071 992
0 994 5 2 1 2205
0 995 7 1 2 2065 2207
0 996 5 1 1 995
0 997 7 4 2 2063 996
0 998 7 1 2 1433 2209
0 999 5 1 1 998
0 1000 7 1 2 1435 999
0 1001 5 1 1 1000
0 1002 7 1 2 2057 1001
0 1003 5 1 1 1002
0 1004 7 2 2 1436 2054
0 1005 5 1 1 2213
0 1006 7 1 2 2051 2214
0 1007 5 1 1 1006
0 1008 7 1 2 2210 1007
0 1009 5 1 1 1008
0 1010 7 1 2 1405 1009
0 1011 5 1 1 1010
0 1012 7 1 2 1397 2198
0 1013 5 1 1 1012
0 1014 7 1 2 1428 2200
0 1015 5 1 1 1014
0 1016 7 2 2 1013 1015
0 1017 5 1 1 2215
0 1018 7 1 2 2078 2216
0 1019 5 1 1 1018
0 1020 7 1 2 1426 2194
0 1021 5 1 1 1020
0 1022 7 1 2 1394 2196
0 1023 5 1 1 1022
0 1024 7 2 2 1021 1023
0 1025 5 1 1 2217
0 1026 7 1 2 1391 2190
0 1027 5 1 1 1026
0 1028 7 1 2 1424 2192
0 1029 5 1 1 1028
0 1030 7 2 2 1027 1029
0 1031 5 1 1 2219
0 1032 7 1 2 1388 2186
0 1033 5 1 1 1032
0 1034 7 1 2 1422 2188
0 1035 5 1 1 1034
0 1036 7 2 2 1033 1035
0 1037 5 1 1 2221
0 1038 7 1 2 2100 2222
0 1039 5 1 1 1038
0 1040 7 1 2 1420 2184
0 1041 5 1 1 1040
0 1042 7 1 2 1385 970
0 1043 5 1 1 1042
0 1044 7 2 2 1041 1043
0 1045 5 1 1 2223
0 1046 7 2 2 2176 2178
0 1047 5 1 1 2225
0 1048 7 2 2 2165 2167
0 1049 5 1 1 2227
0 1050 7 1 2 2171 1049
0 1051 5 1 1 1050
0 1052 7 1 2 1376 2159
0 1053 5 1 1 1052
0 1054 7 1 2 1414 2161
0 1055 5 1 1 1054
0 1056 7 2 2 1053 1055
0 1057 5 1 1 2229
0 1058 7 1 2 1373 2155
0 1059 5 1 1 1058
0 1060 7 1 2 1412 2157
0 1061 5 1 1 1060
0 1062 7 2 2 1059 1061
0 1063 5 1 1 2231
0 1064 7 1 2 2123 2232
0 1065 5 1 1 1064
0 1066 7 1 2 1370 2151
0 1067 5 1 1 1066
0 1068 7 1 2 1410 2153
0 1069 5 1 1 1068
0 1070 7 2 2 1067 1069
0 1071 5 1 1 2233
0 1072 7 2 2 1364 928
0 1073 5 1 1 2235
0 1074 7 1 2 2139 1073
0 1075 5 2 1 1074
0 1076 7 2 2 2141 2143
0 1077 5 1 1 2239
0 1078 7 1 2 2147 2240
0 1079 5 1 1 1078
0 1080 7 1 2 2149 1077
0 1081 5 1 1 1080
0 1082 7 1 2 2136 2236
0 1083 5 2 1 1082
0 1084 7 1 2 1081 2241
0 1085 7 1 2 1079 1084
0 1086 5 1 1 1085
0 1087 7 1 2 2237 1086
0 1088 5 1 1 1087
0 1089 7 1 2 1071 1088
0 1090 5 1 1 1089
0 1091 7 1 2 2130 2234
0 1092 5 1 1 1091
0 1093 7 1 2 1090 1092
0 1094 7 1 2 1063 1093
0 1095 5 1 1 1094
0 1096 7 1 2 1065 1095
0 1097 7 1 2 1057 1096
0 1098 5 1 1 1097
0 1099 7 1 2 2115 2230
0 1100 5 1 1 1099
0 1101 7 1 2 1098 1100
0 1102 7 1 2 2228 1101
0 1103 5 1 1 1102
0 1104 7 1 2 1051 1103
0 1105 7 1 2 2226 1104
0 1106 5 1 1 1105
0 1107 7 1 2 2181 1047
0 1108 5 1 1 1107
0 1109 7 1 2 1106 1108
0 1110 7 1 2 1045 1109
0 1111 5 1 1 1110
0 1112 7 1 2 2108 2224
0 1113 5 1 1 1112
0 1114 7 1 2 1111 1113
0 1115 7 1 2 1037 1114
0 1116 5 1 1 1115
0 1117 7 1 2 1039 1116
0 1118 7 1 2 1031 1117
0 1119 5 1 1 1118
0 1120 7 1 2 2093 2220
0 1121 5 1 1 1120
0 1122 7 1 2 1119 1121
0 1123 7 1 2 2218 1122
0 1124 5 1 1 1123
0 1125 7 1 2 2085 1025
0 1126 5 1 1 1125
0 1127 7 1 2 1124 1126
0 1128 7 1 2 1017 1127
0 1129 5 1 1 1128
0 1130 7 1 2 1019 1129
0 1131 5 1 1 1130
0 1132 7 1 2 1400 2204
0 1133 5 1 1 1132
0 1134 7 1 2 1430 2202
0 1135 5 1 1 1134
0 1136 7 2 2 1133 1135
0 1137 5 1 1 2243
0 1138 7 1 2 1131 2244
0 1139 5 1 1 1138
0 1140 7 1 2 2070 1137
0 1141 5 1 1 1140
0 1142 7 1 2 1139 1141
0 1143 5 1 1 1142
0 1144 7 1 2 1403 2208
0 1145 5 1 1 1144
0 1146 7 1 2 1432 2206
0 1147 5 1 1 1146
0 1148 7 2 2 1145 1147
0 1149 5 1 1 2245
0 1150 7 1 2 1143 2246
0 1151 5 1 1 1150
0 1152 7 1 2 2062 1149
0 1153 5 1 1 1152
0 1154 7 1 2 1151 1153
0 1155 7 1 2 1011 1154
0 1156 7 1 2 1003 1155
0 1157 5 1 1 1156
0 1158 7 1 2 2056 2211
0 1159 5 1 1 1158
0 1160 7 1 2 1416 2170
0 1161 5 1 1 1160
0 1162 7 1 2 1379 2172
0 1163 5 1 1 1162
0 1164 7 1 2 1367 2238
0 1165 5 1 1 1164
0 1166 7 1 2 2242 1165
0 1167 7 1 2 2132 1166
0 1168 5 1 1 1167
0 1169 7 1 2 2134 1168
0 1170 7 1 2 2127 1169
0 1171 5 1 1 1170
0 1172 7 1 2 2125 1171
0 1173 7 1 2 2117 1172
0 1174 5 1 1 1173
0 1175 7 1 2 2119 1174
0 1176 5 1 1 1175
0 1177 7 1 2 1163 1176
0 1178 5 1 1 1177
0 1179 7 2 2 1161 1178
0 1180 5 1 1 2247
0 1181 7 1 2 1418 1180
0 1182 5 1 1 1181
0 1183 7 1 2 966 1182
0 1184 5 1 1 1183
0 1185 7 1 2 1382 2248
0 1186 5 1 1 1185
0 1187 7 1 2 2110 1186
0 1188 7 1 2 1184 1187
0 1189 5 1 1 1188
0 1190 7 1 2 2104 2112
0 1191 7 1 2 1189 1190
0 1192 5 1 1 1191
0 1193 7 1 2 2095 2102
0 1194 7 1 2 1192 1193
0 1195 5 1 1 1194
0 1196 7 1 2 2089 2097
0 1197 7 1 2 1195 1196
0 1198 5 1 1 1197
0 1199 7 1 2 2080 2087
0 1200 7 1 2 1198 1199
0 1201 5 1 1 1200
0 1202 7 1 2 2082 1201
0 1203 5 1 1 1202
0 1204 7 1 2 2072 1203
0 1205 5 1 1 1204
0 1206 7 1 2 2066 2074
0 1207 7 2 2 1205 1206
0 1208 5 1 1 2249
0 1209 7 1 2 1437 2064
0 1210 7 1 2 1208 1209
0 1211 5 1 1 1210
0 1212 7 1 2 1159 1211
0 1213 5 1 1 1212
0 1214 7 1 2 1434 1213
0 1215 5 1 1 1214
0 1216 7 2 2 2047 2052
0 1217 5 1 1 2251
0 1218 7 1 2 1005 2252
0 1219 5 1 1 1218
0 1220 7 1 2 2212 2250
0 1221 5 1 1 1220
0 1222 7 1 2 1219 1221
0 1223 5 1 1 1222
0 1224 7 1 2 1406 2058
0 1225 5 1 1 1224
0 1226 7 1 2 1408 1225
0 1227 5 1 1 1226
0 1228 7 1 2 1217 1227
0 1229 5 1 1 1228
0 1230 7 1 2 1223 1229
0 1231 7 1 2 1215 1230
0 1232 7 1 2 1157 1231
3 4299 5 0 1 1232
