1 0 0 2 0
2 49 1 0
2 715 1 0
1 1 0 2 0
2 716 1 1
2 717 1 1
1 2 0 2 0
2 718 1 2
2 719 1 2
1 3 0 2 0
2 720 1 3
2 721 1 3
1 4 0 2 0
2 722 1 4
2 723 1 4
1 5 0 2 0
2 724 1 5
2 725 1 5
1 6 0 2 0
2 726 1 6
2 727 1 6
1 7 0 2 0
2 728 1 7
2 729 1 7
1 8 0 2 0
2 730 1 8
2 731 1 8
1 9 0 2 0
2 732 1 9
2 733 1 9
1 10 0 2 0
2 734 1 10
2 735 1 10
1 11 0 2 0
2 736 1 11
2 737 1 11
1 12 0 2 0
2 738 1 12
2 739 1 12
1 13 0 2 0
2 740 1 13
2 741 1 13
1 14 0 2 0
2 742 1 14
2 743 1 14
1 15 0 2 0
2 744 1 15
2 745 1 15
1 16 0 2 0
2 746 1 16
2 747 1 16
1 17 0 2 0
2 748 1 17
2 749 1 17
1 18 0 2 0
2 750 1 18
2 751 1 18
1 19 0 2 0
2 752 1 19
2 753 1 19
1 20 0 2 0
2 754 1 20
2 755 1 20
1 21 0 2 0
2 756 1 21
2 757 1 21
1 22 0 2 0
2 758 1 22
2 759 1 22
1 23 0 2 0
2 760 1 23
2 761 1 23
1 24 0 2 0
2 762 1 24
2 763 1 24
1 25 0 2 0
2 764 1 25
2 765 1 25
1 26 0 2 0
2 766 1 26
2 767 1 26
1 27 0 2 0
2 768 1 27
2 769 1 27
1 28 0 2 0
2 770 1 28
2 771 1 28
1 29 0 2 0
2 772 1 29
2 773 1 29
1 30 0 2 0
2 774 1 30
2 775 1 30
1 31 0 2 0
2 776 1 31
2 777 1 31
1 32 0 2 0
2 778 1 32
2 779 1 32
1 33 0 3 0
2 780 1 33
2 781 1 33
2 782 1 33
1 34 0 2 0
2 783 1 34
2 784 1 34
1 35 0 2 0
2 785 1 35
2 786 1 35
1 36 0 2 0
2 787 1 36
2 788 1 36
1 37 0 2 0
2 789 1 37
2 790 1 37
1 38 0 2 0
2 791 1 38
2 792 1 38
1 39 0 2 0
2 793 1 39
2 794 1 39
1 40 0 2 0
2 795 1 40
2 796 1 40
1 41 0 2 0
2 797 1 41
2 798 1 41
1 42 0 2 0
2 799 1 42
2 800 1 42
1 43 0 2 0
2 801 1 43
2 802 1 43
1 44 0 2 0
2 803 1 44
2 804 1 44
1 45 0 2 0
2 805 1 45
2 806 1 45
1 46 0 2 0
2 807 1 46
2 808 1 46
1 47 0 2 0
2 809 1 47
2 810 1 47
1 48 0 2 0
2 811 1 48
2 812 1 48
2 813 1 69
2 814 1 69
2 815 1 70
2 816 1 70
2 817 1 71
2 818 1 71
2 819 1 72
2 820 1 72
2 821 1 73
2 822 1 73
2 823 1 74
2 824 1 74
2 825 1 75
2 826 1 75
2 827 1 76
2 828 1 76
2 829 1 77
2 830 1 77
2 831 1 78
2 832 1 78
2 833 1 79
2 834 1 79
2 835 1 80
2 836 1 80
2 837 1 100
2 838 1 100
2 839 1 102
2 840 1 102
2 841 1 104
2 842 1 104
2 843 1 106
2 844 1 106
2 845 1 108
2 846 1 108
2 847 1 110
2 848 1 110
2 849 1 111
2 850 1 111
2 851 1 112
2 852 1 112
2 853 1 112
2 854 1 115
2 855 1 115
2 856 1 116
2 857 1 116
2 858 1 119
2 859 1 119
2 860 1 122
2 861 1 122
2 862 1 124
2 863 1 124
2 864 1 127
2 865 1 127
2 866 1 130
2 867 1 130
2 868 1 132
2 869 1 132
2 870 1 135
2 871 1 135
2 872 1 138
2 873 1 138
2 874 1 140
2 875 1 140
2 876 1 143
2 877 1 143
2 878 1 146
2 879 1 146
2 880 1 148
2 881 1 148
2 882 1 151
2 883 1 151
2 884 1 154
2 885 1 154
2 886 1 156
2 887 1 156
2 888 1 159
2 889 1 159
2 890 1 162
2 891 1 162
2 892 1 164
2 893 1 164
2 894 1 167
2 895 1 167
2 896 1 170
2 897 1 170
2 898 1 172
2 899 1 172
2 900 1 175
2 901 1 175
2 902 1 178
2 903 1 178
2 904 1 180
2 905 1 180
2 906 1 183
2 907 1 183
2 908 1 186
2 909 1 186
2 910 1 188
2 911 1 188
2 912 1 191
2 913 1 191
2 914 1 194
2 915 1 194
2 916 1 196
2 917 1 196
2 918 1 199
2 919 1 199
2 920 1 202
2 921 1 202
2 922 1 204
2 923 1 204
2 924 1 207
2 925 1 207
2 926 1 210
2 927 1 210
2 928 1 212
2 929 1 212
2 930 1 215
2 931 1 215
2 932 1 216
2 933 1 216
2 934 1 219
2 935 1 219
2 936 1 221
2 937 1 221
2 938 1 222
2 939 1 222
2 940 1 223
2 941 1 223
2 942 1 223
2 943 1 224
2 944 1 224
2 945 1 225
2 946 1 225
2 947 1 231
2 948 1 231
2 949 1 233
2 950 1 233
2 951 1 234
2 952 1 234
2 953 1 236
2 954 1 236
2 955 1 236
2 956 1 237
2 957 1 237
2 958 1 243
2 959 1 243
2 960 1 246
2 961 1 246
2 962 1 246
2 963 1 247
2 964 1 247
2 965 1 253
2 966 1 253
2 967 1 256
2 968 1 256
2 969 1 256
2 970 1 258
2 971 1 258
2 972 1 258
2 973 1 258
2 974 1 259
2 975 1 259
2 976 1 265
2 977 1 265
2 978 1 268
2 979 1 268
2 980 1 268
2 981 1 270
2 982 1 270
2 983 1 270
2 984 1 270
2 985 1 271
2 986 1 271
2 987 1 277
2 988 1 277
2 989 1 280
2 990 1 280
2 991 1 280
2 992 1 280
2 993 1 282
2 994 1 282
2 995 1 282
2 996 1 282
2 997 1 283
2 998 1 283
2 999 1 289
2 1000 1 289
2 1001 1 291
2 1002 1 291
2 1003 1 291
2 1004 1 292
2 1005 1 292
2 1006 1 293
2 1007 1 293
2 1008 1 293
2 1009 1 294
2 1010 1 294
2 1011 1 295
2 1012 1 295
2 1013 1 301
2 1014 1 301
2 1015 1 304
2 1016 1 304
2 1017 1 304
2 1018 1 306
2 1019 1 306
2 1020 1 306
2 1021 1 307
2 1022 1 307
2 1023 1 313
2 1024 1 313
2 1025 1 316
2 1026 1 316
2 1027 1 316
2 1028 1 316
2 1029 1 317
2 1030 1 317
2 1031 1 323
2 1032 1 323
2 1033 1 326
2 1034 1 326
2 1035 1 326
2 1036 1 326
2 1037 1 328
2 1038 1 328
2 1039 1 328
2 1040 1 329
2 1041 1 329
2 1042 1 335
2 1043 1 335
2 1044 1 338
2 1045 1 338
2 1046 1 338
2 1047 1 338
2 1048 1 339
2 1049 1 339
2 1050 1 345
2 1051 1 345
2 1052 1 348
2 1053 1 348
2 1054 1 348
2 1055 1 348
2 1056 1 350
2 1057 1 350
2 1058 1 350
2 1059 1 351
2 1060 1 351
2 1061 1 357
2 1062 1 357
2 1063 1 360
2 1064 1 360
2 1065 1 360
2 1066 1 361
2 1067 1 361
2 1068 1 367
2 1069 1 367
2 1070 1 370
2 1071 1 370
2 1072 1 370
2 1073 1 372
2 1074 1 372
2 1075 1 372
2 1076 1 373
2 1077 1 373
2 1078 1 379
2 1079 1 379
2 1080 1 382
2 1081 1 382
2 1082 1 383
2 1083 1 383
2 1084 1 384
2 1085 1 384
2 1086 1 389
2 1087 1 389
2 1088 1 394
2 1089 1 394
2 1090 1 397
2 1091 1 397
2 1092 1 407
2 1093 1 407
2 1094 1 408
2 1095 1 408
2 1096 1 409
2 1097 1 409
2 1098 1 412
2 1099 1 412
2 1100 1 413
2 1101 1 413
2 1102 1 415
2 1103 1 415
2 1104 1 415
2 1105 1 418
2 1106 1 418
2 1107 1 419
2 1108 1 419
2 1109 1 422
2 1110 1 422
2 1111 1 423
2 1112 1 423
2 1113 1 425
2 1114 1 425
2 1115 1 425
2 1116 1 428
2 1117 1 428
2 1118 1 429
2 1119 1 429
2 1120 1 432
2 1121 1 432
2 1122 1 435
2 1123 1 435
2 1124 1 435
2 1125 1 436
2 1126 1 436
2 1127 1 438
2 1128 1 438
2 1129 1 439
2 1130 1 439
2 1131 1 442
2 1132 1 442
2 1133 1 442
2 1134 1 450
2 1135 1 450
2 1136 1 453
2 1137 1 453
2 1138 1 454
2 1139 1 454
2 1140 1 457
2 1141 1 457
2 1142 1 458
2 1143 1 458
2 1144 1 460
2 1145 1 460
2 1146 1 460
2 1147 1 463
2 1148 1 463
2 1149 1 463
2 1150 1 468
2 1151 1 468
2 1152 1 471
2 1153 1 471
2 1154 1 475
2 1155 1 475
2 1156 1 476
2 1157 1 476
2 1158 1 483
2 1159 1 483
2 1160 1 483
2 1161 1 484
2 1162 1 484
2 1163 1 489
2 1164 1 489
2 1165 1 490
2 1166 1 490
2 1167 1 497
2 1168 1 497
2 1169 1 498
2 1170 1 498
2 1171 1 504
2 1172 1 504
2 1173 1 511
2 1174 1 511
2 1175 1 511
2 1176 1 512
2 1177 1 512
2 1178 1 519
2 1179 1 519
2 1180 1 520
2 1181 1 520
2 1182 1 525
2 1183 1 525
2 1184 1 526
2 1185 1 526
2 1186 1 531
2 1187 1 531
2 1188 1 531
2 1189 1 537
2 1190 1 537
2 1191 1 538
2 1192 1 538
2 1193 1 545
2 1194 1 545
2 1195 1 545
2 1196 1 546
2 1197 1 546
2 1198 1 551
2 1199 1 551
2 1200 1 551
2 1201 1 552
2 1202 1 552
2 1203 1 591
2 1204 1 591
2 1205 1 591
2 1206 1 595
2 1207 1 595
2 1208 1 595
2 1209 1 599
2 1210 1 599
2 1211 1 602
2 1212 1 602
2 1213 1 610
2 1214 1 610
2 1215 1 613
2 1216 1 613
2 1217 1 614
2 1218 1 614
2 1219 1 617
2 1220 1 617
2 1221 1 618
2 1222 1 618
2 1223 1 630
2 1224 1 630
2 1225 1 632
2 1226 1 632
2 1227 1 633
2 1228 1 633
2 1229 1 642
2 1230 1 642
2 1231 1 702
2 1232 1 702
0 50 5 1 1 49
0 51 5 1 1 716
0 52 5 1 1 718
0 53 5 1 1 720
0 54 5 1 1 722
0 55 5 1 1 724
0 56 5 1 1 726
0 57 5 1 1 728
0 58 5 1 1 730
0 59 5 1 1 732
0 60 5 1 1 734
0 61 5 1 1 736
0 62 5 1 1 738
0 63 5 1 1 740
0 64 5 1 1 742
0 65 5 1 1 744
0 66 5 1 1 746
0 67 5 1 1 748
0 68 5 1 1 750
0 69 5 2 1 752
0 70 5 2 1 754
0 71 5 2 1 756
0 72 5 2 1 758
0 73 5 2 1 760
0 74 5 2 1 762
0 75 5 2 1 764
0 76 5 2 1 766
0 77 5 2 1 768
0 78 5 2 1 770
0 79 5 2 1 772
0 80 5 2 1 774
0 81 5 1 1 776
0 82 5 1 1 778
0 83 5 1 1 780
0 84 5 1 1 783
0 85 5 1 1 785
0 86 5 1 1 787
0 87 5 1 1 789
0 88 5 1 1 791
0 89 5 1 1 793
0 90 5 1 1 795
0 91 5 1 1 797
0 92 5 1 1 799
0 93 5 1 1 801
0 94 5 1 1 803
0 95 5 1 1 805
0 96 5 1 1 807
0 97 5 1 1 809
0 98 5 1 1 811
0 99 7 1 2 65 81
0 100 5 2 1 99
0 101 7 1 2 745 777
0 102 5 2 1 101
0 103 7 1 2 52 68
0 104 5 2 1 103
0 105 7 1 2 719 751
0 106 5 2 1 105
0 107 7 1 2 51 67
0 108 5 2 1 107
0 109 7 1 2 717 749
0 110 5 2 1 109
0 111 7 2 2 715 747
0 112 5 3 1 849
0 113 7 1 2 847 851
0 114 5 1 1 113
0 115 7 2 2 845 114
0 116 5 2 1 854
0 117 7 1 2 843 856
0 118 5 1 1 117
0 119 7 2 2 841 118
0 120 5 1 1 858
0 121 7 1 2 53 120
0 122 5 2 1 121
0 123 7 1 2 721 859
0 124 5 2 1 123
0 125 7 1 2 813 862
0 126 5 1 1 125
0 127 7 2 2 860 126
0 128 5 1 1 864
0 129 7 1 2 54 128
0 130 5 2 1 129
0 131 7 1 2 723 865
0 132 5 2 1 131
0 133 7 1 2 815 868
0 134 5 1 1 133
0 135 7 2 2 866 134
0 136 5 1 1 870
0 137 7 1 2 55 136
0 138 5 2 1 137
0 139 7 1 2 725 871
0 140 5 2 1 139
0 141 7 1 2 817 874
0 142 5 1 1 141
0 143 7 2 2 872 142
0 144 5 1 1 876
0 145 7 1 2 56 144
0 146 5 2 1 145
0 147 7 1 2 727 877
0 148 5 2 1 147
0 149 7 1 2 819 880
0 150 5 1 1 149
0 151 7 2 2 878 150
0 152 5 1 1 882
0 153 7 1 2 57 152
0 154 5 2 1 153
0 155 7 1 2 729 883
0 156 5 2 1 155
0 157 7 1 2 821 886
0 158 5 1 1 157
0 159 7 2 2 884 158
0 160 5 1 1 888
0 161 7 1 2 58 160
0 162 5 2 1 161
0 163 7 1 2 731 889
0 164 5 2 1 163
0 165 7 1 2 823 892
0 166 5 1 1 165
0 167 7 2 2 890 166
0 168 5 1 1 894
0 169 7 1 2 59 168
0 170 5 2 1 169
0 171 7 1 2 733 895
0 172 5 2 1 171
0 173 7 1 2 825 898
0 174 5 1 1 173
0 175 7 2 2 896 174
0 176 5 1 1 900
0 177 7 1 2 60 176
0 178 5 2 1 177
0 179 7 1 2 735 901
0 180 5 2 1 179
0 181 7 1 2 827 904
0 182 5 1 1 181
0 183 7 2 2 902 182
0 184 5 1 1 906
0 185 7 1 2 61 184
0 186 5 2 1 185
0 187 7 1 2 737 907
0 188 5 2 1 187
0 189 7 1 2 829 910
0 190 5 1 1 189
0 191 7 2 2 908 190
0 192 5 1 1 912
0 193 7 1 2 62 192
0 194 5 2 1 193
0 195 7 1 2 739 913
0 196 5 2 1 195
0 197 7 1 2 831 916
0 198 5 1 1 197
0 199 7 2 2 914 198
0 200 5 1 1 918
0 201 7 1 2 63 200
0 202 5 2 1 201
0 203 7 1 2 741 919
0 204 5 2 1 203
0 205 7 1 2 833 922
0 206 5 1 1 205
0 207 7 2 2 920 206
0 208 5 1 1 924
0 209 7 1 2 64 208
0 210 5 2 1 209
0 211 7 1 2 743 925
0 212 5 2 1 211
0 213 7 1 2 835 928
0 214 5 1 1 213
0 215 7 2 2 926 214
0 216 5 2 1 930
0 217 7 1 2 839 932
0 218 5 1 1 217
0 219 7 2 2 837 218
0 220 5 1 1 934
0 221 7 2 2 98 935
0 222 5 2 1 936
0 223 7 3 2 812 220
0 224 5 2 1 940
0 225 7 2 2 838 840
0 226 5 1 1 945
0 227 7 1 2 931 226
0 228 5 1 1 227
0 229 7 1 2 933 946
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 947
0 233 7 2 2 97 232
0 234 5 2 1 949
0 235 7 1 2 810 948
0 236 5 3 1 235
0 237 7 2 2 927 929
0 238 5 1 1 956
0 239 7 1 2 775 957
0 240 5 1 1 239
0 241 7 1 2 836 238
0 242 5 1 1 241
0 243 7 2 2 240 242
0 244 5 1 1 958
0 245 7 1 2 808 244
0 246 5 3 1 245
0 247 7 2 2 921 923
0 248 5 1 1 963
0 249 7 1 2 773 964
0 250 5 1 1 249
0 251 7 1 2 834 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 965
0 255 7 1 2 806 254
0 256 5 3 1 255
0 257 7 1 2 95 966
0 258 5 4 1 257
0 259 7 2 2 915 917
0 260 5 1 1 974
0 261 7 1 2 771 975
0 262 5 1 1 261
0 263 7 1 2 832 260
0 264 5 1 1 263
0 265 7 2 2 262 264
0 266 5 1 1 976
0 267 7 1 2 804 266
0 268 5 3 1 267
0 269 7 1 2 94 977
0 270 5 4 1 269
0 271 7 2 2 909 911
0 272 5 1 1 985
0 273 7 1 2 769 986
0 274 5 1 1 273
0 275 7 1 2 830 272
0 276 5 1 1 275
0 277 7 2 2 274 276
0 278 5 1 1 987
0 279 7 1 2 802 278
0 280 5 4 1 279
0 281 7 1 2 93 988
0 282 5 4 1 281
0 283 7 2 2 903 905
0 284 5 1 1 997
0 285 7 1 2 767 998
0 286 5 1 1 285
0 287 7 1 2 828 284
0 288 5 1 1 287
0 289 7 2 2 286 288
0 290 5 1 1 999
0 291 7 3 2 92 1000
0 292 5 2 1 1001
0 293 7 3 2 800 290
0 294 5 2 1 1006
0 295 7 2 2 897 899
0 296 5 1 1 1011
0 297 7 1 2 765 1012
0 298 5 1 1 297
0 299 7 1 2 826 296
0 300 5 1 1 299
0 301 7 2 2 298 300
0 302 5 1 1 1013
0 303 7 1 2 798 302
0 304 5 3 1 303
0 305 7 1 2 91 1014
0 306 5 3 1 305
0 307 7 2 2 891 893
0 308 5 1 1 1021
0 309 7 1 2 763 1022
0 310 5 1 1 309
0 311 7 1 2 824 308
0 312 5 1 1 311
0 313 7 2 2 310 312
0 314 5 1 1 1023
0 315 7 1 2 796 314
0 316 5 4 1 315
0 317 7 2 2 885 887
0 318 5 1 1 1029
0 319 7 1 2 761 1030
0 320 5 1 1 319
0 321 7 1 2 822 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1031
0 325 7 1 2 794 324
0 326 5 4 1 325
0 327 7 1 2 89 1032
0 328 5 3 1 327
0 329 7 2 2 879 881
0 330 5 1 1 1040
0 331 7 1 2 759 1041
0 332 5 1 1 331
0 333 7 1 2 820 330
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 1042
0 337 7 1 2 792 336
0 338 5 4 1 337
0 339 7 2 2 873 875
0 340 5 1 1 1048
0 341 7 1 2 757 1049
0 342 5 1 1 341
0 343 7 1 2 818 340
0 344 5 1 1 343
0 345 7 2 2 342 344
0 346 5 1 1 1050
0 347 7 1 2 790 346
0 348 5 4 1 347
0 349 7 1 2 87 1051
0 350 5 3 1 349
0 351 7 2 2 867 869
0 352 5 1 1 1059
0 353 7 1 2 755 1060
0 354 5 1 1 353
0 355 7 1 2 816 352
0 356 5 1 1 355
0 357 7 2 2 354 356
0 358 5 1 1 1061
0 359 7 1 2 788 358
0 360 5 3 1 359
0 361 7 2 2 861 863
0 362 5 1 1 1066
0 363 7 1 2 753 1067
0 364 5 1 1 363
0 365 7 1 2 814 362
0 366 5 1 1 365
0 367 7 2 2 364 366
0 368 5 1 1 1068
0 369 7 1 2 786 368
0 370 5 3 1 369
0 371 7 1 2 85 1069
0 372 5 3 1 371
0 373 7 2 2 842 844
0 374 5 1 1 1076
0 375 7 1 2 855 374
0 376 5 1 1 375
0 377 7 1 2 857 1077
0 378 5 1 1 377
0 379 7 2 2 376 378
0 380 5 1 1 1078
0 381 7 1 2 84 380
0 382 5 2 1 381
0 383 7 2 2 846 848
0 384 5 2 1 1082
0 385 7 1 2 850 1084
0 386 5 1 1 385
0 387 7 1 2 852 1083
0 388 5 1 1 387
0 389 7 2 2 386 388
0 390 5 1 1 1086
0 391 7 1 2 781 1087
0 392 5 1 1 391
0 393 7 1 2 83 390
0 394 5 2 1 393
0 395 7 1 2 50 66
0 396 5 1 1 395
0 397 7 2 2 853 396
0 398 5 1 1 1090
0 399 7 1 2 779 398
0 400 7 1 2 1088 399
0 401 5 1 1 400
0 402 7 1 2 392 401
0 403 5 1 1 402
0 404 7 1 2 1080 403
0 405 5 1 1 404
0 406 7 1 2 784 1079
0 407 5 2 1 406
0 408 7 2 2 405 1092
0 409 5 2 1 1094
0 410 7 1 2 1073 1096
0 411 5 1 1 410
0 412 7 2 2 1070 411
0 413 5 2 1 1098
0 414 7 1 2 86 1062
0 415 5 3 1 414
0 416 7 1 2 1100 1102
0 417 5 1 1 416
0 418 7 2 2 1063 417
0 419 5 2 1 1105
0 420 7 1 2 1056 1107
0 421 5 1 1 420
0 422 7 2 2 1052 421
0 423 5 2 1 1109
0 424 7 1 2 88 1043
0 425 5 3 1 424
0 426 7 1 2 1111 1113
0 427 5 1 1 426
0 428 7 2 2 1044 427
0 429 5 2 1 1116
0 430 7 1 2 1037 1118
0 431 5 1 1 430
0 432 7 2 2 1033 431
0 433 5 1 1 1120
0 434 7 1 2 90 1024
0 435 5 3 1 434
0 436 7 2 2 433 1122
0 437 5 1 1 1125
0 438 7 2 2 1025 437
0 439 5 2 1 1127
0 440 7 1 2 1018 1129
0 441 5 1 1 440
0 442 7 3 2 1015 441
0 443 5 1 1 1131
0 444 7 1 2 1009 1132
0 445 5 1 1 444
0 446 7 1 2 1004 445
0 447 7 1 2 993 446
0 448 5 1 1 447
0 449 7 1 2 989 448
0 450 5 2 1 449
0 451 7 1 2 981 1134
0 452 5 1 1 451
0 453 7 2 2 978 452
0 454 5 2 1 1136
0 455 7 1 2 970 1138
0 456 5 1 1 455
0 457 7 2 2 967 456
0 458 5 2 1 1140
0 459 7 1 2 96 959
0 460 5 3 1 459
0 461 7 1 2 1142 1144
0 462 5 1 1 461
0 463 7 3 2 960 462
0 464 5 1 1 1147
0 465 7 1 2 953 1148
0 466 5 1 1 465
0 467 7 1 2 951 466
0 468 5 2 1 467
0 469 7 1 2 943 1150
0 470 5 1 1 469
0 471 7 2 2 938 470
0 472 5 1 1 1152
0 473 7 1 2 937 1151
0 474 5 1 1 473
0 475 7 2 2 952 954
0 476 5 2 1 1154
0 477 7 1 2 464 1156
0 478 5 1 1 477
0 479 7 1 2 1149 1155
0 480 5 1 1 479
0 481 7 1 2 478 480
0 482 5 1 1 481
0 483 7 3 2 961 1145
0 484 5 2 1 1158
0 485 7 1 2 1143 1159
0 486 5 1 1 485
0 487 7 1 2 1141 1161
0 488 5 1 1 487
0 489 7 2 2 968 971
0 490 5 2 1 1163
0 491 7 1 2 1139 1165
0 492 5 1 1 491
0 493 7 1 2 1137 1164
0 494 5 1 1 493
0 495 7 1 2 492 494
0 496 5 1 1 495
0 497 7 2 2 979 982
0 498 5 2 1 1167
0 499 7 1 2 1135 1168
0 500 5 1 1 499
0 501 7 1 2 990 1169
0 502 5 1 1 501
0 503 7 1 2 991 994
0 504 5 2 1 503
0 505 7 1 2 1007 443
0 506 5 1 1 505
0 507 7 1 2 1171 506
0 508 5 1 1 507
0 509 7 1 2 1002 1133
0 510 5 1 1 509
0 511 7 3 2 1016 1019
0 512 5 2 1 1173
0 513 7 1 2 1128 1174
0 514 5 1 1 513
0 515 7 1 2 1130 1176
0 516 5 1 1 515
0 517 7 1 2 1026 1126
0 518 5 1 1 517
0 519 7 2 2 1027 1123
0 520 5 2 1 1178
0 521 7 1 2 1121 1180
0 522 5 1 1 521
0 523 7 1 2 518 522
0 524 5 1 1 523
0 525 7 2 2 1034 1038
0 526 5 2 1 1182
0 527 7 1 2 1119 1184
0 528 5 1 1 527
0 529 7 1 2 1117 1183
0 530 5 1 1 529
0 531 7 3 2 1045 1114
0 532 5 1 1 1186
0 533 7 1 2 1112 532
0 534 5 1 1 533
0 535 7 1 2 1110 1187
0 536 5 1 1 535
0 537 7 2 2 1053 1057
0 538 5 2 1 1189
0 539 7 1 2 1106 1191
0 540 5 1 1 539
0 541 7 1 2 1108 1190
0 542 5 1 1 541
0 543 7 1 2 540 542
0 544 5 1 1 543
0 545 7 3 2 1064 1103
0 546 5 2 1 1193
0 547 7 1 2 1099 1196
0 548 5 1 1 547
0 549 7 1 2 1101 1194
0 550 5 1 1 549
0 551 7 3 2 1071 1074
0 552 5 2 1 1198
0 553 7 1 2 1095 1201
0 554 5 1 1 553
0 555 7 1 2 1097 1199
0 556 5 1 1 555
0 557 7 1 2 554 556
0 558 7 1 2 550 557
0 559 7 1 2 548 558
0 560 5 1 1 559
0 561 7 1 2 544 560
0 562 7 1 2 536 561
0 563 7 1 2 534 562
0 564 7 1 2 530 563
0 565 7 1 2 528 564
0 566 7 1 2 524 565
0 567 7 1 2 516 566
0 568 7 1 2 514 567
0 569 5 1 1 568
0 570 7 1 2 510 569
0 571 7 1 2 508 570
0 572 7 1 2 502 571
0 573 7 1 2 500 572
0 574 7 1 2 496 573
0 575 7 1 2 944 574
0 576 7 1 2 488 575
0 577 7 1 2 486 576
0 578 7 1 2 482 577
0 579 7 1 2 474 578
0 580 7 1 2 472 579
0 581 5 1 1 580
0 582 7 1 2 782 1085
0 583 5 1 1 582
0 584 7 1 2 82 1091
0 585 7 1 2 583 584
0 586 5 1 1 585
0 587 7 1 2 1089 586
0 588 5 1 1 587
0 589 7 1 2 1093 588
0 590 5 1 1 589
0 591 7 3 2 1081 590
0 592 5 1 1 1203
0 593 7 1 2 1075 1204
0 594 5 1 1 593
0 595 7 3 2 1072 594
0 596 5 1 1 1206
0 597 7 1 2 1065 1207
0 598 5 1 1 597
0 599 7 2 2 1104 598
0 600 5 1 1 1209
0 601 7 1 2 1058 1210
0 602 5 2 1 601
0 603 7 1 2 1054 1211
0 604 7 1 2 1046 603
0 605 5 1 1 604
0 606 7 1 2 1115 605
0 607 7 1 2 1039 606
0 608 5 1 1 607
0 609 7 1 2 1035 608
0 610 5 2 1 609
0 611 7 1 2 1124 1213
0 612 5 1 1 611
0 613 7 2 2 1028 612
0 614 5 2 1 1215
0 615 7 1 2 1020 1217
0 616 5 1 1 615
0 617 7 2 2 1017 616
0 618 5 2 1 1219
0 619 7 1 2 1005 1221
0 620 5 1 1 619
0 621 7 1 2 1010 620
0 622 7 1 2 992 621
0 623 5 1 1 622
0 624 7 1 2 995 623
0 625 5 1 1 624
0 626 7 1 2 980 625
0 627 5 1 1 626
0 628 7 1 2 983 627
0 629 5 1 1 628
0 630 7 2 2 969 629
0 631 5 1 1 1223
0 632 7 2 2 972 631
0 633 5 2 1 1225
0 634 7 1 2 1162 1227
0 635 5 1 1 634
0 636 7 1 2 1160 1226
0 637 5 1 1 636
0 638 7 1 2 635 637
0 639 5 1 1 638
0 640 7 1 2 962 1228
0 641 5 1 1 640
0 642 7 2 2 1146 641
0 643 5 1 1 1229
0 644 7 1 2 1157 1230
0 645 5 1 1 644
0 646 7 1 2 973 1224
0 647 5 1 1 646
0 648 7 1 2 984 1166
0 649 5 1 1 648
0 650 7 1 2 996 1170
0 651 5 1 1 650
0 652 7 1 2 1003 1220
0 653 5 1 1 652
0 654 7 1 2 1172 653
0 655 5 1 1 654
0 656 7 1 2 1008 1222
0 657 5 1 1 656
0 658 7 1 2 1177 1216
0 659 5 1 1 658
0 660 7 1 2 1175 1218
0 661 5 1 1 660
0 662 7 1 2 1036 1181
0 663 5 1 1 662
0 664 7 1 2 1179 1214
0 665 5 1 1 664
0 666 7 1 2 1047 1185
0 667 5 1 1 666
0 668 7 1 2 1188 1212
0 669 5 1 1 668
0 670 7 1 2 1055 669
0 671 5 1 1 670
0 672 7 1 2 1192 600
0 673 5 1 1 672
0 674 7 1 2 1195 1208
0 675 5 1 1 674
0 676 7 1 2 1197 596
0 677 5 1 1 676
0 678 7 1 2 1202 1205
0 679 5 1 1 678
0 680 7 1 2 1200 592
0 681 5 1 1 680
0 682 7 1 2 679 681
0 683 7 1 2 677 682
0 684 7 1 2 675 683
0 685 5 1 1 684
0 686 7 1 2 673 685
0 687 7 1 2 671 686
0 688 7 1 2 667 687
0 689 7 1 2 665 688
0 690 7 1 2 663 689
0 691 7 1 2 661 690
0 692 7 1 2 659 691
0 693 5 1 1 692
0 694 7 1 2 657 693
0 695 7 1 2 655 694
0 696 7 1 2 651 695
0 697 7 1 2 649 696
0 698 7 1 2 647 697
0 699 7 1 2 939 698
0 700 7 1 2 645 699
0 701 7 1 2 639 700
0 702 7 2 2 955 643
0 703 5 1 1 1231
0 704 7 1 2 941 703
0 705 5 1 1 704
0 706 7 1 2 942 950
0 707 5 1 1 706
0 708 7 1 2 1232 707
0 709 5 1 1 708
0 710 7 1 2 705 709
0 711 7 1 2 701 710
0 712 7 1 2 1153 711
0 713 5 1 1 712
0 714 7 1 2 581 713
3 1499 5 0 1 714
