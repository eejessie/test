1 0 0 2 0
2 49 1 0
2 723 1 0
1 1 0 2 0
2 724 1 1
2 725 1 1
1 2 0 2 0
2 726 1 2
2 727 1 2
1 3 0 2 0
2 728 1 3
2 729 1 3
1 4 0 2 0
2 730 1 4
2 731 1 4
1 5 0 2 0
2 732 1 5
2 733 1 5
1 6 0 2 0
2 734 1 6
2 735 1 6
1 7 0 2 0
2 736 1 7
2 737 1 7
1 8 0 2 0
2 738 1 8
2 739 1 8
1 9 0 2 0
2 740 1 9
2 741 1 9
1 10 0 2 0
2 742 1 10
2 743 1 10
1 11 0 2 0
2 744 1 11
2 745 1 11
1 12 0 2 0
2 746 1 12
2 747 1 12
1 13 0 2 0
2 748 1 13
2 749 1 13
1 14 0 2 0
2 750 1 14
2 751 1 14
1 15 0 2 0
2 752 1 15
2 753 1 15
1 16 0 2 0
2 754 1 16
2 755 1 16
1 17 0 2 0
2 756 1 17
2 757 1 17
1 18 0 2 0
2 758 1 18
2 759 1 18
1 19 0 2 0
2 760 1 19
2 761 1 19
1 20 0 2 0
2 762 1 20
2 763 1 20
1 21 0 2 0
2 764 1 21
2 765 1 21
1 22 0 2 0
2 766 1 22
2 767 1 22
1 23 0 2 0
2 768 1 23
2 769 1 23
1 24 0 2 0
2 770 1 24
2 771 1 24
1 25 0 2 0
2 772 1 25
2 773 1 25
1 26 0 2 0
2 774 1 26
2 775 1 26
1 27 0 2 0
2 776 1 27
2 777 1 27
1 28 0 2 0
2 778 1 28
2 779 1 28
1 29 0 2 0
2 780 1 29
2 781 1 29
1 30 0 2 0
2 782 1 30
2 783 1 30
1 31 0 2 0
2 784 1 31
2 785 1 31
1 32 0 2 0
2 786 1 32
2 787 1 32
1 33 0 2 0
2 788 1 33
2 789 1 33
1 34 0 2 0
2 790 1 34
2 791 1 34
1 35 0 2 0
2 792 1 35
2 793 1 35
1 36 0 2 0
2 794 1 36
2 795 1 36
1 37 0 2 0
2 796 1 37
2 797 1 37
1 38 0 2 0
2 798 1 38
2 799 1 38
1 39 0 2 0
2 800 1 39
2 801 1 39
1 40 0 2 0
2 802 1 40
2 803 1 40
1 41 0 2 0
2 804 1 41
2 805 1 41
1 42 0 2 0
2 806 1 42
2 807 1 42
1 43 0 2 0
2 808 1 43
2 809 1 43
1 44 0 2 0
2 810 1 44
2 811 1 44
1 45 0 2 0
2 812 1 45
2 813 1 45
1 46 0 2 0
2 814 1 46
2 815 1 46
1 47 0 2 0
2 816 1 47
2 817 1 47
1 48 0 2 0
2 818 1 48
2 819 1 48
2 820 1 69
2 821 1 69
2 822 1 70
2 823 1 70
2 824 1 71
2 825 1 71
2 826 1 72
2 827 1 72
2 828 1 73
2 829 1 73
2 830 1 74
2 831 1 74
2 832 1 75
2 833 1 75
2 834 1 76
2 835 1 76
2 836 1 77
2 837 1 77
2 838 1 78
2 839 1 78
2 840 1 79
2 841 1 79
2 842 1 80
2 843 1 80
2 844 1 81
2 845 1 81
2 846 1 100
2 847 1 100
2 848 1 102
2 849 1 102
2 850 1 104
2 851 1 104
2 852 1 106
2 853 1 106
2 854 1 107
2 855 1 107
2 856 1 108
2 857 1 108
2 858 1 108
2 859 1 111
2 860 1 111
2 861 1 112
2 862 1 112
2 863 1 115
2 864 1 115
2 865 1 118
2 866 1 118
2 867 1 120
2 868 1 120
2 869 1 123
2 870 1 123
2 871 1 126
2 872 1 126
2 873 1 128
2 874 1 128
2 875 1 131
2 876 1 131
2 877 1 134
2 878 1 134
2 879 1 136
2 880 1 136
2 881 1 139
2 882 1 139
2 883 1 142
2 884 1 142
2 885 1 144
2 886 1 144
2 887 1 147
2 888 1 147
2 889 1 150
2 890 1 150
2 891 1 152
2 892 1 152
2 893 1 155
2 894 1 155
2 895 1 158
2 896 1 158
2 897 1 160
2 898 1 160
2 899 1 163
2 900 1 163
2 901 1 166
2 902 1 166
2 903 1 168
2 904 1 168
2 905 1 171
2 906 1 171
2 907 1 174
2 908 1 174
2 909 1 176
2 910 1 176
2 911 1 179
2 912 1 179
2 913 1 182
2 914 1 182
2 915 1 184
2 916 1 184
2 917 1 187
2 918 1 187
2 919 1 190
2 920 1 190
2 921 1 192
2 922 1 192
2 923 1 195
2 924 1 195
2 925 1 198
2 926 1 198
2 927 1 200
2 928 1 200
2 929 1 203
2 930 1 203
2 931 1 206
2 932 1 206
2 933 1 208
2 934 1 208
2 935 1 211
2 936 1 211
2 937 1 214
2 938 1 214
2 939 1 216
2 940 1 216
2 941 1 219
2 942 1 219
2 943 1 221
2 944 1 221
2 945 1 222
2 946 1 222
2 947 1 223
2 948 1 223
2 949 1 224
2 950 1 224
2 951 1 225
2 952 1 225
2 953 1 231
2 954 1 231
2 955 1 233
2 956 1 233
2 957 1 234
2 958 1 234
2 959 1 234
2 960 1 235
2 961 1 235
2 962 1 241
2 963 1 241
2 964 1 244
2 965 1 244
2 966 1 244
2 967 1 244
2 968 1 246
2 969 1 246
2 970 1 246
2 971 1 247
2 972 1 247
2 973 1 253
2 974 1 253
2 975 1 256
2 976 1 256
2 977 1 256
2 978 1 256
2 979 1 258
2 980 1 258
2 981 1 258
2 982 1 258
2 983 1 259
2 984 1 259
2 985 1 265
2 986 1 265
2 987 1 268
2 988 1 268
2 989 1 268
2 990 1 268
2 991 1 270
2 992 1 270
2 993 1 270
2 994 1 270
2 995 1 271
2 996 1 271
2 997 1 277
2 998 1 277
2 999 1 280
2 1000 1 280
2 1001 1 280
2 1002 1 280
2 1003 1 282
2 1004 1 282
2 1005 1 282
2 1006 1 282
2 1007 1 283
2 1008 1 283
2 1009 1 289
2 1010 1 289
2 1011 1 292
2 1012 1 292
2 1013 1 292
2 1014 1 292
2 1015 1 294
2 1016 1 294
2 1017 1 294
2 1018 1 295
2 1019 1 295
2 1020 1 301
2 1021 1 301
2 1022 1 304
2 1023 1 304
2 1024 1 304
2 1025 1 304
2 1026 1 305
2 1027 1 305
2 1028 1 311
2 1029 1 311
2 1030 1 314
2 1031 1 314
2 1032 1 314
2 1033 1 314
2 1034 1 316
2 1035 1 316
2 1036 1 316
2 1037 1 316
2 1038 1 317
2 1039 1 317
2 1040 1 323
2 1041 1 323
2 1042 1 326
2 1043 1 326
2 1044 1 326
2 1045 1 328
2 1046 1 328
2 1047 1 328
2 1048 1 329
2 1049 1 329
2 1050 1 335
2 1051 1 335
2 1052 1 338
2 1053 1 338
2 1054 1 338
2 1055 1 340
2 1056 1 340
2 1057 1 340
2 1058 1 341
2 1059 1 341
2 1060 1 347
2 1061 1 347
2 1062 1 349
2 1063 1 349
2 1064 1 350
2 1065 1 350
2 1066 1 350
2 1067 1 351
2 1068 1 351
2 1069 1 352
2 1070 1 352
2 1071 1 352
2 1072 1 353
2 1073 1 353
2 1074 1 359
2 1075 1 359
2 1076 1 362
2 1077 1 362
2 1078 1 362
2 1079 1 364
2 1080 1 364
2 1081 1 364
2 1082 1 365
2 1083 1 365
2 1084 1 371
2 1085 1 371
2 1086 1 374
2 1087 1 374
2 1088 1 374
2 1089 1 376
2 1090 1 376
2 1091 1 376
2 1092 1 377
2 1093 1 377
2 1094 1 383
2 1095 1 383
2 1096 1 386
2 1097 1 386
2 1098 1 386
2 1099 1 388
2 1100 1 388
2 1101 1 388
2 1102 1 389
2 1103 1 389
2 1104 1 395
2 1105 1 395
2 1106 1 398
2 1107 1 398
2 1108 1 400
2 1109 1 400
2 1110 1 403
2 1111 1 403
2 1112 1 409
2 1113 1 409
2 1114 1 410
2 1115 1 410
2 1116 1 413
2 1117 1 413
2 1118 1 413
2 1119 1 417
2 1120 1 417
2 1121 1 418
2 1122 1 418
2 1123 1 422
2 1124 1 422
2 1125 1 425
2 1126 1 425
2 1127 1 429
2 1128 1 429
2 1129 1 430
2 1130 1 430
2 1131 1 433
2 1132 1 433
2 1133 1 436
2 1134 1 436
2 1135 1 441
2 1136 1 441
2 1137 1 441
2 1138 1 441
2 1139 1 444
2 1140 1 444
2 1141 1 448
2 1142 1 448
2 1143 1 452
2 1144 1 452
2 1145 1 456
2 1146 1 456
2 1147 1 462
2 1148 1 462
2 1149 1 463
2 1150 1 463
2 1151 1 464
2 1152 1 464
2 1153 1 464
2 1154 1 467
2 1155 1 467
2 1156 1 471
2 1157 1 471
2 1158 1 475
2 1159 1 475
2 1160 1 481
2 1161 1 481
2 1162 1 481
2 1163 1 487
2 1164 1 487
2 1165 1 493
2 1166 1 493
2 1167 1 498
2 1168 1 498
2 1169 1 504
2 1170 1 504
2 1171 1 505
2 1172 1 505
2 1173 1 508
2 1174 1 508
2 1175 1 514
2 1176 1 514
2 1177 1 517
2 1178 1 517
2 1179 1 517
2 1180 1 518
2 1181 1 518
2 1182 1 525
2 1183 1 525
2 1184 1 525
2 1185 1 525
2 1186 1 526
2 1187 1 526
2 1188 1 535
2 1189 1 535
2 1190 1 535
2 1191 1 536
2 1192 1 536
2 1193 1 541
2 1194 1 541
2 1195 1 541
2 1196 1 542
2 1197 1 542
2 1198 1 545
2 1199 1 545
2 1200 1 546
2 1201 1 546
2 1202 1 548
2 1203 1 548
2 1204 1 552
2 1205 1 552
2 1206 1 583
2 1207 1 583
2 1208 1 586
2 1209 1 586
2 1210 1 587
2 1211 1 587
2 1212 1 590
2 1213 1 590
2 1214 1 591
2 1215 1 591
2 1216 1 594
2 1217 1 594
2 1218 1 595
2 1219 1 595
2 1220 1 598
2 1221 1 598
2 1222 1 602
2 1223 1 602
2 1224 1 603
2 1225 1 603
2 1226 1 606
2 1227 1 606
2 1228 1 609
2 1229 1 609
2 1230 1 614
2 1231 1 614
2 1232 1 618
2 1233 1 618
2 1234 1 621
2 1235 1 621
2 1236 1 626
2 1237 1 626
2 1238 1 628
2 1239 1 628
2 1240 1 628
2 1241 1 632
2 1242 1 632
2 1243 1 632
0 50 5 1 1 49
0 51 5 1 1 724
0 52 5 1 1 726
0 53 5 1 1 728
0 54 5 1 1 730
0 55 5 1 1 732
0 56 5 1 1 734
0 57 5 1 1 736
0 58 5 1 1 738
0 59 5 1 1 740
0 60 5 1 1 742
0 61 5 1 1 744
0 62 5 1 1 746
0 63 5 1 1 748
0 64 5 1 1 750
0 65 5 1 1 752
0 66 5 1 1 754
0 67 5 1 1 756
0 68 5 1 1 758
0 69 5 2 1 760
0 70 5 2 1 762
0 71 5 2 1 764
0 72 5 2 1 766
0 73 5 2 1 768
0 74 5 2 1 770
0 75 5 2 1 772
0 76 5 2 1 774
0 77 5 2 1 776
0 78 5 2 1 778
0 79 5 2 1 780
0 80 5 2 1 782
0 81 5 2 1 784
0 82 5 1 1 786
0 83 5 1 1 788
0 84 5 1 1 790
0 85 5 1 1 792
0 86 5 1 1 794
0 87 5 1 1 796
0 88 5 1 1 798
0 89 5 1 1 800
0 90 5 1 1 802
0 91 5 1 1 804
0 92 5 1 1 806
0 93 5 1 1 808
0 94 5 1 1 810
0 95 5 1 1 812
0 96 5 1 1 814
0 97 5 1 1 816
0 98 5 1 1 818
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 727 759
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 725 757
0 106 5 2 1 105
0 107 7 2 2 723 755
0 108 5 3 1 854
0 109 7 1 2 852 856
0 110 5 1 1 109
0 111 7 2 2 850 110
0 112 5 2 1 859
0 113 7 1 2 848 861
0 114 5 1 1 113
0 115 7 2 2 846 114
0 116 5 1 1 863
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 729 864
0 120 5 2 1 119
0 121 7 1 2 820 867
0 122 5 1 1 121
0 123 7 2 2 865 122
0 124 5 1 1 869
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 731 870
0 128 5 2 1 127
0 129 7 1 2 822 873
0 130 5 1 1 129
0 131 7 2 2 871 130
0 132 5 1 1 875
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 733 876
0 136 5 2 1 135
0 137 7 1 2 824 879
0 138 5 1 1 137
0 139 7 2 2 877 138
0 140 5 1 1 881
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 735 882
0 144 5 2 1 143
0 145 7 1 2 826 885
0 146 5 1 1 145
0 147 7 2 2 883 146
0 148 5 1 1 887
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 737 888
0 152 5 2 1 151
0 153 7 1 2 828 891
0 154 5 1 1 153
0 155 7 2 2 889 154
0 156 5 1 1 893
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 739 894
0 160 5 2 1 159
0 161 7 1 2 830 897
0 162 5 1 1 161
0 163 7 2 2 895 162
0 164 5 1 1 899
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 741 900
0 168 5 2 1 167
0 169 7 1 2 832 903
0 170 5 1 1 169
0 171 7 2 2 901 170
0 172 5 1 1 905
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 743 906
0 176 5 2 1 175
0 177 7 1 2 834 909
0 178 5 1 1 177
0 179 7 2 2 907 178
0 180 5 1 1 911
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 745 912
0 184 5 2 1 183
0 185 7 1 2 836 915
0 186 5 1 1 185
0 187 7 2 2 913 186
0 188 5 1 1 917
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 747 918
0 192 5 2 1 191
0 193 7 1 2 838 921
0 194 5 1 1 193
0 195 7 2 2 919 194
0 196 5 1 1 923
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 749 924
0 200 5 2 1 199
0 201 7 1 2 840 927
0 202 5 1 1 201
0 203 7 2 2 925 202
0 204 5 1 1 929
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 751 930
0 208 5 2 1 207
0 209 7 1 2 842 933
0 210 5 1 1 209
0 211 7 2 2 931 210
0 212 5 1 1 935
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 753 936
0 216 5 2 1 215
0 217 7 1 2 844 939
0 218 5 1 1 217
0 219 7 2 2 937 218
0 220 5 1 1 941
0 221 7 2 2 819 220
0 222 5 2 1 943
0 223 7 2 2 98 942
0 224 5 2 1 947
0 225 7 2 2 938 940
0 226 5 1 1 951
0 227 7 1 2 785 226
0 228 5 1 1 227
0 229 7 1 2 845 952
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 953
0 233 7 2 2 817 954
0 234 5 3 1 955
0 235 7 2 2 932 934
0 236 5 1 1 960
0 237 7 1 2 783 961
0 238 5 1 1 237
0 239 7 1 2 843 236
0 240 5 1 1 239
0 241 7 2 2 238 240
0 242 5 1 1 962
0 243 7 1 2 815 242
0 244 5 4 1 243
0 245 7 1 2 96 963
0 246 5 3 1 245
0 247 7 2 2 926 928
0 248 5 1 1 971
0 249 7 1 2 781 972
0 250 5 1 1 249
0 251 7 1 2 841 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 973
0 255 7 1 2 813 254
0 256 5 4 1 255
0 257 7 1 2 95 974
0 258 5 4 1 257
0 259 7 2 2 920 922
0 260 5 1 1 983
0 261 7 1 2 779 984
0 262 5 1 1 261
0 263 7 1 2 839 260
0 264 5 1 1 263
0 265 7 2 2 262 264
0 266 5 1 1 985
0 267 7 1 2 811 266
0 268 5 4 1 267
0 269 7 1 2 94 986
0 270 5 4 1 269
0 271 7 2 2 914 916
0 272 5 1 1 995
0 273 7 1 2 777 996
0 274 5 1 1 273
0 275 7 1 2 837 272
0 276 5 1 1 275
0 277 7 2 2 274 276
0 278 5 1 1 997
0 279 7 1 2 809 278
0 280 5 4 1 279
0 281 7 1 2 93 998
0 282 5 4 1 281
0 283 7 2 2 908 910
0 284 5 1 1 1007
0 285 7 1 2 775 1008
0 286 5 1 1 285
0 287 7 1 2 835 284
0 288 5 1 1 287
0 289 7 2 2 286 288
0 290 5 1 1 1009
0 291 7 1 2 807 290
0 292 5 4 1 291
0 293 7 1 2 92 1010
0 294 5 3 1 293
0 295 7 2 2 902 904
0 296 5 1 1 1018
0 297 7 1 2 773 1019
0 298 5 1 1 297
0 299 7 1 2 833 296
0 300 5 1 1 299
0 301 7 2 2 298 300
0 302 5 1 1 1020
0 303 7 1 2 805 302
0 304 5 4 1 303
0 305 7 2 2 896 898
0 306 5 1 1 1026
0 307 7 1 2 771 1027
0 308 5 1 1 307
0 309 7 1 2 831 306
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 1028
0 313 7 1 2 803 312
0 314 5 4 1 313
0 315 7 1 2 90 1029
0 316 5 4 1 315
0 317 7 2 2 890 892
0 318 5 1 1 1038
0 319 7 1 2 769 1039
0 320 5 1 1 319
0 321 7 1 2 829 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1040
0 325 7 1 2 801 324
0 326 5 3 1 325
0 327 7 1 2 89 1041
0 328 5 3 1 327
0 329 7 2 2 884 886
0 330 5 1 1 1048
0 331 7 1 2 767 1049
0 332 5 1 1 331
0 333 7 1 2 827 330
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 1050
0 337 7 1 2 799 336
0 338 5 3 1 337
0 339 7 1 2 88 1051
0 340 5 3 1 339
0 341 7 2 2 878 880
0 342 5 1 1 1058
0 343 7 1 2 765 1059
0 344 5 1 1 343
0 345 7 1 2 825 342
0 346 5 1 1 345
0 347 7 2 2 344 346
0 348 5 1 1 1060
0 349 7 2 2 797 348
0 350 5 3 1 1062
0 351 7 2 2 87 1061
0 352 5 3 1 1067
0 353 7 2 2 872 874
0 354 5 1 1 1072
0 355 7 1 2 763 1073
0 356 5 1 1 355
0 357 7 1 2 823 354
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 1074
0 361 7 1 2 795 360
0 362 5 3 1 361
0 363 7 1 2 86 1075
0 364 5 3 1 363
0 365 7 2 2 866 868
0 366 5 1 1 1082
0 367 7 1 2 761 1083
0 368 5 1 1 367
0 369 7 1 2 821 366
0 370 5 1 1 369
0 371 7 2 2 368 370
0 372 5 1 1 1084
0 373 7 1 2 793 372
0 374 5 3 1 373
0 375 7 1 2 85 1085
0 376 5 3 1 375
0 377 7 2 2 847 849
0 378 5 1 1 1092
0 379 7 1 2 860 378
0 380 5 1 1 379
0 381 7 1 2 862 1093
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 1094
0 385 7 1 2 84 384
0 386 5 3 1 385
0 387 7 1 2 791 1095
0 388 5 3 1 387
0 389 7 2 2 851 853
0 390 5 1 1 1102
0 391 7 1 2 855 390
0 392 5 1 1 391
0 393 7 1 2 857 1103
0 394 5 1 1 393
0 395 7 2 2 392 394
0 396 5 1 1 1104
0 397 7 1 2 83 396
0 398 5 2 1 397
0 399 7 1 2 789 1105
0 400 5 2 1 399
0 401 7 1 2 50 66
0 402 5 1 1 401
0 403 7 2 2 858 402
0 404 5 1 1 1110
0 405 7 1 2 787 404
0 406 5 1 1 405
0 407 7 1 2 1108 406
0 408 5 1 1 407
0 409 7 2 2 1106 408
0 410 5 2 1 1112
0 411 7 1 2 1099 1114
0 412 5 1 1 411
0 413 7 3 2 1096 412
0 414 5 1 1 1116
0 415 7 1 2 1089 1117
0 416 5 1 1 415
0 417 7 2 2 1086 416
0 418 5 2 1 1119
0 419 7 1 2 1079 1121
0 420 5 1 1 419
0 421 7 1 2 1076 420
0 422 5 2 1 421
0 423 7 1 2 1069 1123
0 424 5 1 1 423
0 425 7 2 2 1064 424
0 426 5 1 1 1125
0 427 7 1 2 1055 426
0 428 5 1 1 427
0 429 7 2 2 1052 428
0 430 5 2 1 1127
0 431 7 1 2 1045 1129
0 432 5 1 1 431
0 433 7 2 2 1042 432
0 434 5 1 1 1131
0 435 7 1 2 1034 434
0 436 5 2 1 435
0 437 7 1 2 1030 1133
0 438 7 1 2 1022 437
0 439 5 1 1 438
0 440 7 1 2 91 1021
0 441 5 4 1 440
0 442 7 1 2 439 1135
0 443 7 1 2 1015 442
0 444 5 2 1 443
0 445 7 1 2 1011 1139
0 446 5 1 1 445
0 447 7 1 2 1003 446
0 448 5 2 1 447
0 449 7 1 2 999 1141
0 450 5 1 1 449
0 451 7 1 2 991 450
0 452 5 2 1 451
0 453 7 1 2 987 1143
0 454 5 1 1 453
0 455 7 1 2 979 454
0 456 5 2 1 455
0 457 7 1 2 975 1145
0 458 5 1 1 457
0 459 7 1 2 968 458
0 460 5 1 1 459
0 461 7 1 2 964 460
0 462 5 2 1 461
0 463 7 2 2 97 232
0 464 5 3 1 1149
0 465 7 1 2 1147 1151
0 466 5 1 1 465
0 467 7 2 2 957 466
0 468 5 1 1 1154
0 469 7 1 2 949 468
0 470 5 1 1 469
0 471 7 2 2 945 470
0 472 5 1 1 1156
0 473 7 1 2 948 1155
0 474 5 1 1 473
0 475 7 2 2 1152 958
0 476 5 1 1 1158
0 477 7 1 2 965 476
0 478 5 1 1 477
0 479 7 1 2 1148 1159
0 480 5 1 1 479
0 481 7 3 2 966 969
0 482 5 1 1 1160
0 483 7 1 2 1146 1161
0 484 5 1 1 483
0 485 7 1 2 976 484
0 486 5 1 1 485
0 487 7 2 2 977 980
0 488 5 1 1 1163
0 489 7 1 2 1144 1164
0 490 5 1 1 489
0 491 7 1 2 988 490
0 492 5 1 1 491
0 493 7 2 2 989 992
0 494 7 1 2 1142 1165
0 495 5 1 1 494
0 496 7 1 2 1000 495
0 497 5 1 1 496
0 498 7 2 2 1001 1004
0 499 5 1 1 1167
0 500 7 1 2 1140 1168
0 501 5 1 1 500
0 502 7 1 2 1012 501
0 503 5 1 1 502
0 504 7 2 2 1013 1016
0 505 5 2 1 1169
0 506 7 1 2 1023 1171
0 507 5 1 1 506
0 508 7 2 2 1024 1136
0 509 7 1 2 1134 1173
0 510 5 1 1 509
0 511 7 1 2 1031 510
0 512 5 1 1 511
0 513 7 1 2 1032 1035
0 514 5 2 1 513
0 515 7 1 2 1132 1175
0 516 5 1 1 515
0 517 7 3 2 1043 1046
0 518 5 2 1 1177
0 519 7 1 2 1130 1180
0 520 5 1 1 519
0 521 7 1 2 1128 1178
0 522 5 1 1 521
0 523 7 1 2 520 522
0 524 5 1 1 523
0 525 7 4 2 1053 1056
0 526 5 2 1 1182
0 527 7 1 2 1065 1183
0 528 5 1 1 527
0 529 7 1 2 1124 528
0 530 5 1 1 529
0 531 7 1 2 1126 1184
0 532 5 1 1 531
0 533 7 1 2 1070 1186
0 534 5 1 1 533
0 535 7 3 2 1077 1080
0 536 5 2 1 1188
0 537 7 1 2 1122 1189
0 538 5 1 1 537
0 539 7 1 2 1120 1191
0 540 5 1 1 539
0 541 7 3 2 1087 1090
0 542 5 2 1 1193
0 543 7 1 2 1118 1194
0 544 5 1 1 543
0 545 7 2 2 1097 1100
0 546 5 2 1 1198
0 547 7 1 2 1113 1200
0 548 5 2 1 547
0 549 7 1 2 82 1111
0 550 5 1 1 549
0 551 7 1 2 1107 550
0 552 5 2 1 551
0 553 7 1 2 1201 1204
0 554 5 1 1 553
0 555 7 1 2 1115 554
0 556 5 1 1 555
0 557 7 1 2 1202 556
0 558 5 1 1 557
0 559 7 1 2 414 1196
0 560 5 1 1 559
0 561 7 1 2 558 560
0 562 7 1 2 544 561
0 563 7 1 2 540 562
0 564 7 1 2 538 563
0 565 5 1 1 564
0 566 7 1 2 534 565
0 567 7 1 2 532 566
0 568 7 1 2 530 567
0 569 5 1 1 568
0 570 7 1 2 524 569
0 571 7 1 2 516 570
0 572 7 1 2 512 571
0 573 7 1 2 507 572
0 574 7 1 2 503 573
0 575 7 1 2 497 574
0 576 7 1 2 492 575
0 577 7 1 2 486 576
0 578 7 1 2 480 577
0 579 7 1 2 478 578
0 580 7 1 2 474 579
0 581 7 1 2 1157 580
0 582 5 1 1 581
0 583 7 2 2 1109 1205
0 584 7 1 2 1101 1206
0 585 5 1 1 584
0 586 7 2 2 1098 585
0 587 5 2 1 1208
0 588 7 1 2 1088 1210
0 589 5 1 1 588
0 590 7 2 2 1091 589
0 591 5 2 1 1212
0 592 7 1 2 1078 1214
0 593 5 1 1 592
0 594 7 2 2 1081 593
0 595 5 2 1 1216
0 596 7 1 2 1066 1218
0 597 5 1 1 596
0 598 7 2 2 1071 597
0 599 5 1 1 1220
0 600 7 1 2 1054 599
0 601 5 1 1 600
0 602 7 2 2 1057 601
0 603 5 2 1 1222
0 604 7 1 2 1044 1224
0 605 5 1 1 604
0 606 7 2 2 1047 605
0 607 5 1 1 1226
0 608 7 1 2 1033 607
0 609 5 2 1 608
0 610 7 1 2 1036 1228
0 611 5 1 1 610
0 612 7 1 2 1025 611
0 613 5 1 1 612
0 614 7 2 2 1137 613
0 615 5 1 1 1230
0 616 7 1 2 1017 1231
0 617 5 1 1 616
0 618 7 2 2 1014 617
0 619 5 1 1 1232
0 620 7 1 2 1002 1233
0 621 5 2 1 620
0 622 7 1 2 1005 1234
0 623 7 1 2 993 622
0 624 5 1 1 623
0 625 7 1 2 990 624
0 626 7 2 2 978 625
0 627 5 1 1 1236
0 628 7 3 2 981 627
0 629 5 1 1 1238
0 630 7 1 2 970 1239
0 631 5 1 1 630
0 632 7 3 2 967 631
0 633 5 1 1 1241
0 634 7 1 2 959 1242
0 635 5 1 1 634
0 636 7 1 2 946 635
0 637 5 1 1 636
0 638 7 1 2 1153 637
0 639 5 1 1 638
0 640 7 1 2 956 633
0 641 5 1 1 640
0 642 7 1 2 944 1243
0 643 5 1 1 642
0 644 7 1 2 1150 643
0 645 5 1 1 644
0 646 7 1 2 994 488
0 647 5 1 1 646
0 648 7 1 2 982 1237
0 649 5 1 1 648
0 650 7 1 2 1166 1235
0 651 5 1 1 650
0 652 7 1 2 1006 651
0 653 5 1 1 652
0 654 7 1 2 499 619
0 655 5 1 1 654
0 656 7 1 2 1170 615
0 657 5 1 1 656
0 658 7 1 2 1138 1172
0 659 5 1 1 658
0 660 7 1 2 1174 1229
0 661 5 1 1 660
0 662 7 1 2 1037 661
0 663 5 1 1 662
0 664 7 1 2 1176 1227
0 665 5 1 1 664
0 666 7 1 2 1181 1225
0 667 5 1 1 666
0 668 7 1 2 1179 1223
0 669 5 1 1 668
0 670 7 1 2 667 669
0 671 5 1 1 670
0 672 7 1 2 1063 1217
0 673 5 1 1 672
0 674 7 1 2 1187 673
0 675 5 1 1 674
0 676 7 1 2 1185 1221
0 677 5 1 1 676
0 678 7 1 2 1068 1219
0 679 5 1 1 678
0 680 7 1 2 1192 1215
0 681 5 1 1 680
0 682 7 1 2 1190 1213
0 683 5 1 1 682
0 684 7 1 2 681 683
0 685 5 1 1 684
0 686 7 1 2 1197 1209
0 687 5 1 1 686
0 688 7 1 2 1195 1211
0 689 5 1 1 688
0 690 7 1 2 1199 1207
0 691 5 1 1 690
0 692 7 1 2 1203 691
0 693 7 1 2 689 692
0 694 7 1 2 687 693
0 695 7 1 2 685 694
0 696 5 1 1 695
0 697 7 1 2 679 696
0 698 7 1 2 677 697
0 699 7 1 2 675 698
0 700 5 1 1 699
0 701 7 1 2 671 700
0 702 7 1 2 665 701
0 703 7 1 2 663 702
0 704 7 1 2 659 703
0 705 7 1 2 657 704
0 706 7 1 2 655 705
0 707 7 1 2 653 706
0 708 7 1 2 649 707
0 709 7 1 2 647 708
0 710 7 1 2 950 709
0 711 7 1 2 1162 629
0 712 5 1 1 711
0 713 7 1 2 482 1240
0 714 5 1 1 713
0 715 7 1 2 712 714
0 716 7 1 2 710 715
0 717 7 1 2 645 716
0 718 7 1 2 641 717
0 719 7 1 2 639 718
0 720 7 1 2 472 719
0 721 5 1 1 720
0 722 7 1 2 582 721
3 3499 5 0 1 722
