1 0 0 6 0
2 49 1 0
2 4788 1 0
2 4789 1 0
2 4790 1 0
2 4791 1 0
2 4792 1 0
1 1 0 8 0
2 4793 1 1
2 4794 1 1
2 4795 1 1
2 4796 1 1
2 4797 1 1
2 4798 1 1
2 4799 1 1
2 4800 1 1
1 2 0 9 0
2 4801 1 2
2 4802 1 2
2 4803 1 2
2 4804 1 2
2 4805 1 2
2 4806 1 2
2 4807 1 2
2 4808 1 2
2 4809 1 2
1 3 0 8 0
2 4810 1 3
2 4811 1 3
2 4812 1 3
2 4813 1 3
2 4814 1 3
2 4815 1 3
2 4816 1 3
2 4817 1 3
1 4 0 8 0
2 4818 1 4
2 4819 1 4
2 4820 1 4
2 4821 1 4
2 4822 1 4
2 4823 1 4
2 4824 1 4
2 4825 1 4
1 5 0 8 0
2 4826 1 5
2 4827 1 5
2 4828 1 5
2 4829 1 5
2 4830 1 5
2 4831 1 5
2 4832 1 5
2 4833 1 5
1 6 0 8 0
2 4834 1 6
2 4835 1 6
2 4836 1 6
2 4837 1 6
2 4838 1 6
2 4839 1 6
2 4840 1 6
2 4841 1 6
1 7 0 8 0
2 4842 1 7
2 4843 1 7
2 4844 1 7
2 4845 1 7
2 4846 1 7
2 4847 1 7
2 4848 1 7
2 4849 1 7
1 8 0 8 0
2 4850 1 8
2 4851 1 8
2 4852 1 8
2 4853 1 8
2 4854 1 8
2 4855 1 8
2 4856 1 8
2 4857 1 8
1 9 0 8 0
2 4858 1 9
2 4859 1 9
2 4860 1 9
2 4861 1 9
2 4862 1 9
2 4863 1 9
2 4864 1 9
2 4865 1 9
1 10 0 8 0
2 4866 1 10
2 4867 1 10
2 4868 1 10
2 4869 1 10
2 4870 1 10
2 4871 1 10
2 4872 1 10
2 4873 1 10
1 11 0 8 0
2 4874 1 11
2 4875 1 11
2 4876 1 11
2 4877 1 11
2 4878 1 11
2 4879 1 11
2 4880 1 11
2 4881 1 11
1 12 0 8 0
2 4882 1 12
2 4883 1 12
2 4884 1 12
2 4885 1 12
2 4886 1 12
2 4887 1 12
2 4888 1 12
2 4889 1 12
1 13 0 8 0
2 4890 1 13
2 4891 1 13
2 4892 1 13
2 4893 1 13
2 4894 1 13
2 4895 1 13
2 4896 1 13
2 4897 1 13
1 14 0 8 0
2 4898 1 14
2 4899 1 14
2 4900 1 14
2 4901 1 14
2 4902 1 14
2 4903 1 14
2 4904 1 14
2 4905 1 14
1 15 0 8 0
2 4906 1 15
2 4907 1 15
2 4908 1 15
2 4909 1 15
2 4910 1 15
2 4911 1 15
2 4912 1 15
2 4913 1 15
1 16 0 8 0
2 4914 1 16
2 4915 1 16
2 4916 1 16
2 4917 1 16
2 4918 1 16
2 4919 1 16
2 4920 1 16
2 4921 1 16
1 17 0 8 0
2 4922 1 17
2 4923 1 17
2 4924 1 17
2 4925 1 17
2 4926 1 17
2 4927 1 17
2 4928 1 17
2 4929 1 17
1 18 0 8 0
2 4930 1 18
2 4931 1 18
2 4932 1 18
2 4933 1 18
2 4934 1 18
2 4935 1 18
2 4936 1 18
2 4937 1 18
1 19 0 8 0
2 4938 1 19
2 4939 1 19
2 4940 1 19
2 4941 1 19
2 4942 1 19
2 4943 1 19
2 4944 1 19
2 4945 1 19
1 20 0 8 0
2 4946 1 20
2 4947 1 20
2 4948 1 20
2 4949 1 20
2 4950 1 20
2 4951 1 20
2 4952 1 20
2 4953 1 20
1 21 0 8 0
2 4954 1 21
2 4955 1 21
2 4956 1 21
2 4957 1 21
2 4958 1 21
2 4959 1 21
2 4960 1 21
2 4961 1 21
1 22 0 8 0
2 4962 1 22
2 4963 1 22
2 4964 1 22
2 4965 1 22
2 4966 1 22
2 4967 1 22
2 4968 1 22
2 4969 1 22
1 23 0 8 0
2 4970 1 23
2 4971 1 23
2 4972 1 23
2 4973 1 23
2 4974 1 23
2 4975 1 23
2 4976 1 23
2 4977 1 23
1 24 0 8 0
2 4978 1 24
2 4979 1 24
2 4980 1 24
2 4981 1 24
2 4982 1 24
2 4983 1 24
2 4984 1 24
2 4985 1 24
1 25 0 8 0
2 4986 1 25
2 4987 1 25
2 4988 1 25
2 4989 1 25
2 4990 1 25
2 4991 1 25
2 4992 1 25
2 4993 1 25
1 26 0 8 0
2 4994 1 26
2 4995 1 26
2 4996 1 26
2 4997 1 26
2 4998 1 26
2 4999 1 26
2 5000 1 26
2 5001 1 26
1 27 0 8 0
2 5002 1 27
2 5003 1 27
2 5004 1 27
2 5005 1 27
2 5006 1 27
2 5007 1 27
2 5008 1 27
2 5009 1 27
1 28 0 8 0
2 5010 1 28
2 5011 1 28
2 5012 1 28
2 5013 1 28
2 5014 1 28
2 5015 1 28
2 5016 1 28
2 5017 1 28
1 29 0 8 0
2 5018 1 29
2 5019 1 29
2 5020 1 29
2 5021 1 29
2 5022 1 29
2 5023 1 29
2 5024 1 29
2 5025 1 29
1 30 0 8 0
2 5026 1 30
2 5027 1 30
2 5028 1 30
2 5029 1 30
2 5030 1 30
2 5031 1 30
2 5032 1 30
2 5033 1 30
1 31 0 8 0
2 5034 1 31
2 5035 1 31
2 5036 1 31
2 5037 1 31
2 5038 1 31
2 5039 1 31
2 5040 1 31
2 5041 1 31
1 32 0 8 0
2 5042 1 32
2 5043 1 32
2 5044 1 32
2 5045 1 32
2 5046 1 32
2 5047 1 32
2 5048 1 32
2 5049 1 32
1 33 0 8 0
2 5050 1 33
2 5051 1 33
2 5052 1 33
2 5053 1 33
2 5054 1 33
2 5055 1 33
2 5056 1 33
2 5057 1 33
1 34 0 8 0
2 5058 1 34
2 5059 1 34
2 5060 1 34
2 5061 1 34
2 5062 1 34
2 5063 1 34
2 5064 1 34
2 5065 1 34
1 35 0 8 0
2 5066 1 35
2 5067 1 35
2 5068 1 35
2 5069 1 35
2 5070 1 35
2 5071 1 35
2 5072 1 35
2 5073 1 35
1 36 0 8 0
2 5074 1 36
2 5075 1 36
2 5076 1 36
2 5077 1 36
2 5078 1 36
2 5079 1 36
2 5080 1 36
2 5081 1 36
1 37 0 8 0
2 5082 1 37
2 5083 1 37
2 5084 1 37
2 5085 1 37
2 5086 1 37
2 5087 1 37
2 5088 1 37
2 5089 1 37
1 38 0 8 0
2 5090 1 38
2 5091 1 38
2 5092 1 38
2 5093 1 38
2 5094 1 38
2 5095 1 38
2 5096 1 38
2 5097 1 38
1 39 0 8 0
2 5098 1 39
2 5099 1 39
2 5100 1 39
2 5101 1 39
2 5102 1 39
2 5103 1 39
2 5104 1 39
2 5105 1 39
1 40 0 8 0
2 5106 1 40
2 5107 1 40
2 5108 1 40
2 5109 1 40
2 5110 1 40
2 5111 1 40
2 5112 1 40
2 5113 1 40
1 41 0 8 0
2 5114 1 41
2 5115 1 41
2 5116 1 41
2 5117 1 41
2 5118 1 41
2 5119 1 41
2 5120 1 41
2 5121 1 41
1 42 0 8 0
2 5122 1 42
2 5123 1 42
2 5124 1 42
2 5125 1 42
2 5126 1 42
2 5127 1 42
2 5128 1 42
2 5129 1 42
1 43 0 8 0
2 5130 1 43
2 5131 1 43
2 5132 1 43
2 5133 1 43
2 5134 1 43
2 5135 1 43
2 5136 1 43
2 5137 1 43
1 44 0 8 0
2 5138 1 44
2 5139 1 44
2 5140 1 44
2 5141 1 44
2 5142 1 44
2 5143 1 44
2 5144 1 44
2 5145 1 44
1 45 0 10 0
2 5146 1 45
2 5147 1 45
2 5148 1 45
2 5149 1 45
2 5150 1 45
2 5151 1 45
2 5152 1 45
2 5153 1 45
2 5154 1 45
2 5155 1 45
1 46 0 9 0
2 5156 1 46
2 5157 1 46
2 5158 1 46
2 5159 1 46
2 5160 1 46
2 5161 1 46
2 5162 1 46
2 5163 1 46
2 5164 1 46
1 47 0 8 0
2 5165 1 47
2 5166 1 47
2 5167 1 47
2 5168 1 47
2 5169 1 47
2 5170 1 47
2 5171 1 47
2 5172 1 47
1 48 0 7 0
2 5173 1 48
2 5174 1 48
2 5175 1 48
2 5176 1 48
2 5177 1 48
2 5178 1 48
2 5179 1 48
2 5180 1 50
2 5181 1 50
2 5182 1 50
2 5183 1 50
2 5184 1 50
2 5185 1 50
2 5186 1 50
2 5187 1 51
2 5188 1 51
2 5189 1 51
2 5190 1 51
2 5191 1 51
2 5192 1 51
2 5193 1 52
2 5194 1 52
2 5195 1 52
2 5196 1 52
2 5197 1 52
2 5198 1 52
2 5199 1 52
2 5200 1 53
2 5201 1 53
2 5202 1 53
2 5203 1 53
2 5204 1 53
2 5205 1 53
2 5206 1 53
2 5207 1 54
2 5208 1 54
2 5209 1 54
2 5210 1 54
2 5211 1 54
2 5212 1 54
2 5213 1 54
2 5214 1 55
2 5215 1 55
2 5216 1 55
2 5217 1 55
2 5218 1 55
2 5219 1 55
2 5220 1 55
2 5221 1 56
2 5222 1 56
2 5223 1 56
2 5224 1 56
2 5225 1 56
2 5226 1 56
2 5227 1 56
2 5228 1 57
2 5229 1 57
2 5230 1 57
2 5231 1 57
2 5232 1 57
2 5233 1 57
2 5234 1 57
2 5235 1 58
2 5236 1 58
2 5237 1 58
2 5238 1 58
2 5239 1 58
2 5240 1 58
2 5241 1 58
2 5242 1 59
2 5243 1 59
2 5244 1 59
2 5245 1 59
2 5246 1 59
2 5247 1 59
2 5248 1 59
2 5249 1 60
2 5250 1 60
2 5251 1 60
2 5252 1 60
2 5253 1 60
2 5254 1 60
2 5255 1 60
2 5256 1 61
2 5257 1 61
2 5258 1 61
2 5259 1 61
2 5260 1 61
2 5261 1 61
2 5262 1 61
2 5263 1 62
2 5264 1 62
2 5265 1 62
2 5266 1 62
2 5267 1 62
2 5268 1 62
2 5269 1 62
2 5270 1 63
2 5271 1 63
2 5272 1 63
2 5273 1 63
2 5274 1 63
2 5275 1 63
2 5276 1 63
2 5277 1 64
2 5278 1 64
2 5279 1 64
2 5280 1 64
2 5281 1 64
2 5282 1 64
2 5283 1 64
2 5284 1 65
2 5285 1 65
2 5286 1 65
2 5287 1 65
2 5288 1 65
2 5289 1 65
2 5290 1 65
2 5291 1 66
2 5292 1 66
2 5293 1 66
2 5294 1 66
2 5295 1 66
2 5296 1 66
2 5297 1 66
2 5298 1 67
2 5299 1 67
2 5300 1 67
2 5301 1 67
2 5302 1 67
2 5303 1 67
2 5304 1 67
2 5305 1 68
2 5306 1 68
2 5307 1 68
2 5308 1 68
2 5309 1 68
2 5310 1 68
2 5311 1 68
2 5312 1 69
2 5313 1 69
2 5314 1 69
2 5315 1 69
2 5316 1 69
2 5317 1 69
2 5318 1 69
2 5319 1 69
2 5320 1 70
2 5321 1 70
2 5322 1 70
2 5323 1 70
2 5324 1 70
2 5325 1 70
2 5326 1 70
2 5327 1 70
2 5328 1 71
2 5329 1 71
2 5330 1 71
2 5331 1 71
2 5332 1 71
2 5333 1 71
2 5334 1 71
2 5335 1 71
2 5336 1 72
2 5337 1 72
2 5338 1 72
2 5339 1 72
2 5340 1 72
2 5341 1 72
2 5342 1 72
2 5343 1 72
2 5344 1 73
2 5345 1 73
2 5346 1 73
2 5347 1 73
2 5348 1 73
2 5349 1 73
2 5350 1 73
2 5351 1 73
2 5352 1 74
2 5353 1 74
2 5354 1 74
2 5355 1 74
2 5356 1 74
2 5357 1 74
2 5358 1 74
2 5359 1 74
2 5360 1 75
2 5361 1 75
2 5362 1 75
2 5363 1 75
2 5364 1 75
2 5365 1 75
2 5366 1 75
2 5367 1 75
2 5368 1 76
2 5369 1 76
2 5370 1 76
2 5371 1 76
2 5372 1 76
2 5373 1 76
2 5374 1 76
2 5375 1 76
2 5376 1 77
2 5377 1 77
2 5378 1 77
2 5379 1 77
2 5380 1 77
2 5381 1 77
2 5382 1 77
2 5383 1 77
2 5384 1 78
2 5385 1 78
2 5386 1 78
2 5387 1 78
2 5388 1 78
2 5389 1 78
2 5390 1 78
2 5391 1 78
2 5392 1 79
2 5393 1 79
2 5394 1 79
2 5395 1 79
2 5396 1 79
2 5397 1 79
2 5398 1 79
2 5399 1 79
2 5400 1 80
2 5401 1 80
2 5402 1 80
2 5403 1 80
2 5404 1 80
2 5405 1 80
2 5406 1 80
2 5407 1 80
2 5408 1 81
2 5409 1 81
2 5410 1 81
2 5411 1 81
2 5412 1 81
2 5413 1 81
2 5414 1 81
2 5415 1 81
2 5416 1 82
2 5417 1 82
2 5418 1 82
2 5419 1 82
2 5420 1 82
2 5421 1 82
2 5422 1 82
2 5423 1 83
2 5424 1 83
2 5425 1 83
2 5426 1 83
2 5427 1 83
2 5428 1 83
2 5429 1 83
2 5430 1 84
2 5431 1 84
2 5432 1 84
2 5433 1 84
2 5434 1 84
2 5435 1 84
2 5436 1 84
2 5437 1 85
2 5438 1 85
2 5439 1 85
2 5440 1 85
2 5441 1 85
2 5442 1 85
2 5443 1 85
2 5444 1 86
2 5445 1 86
2 5446 1 86
2 5447 1 86
2 5448 1 86
2 5449 1 86
2 5450 1 86
2 5451 1 87
2 5452 1 87
2 5453 1 87
2 5454 1 87
2 5455 1 87
2 5456 1 87
2 5457 1 87
2 5458 1 88
2 5459 1 88
2 5460 1 88
2 5461 1 88
2 5462 1 88
2 5463 1 88
2 5464 1 88
2 5465 1 89
2 5466 1 89
2 5467 1 89
2 5468 1 89
2 5469 1 89
2 5470 1 89
2 5471 1 89
2 5472 1 90
2 5473 1 90
2 5474 1 90
2 5475 1 90
2 5476 1 90
2 5477 1 90
2 5478 1 90
2 5479 1 91
2 5480 1 91
2 5481 1 91
2 5482 1 91
2 5483 1 91
2 5484 1 91
2 5485 1 91
2 5486 1 92
2 5487 1 92
2 5488 1 92
2 5489 1 92
2 5490 1 92
2 5491 1 92
2 5492 1 92
2 5493 1 93
2 5494 1 93
2 5495 1 93
2 5496 1 93
2 5497 1 93
2 5498 1 93
2 5499 1 93
2 5500 1 94
2 5501 1 94
2 5502 1 94
2 5503 1 94
2 5504 1 94
2 5505 1 94
2 5506 1 94
2 5507 1 94
2 5508 1 95
2 5509 1 95
2 5510 1 95
2 5511 1 95
2 5512 1 95
2 5513 1 95
2 5514 1 95
2 5515 1 96
2 5516 1 96
2 5517 1 96
2 5518 1 96
2 5519 1 96
2 5520 1 97
2 5521 1 97
2 5522 1 97
2 5523 1 97
2 5524 1 98
2 5525 1 98
2 5526 1 98
2 5527 1 98
2 5528 1 98
2 5529 1 98
2 5530 1 99
2 5531 1 99
2 5532 1 100
2 5533 1 100
2 5534 1 104
2 5535 1 104
2 5536 1 105
2 5537 1 105
2 5538 1 108
2 5539 1 108
2 5540 1 110
2 5541 1 110
2 5542 1 112
2 5543 1 112
2 5544 1 113
2 5545 1 113
2 5546 1 113
2 5547 1 118
2 5548 1 118
2 5549 1 119
2 5550 1 119
2 5551 1 120
2 5552 1 120
2 5553 1 120
2 5554 1 122
2 5555 1 122
2 5556 1 123
2 5557 1 123
2 5558 1 125
2 5559 1 125
2 5560 1 129
2 5561 1 129
2 5562 1 130
2 5563 1 130
2 5564 1 131
2 5565 1 131
2 5566 1 132
2 5567 1 132
2 5568 1 134
2 5569 1 134
2 5570 1 139
2 5571 1 139
2 5572 1 142
2 5573 1 142
2 5574 1 145
2 5575 1 145
2 5576 1 145
2 5577 1 147
2 5578 1 147
2 5579 1 148
2 5580 1 148
2 5581 1 149
2 5582 1 149
2 5583 1 151
2 5584 1 151
2 5585 1 156
2 5586 1 156
2 5587 1 156
2 5588 1 158
2 5589 1 158
2 5590 1 159
2 5591 1 159
2 5592 1 161
2 5593 1 161
2 5594 1 164
2 5595 1 164
2 5596 1 164
2 5597 1 171
2 5598 1 171
2 5599 1 176
2 5600 1 176
2 5601 1 178
2 5602 1 178
2 5603 1 179
2 5604 1 179
2 5605 1 180
2 5606 1 180
2 5607 1 182
2 5608 1 182
2 5609 1 187
2 5610 1 187
2 5611 1 187
2 5612 1 189
2 5613 1 189
2 5614 1 190
2 5615 1 190
2 5616 1 192
2 5617 1 192
2 5618 1 196
2 5619 1 196
2 5620 1 201
2 5621 1 201
2 5622 1 201
2 5623 1 203
2 5624 1 203
2 5625 1 212
2 5626 1 212
2 5627 1 214
2 5628 1 214
2 5629 1 215
2 5630 1 215
2 5631 1 217
2 5632 1 217
2 5633 1 222
2 5634 1 222
2 5635 1 222
2 5636 1 224
2 5637 1 224
2 5638 1 225
2 5639 1 225
2 5640 1 227
2 5641 1 227
2 5642 1 232
2 5643 1 232
2 5644 1 235
2 5645 1 235
2 5646 1 238
2 5647 1 238
2 5648 1 238
2 5649 1 240
2 5650 1 240
2 5651 1 241
2 5652 1 241
2 5653 1 242
2 5654 1 242
2 5655 1 244
2 5656 1 244
2 5657 1 249
2 5658 1 249
2 5659 1 249
2 5660 1 251
2 5661 1 251
2 5662 1 252
2 5663 1 252
2 5664 1 254
2 5665 1 254
2 5666 1 257
2 5667 1 257
2 5668 1 257
2 5669 1 264
2 5670 1 264
2 5671 1 269
2 5672 1 269
2 5673 1 271
2 5674 1 271
2 5675 1 272
2 5676 1 272
2 5677 1 273
2 5678 1 273
2 5679 1 275
2 5680 1 275
2 5681 1 280
2 5682 1 280
2 5683 1 280
2 5684 1 282
2 5685 1 282
2 5686 1 283
2 5687 1 283
2 5688 1 285
2 5689 1 285
2 5690 1 289
2 5691 1 289
2 5692 1 294
2 5693 1 294
2 5694 1 294
2 5695 1 296
2 5696 1 296
2 5697 1 305
2 5698 1 305
2 5699 1 307
2 5700 1 307
2 5701 1 308
2 5702 1 308
2 5703 1 310
2 5704 1 310
2 5705 1 315
2 5706 1 315
2 5707 1 315
2 5708 1 317
2 5709 1 317
2 5710 1 318
2 5711 1 318
2 5712 1 320
2 5713 1 320
2 5714 1 325
2 5715 1 325
2 5716 1 328
2 5717 1 328
2 5718 1 331
2 5719 1 331
2 5720 1 331
2 5721 1 333
2 5722 1 333
2 5723 1 334
2 5724 1 334
2 5725 1 335
2 5726 1 335
2 5727 1 337
2 5728 1 337
2 5729 1 342
2 5730 1 342
2 5731 1 342
2 5732 1 344
2 5733 1 344
2 5734 1 345
2 5735 1 345
2 5736 1 347
2 5737 1 347
2 5738 1 350
2 5739 1 350
2 5740 1 350
2 5741 1 357
2 5742 1 357
2 5743 1 362
2 5744 1 362
2 5745 1 364
2 5746 1 364
2 5747 1 365
2 5748 1 365
2 5749 1 366
2 5750 1 366
2 5751 1 368
2 5752 1 368
2 5753 1 373
2 5754 1 373
2 5755 1 373
2 5756 1 375
2 5757 1 375
2 5758 1 376
2 5759 1 376
2 5760 1 378
2 5761 1 378
2 5762 1 382
2 5763 1 382
2 5764 1 387
2 5765 1 387
2 5766 1 387
2 5767 1 389
2 5768 1 389
2 5769 1 398
2 5770 1 398
2 5771 1 400
2 5772 1 400
2 5773 1 401
2 5774 1 401
2 5775 1 403
2 5776 1 403
2 5777 1 408
2 5778 1 408
2 5779 1 408
2 5780 1 410
2 5781 1 410
2 5782 1 411
2 5783 1 411
2 5784 1 413
2 5785 1 413
2 5786 1 418
2 5787 1 418
2 5788 1 421
2 5789 1 421
2 5790 1 424
2 5791 1 424
2 5792 1 424
2 5793 1 426
2 5794 1 426
2 5795 1 427
2 5796 1 427
2 5797 1 428
2 5798 1 428
2 5799 1 430
2 5800 1 430
2 5801 1 435
2 5802 1 435
2 5803 1 435
2 5804 1 437
2 5805 1 437
2 5806 1 438
2 5807 1 438
2 5808 1 440
2 5809 1 440
2 5810 1 443
2 5811 1 443
2 5812 1 443
2 5813 1 450
2 5814 1 450
2 5815 1 455
2 5816 1 455
2 5817 1 457
2 5818 1 457
2 5819 1 458
2 5820 1 458
2 5821 1 459
2 5822 1 459
2 5823 1 461
2 5824 1 461
2 5825 1 466
2 5826 1 466
2 5827 1 466
2 5828 1 468
2 5829 1 468
2 5830 1 469
2 5831 1 469
2 5832 1 471
2 5833 1 471
2 5834 1 475
2 5835 1 475
2 5836 1 480
2 5837 1 480
2 5838 1 480
2 5839 1 482
2 5840 1 482
2 5841 1 491
2 5842 1 491
2 5843 1 493
2 5844 1 493
2 5845 1 494
2 5846 1 494
2 5847 1 496
2 5848 1 496
2 5849 1 501
2 5850 1 501
2 5851 1 501
2 5852 1 503
2 5853 1 503
2 5854 1 504
2 5855 1 504
2 5856 1 506
2 5857 1 506
2 5858 1 511
2 5859 1 511
2 5860 1 514
2 5861 1 514
2 5862 1 517
2 5863 1 517
2 5864 1 517
2 5865 1 519
2 5866 1 519
2 5867 1 520
2 5868 1 520
2 5869 1 521
2 5870 1 521
2 5871 1 523
2 5872 1 523
2 5873 1 528
2 5874 1 528
2 5875 1 528
2 5876 1 530
2 5877 1 530
2 5878 1 531
2 5879 1 531
2 5880 1 533
2 5881 1 533
2 5882 1 536
2 5883 1 536
2 5884 1 536
2 5885 1 543
2 5886 1 543
2 5887 1 548
2 5888 1 548
2 5889 1 550
2 5890 1 550
2 5891 1 551
2 5892 1 551
2 5893 1 552
2 5894 1 552
2 5895 1 554
2 5896 1 554
2 5897 1 559
2 5898 1 559
2 5899 1 559
2 5900 1 561
2 5901 1 561
2 5902 1 562
2 5903 1 562
2 5904 1 564
2 5905 1 564
2 5906 1 568
2 5907 1 568
2 5908 1 573
2 5909 1 573
2 5910 1 573
2 5911 1 575
2 5912 1 575
2 5913 1 584
2 5914 1 584
2 5915 1 586
2 5916 1 586
2 5917 1 587
2 5918 1 587
2 5919 1 589
2 5920 1 589
2 5921 1 594
2 5922 1 594
2 5923 1 594
2 5924 1 596
2 5925 1 596
2 5926 1 597
2 5927 1 597
2 5928 1 599
2 5929 1 599
2 5930 1 604
2 5931 1 604
2 5932 1 607
2 5933 1 607
2 5934 1 610
2 5935 1 610
2 5936 1 610
2 5937 1 612
2 5938 1 612
2 5939 1 613
2 5940 1 613
2 5941 1 614
2 5942 1 614
2 5943 1 616
2 5944 1 616
2 5945 1 621
2 5946 1 621
2 5947 1 621
2 5948 1 623
2 5949 1 623
2 5950 1 624
2 5951 1 624
2 5952 1 626
2 5953 1 626
2 5954 1 629
2 5955 1 629
2 5956 1 629
2 5957 1 636
2 5958 1 636
2 5959 1 641
2 5960 1 641
2 5961 1 643
2 5962 1 643
2 5963 1 644
2 5964 1 644
2 5965 1 645
2 5966 1 645
2 5967 1 647
2 5968 1 647
2 5969 1 652
2 5970 1 652
2 5971 1 652
2 5972 1 654
2 5973 1 654
2 5974 1 655
2 5975 1 655
2 5976 1 657
2 5977 1 657
2 5978 1 661
2 5979 1 661
2 5980 1 666
2 5981 1 666
2 5982 1 666
2 5983 1 668
2 5984 1 668
2 5985 1 677
2 5986 1 677
2 5987 1 679
2 5988 1 679
2 5989 1 680
2 5990 1 680
2 5991 1 682
2 5992 1 682
2 5993 1 687
2 5994 1 687
2 5995 1 687
2 5996 1 689
2 5997 1 689
2 5998 1 690
2 5999 1 690
2 6000 1 692
2 6001 1 692
2 6002 1 697
2 6003 1 697
2 6004 1 700
2 6005 1 700
2 6006 1 703
2 6007 1 703
2 6008 1 703
2 6009 1 705
2 6010 1 705
2 6011 1 706
2 6012 1 706
2 6013 1 707
2 6014 1 707
2 6015 1 709
2 6016 1 709
2 6017 1 714
2 6018 1 714
2 6019 1 714
2 6020 1 716
2 6021 1 716
2 6022 1 717
2 6023 1 717
2 6024 1 719
2 6025 1 719
2 6026 1 722
2 6027 1 722
2 6028 1 722
2 6029 1 729
2 6030 1 729
2 6031 1 734
2 6032 1 734
2 6033 1 736
2 6034 1 736
2 6035 1 737
2 6036 1 737
2 6037 1 738
2 6038 1 738
2 6039 1 740
2 6040 1 740
2 6041 1 745
2 6042 1 745
2 6043 1 745
2 6044 1 747
2 6045 1 747
2 6046 1 748
2 6047 1 748
2 6048 1 750
2 6049 1 750
2 6050 1 754
2 6051 1 754
2 6052 1 759
2 6053 1 759
2 6054 1 759
2 6055 1 761
2 6056 1 761
2 6057 1 770
2 6058 1 770
2 6059 1 772
2 6060 1 772
2 6061 1 773
2 6062 1 773
2 6063 1 775
2 6064 1 775
2 6065 1 780
2 6066 1 780
2 6067 1 780
2 6068 1 782
2 6069 1 782
2 6070 1 783
2 6071 1 783
2 6072 1 785
2 6073 1 785
2 6074 1 790
2 6075 1 790
2 6076 1 793
2 6077 1 793
2 6078 1 796
2 6079 1 796
2 6080 1 796
2 6081 1 798
2 6082 1 798
2 6083 1 799
2 6084 1 799
2 6085 1 800
2 6086 1 800
2 6087 1 802
2 6088 1 802
2 6089 1 807
2 6090 1 807
2 6091 1 807
2 6092 1 809
2 6093 1 809
2 6094 1 810
2 6095 1 810
2 6096 1 812
2 6097 1 812
2 6098 1 815
2 6099 1 815
2 6100 1 815
2 6101 1 822
2 6102 1 822
2 6103 1 827
2 6104 1 827
2 6105 1 829
2 6106 1 829
2 6107 1 830
2 6108 1 830
2 6109 1 831
2 6110 1 831
2 6111 1 833
2 6112 1 833
2 6113 1 838
2 6114 1 838
2 6115 1 838
2 6116 1 840
2 6117 1 840
2 6118 1 841
2 6119 1 841
2 6120 1 843
2 6121 1 843
2 6122 1 847
2 6123 1 847
2 6124 1 852
2 6125 1 852
2 6126 1 852
2 6127 1 854
2 6128 1 854
2 6129 1 863
2 6130 1 863
2 6131 1 865
2 6132 1 865
2 6133 1 866
2 6134 1 866
2 6135 1 868
2 6136 1 868
2 6137 1 873
2 6138 1 873
2 6139 1 873
2 6140 1 875
2 6141 1 875
2 6142 1 876
2 6143 1 876
2 6144 1 878
2 6145 1 878
2 6146 1 883
2 6147 1 883
2 6148 1 886
2 6149 1 886
2 6150 1 889
2 6151 1 889
2 6152 1 889
2 6153 1 891
2 6154 1 891
2 6155 1 892
2 6156 1 892
2 6157 1 893
2 6158 1 893
2 6159 1 895
2 6160 1 895
2 6161 1 900
2 6162 1 900
2 6163 1 900
2 6164 1 902
2 6165 1 902
2 6166 1 903
2 6167 1 903
2 6168 1 905
2 6169 1 905
2 6170 1 908
2 6171 1 908
2 6172 1 908
2 6173 1 915
2 6174 1 915
2 6175 1 920
2 6176 1 920
2 6177 1 922
2 6178 1 922
2 6179 1 923
2 6180 1 923
2 6181 1 924
2 6182 1 924
2 6183 1 926
2 6184 1 926
2 6185 1 931
2 6186 1 931
2 6187 1 931
2 6188 1 933
2 6189 1 933
2 6190 1 934
2 6191 1 934
2 6192 1 936
2 6193 1 936
2 6194 1 940
2 6195 1 940
2 6196 1 945
2 6197 1 945
2 6198 1 945
2 6199 1 947
2 6200 1 947
2 6201 1 956
2 6202 1 956
2 6203 1 958
2 6204 1 958
2 6205 1 959
2 6206 1 959
2 6207 1 961
2 6208 1 961
2 6209 1 966
2 6210 1 966
2 6211 1 966
2 6212 1 968
2 6213 1 968
2 6214 1 969
2 6215 1 969
2 6216 1 971
2 6217 1 971
2 6218 1 976
2 6219 1 976
2 6220 1 979
2 6221 1 979
2 6222 1 982
2 6223 1 982
2 6224 1 982
2 6225 1 984
2 6226 1 984
2 6227 1 985
2 6228 1 985
2 6229 1 986
2 6230 1 986
2 6231 1 988
2 6232 1 988
2 6233 1 993
2 6234 1 993
2 6235 1 993
2 6236 1 995
2 6237 1 995
2 6238 1 996
2 6239 1 996
2 6240 1 998
2 6241 1 998
2 6242 1 1001
2 6243 1 1001
2 6244 1 1001
2 6245 1 1008
2 6246 1 1008
2 6247 1 1013
2 6248 1 1013
2 6249 1 1015
2 6250 1 1015
2 6251 1 1016
2 6252 1 1016
2 6253 1 1017
2 6254 1 1017
2 6255 1 1019
2 6256 1 1019
2 6257 1 1024
2 6258 1 1024
2 6259 1 1024
2 6260 1 1026
2 6261 1 1026
2 6262 1 1027
2 6263 1 1027
2 6264 1 1029
2 6265 1 1029
2 6266 1 1033
2 6267 1 1033
2 6268 1 1038
2 6269 1 1038
2 6270 1 1038
2 6271 1 1040
2 6272 1 1040
2 6273 1 1049
2 6274 1 1049
2 6275 1 1051
2 6276 1 1051
2 6277 1 1052
2 6278 1 1052
2 6279 1 1054
2 6280 1 1054
2 6281 1 1059
2 6282 1 1059
2 6283 1 1059
2 6284 1 1061
2 6285 1 1061
2 6286 1 1062
2 6287 1 1062
2 6288 1 1064
2 6289 1 1064
2 6290 1 1069
2 6291 1 1069
2 6292 1 1072
2 6293 1 1072
2 6294 1 1075
2 6295 1 1075
2 6296 1 1075
2 6297 1 1077
2 6298 1 1077
2 6299 1 1078
2 6300 1 1078
2 6301 1 1079
2 6302 1 1079
2 6303 1 1081
2 6304 1 1081
2 6305 1 1086
2 6306 1 1086
2 6307 1 1086
2 6308 1 1088
2 6309 1 1088
2 6310 1 1089
2 6311 1 1089
2 6312 1 1091
2 6313 1 1091
2 6314 1 1094
2 6315 1 1094
2 6316 1 1094
2 6317 1 1101
2 6318 1 1101
2 6319 1 1106
2 6320 1 1106
2 6321 1 1108
2 6322 1 1108
2 6323 1 1109
2 6324 1 1109
2 6325 1 1110
2 6326 1 1110
2 6327 1 1112
2 6328 1 1112
2 6329 1 1117
2 6330 1 1117
2 6331 1 1117
2 6332 1 1119
2 6333 1 1119
2 6334 1 1120
2 6335 1 1120
2 6336 1 1122
2 6337 1 1122
2 6338 1 1126
2 6339 1 1126
2 6340 1 1131
2 6341 1 1131
2 6342 1 1131
2 6343 1 1133
2 6344 1 1133
2 6345 1 1142
2 6346 1 1142
2 6347 1 1144
2 6348 1 1144
2 6349 1 1145
2 6350 1 1145
2 6351 1 1147
2 6352 1 1147
2 6353 1 1152
2 6354 1 1152
2 6355 1 1152
2 6356 1 1154
2 6357 1 1154
2 6358 1 1155
2 6359 1 1155
2 6360 1 1157
2 6361 1 1157
2 6362 1 1162
2 6363 1 1162
2 6364 1 1165
2 6365 1 1165
2 6366 1 1168
2 6367 1 1168
2 6368 1 1168
2 6369 1 1170
2 6370 1 1170
2 6371 1 1171
2 6372 1 1171
2 6373 1 1172
2 6374 1 1172
2 6375 1 1174
2 6376 1 1174
2 6377 1 1179
2 6378 1 1179
2 6379 1 1179
2 6380 1 1181
2 6381 1 1181
2 6382 1 1182
2 6383 1 1182
2 6384 1 1184
2 6385 1 1184
2 6386 1 1187
2 6387 1 1187
2 6388 1 1187
2 6389 1 1194
2 6390 1 1194
2 6391 1 1199
2 6392 1 1199
2 6393 1 1201
2 6394 1 1201
2 6395 1 1202
2 6396 1 1202
2 6397 1 1203
2 6398 1 1203
2 6399 1 1205
2 6400 1 1205
2 6401 1 1210
2 6402 1 1210
2 6403 1 1210
2 6404 1 1212
2 6405 1 1212
2 6406 1 1213
2 6407 1 1213
2 6408 1 1215
2 6409 1 1215
2 6410 1 1219
2 6411 1 1219
2 6412 1 1224
2 6413 1 1224
2 6414 1 1224
2 6415 1 1226
2 6416 1 1226
2 6417 1 1235
2 6418 1 1235
2 6419 1 1237
2 6420 1 1237
2 6421 1 1238
2 6422 1 1238
2 6423 1 1240
2 6424 1 1240
2 6425 1 1245
2 6426 1 1245
2 6427 1 1245
2 6428 1 1247
2 6429 1 1247
2 6430 1 1248
2 6431 1 1248
2 6432 1 1250
2 6433 1 1250
2 6434 1 1255
2 6435 1 1255
2 6436 1 1258
2 6437 1 1258
2 6438 1 1261
2 6439 1 1261
2 6440 1 1261
2 6441 1 1263
2 6442 1 1263
2 6443 1 1264
2 6444 1 1264
2 6445 1 1265
2 6446 1 1265
2 6447 1 1267
2 6448 1 1267
2 6449 1 1272
2 6450 1 1272
2 6451 1 1272
2 6452 1 1274
2 6453 1 1274
2 6454 1 1275
2 6455 1 1275
2 6456 1 1277
2 6457 1 1277
2 6458 1 1280
2 6459 1 1280
2 6460 1 1280
2 6461 1 1287
2 6462 1 1287
2 6463 1 1292
2 6464 1 1292
2 6465 1 1294
2 6466 1 1294
2 6467 1 1295
2 6468 1 1295
2 6469 1 1296
2 6470 1 1296
2 6471 1 1298
2 6472 1 1298
2 6473 1 1303
2 6474 1 1303
2 6475 1 1303
2 6476 1 1305
2 6477 1 1305
2 6478 1 1306
2 6479 1 1306
2 6480 1 1308
2 6481 1 1308
2 6482 1 1312
2 6483 1 1312
2 6484 1 1317
2 6485 1 1317
2 6486 1 1317
2 6487 1 1319
2 6488 1 1319
2 6489 1 1328
2 6490 1 1328
2 6491 1 1330
2 6492 1 1330
2 6493 1 1331
2 6494 1 1331
2 6495 1 1333
2 6496 1 1333
2 6497 1 1338
2 6498 1 1338
2 6499 1 1338
2 6500 1 1340
2 6501 1 1340
2 6502 1 1341
2 6503 1 1341
2 6504 1 1343
2 6505 1 1343
2 6506 1 1348
2 6507 1 1348
2 6508 1 1351
2 6509 1 1351
2 6510 1 1354
2 6511 1 1354
2 6512 1 1354
2 6513 1 1356
2 6514 1 1356
2 6515 1 1357
2 6516 1 1357
2 6517 1 1358
2 6518 1 1358
2 6519 1 1360
2 6520 1 1360
2 6521 1 1365
2 6522 1 1365
2 6523 1 1365
2 6524 1 1367
2 6525 1 1367
2 6526 1 1368
2 6527 1 1368
2 6528 1 1370
2 6529 1 1370
2 6530 1 1373
2 6531 1 1373
2 6532 1 1373
2 6533 1 1380
2 6534 1 1380
2 6535 1 1385
2 6536 1 1385
2 6537 1 1387
2 6538 1 1387
2 6539 1 1388
2 6540 1 1388
2 6541 1 1389
2 6542 1 1389
2 6543 1 1391
2 6544 1 1391
2 6545 1 1396
2 6546 1 1396
2 6547 1 1396
2 6548 1 1398
2 6549 1 1398
2 6550 1 1399
2 6551 1 1399
2 6552 1 1401
2 6553 1 1401
2 6554 1 1404
2 6555 1 1404
2 6556 1 1404
2 6557 1 1406
2 6558 1 1406
2 6559 1 1408
2 6560 1 1408
2 6561 1 1414
2 6562 1 1414
2 6563 1 1419
2 6564 1 1419
2 6565 1 1422
2 6566 1 1422
2 6567 1 1427
2 6568 1 1427
2 6569 1 1433
2 6570 1 1433
2 6571 1 1434
2 6572 1 1434
2 6573 1 1437
2 6574 1 1437
2 6575 1 1439
2 6576 1 1439
2 6577 1 1440
2 6578 1 1440
2 6579 1 1441
2 6580 1 1441
2 6581 1 1448
2 6582 1 1448
2 6583 1 1476
2 6584 1 1476
2 6585 1 1476
2 6586 1 1479
2 6587 1 1479
2 6588 1 1482
2 6589 1 1482
2 6590 1 1486
2 6591 1 1486
2 6592 1 1487
2 6593 1 1487
2 6594 1 1488
2 6595 1 1488
2 6596 1 1488
2 6597 1 1488
2 6598 1 1491
2 6599 1 1491
2 6600 1 1498
2 6601 1 1498
2 6602 1 1502
2 6603 1 1502
2 6604 1 1503
2 6605 1 1503
2 6606 1 1511
2 6607 1 1511
2 6608 1 1514
2 6609 1 1514
2 6610 1 1515
2 6611 1 1515
2 6612 1 1518
2 6613 1 1518
2 6614 1 1518
2 6615 1 1520
2 6616 1 1520
2 6617 1 1522
2 6618 1 1522
2 6619 1 1524
2 6620 1 1524
2 6621 1 1531
2 6622 1 1531
2 6623 1 1532
2 6624 1 1532
2 6625 1 1538
2 6626 1 1538
2 6627 1 1541
2 6628 1 1541
2 6629 1 1542
2 6630 1 1542
2 6631 1 1547
2 6632 1 1547
2 6633 1 1551
2 6634 1 1551
2 6635 1 1551
2 6636 1 1551
2 6637 1 1555
2 6638 1 1555
2 6639 1 1558
2 6640 1 1558
2 6641 1 1559
2 6642 1 1559
2 6643 1 1562
2 6644 1 1562
2 6645 1 1562
2 6646 1 1565
2 6647 1 1565
2 6648 1 1569
2 6649 1 1569
2 6650 1 1570
2 6651 1 1570
2 6652 1 1572
2 6653 1 1572
2 6654 1 1574
2 6655 1 1574
2 6656 1 1576
2 6657 1 1576
2 6658 1 1579
2 6659 1 1579
2 6660 1 1579
2 6661 1 1579
2 6662 1 1581
2 6663 1 1581
2 6664 1 1583
2 6665 1 1583
2 6666 1 1587
2 6667 1 1587
2 6668 1 1596
2 6669 1 1596
2 6670 1 1597
2 6671 1 1597
2 6672 1 1603
2 6673 1 1603
2 6674 1 1606
2 6675 1 1606
2 6676 1 1607
2 6677 1 1607
2 6678 1 1610
2 6679 1 1610
2 6680 1 1612
2 6681 1 1612
2 6682 1 1614
2 6683 1 1614
2 6684 1 1616
2 6685 1 1616
2 6686 1 1618
2 6687 1 1618
2 6688 1 1621
2 6689 1 1621
2 6690 1 1621
2 6691 1 1621
2 6692 1 1626
2 6693 1 1626
2 6694 1 1627
2 6695 1 1627
2 6696 1 1631
2 6697 1 1631
2 6698 1 1640
2 6699 1 1640
2 6700 1 1643
2 6701 1 1643
2 6702 1 1644
2 6703 1 1644
2 6704 1 1647
2 6705 1 1647
2 6706 1 1647
2 6707 1 1649
2 6708 1 1649
2 6709 1 1651
2 6710 1 1651
2 6711 1 1653
2 6712 1 1653
2 6713 1 1660
2 6714 1 1660
2 6715 1 1661
2 6716 1 1661
2 6717 1 1667
2 6718 1 1667
2 6719 1 1670
2 6720 1 1670
2 6721 1 1671
2 6722 1 1671
2 6723 1 1676
2 6724 1 1676
2 6725 1 1680
2 6726 1 1680
2 6727 1 1680
2 6728 1 1680
2 6729 1 1684
2 6730 1 1684
2 6731 1 1687
2 6732 1 1687
2 6733 1 1688
2 6734 1 1688
2 6735 1 1691
2 6736 1 1691
2 6737 1 1691
2 6738 1 1694
2 6739 1 1694
2 6740 1 1698
2 6741 1 1698
2 6742 1 1699
2 6743 1 1699
2 6744 1 1701
2 6745 1 1701
2 6746 1 1703
2 6747 1 1703
2 6748 1 1705
2 6749 1 1705
2 6750 1 1708
2 6751 1 1708
2 6752 1 1708
2 6753 1 1708
2 6754 1 1710
2 6755 1 1710
2 6756 1 1712
2 6757 1 1712
2 6758 1 1716
2 6759 1 1716
2 6760 1 1725
2 6761 1 1725
2 6762 1 1726
2 6763 1 1726
2 6764 1 1732
2 6765 1 1732
2 6766 1 1735
2 6767 1 1735
2 6768 1 1736
2 6769 1 1736
2 6770 1 1739
2 6771 1 1739
2 6772 1 1741
2 6773 1 1741
2 6774 1 1743
2 6775 1 1743
2 6776 1 1745
2 6777 1 1745
2 6778 1 1747
2 6779 1 1747
2 6780 1 1750
2 6781 1 1750
2 6782 1 1750
2 6783 1 1750
2 6784 1 1755
2 6785 1 1755
2 6786 1 1756
2 6787 1 1756
2 6788 1 1760
2 6789 1 1760
2 6790 1 1769
2 6791 1 1769
2 6792 1 1772
2 6793 1 1772
2 6794 1 1773
2 6795 1 1773
2 6796 1 1776
2 6797 1 1776
2 6798 1 1776
2 6799 1 1778
2 6800 1 1778
2 6801 1 1780
2 6802 1 1780
2 6803 1 1782
2 6804 1 1782
2 6805 1 1789
2 6806 1 1789
2 6807 1 1790
2 6808 1 1790
2 6809 1 1796
2 6810 1 1796
2 6811 1 1799
2 6812 1 1799
2 6813 1 1800
2 6814 1 1800
2 6815 1 1805
2 6816 1 1805
2 6817 1 1809
2 6818 1 1809
2 6819 1 1809
2 6820 1 1809
2 6821 1 1813
2 6822 1 1813
2 6823 1 1816
2 6824 1 1816
2 6825 1 1817
2 6826 1 1817
2 6827 1 1820
2 6828 1 1820
2 6829 1 1820
2 6830 1 1823
2 6831 1 1823
2 6832 1 1827
2 6833 1 1827
2 6834 1 1828
2 6835 1 1828
2 6836 1 1830
2 6837 1 1830
2 6838 1 1832
2 6839 1 1832
2 6840 1 1834
2 6841 1 1834
2 6842 1 1837
2 6843 1 1837
2 6844 1 1837
2 6845 1 1837
2 6846 1 1839
2 6847 1 1839
2 6848 1 1841
2 6849 1 1841
2 6850 1 1845
2 6851 1 1845
2 6852 1 1854
2 6853 1 1854
2 6854 1 1855
2 6855 1 1855
2 6856 1 1861
2 6857 1 1861
2 6858 1 1864
2 6859 1 1864
2 6860 1 1865
2 6861 1 1865
2 6862 1 1868
2 6863 1 1868
2 6864 1 1870
2 6865 1 1870
2 6866 1 1872
2 6867 1 1872
2 6868 1 1874
2 6869 1 1874
2 6870 1 1876
2 6871 1 1876
2 6872 1 1879
2 6873 1 1879
2 6874 1 1879
2 6875 1 1879
2 6876 1 1884
2 6877 1 1884
2 6878 1 1885
2 6879 1 1885
2 6880 1 1889
2 6881 1 1889
2 6882 1 1898
2 6883 1 1898
2 6884 1 1901
2 6885 1 1901
2 6886 1 1902
2 6887 1 1902
2 6888 1 1905
2 6889 1 1905
2 6890 1 1905
2 6891 1 1907
2 6892 1 1907
2 6893 1 1909
2 6894 1 1909
2 6895 1 1911
2 6896 1 1911
2 6897 1 1918
2 6898 1 1918
2 6899 1 1919
2 6900 1 1919
2 6901 1 1925
2 6902 1 1925
2 6903 1 1928
2 6904 1 1928
2 6905 1 1929
2 6906 1 1929
2 6907 1 1934
2 6908 1 1934
2 6909 1 1938
2 6910 1 1938
2 6911 1 1938
2 6912 1 1938
2 6913 1 1942
2 6914 1 1942
2 6915 1 1945
2 6916 1 1945
2 6917 1 1946
2 6918 1 1946
2 6919 1 1949
2 6920 1 1949
2 6921 1 1949
2 6922 1 1952
2 6923 1 1952
2 6924 1 1956
2 6925 1 1956
2 6926 1 1957
2 6927 1 1957
2 6928 1 1959
2 6929 1 1959
2 6930 1 1961
2 6931 1 1961
2 6932 1 1963
2 6933 1 1963
2 6934 1 1966
2 6935 1 1966
2 6936 1 1966
2 6937 1 1966
2 6938 1 1968
2 6939 1 1968
2 6940 1 1970
2 6941 1 1970
2 6942 1 1974
2 6943 1 1974
2 6944 1 1983
2 6945 1 1983
2 6946 1 1984
2 6947 1 1984
2 6948 1 1990
2 6949 1 1990
2 6950 1 1993
2 6951 1 1993
2 6952 1 1994
2 6953 1 1994
2 6954 1 1997
2 6955 1 1997
2 6956 1 1999
2 6957 1 1999
2 6958 1 2001
2 6959 1 2001
2 6960 1 2003
2 6961 1 2003
2 6962 1 2005
2 6963 1 2005
2 6964 1 2008
2 6965 1 2008
2 6966 1 2008
2 6967 1 2008
2 6968 1 2013
2 6969 1 2013
2 6970 1 2014
2 6971 1 2014
2 6972 1 2018
2 6973 1 2018
2 6974 1 2027
2 6975 1 2027
2 6976 1 2030
2 6977 1 2030
2 6978 1 2031
2 6979 1 2031
2 6980 1 2034
2 6981 1 2034
2 6982 1 2034
2 6983 1 2036
2 6984 1 2036
2 6985 1 2038
2 6986 1 2038
2 6987 1 2040
2 6988 1 2040
2 6989 1 2047
2 6990 1 2047
2 6991 1 2048
2 6992 1 2048
2 6993 1 2054
2 6994 1 2054
2 6995 1 2057
2 6996 1 2057
2 6997 1 2058
2 6998 1 2058
2 6999 1 2063
2 7000 1 2063
2 7001 1 2067
2 7002 1 2067
2 7003 1 2067
2 7004 1 2067
2 7005 1 2071
2 7006 1 2071
2 7007 1 2074
2 7008 1 2074
2 7009 1 2075
2 7010 1 2075
2 7011 1 2078
2 7012 1 2078
2 7013 1 2078
2 7014 1 2081
2 7015 1 2081
2 7016 1 2085
2 7017 1 2085
2 7018 1 2086
2 7019 1 2086
2 7020 1 2088
2 7021 1 2088
2 7022 1 2090
2 7023 1 2090
2 7024 1 2092
2 7025 1 2092
2 7026 1 2095
2 7027 1 2095
2 7028 1 2095
2 7029 1 2095
2 7030 1 2097
2 7031 1 2097
2 7032 1 2099
2 7033 1 2099
2 7034 1 2103
2 7035 1 2103
2 7036 1 2112
2 7037 1 2112
2 7038 1 2113
2 7039 1 2113
2 7040 1 2119
2 7041 1 2119
2 7042 1 2122
2 7043 1 2122
2 7044 1 2123
2 7045 1 2123
2 7046 1 2126
2 7047 1 2126
2 7048 1 2128
2 7049 1 2128
2 7050 1 2130
2 7051 1 2130
2 7052 1 2132
2 7053 1 2132
2 7054 1 2134
2 7055 1 2134
2 7056 1 2137
2 7057 1 2137
2 7058 1 2137
2 7059 1 2137
2 7060 1 2142
2 7061 1 2142
2 7062 1 2143
2 7063 1 2143
2 7064 1 2147
2 7065 1 2147
2 7066 1 2156
2 7067 1 2156
2 7068 1 2159
2 7069 1 2159
2 7070 1 2160
2 7071 1 2160
2 7072 1 2163
2 7073 1 2163
2 7074 1 2163
2 7075 1 2165
2 7076 1 2165
2 7077 1 2167
2 7078 1 2167
2 7079 1 2169
2 7080 1 2169
2 7081 1 2176
2 7082 1 2176
2 7083 1 2177
2 7084 1 2177
2 7085 1 2183
2 7086 1 2183
2 7087 1 2186
2 7088 1 2186
2 7089 1 2187
2 7090 1 2187
2 7091 1 2192
2 7092 1 2192
2 7093 1 2196
2 7094 1 2196
2 7095 1 2196
2 7096 1 2196
2 7097 1 2200
2 7098 1 2200
2 7099 1 2203
2 7100 1 2203
2 7101 1 2204
2 7102 1 2204
2 7103 1 2207
2 7104 1 2207
2 7105 1 2207
2 7106 1 2210
2 7107 1 2210
2 7108 1 2214
2 7109 1 2214
2 7110 1 2215
2 7111 1 2215
2 7112 1 2217
2 7113 1 2217
2 7114 1 2219
2 7115 1 2219
2 7116 1 2221
2 7117 1 2221
2 7118 1 2224
2 7119 1 2224
2 7120 1 2224
2 7121 1 2224
2 7122 1 2226
2 7123 1 2226
2 7124 1 2228
2 7125 1 2228
2 7126 1 2232
2 7127 1 2232
2 7128 1 2241
2 7129 1 2241
2 7130 1 2242
2 7131 1 2242
2 7132 1 2248
2 7133 1 2248
2 7134 1 2251
2 7135 1 2251
2 7136 1 2252
2 7137 1 2252
2 7138 1 2255
2 7139 1 2255
2 7140 1 2257
2 7141 1 2257
2 7142 1 2259
2 7143 1 2259
2 7144 1 2261
2 7145 1 2261
2 7146 1 2263
2 7147 1 2263
2 7148 1 2266
2 7149 1 2266
2 7150 1 2266
2 7151 1 2266
2 7152 1 2271
2 7153 1 2271
2 7154 1 2272
2 7155 1 2272
2 7156 1 2276
2 7157 1 2276
2 7158 1 2285
2 7159 1 2285
2 7160 1 2288
2 7161 1 2288
2 7162 1 2289
2 7163 1 2289
2 7164 1 2292
2 7165 1 2292
2 7166 1 2292
2 7167 1 2294
2 7168 1 2294
2 7169 1 2296
2 7170 1 2296
2 7171 1 2298
2 7172 1 2298
2 7173 1 2305
2 7174 1 2305
2 7175 1 2306
2 7176 1 2306
2 7177 1 2312
2 7178 1 2312
2 7179 1 2315
2 7180 1 2315
2 7181 1 2316
2 7182 1 2316
2 7183 1 2321
2 7184 1 2321
2 7185 1 2325
2 7186 1 2325
2 7187 1 2325
2 7188 1 2325
2 7189 1 2329
2 7190 1 2329
2 7191 1 2332
2 7192 1 2332
2 7193 1 2333
2 7194 1 2333
2 7195 1 2336
2 7196 1 2336
2 7197 1 2336
2 7198 1 2339
2 7199 1 2339
2 7200 1 2343
2 7201 1 2343
2 7202 1 2344
2 7203 1 2344
2 7204 1 2346
2 7205 1 2346
2 7206 1 2348
2 7207 1 2348
2 7208 1 2350
2 7209 1 2350
2 7210 1 2353
2 7211 1 2353
2 7212 1 2353
2 7213 1 2353
2 7214 1 2355
2 7215 1 2355
2 7216 1 2357
2 7217 1 2357
2 7218 1 2359
2 7219 1 2359
2 7220 1 2366
2 7221 1 2366
2 7222 1 2367
2 7223 1 2367
2 7224 1 2370
2 7225 1 2370
2 7226 1 2371
2 7227 1 2371
2 7228 1 2374
2 7229 1 2374
2 7230 1 2385
2 7231 1 2385
2 7232 1 2386
2 7233 1 2386
2 7234 1 2388
2 7235 1 2388
2 7236 1 2390
2 7237 1 2390
2 7238 1 2392
2 7239 1 2392
2 7240 1 2396
2 7241 1 2396
2 7242 1 2397
2 7243 1 2397
2 7244 1 2401
2 7245 1 2401
2 7246 1 2401
2 7247 1 2401
2 7248 1 2405
2 7249 1 2405
2 7250 1 2414
2 7251 1 2414
2 7252 1 2417
2 7253 1 2417
2 7254 1 2418
2 7255 1 2418
2 7256 1 2421
2 7257 1 2421
2 7258 1 2421
2 7259 1 2424
2 7260 1 2424
2 7261 1 2427
2 7262 1 2427
2 7263 1 2428
2 7264 1 2428
2 7265 1 2429
2 7266 1 2429
2 7267 1 2431
2 7268 1 2431
2 7269 1 2434
2 7270 1 2434
2 7271 1 2435
2 7272 1 2435
2 7273 1 2440
2 7274 1 2440
2 7275 1 2458
2 7276 1 2458
2 7277 1 2469
2 7278 1 2469
2 7279 1 2470
2 7280 1 2470
2 7281 1 2475
2 7282 1 2475
2 7283 1 2478
2 7284 1 2478
2 7285 1 2481
2 7286 1 2481
2 7287 1 2483
2 7288 1 2483
2 7289 1 2484
2 7290 1 2484
2 7291 1 2489
2 7292 1 2489
2 7293 1 2492
2 7294 1 2492
2 7295 1 2497
2 7296 1 2497
2 7297 1 2498
2 7298 1 2498
2 7299 1 2499
2 7300 1 2499
2 7301 1 2502
2 7302 1 2502
2 7303 1 2505
2 7304 1 2505
2 7305 1 2507
2 7306 1 2507
2 7307 1 2508
2 7308 1 2508
2 7309 1 2513
2 7310 1 2513
2 7311 1 2516
2 7312 1 2516
2 7313 1 2521
2 7314 1 2521
2 7315 1 2521
2 7316 1 2527
2 7317 1 2527
2 7318 1 2527
2 7319 1 2529
2 7320 1 2529
2 7321 1 2532
2 7322 1 2532
2 7323 1 2535
2 7324 1 2535
2 7325 1 2537
2 7326 1 2537
2 7327 1 2538
2 7328 1 2538
2 7329 1 2543
2 7330 1 2543
2 7331 1 2546
2 7332 1 2546
2 7333 1 2547
2 7334 1 2547
2 7335 1 2550
2 7336 1 2550
2 7337 1 2553
2 7338 1 2553
2 7339 1 2555
2 7340 1 2555
2 7341 1 2556
2 7342 1 2556
2 7343 1 2561
2 7344 1 2561
2 7345 1 2564
2 7346 1 2564
2 7347 1 2569
2 7348 1 2569
2 7349 1 2569
2 7350 1 2575
2 7351 1 2575
2 7352 1 2575
2 7353 1 2577
2 7354 1 2577
2 7355 1 2580
2 7356 1 2580
2 7357 1 2583
2 7358 1 2583
2 7359 1 2585
2 7360 1 2585
2 7361 1 2586
2 7362 1 2586
2 7363 1 2591
2 7364 1 2591
2 7365 1 2594
2 7366 1 2594
2 7367 1 2595
2 7368 1 2595
2 7369 1 2598
2 7370 1 2598
2 7371 1 2601
2 7372 1 2601
2 7373 1 2603
2 7374 1 2603
2 7375 1 2604
2 7376 1 2604
2 7377 1 2609
2 7378 1 2609
2 7379 1 2612
2 7380 1 2612
2 7381 1 2617
2 7382 1 2617
2 7383 1 2617
2 7384 1 2623
2 7385 1 2623
2 7386 1 2623
2 7387 1 2625
2 7388 1 2625
2 7389 1 2628
2 7390 1 2628
2 7391 1 2631
2 7392 1 2631
2 7393 1 2633
2 7394 1 2633
2 7395 1 2634
2 7396 1 2634
2 7397 1 2639
2 7398 1 2639
2 7399 1 2642
2 7400 1 2642
2 7401 1 2643
2 7402 1 2643
2 7403 1 2646
2 7404 1 2646
2 7405 1 2649
2 7406 1 2649
2 7407 1 2651
2 7408 1 2651
2 7409 1 2652
2 7410 1 2652
2 7411 1 2657
2 7412 1 2657
2 7413 1 2660
2 7414 1 2660
2 7415 1 2665
2 7416 1 2665
2 7417 1 2665
2 7418 1 2671
2 7419 1 2671
2 7420 1 2671
2 7421 1 2673
2 7422 1 2673
2 7423 1 2676
2 7424 1 2676
2 7425 1 2679
2 7426 1 2679
2 7427 1 2681
2 7428 1 2681
2 7429 1 2682
2 7430 1 2682
2 7431 1 2687
2 7432 1 2687
2 7433 1 2690
2 7434 1 2690
2 7435 1 2691
2 7436 1 2691
2 7437 1 2694
2 7438 1 2694
2 7439 1 2697
2 7440 1 2697
2 7441 1 2699
2 7442 1 2699
2 7443 1 2700
2 7444 1 2700
2 7445 1 2705
2 7446 1 2705
2 7447 1 2708
2 7448 1 2708
2 7449 1 2713
2 7450 1 2713
2 7451 1 2713
2 7452 1 2719
2 7453 1 2719
2 7454 1 2719
2 7455 1 2721
2 7456 1 2721
2 7457 1 2724
2 7458 1 2724
2 7459 1 2727
2 7460 1 2727
2 7461 1 2729
2 7462 1 2729
2 7463 1 2730
2 7464 1 2730
2 7465 1 2735
2 7466 1 2735
2 7467 1 2738
2 7468 1 2738
2 7469 1 2739
2 7470 1 2739
2 7471 1 2742
2 7472 1 2742
2 7473 1 2745
2 7474 1 2745
2 7475 1 2747
2 7476 1 2747
2 7477 1 2748
2 7478 1 2748
2 7479 1 2753
2 7480 1 2753
2 7481 1 2756
2 7482 1 2756
2 7483 1 2761
2 7484 1 2761
2 7485 1 2761
2 7486 1 2767
2 7487 1 2767
2 7488 1 2767
2 7489 1 2769
2 7490 1 2769
2 7491 1 2772
2 7492 1 2772
2 7493 1 2775
2 7494 1 2775
2 7495 1 2777
2 7496 1 2777
2 7497 1 2778
2 7498 1 2778
2 7499 1 2783
2 7500 1 2783
2 7501 1 2786
2 7502 1 2786
2 7503 1 2787
2 7504 1 2787
2 7505 1 2790
2 7506 1 2790
2 7507 1 2793
2 7508 1 2793
2 7509 1 2795
2 7510 1 2795
2 7511 1 2796
2 7512 1 2796
2 7513 1 2801
2 7514 1 2801
2 7515 1 2804
2 7516 1 2804
2 7517 1 2809
2 7518 1 2809
2 7519 1 2809
2 7520 1 2815
2 7521 1 2815
2 7522 1 2815
2 7523 1 2817
2 7524 1 2817
2 7525 1 2820
2 7526 1 2820
2 7527 1 2823
2 7528 1 2823
2 7529 1 2825
2 7530 1 2825
2 7531 1 2826
2 7532 1 2826
2 7533 1 2831
2 7534 1 2831
2 7535 1 2834
2 7536 1 2834
2 7537 1 2835
2 7538 1 2835
2 7539 1 2838
2 7540 1 2838
2 7541 1 2841
2 7542 1 2841
2 7543 1 2843
2 7544 1 2843
2 7545 1 2844
2 7546 1 2844
2 7547 1 2849
2 7548 1 2849
2 7549 1 2852
2 7550 1 2852
2 7551 1 2857
2 7552 1 2857
2 7553 1 2857
2 7554 1 2863
2 7555 1 2863
2 7556 1 2863
2 7557 1 2865
2 7558 1 2865
2 7559 1 2868
2 7560 1 2868
2 7561 1 2871
2 7562 1 2871
2 7563 1 2873
2 7564 1 2873
2 7565 1 2874
2 7566 1 2874
2 7567 1 2879
2 7568 1 2879
2 7569 1 2882
2 7570 1 2882
2 7571 1 2883
2 7572 1 2883
2 7573 1 2886
2 7574 1 2886
2 7575 1 2889
2 7576 1 2889
2 7577 1 2891
2 7578 1 2891
2 7579 1 2892
2 7580 1 2892
2 7581 1 2897
2 7582 1 2897
2 7583 1 2900
2 7584 1 2900
2 7585 1 2905
2 7586 1 2905
2 7587 1 2905
2 7588 1 2911
2 7589 1 2911
2 7590 1 2911
2 7591 1 2913
2 7592 1 2913
2 7593 1 2916
2 7594 1 2916
2 7595 1 2919
2 7596 1 2919
2 7597 1 2921
2 7598 1 2921
2 7599 1 2922
2 7600 1 2922
2 7601 1 2927
2 7602 1 2927
2 7603 1 2930
2 7604 1 2930
2 7605 1 2931
2 7606 1 2931
2 7607 1 2934
2 7608 1 2934
2 7609 1 2937
2 7610 1 2937
2 7611 1 2939
2 7612 1 2939
2 7613 1 2940
2 7614 1 2940
2 7615 1 2945
2 7616 1 2945
2 7617 1 2948
2 7618 1 2948
2 7619 1 2953
2 7620 1 2953
2 7621 1 2953
2 7622 1 2959
2 7623 1 2959
2 7624 1 2959
2 7625 1 2961
2 7626 1 2961
2 7627 1 2964
2 7628 1 2964
2 7629 1 2967
2 7630 1 2967
2 7631 1 2969
2 7632 1 2969
2 7633 1 2970
2 7634 1 2970
2 7635 1 2975
2 7636 1 2975
2 7637 1 2978
2 7638 1 2978
2 7639 1 2979
2 7640 1 2979
2 7641 1 2982
2 7642 1 2982
2 7643 1 2985
2 7644 1 2985
2 7645 1 2987
2 7646 1 2987
2 7647 1 2988
2 7648 1 2988
2 7649 1 2993
2 7650 1 2993
2 7651 1 2996
2 7652 1 2996
2 7653 1 3001
2 7654 1 3001
2 7655 1 3001
2 7656 1 3007
2 7657 1 3007
2 7658 1 3007
2 7659 1 3009
2 7660 1 3009
2 7661 1 3012
2 7662 1 3012
2 7663 1 3015
2 7664 1 3015
2 7665 1 3017
2 7666 1 3017
2 7667 1 3018
2 7668 1 3018
2 7669 1 3023
2 7670 1 3023
2 7671 1 3026
2 7672 1 3026
2 7673 1 3027
2 7674 1 3027
2 7675 1 3030
2 7676 1 3030
2 7677 1 3033
2 7678 1 3033
2 7679 1 3035
2 7680 1 3035
2 7681 1 3036
2 7682 1 3036
2 7683 1 3041
2 7684 1 3041
2 7685 1 3044
2 7686 1 3044
2 7687 1 3049
2 7688 1 3049
2 7689 1 3049
2 7690 1 3055
2 7691 1 3055
2 7692 1 3055
2 7693 1 3057
2 7694 1 3057
2 7695 1 3060
2 7696 1 3060
2 7697 1 3063
2 7698 1 3063
2 7699 1 3065
2 7700 1 3065
2 7701 1 3066
2 7702 1 3066
2 7703 1 3071
2 7704 1 3071
2 7705 1 3074
2 7706 1 3074
2 7707 1 3075
2 7708 1 3075
2 7709 1 3078
2 7710 1 3078
2 7711 1 3081
2 7712 1 3081
2 7713 1 3083
2 7714 1 3083
2 7715 1 3084
2 7716 1 3084
2 7717 1 3089
2 7718 1 3089
2 7719 1 3092
2 7720 1 3092
2 7721 1 3097
2 7722 1 3097
2 7723 1 3097
2 7724 1 3103
2 7725 1 3103
2 7726 1 3103
2 7727 1 3105
2 7728 1 3105
2 7729 1 3108
2 7730 1 3108
2 7731 1 3111
2 7732 1 3111
2 7733 1 3113
2 7734 1 3113
2 7735 1 3114
2 7736 1 3114
2 7737 1 3119
2 7738 1 3119
2 7739 1 3122
2 7740 1 3122
2 7741 1 3123
2 7742 1 3123
2 7743 1 3126
2 7744 1 3126
2 7745 1 3129
2 7746 1 3129
2 7747 1 3131
2 7748 1 3131
2 7749 1 3132
2 7750 1 3132
2 7751 1 3137
2 7752 1 3137
2 7753 1 3140
2 7754 1 3140
2 7755 1 3145
2 7756 1 3145
2 7757 1 3145
2 7758 1 3151
2 7759 1 3151
2 7760 1 3151
2 7761 1 3153
2 7762 1 3153
2 7763 1 3156
2 7764 1 3156
2 7765 1 3159
2 7766 1 3159
2 7767 1 3161
2 7768 1 3161
2 7769 1 3162
2 7770 1 3162
2 7771 1 3167
2 7772 1 3167
2 7773 1 3170
2 7774 1 3170
2 7775 1 3171
2 7776 1 3171
2 7777 1 3174
2 7778 1 3174
2 7779 1 3177
2 7780 1 3177
2 7781 1 3179
2 7782 1 3179
2 7783 1 3180
2 7784 1 3180
2 7785 1 3185
2 7786 1 3185
2 7787 1 3188
2 7788 1 3188
2 7789 1 3193
2 7790 1 3193
2 7791 1 3193
2 7792 1 3199
2 7793 1 3199
2 7794 1 3199
2 7795 1 3201
2 7796 1 3201
2 7797 1 3204
2 7798 1 3204
2 7799 1 3207
2 7800 1 3207
2 7801 1 3209
2 7802 1 3209
2 7803 1 3210
2 7804 1 3210
2 7805 1 3215
2 7806 1 3215
2 7807 1 3218
2 7808 1 3218
2 7809 1 3219
2 7810 1 3219
2 7811 1 3222
2 7812 1 3222
2 7813 1 3225
2 7814 1 3225
2 7815 1 3227
2 7816 1 3227
2 7817 1 3228
2 7818 1 3228
2 7819 1 3233
2 7820 1 3233
2 7821 1 3236
2 7822 1 3236
2 7823 1 3241
2 7824 1 3241
2 7825 1 3241
2 7826 1 3247
2 7827 1 3247
2 7828 1 3247
2 7829 1 3249
2 7830 1 3249
2 7831 1 3252
2 7832 1 3252
2 7833 1 3255
2 7834 1 3255
2 7835 1 3257
2 7836 1 3257
2 7837 1 3258
2 7838 1 3258
2 7839 1 3263
2 7840 1 3263
2 7841 1 3266
2 7842 1 3266
2 7843 1 3267
2 7844 1 3267
2 7845 1 3270
2 7846 1 3270
2 7847 1 3273
2 7848 1 3273
2 7849 1 3275
2 7850 1 3275
2 7851 1 3276
2 7852 1 3276
2 7853 1 3281
2 7854 1 3281
2 7855 1 3284
2 7856 1 3284
2 7857 1 3289
2 7858 1 3289
2 7859 1 3289
2 7860 1 3295
2 7861 1 3295
2 7862 1 3295
2 7863 1 3297
2 7864 1 3297
2 7865 1 3300
2 7866 1 3300
2 7867 1 3303
2 7868 1 3303
2 7869 1 3305
2 7870 1 3305
2 7871 1 3306
2 7872 1 3306
2 7873 1 3311
2 7874 1 3311
2 7875 1 3314
2 7876 1 3314
2 7877 1 3315
2 7878 1 3315
2 7879 1 3318
2 7880 1 3318
2 7881 1 3321
2 7882 1 3321
2 7883 1 3323
2 7884 1 3323
2 7885 1 3324
2 7886 1 3324
2 7887 1 3329
2 7888 1 3329
2 7889 1 3332
2 7890 1 3332
2 7891 1 3337
2 7892 1 3337
2 7893 1 3337
2 7894 1 3343
2 7895 1 3343
2 7896 1 3343
2 7897 1 3345
2 7898 1 3345
2 7899 1 3348
2 7900 1 3348
2 7901 1 3351
2 7902 1 3351
2 7903 1 3353
2 7904 1 3353
2 7905 1 3354
2 7906 1 3354
2 7907 1 3359
2 7908 1 3359
2 7909 1 3362
2 7910 1 3362
2 7911 1 3363
2 7912 1 3363
2 7913 1 3366
2 7914 1 3366
2 7915 1 3369
2 7916 1 3369
2 7917 1 3371
2 7918 1 3371
2 7919 1 3372
2 7920 1 3372
2 7921 1 3377
2 7922 1 3377
2 7923 1 3380
2 7924 1 3380
2 7925 1 3385
2 7926 1 3385
2 7927 1 3385
2 7928 1 3391
2 7929 1 3391
2 7930 1 3391
2 7931 1 3393
2 7932 1 3393
2 7933 1 3396
2 7934 1 3396
2 7935 1 3399
2 7936 1 3399
2 7937 1 3401
2 7938 1 3401
2 7939 1 3402
2 7940 1 3402
2 7941 1 3407
2 7942 1 3407
2 7943 1 3410
2 7944 1 3410
2 7945 1 3411
2 7946 1 3411
2 7947 1 3414
2 7948 1 3414
2 7949 1 3417
2 7950 1 3417
2 7951 1 3419
2 7952 1 3419
2 7953 1 3420
2 7954 1 3420
2 7955 1 3425
2 7956 1 3425
2 7957 1 3428
2 7958 1 3428
2 7959 1 3433
2 7960 1 3433
2 7961 1 3433
2 7962 1 3439
2 7963 1 3439
2 7964 1 3439
2 7965 1 3441
2 7966 1 3441
2 7967 1 3444
2 7968 1 3444
2 7969 1 3447
2 7970 1 3447
2 7971 1 3449
2 7972 1 3449
2 7973 1 3450
2 7974 1 3450
2 7975 1 3455
2 7976 1 3455
2 7977 1 3458
2 7978 1 3458
2 7979 1 3459
2 7980 1 3459
2 7981 1 3462
2 7982 1 3462
2 7983 1 3465
2 7984 1 3465
2 7985 1 3467
2 7986 1 3467
2 7987 1 3468
2 7988 1 3468
2 7989 1 3473
2 7990 1 3473
2 7991 1 3476
2 7992 1 3476
2 7993 1 3481
2 7994 1 3481
2 7995 1 3481
2 7996 1 3483
2 7997 1 3483
2 7998 1 3486
2 7999 1 3486
2 8000 1 3489
2 8001 1 3489
2 8002 1 3489
2 8003 1 3491
2 8004 1 3491
2 8005 1 3492
2 8006 1 3492
2 8007 1 3497
2 8008 1 3497
2 8009 1 3500
2 8010 1 3500
2 8011 1 3505
2 8012 1 3505
2 8013 1 3505
2 8014 1 3511
2 8015 1 3511
2 8016 1 3514
2 8017 1 3514
2 8018 1 3516
2 8019 1 3516
2 8020 1 3517
2 8021 1 3517
2 8022 1 3530
2 8023 1 3530
2 8024 1 3536
2 8025 1 3536
2 8026 1 3541
2 8027 1 3541
2 8028 1 3544
2 8029 1 3544
2 8030 1 3547
2 8031 1 3547
2 8032 1 3550
2 8033 1 3550
2 8034 1 3553
2 8035 1 3553
2 8036 1 3553
2 8037 1 3559
2 8038 1 3559
2 8039 1 3561
2 8040 1 3561
2 8041 1 3567
2 8042 1 3567
2 8043 1 3568
2 8044 1 3568
2 8045 1 3573
2 8046 1 3573
2 8047 1 3576
2 8048 1 3576
2 8049 1 3581
2 8050 1 3581
2 8051 1 3584
2 8052 1 3584
2 8053 1 3587
2 8054 1 3587
2 8055 1 3594
2 8056 1 3594
2 8057 1 3597
2 8058 1 3597
2 8059 1 3599
2 8060 1 3599
2 8061 1 3601
2 8062 1 3601
2 8063 1 3604
2 8064 1 3604
2 8065 1 3607
2 8066 1 3607
2 8067 1 3610
2 8068 1 3610
2 8069 1 3613
2 8070 1 3613
2 8071 1 3620
2 8072 1 3620
2 8073 1 3623
2 8074 1 3623
2 8075 1 3625
2 8076 1 3625
2 8077 1 3627
2 8078 1 3627
2 8079 1 3630
2 8080 1 3630
2 8081 1 3633
2 8082 1 3633
2 8083 1 3636
2 8084 1 3636
2 8085 1 3639
2 8086 1 3639
2 8087 1 3646
2 8088 1 3646
2 8089 1 3649
2 8090 1 3649
2 8091 1 3651
2 8092 1 3651
2 8093 1 3653
2 8094 1 3653
2 8095 1 3656
2 8096 1 3656
2 8097 1 3659
2 8098 1 3659
2 8099 1 3662
2 8100 1 3662
2 8101 1 3665
2 8102 1 3665
2 8103 1 3672
2 8104 1 3672
2 8105 1 3675
2 8106 1 3675
2 8107 1 3677
2 8108 1 3677
2 8109 1 3679
2 8110 1 3679
2 8111 1 3682
2 8112 1 3682
2 8113 1 3685
2 8114 1 3685
2 8115 1 3688
2 8116 1 3688
2 8117 1 3691
2 8118 1 3691
2 8119 1 3698
2 8120 1 3698
2 8121 1 3701
2 8122 1 3701
2 8123 1 3703
2 8124 1 3703
2 8125 1 3705
2 8126 1 3705
2 8127 1 3708
2 8128 1 3708
2 8129 1 3711
2 8130 1 3711
2 8131 1 3714
2 8132 1 3714
2 8133 1 3717
2 8134 1 3717
2 8135 1 3724
2 8136 1 3724
2 8137 1 3727
2 8138 1 3727
2 8139 1 3729
2 8140 1 3729
2 8141 1 3731
2 8142 1 3731
2 8143 1 3734
2 8144 1 3734
2 8145 1 3737
2 8146 1 3737
2 8147 1 3740
2 8148 1 3740
2 8149 1 3743
2 8150 1 3743
2 8151 1 3750
2 8152 1 3750
2 8153 1 3753
2 8154 1 3753
2 8155 1 3755
2 8156 1 3755
2 8157 1 3757
2 8158 1 3757
2 8159 1 3760
2 8160 1 3760
2 8161 1 3763
2 8162 1 3763
2 8163 1 3766
2 8164 1 3766
2 8165 1 3769
2 8166 1 3769
2 8167 1 3776
2 8168 1 3776
2 8169 1 3779
2 8170 1 3779
2 8171 1 3781
2 8172 1 3781
2 8173 1 3783
2 8174 1 3783
2 8175 1 3786
2 8176 1 3786
2 8177 1 3789
2 8178 1 3789
2 8179 1 3792
2 8180 1 3792
2 8181 1 3795
2 8182 1 3795
2 8183 1 3802
2 8184 1 3802
2 8185 1 3805
2 8186 1 3805
2 8187 1 3807
2 8188 1 3807
2 8189 1 3809
2 8190 1 3809
2 8191 1 3812
2 8192 1 3812
2 8193 1 3815
2 8194 1 3815
2 8195 1 3818
2 8196 1 3818
2 8197 1 3821
2 8198 1 3821
2 8199 1 3828
2 8200 1 3828
2 8201 1 3831
2 8202 1 3831
2 8203 1 3833
2 8204 1 3833
2 8205 1 3835
2 8206 1 3835
2 8207 1 3838
2 8208 1 3838
2 8209 1 3841
2 8210 1 3841
2 8211 1 3844
2 8212 1 3844
2 8213 1 3847
2 8214 1 3847
2 8215 1 3854
2 8216 1 3854
2 8217 1 3857
2 8218 1 3857
2 8219 1 3859
2 8220 1 3859
2 8221 1 3861
2 8222 1 3861
2 8223 1 3864
2 8224 1 3864
2 8225 1 3867
2 8226 1 3867
2 8227 1 3870
2 8228 1 3870
2 8229 1 3873
2 8230 1 3873
2 8231 1 3880
2 8232 1 3880
2 8233 1 3883
2 8234 1 3883
2 8235 1 3885
2 8236 1 3885
2 8237 1 3887
2 8238 1 3887
2 8239 1 3890
2 8240 1 3890
2 8241 1 3893
2 8242 1 3893
2 8243 1 3896
2 8244 1 3896
2 8245 1 3899
2 8246 1 3899
2 8247 1 3906
2 8248 1 3906
2 8249 1 3909
2 8250 1 3909
2 8251 1 3911
2 8252 1 3911
2 8253 1 3913
2 8254 1 3913
2 8255 1 3916
2 8256 1 3916
2 8257 1 3919
2 8258 1 3919
2 8259 1 3922
2 8260 1 3922
2 8261 1 3925
2 8262 1 3925
2 8263 1 3932
2 8264 1 3932
2 8265 1 3935
2 8266 1 3935
2 8267 1 3937
2 8268 1 3937
2 8269 1 3939
2 8270 1 3939
2 8271 1 3942
2 8272 1 3942
2 8273 1 3945
2 8274 1 3945
2 8275 1 3948
2 8276 1 3948
2 8277 1 3951
2 8278 1 3951
2 8279 1 3958
2 8280 1 3958
2 8281 1 3961
2 8282 1 3961
2 8283 1 3963
2 8284 1 3963
2 8285 1 3965
2 8286 1 3965
2 8287 1 3968
2 8288 1 3968
2 8289 1 3971
2 8290 1 3971
2 8291 1 3974
2 8292 1 3974
2 8293 1 3977
2 8294 1 3977
2 8295 1 3984
2 8296 1 3984
2 8297 1 3987
2 8298 1 3987
2 8299 1 3989
2 8300 1 3989
2 8301 1 3991
2 8302 1 3991
2 8303 1 3994
2 8304 1 3994
2 8305 1 3997
2 8306 1 3997
2 8307 1 4000
2 8308 1 4000
2 8309 1 4003
2 8310 1 4003
2 8311 1 4010
2 8312 1 4010
2 8313 1 4013
2 8314 1 4013
2 8315 1 4015
2 8316 1 4015
2 8317 1 4017
2 8318 1 4017
2 8319 1 4020
2 8320 1 4020
2 8321 1 4023
2 8322 1 4023
2 8323 1 4026
2 8324 1 4026
2 8325 1 4029
2 8326 1 4029
2 8327 1 4036
2 8328 1 4036
2 8329 1 4039
2 8330 1 4039
2 8331 1 4041
2 8332 1 4041
2 8333 1 4043
2 8334 1 4043
2 8335 1 4046
2 8336 1 4046
2 8337 1 4049
2 8338 1 4049
2 8339 1 4052
2 8340 1 4052
2 8341 1 4055
2 8342 1 4055
2 8343 1 4062
2 8344 1 4062
2 8345 1 4065
2 8346 1 4065
2 8347 1 4067
2 8348 1 4067
2 8349 1 4069
2 8350 1 4069
2 8351 1 4072
2 8352 1 4072
2 8353 1 4075
2 8354 1 4075
2 8355 1 4078
2 8356 1 4078
2 8357 1 4081
2 8358 1 4081
2 8359 1 4088
2 8360 1 4088
2 8361 1 4091
2 8362 1 4091
2 8363 1 4093
2 8364 1 4093
2 8365 1 4095
2 8366 1 4095
2 8367 1 4098
2 8368 1 4098
2 8369 1 4101
2 8370 1 4101
2 8371 1 4104
2 8372 1 4104
2 8373 1 4107
2 8374 1 4107
2 8375 1 4114
2 8376 1 4114
2 8377 1 4117
2 8378 1 4117
2 8379 1 4119
2 8380 1 4119
2 8381 1 4121
2 8382 1 4121
2 8383 1 4129
2 8384 1 4129
2 8385 1 4151
2 8386 1 4151
2 8387 1 4154
2 8388 1 4154
2 8389 1 4156
2 8390 1 4156
2 8391 1 4158
2 8392 1 4158
2 8393 1 4160
2 8394 1 4160
2 8395 1 4161
2 8396 1 4161
2 8397 1 4162
2 8398 1 4162
2 8399 1 4162
2 8400 1 4165
2 8401 1 4165
2 8402 1 4166
2 8403 1 4166
2 8404 1 4169
2 8405 1 4169
2 8406 1 4172
2 8407 1 4172
2 8408 1 4174
2 8409 1 4174
2 8410 1 4177
2 8411 1 4177
2 8412 1 4180
2 8413 1 4180
2 8414 1 4182
2 8415 1 4182
2 8416 1 4185
2 8417 1 4185
2 8418 1 4188
2 8419 1 4188
2 8420 1 4190
2 8421 1 4190
2 8422 1 4193
2 8423 1 4193
2 8424 1 4196
2 8425 1 4196
2 8426 1 4198
2 8427 1 4198
2 8428 1 4201
2 8429 1 4201
2 8430 1 4204
2 8431 1 4204
2 8432 1 4206
2 8433 1 4206
2 8434 1 4209
2 8435 1 4209
2 8436 1 4212
2 8437 1 4212
2 8438 1 4214
2 8439 1 4214
2 8440 1 4217
2 8441 1 4217
2 8442 1 4220
2 8443 1 4220
2 8444 1 4222
2 8445 1 4222
2 8446 1 4225
2 8447 1 4225
2 8448 1 4228
2 8449 1 4228
2 8450 1 4230
2 8451 1 4230
2 8452 1 4233
2 8453 1 4233
2 8454 1 4236
2 8455 1 4236
2 8456 1 4238
2 8457 1 4238
2 8458 1 4241
2 8459 1 4241
2 8460 1 4244
2 8461 1 4244
2 8462 1 4246
2 8463 1 4246
2 8464 1 4249
2 8465 1 4249
2 8466 1 4252
2 8467 1 4252
2 8468 1 4254
2 8469 1 4254
2 8470 1 4257
2 8471 1 4257
2 8472 1 4260
2 8473 1 4260
2 8474 1 4262
2 8475 1 4262
2 8476 1 4263
2 8477 1 4263
2 8478 1 4269
2 8479 1 4269
2 8480 1 4272
2 8481 1 4272
2 8482 1 4272
2 8483 1 4273
2 8484 1 4273
2 8485 1 4279
2 8486 1 4279
2 8487 1 4282
2 8488 1 4282
2 8489 1 4282
2 8490 1 4284
2 8491 1 4284
2 8492 1 4284
2 8493 1 4284
2 8494 1 4285
2 8495 1 4285
2 8496 1 4291
2 8497 1 4291
2 8498 1 4294
2 8499 1 4294
2 8500 1 4294
2 8501 1 4296
2 8502 1 4296
2 8503 1 4296
2 8504 1 4296
2 8505 1 4297
2 8506 1 4297
2 8507 1 4303
2 8508 1 4303
2 8509 1 4306
2 8510 1 4306
2 8511 1 4306
2 8512 1 4306
2 8513 1 4307
2 8514 1 4307
2 8515 1 4313
2 8516 1 4313
2 8517 1 4315
2 8518 1 4315
2 8519 1 4315
2 8520 1 4316
2 8521 1 4316
2 8522 1 4318
2 8523 1 4318
2 8524 1 4318
2 8525 1 4318
2 8526 1 4319
2 8527 1 4319
2 8528 1 4320
2 8529 1 4320
2 8530 1 4326
2 8531 1 4326
2 8532 1 4329
2 8533 1 4329
2 8534 1 4329
2 8535 1 4331
2 8536 1 4331
2 8537 1 4331
2 8538 1 4331
2 8539 1 4332
2 8540 1 4332
2 8541 1 4338
2 8542 1 4338
2 8543 1 4341
2 8544 1 4341
2 8545 1 4341
2 8546 1 4343
2 8547 1 4343
2 8548 1 4343
2 8549 1 4343
2 8550 1 4344
2 8551 1 4344
2 8552 1 4350
2 8553 1 4350
2 8554 1 4353
2 8555 1 4353
2 8556 1 4353
2 8557 1 4353
2 8558 1 4355
2 8559 1 4355
2 8560 1 4355
2 8561 1 4355
2 8562 1 4356
2 8563 1 4356
2 8564 1 4362
2 8565 1 4362
2 8566 1 4365
2 8567 1 4365
2 8568 1 4365
2 8569 1 4365
2 8570 1 4366
2 8571 1 4366
2 8572 1 4372
2 8573 1 4372
2 8574 1 4375
2 8575 1 4375
2 8576 1 4375
2 8577 1 4375
2 8578 1 4376
2 8579 1 4376
2 8580 1 4382
2 8581 1 4382
2 8582 1 4385
2 8583 1 4385
2 8584 1 4385
2 8585 1 4385
2 8586 1 4387
2 8587 1 4387
2 8588 1 4387
2 8589 1 4388
2 8590 1 4388
2 8591 1 4394
2 8592 1 4394
2 8593 1 4397
2 8594 1 4397
2 8595 1 4397
2 8596 1 4397
2 8597 1 4399
2 8598 1 4399
2 8599 1 4399
2 8600 1 4402
2 8601 1 4402
2 8602 1 4406
2 8603 1 4406
2 8604 1 4412
2 8605 1 4412
2 8606 1 4415
2 8607 1 4415
2 8608 1 4416
2 8609 1 4416
2 8610 1 4422
2 8611 1 4422
2 8612 1 4426
2 8613 1 4426
2 8614 1 4428
2 8615 1 4428
2 8616 1 4430
2 8617 1 4430
2 8618 1 4435
2 8619 1 4435
2 8620 1 4435
2 8621 1 4437
2 8622 1 4437
2 8623 1 4438
2 8624 1 4438
2 8625 1 4441
2 8626 1 4441
2 8627 1 4442
2 8628 1 4442
2 8629 1 4445
2 8630 1 4445
2 8631 1 4448
2 8632 1 4448
2 8633 1 4450
2 8634 1 4450
2 8635 1 4450
2 8636 1 4450
2 8637 1 4452
2 8638 1 4452
2 8639 1 4452
2 8640 1 4452
2 8641 1 4453
2 8642 1 4453
2 8643 1 4456
2 8644 1 4456
2 8645 1 4460
2 8646 1 4460
2 8647 1 4461
2 8648 1 4461
2 8649 1 4464
2 8650 1 4464
2 8651 1 4465
2 8652 1 4465
2 8653 1 4468
2 8654 1 4468
2 8655 1 4468
2 8656 1 4470
2 8657 1 4470
2 8658 1 4470
2 8659 1 4471
2 8660 1 4471
2 8661 1 4477
2 8662 1 4477
2 8663 1 4480
2 8664 1 4480
2 8665 1 4481
2 8666 1 4481
2 8667 1 4484
2 8668 1 4484
2 8669 1 4485
2 8670 1 4485
2 8671 1 4487
2 8672 1 4487
2 8673 1 4487
2 8674 1 4487
2 8675 1 4490
2 8676 1 4490
2 8677 1 4491
2 8678 1 4491
2 8679 1 4494
2 8680 1 4494
2 8681 1 4497
2 8682 1 4497
2 8683 1 4499
2 8684 1 4499
2 8685 1 4500
2 8686 1 4500
2 8687 1 4506
2 8688 1 4506
2 8689 1 4509
2 8690 1 4509
2 8691 1 4509
2 8692 1 4510
2 8693 1 4510
2 8694 1 4511
2 8695 1 4511
2 8696 1 4511
2 8697 1 4512
2 8698 1 4512
2 8699 1 4517
2 8700 1 4517
2 8701 1 4518
2 8702 1 4518
2 8703 1 4518
2 8704 1 4519
2 8705 1 4519
2 8706 1 4528
2 8707 1 4528
2 8708 1 4530
2 8709 1 4530
2 8710 1 4531
2 8711 1 4531
2 8712 1 4532
2 8713 1 4532
2 8714 1 4532
2 8715 1 4533
2 8716 1 4533
2 8717 1 4538
2 8718 1 4538
2 8719 1 4538
2 8720 1 4539
2 8721 1 4539
2 8722 1 4545
2 8723 1 4545
2 8724 1 4552
2 8725 1 4552
2 8726 1 4552
2 8727 1 4553
2 8728 1 4553
2 8729 1 4560
2 8730 1 4560
2 8731 1 4560
2 8732 1 4561
2 8733 1 4561
2 8734 1 4566
2 8735 1 4566
2 8736 1 4567
2 8737 1 4567
2 8738 1 4572
2 8739 1 4572
2 8740 1 4578
2 8741 1 4578
2 8742 1 4581
2 8743 1 4581
2 8744 1 4581
2 8745 1 4582
2 8746 1 4582
2 8747 1 4585
2 8748 1 4585
2 8749 1 4585
2 8750 1 4586
2 8751 1 4586
2 8752 1 4592
2 8753 1 4592
2 8754 1 4592
2 8755 1 4595
2 8756 1 4595
2 8757 1 4624
2 8758 1 4624
2 8759 1 4625
2 8760 1 4625
2 8761 1 4625
2 8762 1 4628
2 8763 1 4628
2 8764 1 4631
2 8765 1 4631
2 8766 1 4639
2 8767 1 4639
2 8768 1 4640
2 8769 1 4640
2 8770 1 4643
2 8771 1 4643
2 8772 1 4644
2 8773 1 4644
2 8774 1 4647
2 8775 1 4647
2 8776 1 4650
2 8777 1 4650
2 8778 1 4655
2 8779 1 4655
2 8780 1 4657
2 8781 1 4657
2 8782 1 4658
2 8783 1 4658
2 8784 1 4661
2 8785 1 4661
2 8786 1 4662
2 8787 1 4662
2 8788 1 4665
2 8789 1 4665
2 8790 1 4666
2 8791 1 4666
2 8792 1 4672
2 8793 1 4672
2 8794 1 4676
2 8795 1 4676
2 8796 1 4677
2 8797 1 4677
2 8798 1 4680
2 8799 1 4680
2 8800 1 4681
2 8801 1 4681
2 8802 1 4684
2 8803 1 4684
2 8804 1 4684
2 8805 1 4690
2 8806 1 4690
0 50 5 7 1 49
0 51 5 6 1 4793
0 52 5 7 1 4801
0 53 5 7 1 4810
0 54 5 7 1 4818
0 55 5 7 1 4826
0 56 5 7 1 4834
0 57 5 7 1 4842
0 58 5 7 1 4850
0 59 5 7 1 4858
0 60 5 7 1 4866
0 61 5 7 1 4874
0 62 5 7 1 4882
0 63 5 7 1 4890
0 64 5 7 1 4898
0 65 5 7 1 4906
0 66 5 7 1 4914
0 67 5 7 1 4922
0 68 5 7 1 4930
0 69 5 8 1 4938
0 70 5 8 1 4946
0 71 5 8 1 4954
0 72 5 8 1 4962
0 73 5 8 1 4970
0 74 5 8 1 4978
0 75 5 8 1 4986
0 76 5 8 1 4994
0 77 5 8 1 5002
0 78 5 8 1 5010
0 79 5 8 1 5018
0 80 5 8 1 5026
0 81 5 8 1 5034
0 82 5 7 1 5042
0 83 5 7 1 5050
0 84 5 7 1 5058
0 85 5 7 1 5066
0 86 5 7 1 5074
0 87 5 7 1 5082
0 88 5 7 1 5090
0 89 5 7 1 5098
0 90 5 7 1 5106
0 91 5 7 1 5114
0 92 5 7 1 5122
0 93 5 7 1 5130
0 94 5 8 1 5138
0 95 5 7 1 5146
0 96 5 5 1 5156
0 97 5 4 1 5165
0 98 5 6 1 5173
0 99 7 2 2 5508 5174
0 100 5 2 1 5530
0 101 7 1 2 5157 5532
0 102 5 1 1 101
0 103 7 1 2 5515 5166
0 104 7 2 2 5175 103
0 105 5 2 1 5534
0 106 7 1 2 5509 5535
0 107 5 1 1 106
0 108 7 2 2 102 107
0 109 5 1 1 5538
0 110 7 2 2 5520 5176
0 111 5 1 1 5540
0 112 7 2 2 5516 5541
0 113 5 3 1 5542
0 114 7 1 2 5147 5524
0 115 5 1 1 114
0 116 7 1 2 5533 115
0 117 5 1 1 116
0 118 7 2 2 5544 117
0 119 5 2 1 5547
0 120 7 3 2 5500 5549
0 121 7 1 2 5539 5551
0 122 5 2 1 121
0 123 7 2 2 5517 5531
0 124 5 1 1 5556
0 125 7 2 2 5167 124
0 126 5 1 1 5558
0 127 7 1 2 5554 5559
0 128 5 1 1 127
0 129 7 2 2 5521 5557
0 130 5 2 1 5560
0 131 7 2 2 128 5562
0 132 5 2 1 5564
0 133 7 1 2 5552 5566
0 134 5 2 1 133
0 135 7 1 2 109 5568
0 136 5 1 1 135
0 137 7 1 2 5501 5561
0 138 5 1 1 137
0 139 7 2 2 136 138
0 140 5 1 1 5570
0 141 7 1 2 5502 5567
0 142 5 2 1 141
0 143 7 1 2 5139 5565
0 144 5 1 1 143
0 145 7 3 2 5572 144
0 146 5 1 1 5574
0 147 7 2 2 5493 5575
0 148 7 2 2 5550 5577
0 149 5 2 1 5579
0 150 7 1 2 140 5581
0 151 5 2 1 150
0 152 7 1 2 5555 5563
0 153 5 1 1 152
0 154 7 1 2 5553 126
0 155 5 1 1 154
0 156 7 3 2 153 155
0 157 5 1 1 5585
0 158 7 2 2 5583 157
0 159 5 2 1 5588
0 160 7 1 2 5494 5590
0 161 5 2 1 160
0 162 7 1 2 5131 5589
0 163 5 1 1 162
0 164 7 3 2 5592 163
0 165 5 1 1 5594
0 166 7 1 2 5548 5573
0 167 5 1 1 166
0 168 7 1 2 5569 167
0 169 5 1 1 168
0 170 7 1 2 5578 5591
0 171 5 2 1 170
0 172 7 1 2 169 5597
0 173 5 1 1 172
0 174 7 1 2 5580 5586
0 175 5 1 1 174
0 176 7 2 2 173 175
0 177 5 1 1 5599
0 178 7 2 2 5486 5595
0 179 7 2 2 5576 5601
0 180 5 2 1 5603
0 181 7 1 2 177 5605
0 182 5 2 1 181
0 183 7 1 2 5582 5587
0 184 5 1 1 183
0 185 7 1 2 5571 184
0 186 5 1 1 185
0 187 7 3 2 5584 186
0 188 5 1 1 5609
0 189 7 2 2 5607 188
0 190 5 2 1 5612
0 191 7 1 2 5487 5614
0 192 5 2 1 191
0 193 7 1 2 165 5616
0 194 5 1 1 193
0 195 7 1 2 5602 5615
0 196 5 2 1 195
0 197 7 1 2 194 5618
0 198 5 1 1 197
0 199 7 1 2 5123 5613
0 200 5 1 1 199
0 201 7 3 2 5617 200
0 202 5 1 1 5620
0 203 7 2 2 5479 5621
0 204 7 1 2 146 5593
0 205 5 1 1 204
0 206 7 1 2 5598 205
0 207 5 1 1 206
0 208 7 1 2 5619 207
0 209 5 1 1 208
0 210 7 1 2 5604 5610
0 211 5 1 1 210
0 212 7 2 2 209 211
0 213 5 1 1 5625
0 214 7 2 2 5596 5623
0 215 5 2 1 5627
0 216 7 1 2 213 5629
0 217 5 2 1 216
0 218 7 1 2 5606 5611
0 219 5 1 1 218
0 220 7 1 2 5600 219
0 221 5 1 1 220
0 222 7 3 2 5608 221
0 223 5 1 1 5633
0 224 7 2 2 5631 223
0 225 5 2 1 5636
0 226 7 1 2 5624 5638
0 227 5 2 1 226
0 228 7 1 2 198 5640
0 229 5 1 1 228
0 230 7 1 2 5628 5634
0 231 5 1 1 230
0 232 7 2 2 229 231
0 233 5 1 1 5642
0 234 7 1 2 5480 5639
0 235 5 2 1 234
0 236 7 1 2 5115 5637
0 237 5 1 1 236
0 238 7 3 2 5644 237
0 239 5 1 1 5646
0 240 7 2 2 5472 5647
0 241 7 2 2 5622 5649
0 242 5 2 1 5651
0 243 7 1 2 233 5653
0 244 5 2 1 243
0 245 7 1 2 5630 5635
0 246 5 1 1 245
0 247 7 1 2 5626 246
0 248 5 1 1 247
0 249 7 3 2 5632 248
0 250 5 1 1 5657
0 251 7 2 2 5655 250
0 252 5 2 1 5660
0 253 7 1 2 5473 5662
0 254 5 2 1 253
0 255 7 1 2 5107 5661
0 256 5 1 1 255
0 257 7 3 2 5664 256
0 258 5 1 1 5666
0 259 7 1 2 202 5645
0 260 5 1 1 259
0 261 7 1 2 5641 260
0 262 5 1 1 261
0 263 7 1 2 5650 5663
0 264 5 2 1 263
0 265 7 1 2 262 5669
0 266 5 1 1 265
0 267 7 1 2 5652 5658
0 268 5 1 1 267
0 269 7 2 2 266 268
0 270 5 1 1 5671
0 271 7 2 2 5465 5667
0 272 7 2 2 5648 5673
0 273 5 2 1 5675
0 274 7 1 2 270 5677
0 275 5 2 1 274
0 276 7 1 2 5654 5659
0 277 5 1 1 276
0 278 7 1 2 5643 277
0 279 5 1 1 278
0 280 7 3 2 5656 279
0 281 5 1 1 5681
0 282 7 2 2 5679 281
0 283 5 2 1 5684
0 284 7 1 2 5466 5686
0 285 5 2 1 284
0 286 7 1 2 258 5688
0 287 5 1 1 286
0 288 7 1 2 5674 5687
0 289 5 2 1 288
0 290 7 1 2 287 5690
0 291 5 1 1 290
0 292 7 1 2 5099 5685
0 293 5 1 1 292
0 294 7 3 2 5689 293
0 295 5 1 1 5692
0 296 7 2 2 5458 5693
0 297 7 1 2 239 5665
0 298 5 1 1 297
0 299 7 1 2 5670 298
0 300 5 1 1 299
0 301 7 1 2 5691 300
0 302 5 1 1 301
0 303 7 1 2 5676 5682
0 304 5 1 1 303
0 305 7 2 2 302 304
0 306 5 1 1 5697
0 307 7 2 2 5668 5695
0 308 5 2 1 5699
0 309 7 1 2 306 5701
0 310 5 2 1 309
0 311 7 1 2 5678 5683
0 312 5 1 1 311
0 313 7 1 2 5672 312
0 314 5 1 1 313
0 315 7 3 2 5680 314
0 316 5 1 1 5705
0 317 7 2 2 5703 316
0 318 5 2 1 5708
0 319 7 1 2 5696 5710
0 320 5 2 1 319
0 321 7 1 2 291 5712
0 322 5 1 1 321
0 323 7 1 2 5700 5706
0 324 5 1 1 323
0 325 7 2 2 322 324
0 326 5 1 1 5714
0 327 7 1 2 5459 5711
0 328 5 2 1 327
0 329 7 1 2 5091 5709
0 330 5 1 1 329
0 331 7 3 2 5716 330
0 332 5 1 1 5718
0 333 7 2 2 5451 5719
0 334 7 2 2 5694 5721
0 335 5 2 1 5723
0 336 7 1 2 326 5725
0 337 5 2 1 336
0 338 7 1 2 5702 5707
0 339 5 1 1 338
0 340 7 1 2 5698 339
0 341 5 1 1 340
0 342 7 3 2 5704 341
0 343 5 1 1 5729
0 344 7 2 2 5727 343
0 345 5 2 1 5732
0 346 7 1 2 5452 5734
0 347 5 2 1 346
0 348 7 1 2 5083 5733
0 349 5 1 1 348
0 350 7 3 2 5736 349
0 351 5 1 1 5738
0 352 7 1 2 295 5717
0 353 5 1 1 352
0 354 7 1 2 5713 353
0 355 5 1 1 354
0 356 7 1 2 5722 5735
0 357 5 2 1 356
0 358 7 1 2 355 5741
0 359 5 1 1 358
0 360 7 1 2 5724 5730
0 361 5 1 1 360
0 362 7 2 2 359 361
0 363 5 1 1 5743
0 364 7 2 2 5444 5739
0 365 7 2 2 5720 5745
0 366 5 2 1 5747
0 367 7 1 2 363 5749
0 368 5 2 1 367
0 369 7 1 2 5726 5731
0 370 5 1 1 369
0 371 7 1 2 5715 370
0 372 5 1 1 371
0 373 7 3 2 5728 372
0 374 5 1 1 5753
0 375 7 2 2 5751 374
0 376 5 2 1 5756
0 377 7 1 2 5445 5758
0 378 5 2 1 377
0 379 7 1 2 351 5760
0 380 5 1 1 379
0 381 7 1 2 5746 5759
0 382 5 2 1 381
0 383 7 1 2 380 5762
0 384 5 1 1 383
0 385 7 1 2 5075 5757
0 386 5 1 1 385
0 387 7 3 2 5761 386
0 388 5 1 1 5764
0 389 7 2 2 5437 5765
0 390 7 1 2 332 5737
0 391 5 1 1 390
0 392 7 1 2 5742 391
0 393 5 1 1 392
0 394 7 1 2 5763 393
0 395 5 1 1 394
0 396 7 1 2 5748 5754
0 397 5 1 1 396
0 398 7 2 2 395 397
0 399 5 1 1 5769
0 400 7 2 2 5740 5767
0 401 5 2 1 5771
0 402 7 1 2 399 5773
0 403 5 2 1 402
0 404 7 1 2 5750 5755
0 405 5 1 1 404
0 406 7 1 2 5744 405
0 407 5 1 1 406
0 408 7 3 2 5752 407
0 409 5 1 1 5777
0 410 7 2 2 5775 409
0 411 5 2 1 5780
0 412 7 1 2 5768 5782
0 413 5 2 1 412
0 414 7 1 2 384 5784
0 415 5 1 1 414
0 416 7 1 2 5772 5778
0 417 5 1 1 416
0 418 7 2 2 415 417
0 419 5 1 1 5786
0 420 7 1 2 5438 5783
0 421 5 2 1 420
0 422 7 1 2 5067 5781
0 423 5 1 1 422
0 424 7 3 2 5788 423
0 425 5 1 1 5790
0 426 7 2 2 5430 5791
0 427 7 2 2 5766 5793
0 428 5 2 1 5795
0 429 7 1 2 419 5797
0 430 5 2 1 429
0 431 7 1 2 5774 5779
0 432 5 1 1 431
0 433 7 1 2 5770 432
0 434 5 1 1 433
0 435 7 3 2 5776 434
0 436 5 1 1 5801
0 437 7 2 2 5799 436
0 438 5 2 1 5804
0 439 7 1 2 5431 5806
0 440 5 2 1 439
0 441 7 1 2 5059 5805
0 442 5 1 1 441
0 443 7 3 2 5808 442
0 444 5 1 1 5810
0 445 7 1 2 388 5789
0 446 5 1 1 445
0 447 7 1 2 5785 446
0 448 5 1 1 447
0 449 7 1 2 5794 5807
0 450 5 2 1 449
0 451 7 1 2 448 5813
0 452 5 1 1 451
0 453 7 1 2 5796 5802
0 454 5 1 1 453
0 455 7 2 2 452 454
0 456 5 1 1 5815
0 457 7 2 2 5423 5811
0 458 7 2 2 5792 5817
0 459 5 2 1 5819
0 460 7 1 2 456 5821
0 461 5 2 1 460
0 462 7 1 2 5798 5803
0 463 5 1 1 462
0 464 7 1 2 5787 463
0 465 5 1 1 464
0 466 7 3 2 5800 465
0 467 5 1 1 5825
0 468 7 2 2 5823 467
0 469 5 2 1 5828
0 470 7 1 2 5424 5830
0 471 5 2 1 470
0 472 7 1 2 444 5832
0 473 5 1 1 472
0 474 7 1 2 5818 5831
0 475 5 2 1 474
0 476 7 1 2 473 5834
0 477 5 1 1 476
0 478 7 1 2 5051 5829
0 479 5 1 1 478
0 480 7 3 2 5833 479
0 481 5 1 1 5836
0 482 7 2 2 5416 5837
0 483 7 1 2 425 5809
0 484 5 1 1 483
0 485 7 1 2 5814 484
0 486 5 1 1 485
0 487 7 1 2 5835 486
0 488 5 1 1 487
0 489 7 1 2 5820 5826
0 490 5 1 1 489
0 491 7 2 2 488 490
0 492 5 1 1 5841
0 493 7 2 2 5812 5839
0 494 5 2 1 5843
0 495 7 1 2 492 5845
0 496 5 2 1 495
0 497 7 1 2 5822 5827
0 498 5 1 1 497
0 499 7 1 2 5816 498
0 500 5 1 1 499
0 501 7 3 2 5824 500
0 502 5 1 1 5849
0 503 7 2 2 5847 502
0 504 5 2 1 5852
0 505 7 1 2 5840 5854
0 506 5 2 1 505
0 507 7 1 2 477 5856
0 508 5 1 1 507
0 509 7 1 2 5844 5850
0 510 5 1 1 509
0 511 7 2 2 508 510
0 512 5 1 1 5858
0 513 7 1 2 5417 5855
0 514 5 2 1 513
0 515 7 1 2 5043 5853
0 516 5 1 1 515
0 517 7 3 2 5860 516
0 518 5 1 1 5862
0 519 7 2 2 5408 5863
0 520 7 2 2 5838 5865
0 521 5 2 1 5867
0 522 7 1 2 512 5869
0 523 5 2 1 522
0 524 7 1 2 5846 5851
0 525 5 1 1 524
0 526 7 1 2 5842 525
0 527 5 1 1 526
0 528 7 3 2 5848 527
0 529 5 1 1 5873
0 530 7 2 2 5871 529
0 531 5 2 1 5876
0 532 7 1 2 5409 5878
0 533 5 2 1 532
0 534 7 1 2 5035 5877
0 535 5 1 1 534
0 536 7 3 2 5880 535
0 537 5 1 1 5882
0 538 7 1 2 481 5861
0 539 5 1 1 538
0 540 7 1 2 5857 539
0 541 5 1 1 540
0 542 7 1 2 5866 5879
0 543 5 2 1 542
0 544 7 1 2 541 5885
0 545 5 1 1 544
0 546 7 1 2 5868 5874
0 547 5 1 1 546
0 548 7 2 2 545 547
0 549 5 1 1 5887
0 550 7 2 2 5400 5883
0 551 7 2 2 5864 5889
0 552 5 2 1 5891
0 553 7 1 2 549 5893
0 554 5 2 1 553
0 555 7 1 2 5870 5875
0 556 5 1 1 555
0 557 7 1 2 5859 556
0 558 5 1 1 557
0 559 7 3 2 5872 558
0 560 5 1 1 5897
0 561 7 2 2 5895 560
0 562 5 2 1 5900
0 563 7 1 2 5401 5902
0 564 5 2 1 563
0 565 7 1 2 537 5904
0 566 5 1 1 565
0 567 7 1 2 5890 5903
0 568 5 2 1 567
0 569 7 1 2 566 5906
0 570 5 1 1 569
0 571 7 1 2 5027 5901
0 572 5 1 1 571
0 573 7 3 2 5905 572
0 574 5 1 1 5908
0 575 7 2 2 5392 5909
0 576 7 1 2 518 5881
0 577 5 1 1 576
0 578 7 1 2 5886 577
0 579 5 1 1 578
0 580 7 1 2 5907 579
0 581 5 1 1 580
0 582 7 1 2 5892 5898
0 583 5 1 1 582
0 584 7 2 2 581 583
0 585 5 1 1 5913
0 586 7 2 2 5884 5911
0 587 5 2 1 5915
0 588 7 1 2 585 5917
0 589 5 2 1 588
0 590 7 1 2 5894 5899
0 591 5 1 1 590
0 592 7 1 2 5888 591
0 593 5 1 1 592
0 594 7 3 2 5896 593
0 595 5 1 1 5921
0 596 7 2 2 5919 595
0 597 5 2 1 5924
0 598 7 1 2 5912 5926
0 599 5 2 1 598
0 600 7 1 2 570 5928
0 601 5 1 1 600
0 602 7 1 2 5916 5922
0 603 5 1 1 602
0 604 7 2 2 601 603
0 605 5 1 1 5930
0 606 7 1 2 5393 5927
0 607 5 2 1 606
0 608 7 1 2 5019 5925
0 609 5 1 1 608
0 610 7 3 2 5932 609
0 611 5 1 1 5934
0 612 7 2 2 5384 5935
0 613 7 2 2 5910 5937
0 614 5 2 1 5939
0 615 7 1 2 605 5941
0 616 5 2 1 615
0 617 7 1 2 5918 5923
0 618 5 1 1 617
0 619 7 1 2 5914 618
0 620 5 1 1 619
0 621 7 3 2 5920 620
0 622 5 1 1 5945
0 623 7 2 2 5943 622
0 624 5 2 1 5948
0 625 7 1 2 5385 5950
0 626 5 2 1 625
0 627 7 1 2 5011 5949
0 628 5 1 1 627
0 629 7 3 2 5952 628
0 630 5 1 1 5954
0 631 7 1 2 574 5933
0 632 5 1 1 631
0 633 7 1 2 5929 632
0 634 5 1 1 633
0 635 7 1 2 5938 5951
0 636 5 2 1 635
0 637 7 1 2 634 5957
0 638 5 1 1 637
0 639 7 1 2 5940 5946
0 640 5 1 1 639
0 641 7 2 2 638 640
0 642 5 1 1 5959
0 643 7 2 2 5376 5955
0 644 7 2 2 5936 5961
0 645 5 2 1 5963
0 646 7 1 2 642 5965
0 647 5 2 1 646
0 648 7 1 2 5942 5947
0 649 5 1 1 648
0 650 7 1 2 5931 649
0 651 5 1 1 650
0 652 7 3 2 5944 651
0 653 5 1 1 5969
0 654 7 2 2 5967 653
0 655 5 2 1 5972
0 656 7 1 2 5377 5974
0 657 5 2 1 656
0 658 7 1 2 630 5976
0 659 5 1 1 658
0 660 7 1 2 5962 5975
0 661 5 2 1 660
0 662 7 1 2 659 5978
0 663 5 1 1 662
0 664 7 1 2 5003 5973
0 665 5 1 1 664
0 666 7 3 2 5977 665
0 667 5 1 1 5980
0 668 7 2 2 5368 5981
0 669 7 1 2 611 5953
0 670 5 1 1 669
0 671 7 1 2 5958 670
0 672 5 1 1 671
0 673 7 1 2 5979 672
0 674 5 1 1 673
0 675 7 1 2 5964 5970
0 676 5 1 1 675
0 677 7 2 2 674 676
0 678 5 1 1 5985
0 679 7 2 2 5956 5983
0 680 5 2 1 5987
0 681 7 1 2 678 5989
0 682 5 2 1 681
0 683 7 1 2 5966 5971
0 684 5 1 1 683
0 685 7 1 2 5960 684
0 686 5 1 1 685
0 687 7 3 2 5968 686
0 688 5 1 1 5993
0 689 7 2 2 5991 688
0 690 5 2 1 5996
0 691 7 1 2 5984 5998
0 692 5 2 1 691
0 693 7 1 2 663 6000
0 694 5 1 1 693
0 695 7 1 2 5988 5994
0 696 5 1 1 695
0 697 7 2 2 694 696
0 698 5 1 1 6002
0 699 7 1 2 5369 5999
0 700 5 2 1 699
0 701 7 1 2 4995 5997
0 702 5 1 1 701
0 703 7 3 2 6004 702
0 704 5 1 1 6006
0 705 7 2 2 5360 6007
0 706 7 2 2 5982 6009
0 707 5 2 1 6011
0 708 7 1 2 698 6013
0 709 5 2 1 708
0 710 7 1 2 5990 5995
0 711 5 1 1 710
0 712 7 1 2 5986 711
0 713 5 1 1 712
0 714 7 3 2 5992 713
0 715 5 1 1 6017
0 716 7 2 2 6015 715
0 717 5 2 1 6020
0 718 7 1 2 5361 6022
0 719 5 2 1 718
0 720 7 1 2 4987 6021
0 721 5 1 1 720
0 722 7 3 2 6024 721
0 723 5 1 1 6026
0 724 7 1 2 667 6005
0 725 5 1 1 724
0 726 7 1 2 6001 725
0 727 5 1 1 726
0 728 7 1 2 6010 6023
0 729 5 2 1 728
0 730 7 1 2 727 6029
0 731 5 1 1 730
0 732 7 1 2 6012 6018
0 733 5 1 1 732
0 734 7 2 2 731 733
0 735 5 1 1 6031
0 736 7 2 2 5352 6027
0 737 7 2 2 6008 6033
0 738 5 2 1 6035
0 739 7 1 2 735 6037
0 740 5 2 1 739
0 741 7 1 2 6014 6019
0 742 5 1 1 741
0 743 7 1 2 6003 742
0 744 5 1 1 743
0 745 7 3 2 6016 744
0 746 5 1 1 6041
0 747 7 2 2 6039 746
0 748 5 2 1 6044
0 749 7 1 2 5353 6046
0 750 5 2 1 749
0 751 7 1 2 723 6048
0 752 5 1 1 751
0 753 7 1 2 6034 6047
0 754 5 2 1 753
0 755 7 1 2 752 6050
0 756 5 1 1 755
0 757 7 1 2 4979 6045
0 758 5 1 1 757
0 759 7 3 2 6049 758
0 760 5 1 1 6052
0 761 7 2 2 5344 6053
0 762 7 1 2 704 6025
0 763 5 1 1 762
0 764 7 1 2 6030 763
0 765 5 1 1 764
0 766 7 1 2 6051 765
0 767 5 1 1 766
0 768 7 1 2 6036 6042
0 769 5 1 1 768
0 770 7 2 2 767 769
0 771 5 1 1 6057
0 772 7 2 2 6028 6055
0 773 5 2 1 6059
0 774 7 1 2 771 6061
0 775 5 2 1 774
0 776 7 1 2 6038 6043
0 777 5 1 1 776
0 778 7 1 2 6032 777
0 779 5 1 1 778
0 780 7 3 2 6040 779
0 781 5 1 1 6065
0 782 7 2 2 6063 781
0 783 5 2 1 6068
0 784 7 1 2 6056 6070
0 785 5 2 1 784
0 786 7 1 2 756 6072
0 787 5 1 1 786
0 788 7 1 2 6060 6066
0 789 5 1 1 788
0 790 7 2 2 787 789
0 791 5 1 1 6074
0 792 7 1 2 5345 6071
0 793 5 2 1 792
0 794 7 1 2 4971 6069
0 795 5 1 1 794
0 796 7 3 2 6076 795
0 797 5 1 1 6078
0 798 7 2 2 5336 6079
0 799 7 2 2 6054 6081
0 800 5 2 1 6083
0 801 7 1 2 791 6085
0 802 5 2 1 801
0 803 7 1 2 6062 6067
0 804 5 1 1 803
0 805 7 1 2 6058 804
0 806 5 1 1 805
0 807 7 3 2 6064 806
0 808 5 1 1 6089
0 809 7 2 2 6087 808
0 810 5 2 1 6092
0 811 7 1 2 5337 6094
0 812 5 2 1 811
0 813 7 1 2 4963 6093
0 814 5 1 1 813
0 815 7 3 2 6096 814
0 816 5 1 1 6098
0 817 7 1 2 760 6077
0 818 5 1 1 817
0 819 7 1 2 6073 818
0 820 5 1 1 819
0 821 7 1 2 6082 6095
0 822 5 2 1 821
0 823 7 1 2 820 6101
0 824 5 1 1 823
0 825 7 1 2 6084 6090
0 826 5 1 1 825
0 827 7 2 2 824 826
0 828 5 1 1 6103
0 829 7 2 2 5328 6099
0 830 7 2 2 6080 6105
0 831 5 2 1 6107
0 832 7 1 2 828 6109
0 833 5 2 1 832
0 834 7 1 2 6086 6091
0 835 5 1 1 834
0 836 7 1 2 6075 835
0 837 5 1 1 836
0 838 7 3 2 6088 837
0 839 5 1 1 6113
0 840 7 2 2 6111 839
0 841 5 2 1 6116
0 842 7 1 2 5329 6118
0 843 5 2 1 842
0 844 7 1 2 816 6120
0 845 5 1 1 844
0 846 7 1 2 6106 6119
0 847 5 2 1 846
0 848 7 1 2 845 6122
0 849 5 1 1 848
0 850 7 1 2 4955 6117
0 851 5 1 1 850
0 852 7 3 2 6121 851
0 853 5 1 1 6124
0 854 7 2 2 5320 6125
0 855 7 1 2 797 6097
0 856 5 1 1 855
0 857 7 1 2 6102 856
0 858 5 1 1 857
0 859 7 1 2 6123 858
0 860 5 1 1 859
0 861 7 1 2 6108 6114
0 862 5 1 1 861
0 863 7 2 2 860 862
0 864 5 1 1 6129
0 865 7 2 2 6100 6127
0 866 5 2 1 6131
0 867 7 1 2 864 6133
0 868 5 2 1 867
0 869 7 1 2 6110 6115
0 870 5 1 1 869
0 871 7 1 2 6104 870
0 872 5 1 1 871
0 873 7 3 2 6112 872
0 874 5 1 1 6137
0 875 7 2 2 6135 874
0 876 5 2 1 6140
0 877 7 1 2 6128 6142
0 878 5 2 1 877
0 879 7 1 2 849 6144
0 880 5 1 1 879
0 881 7 1 2 6132 6138
0 882 5 1 1 881
0 883 7 2 2 880 882
0 884 5 1 1 6146
0 885 7 1 2 5321 6143
0 886 5 2 1 885
0 887 7 1 2 4947 6141
0 888 5 1 1 887
0 889 7 3 2 6148 888
0 890 5 1 1 6150
0 891 7 2 2 5312 6151
0 892 7 2 2 6126 6153
0 893 5 2 1 6155
0 894 7 1 2 884 6157
0 895 5 2 1 894
0 896 7 1 2 6134 6139
0 897 5 1 1 896
0 898 7 1 2 6130 897
0 899 5 1 1 898
0 900 7 3 2 6136 899
0 901 5 1 1 6161
0 902 7 2 2 6159 901
0 903 5 2 1 6164
0 904 7 1 2 5313 6166
0 905 5 2 1 904
0 906 7 1 2 4939 6165
0 907 5 1 1 906
0 908 7 3 2 6168 907
0 909 5 1 1 6170
0 910 7 1 2 853 6149
0 911 5 1 1 910
0 912 7 1 2 6145 911
0 913 5 1 1 912
0 914 7 1 2 6154 6167
0 915 5 2 1 914
0 916 7 1 2 913 6173
0 917 5 1 1 916
0 918 7 1 2 6156 6162
0 919 5 1 1 918
0 920 7 2 2 917 919
0 921 5 1 1 6175
0 922 7 2 2 5305 6171
0 923 7 2 2 6152 6177
0 924 5 2 1 6179
0 925 7 1 2 921 6181
0 926 5 2 1 925
0 927 7 1 2 6158 6163
0 928 5 1 1 927
0 929 7 1 2 6147 928
0 930 5 1 1 929
0 931 7 3 2 6160 930
0 932 5 1 1 6185
0 933 7 2 2 6183 932
0 934 5 2 1 6188
0 935 7 1 2 5306 6190
0 936 5 2 1 935
0 937 7 1 2 909 6192
0 938 5 1 1 937
0 939 7 1 2 6178 6191
0 940 5 2 1 939
0 941 7 1 2 938 6194
0 942 5 1 1 941
0 943 7 1 2 4931 6189
0 944 5 1 1 943
0 945 7 3 2 6193 944
0 946 5 1 1 6196
0 947 7 2 2 5298 6197
0 948 7 1 2 890 6169
0 949 5 1 1 948
0 950 7 1 2 6174 949
0 951 5 1 1 950
0 952 7 1 2 6195 951
0 953 5 1 1 952
0 954 7 1 2 6180 6186
0 955 5 1 1 954
0 956 7 2 2 953 955
0 957 5 1 1 6201
0 958 7 2 2 6172 6199
0 959 5 2 1 6203
0 960 7 1 2 957 6205
0 961 5 2 1 960
0 962 7 1 2 6182 6187
0 963 5 1 1 962
0 964 7 1 2 6176 963
0 965 5 1 1 964
0 966 7 3 2 6184 965
0 967 5 1 1 6209
0 968 7 2 2 6207 967
0 969 5 2 1 6212
0 970 7 1 2 6200 6214
0 971 5 2 1 970
0 972 7 1 2 942 6216
0 973 5 1 1 972
0 974 7 1 2 6204 6210
0 975 5 1 1 974
0 976 7 2 2 973 975
0 977 5 1 1 6218
0 978 7 1 2 5299 6215
0 979 5 2 1 978
0 980 7 1 2 4923 6213
0 981 5 1 1 980
0 982 7 3 2 6220 981
0 983 5 1 1 6222
0 984 7 2 2 5291 6223
0 985 7 2 2 6198 6225
0 986 5 2 1 6227
0 987 7 1 2 977 6229
0 988 5 2 1 987
0 989 7 1 2 6206 6211
0 990 5 1 1 989
0 991 7 1 2 6202 990
0 992 5 1 1 991
0 993 7 3 2 6208 992
0 994 5 1 1 6233
0 995 7 2 2 6231 994
0 996 5 2 1 6236
0 997 7 1 2 5292 6238
0 998 5 2 1 997
0 999 7 1 2 4915 6237
0 1000 5 1 1 999
0 1001 7 3 2 6240 1000
0 1002 5 1 1 6242
0 1003 7 1 2 946 6221
0 1004 5 1 1 1003
0 1005 7 1 2 6217 1004
0 1006 5 1 1 1005
0 1007 7 1 2 6226 6239
0 1008 5 2 1 1007
0 1009 7 1 2 1006 6245
0 1010 5 1 1 1009
0 1011 7 1 2 6228 6234
0 1012 5 1 1 1011
0 1013 7 2 2 1010 1012
0 1014 5 1 1 6247
0 1015 7 2 2 5284 6243
0 1016 7 2 2 6224 6249
0 1017 5 2 1 6251
0 1018 7 1 2 1014 6253
0 1019 5 2 1 1018
0 1020 7 1 2 6230 6235
0 1021 5 1 1 1020
0 1022 7 1 2 6219 1021
0 1023 5 1 1 1022
0 1024 7 3 2 6232 1023
0 1025 5 1 1 6257
0 1026 7 2 2 6255 1025
0 1027 5 2 1 6260
0 1028 7 1 2 5285 6262
0 1029 5 2 1 1028
0 1030 7 1 2 1002 6264
0 1031 5 1 1 1030
0 1032 7 1 2 6250 6263
0 1033 5 2 1 1032
0 1034 7 1 2 1031 6266
0 1035 5 1 1 1034
0 1036 7 1 2 4907 6261
0 1037 5 1 1 1036
0 1038 7 3 2 6265 1037
0 1039 5 1 1 6268
0 1040 7 2 2 5277 6269
0 1041 7 1 2 983 6241
0 1042 5 1 1 1041
0 1043 7 1 2 6246 1042
0 1044 5 1 1 1043
0 1045 7 1 2 6267 1044
0 1046 5 1 1 1045
0 1047 7 1 2 6252 6258
0 1048 5 1 1 1047
0 1049 7 2 2 1046 1048
0 1050 5 1 1 6273
0 1051 7 2 2 6244 6271
0 1052 5 2 1 6275
0 1053 7 1 2 1050 6277
0 1054 5 2 1 1053
0 1055 7 1 2 6254 6259
0 1056 5 1 1 1055
0 1057 7 1 2 6248 1056
0 1058 5 1 1 1057
0 1059 7 3 2 6256 1058
0 1060 5 1 1 6281
0 1061 7 2 2 6279 1060
0 1062 5 2 1 6284
0 1063 7 1 2 6272 6286
0 1064 5 2 1 1063
0 1065 7 1 2 1035 6288
0 1066 5 1 1 1065
0 1067 7 1 2 6276 6282
0 1068 5 1 1 1067
0 1069 7 2 2 1066 1068
0 1070 5 1 1 6290
0 1071 7 1 2 5278 6287
0 1072 5 2 1 1071
0 1073 7 1 2 4899 6285
0 1074 5 1 1 1073
0 1075 7 3 2 6292 1074
0 1076 5 1 1 6294
0 1077 7 2 2 5270 6295
0 1078 7 2 2 6270 6297
0 1079 5 2 1 6299
0 1080 7 1 2 1070 6301
0 1081 5 2 1 1080
0 1082 7 1 2 6278 6283
0 1083 5 1 1 1082
0 1084 7 1 2 6274 1083
0 1085 5 1 1 1084
0 1086 7 3 2 6280 1085
0 1087 5 1 1 6305
0 1088 7 2 2 6303 1087
0 1089 5 2 1 6308
0 1090 7 1 2 5271 6310
0 1091 5 2 1 1090
0 1092 7 1 2 4891 6309
0 1093 5 1 1 1092
0 1094 7 3 2 6312 1093
0 1095 5 1 1 6314
0 1096 7 1 2 1039 6293
0 1097 5 1 1 1096
0 1098 7 1 2 6289 1097
0 1099 5 1 1 1098
0 1100 7 1 2 6298 6311
0 1101 5 2 1 1100
0 1102 7 1 2 1099 6317
0 1103 5 1 1 1102
0 1104 7 1 2 6300 6306
0 1105 5 1 1 1104
0 1106 7 2 2 1103 1105
0 1107 5 1 1 6319
0 1108 7 2 2 5263 6315
0 1109 7 2 2 6296 6321
0 1110 5 2 1 6323
0 1111 7 1 2 1107 6325
0 1112 5 2 1 1111
0 1113 7 1 2 6302 6307
0 1114 5 1 1 1113
0 1115 7 1 2 6291 1114
0 1116 5 1 1 1115
0 1117 7 3 2 6304 1116
0 1118 5 1 1 6329
0 1119 7 2 2 6327 1118
0 1120 5 2 1 6332
0 1121 7 1 2 5264 6334
0 1122 5 2 1 1121
0 1123 7 1 2 1095 6336
0 1124 5 1 1 1123
0 1125 7 1 2 6322 6335
0 1126 5 2 1 1125
0 1127 7 1 2 1124 6338
0 1128 5 1 1 1127
0 1129 7 1 2 4883 6333
0 1130 5 1 1 1129
0 1131 7 3 2 6337 1130
0 1132 5 1 1 6340
0 1133 7 2 2 5256 6341
0 1134 7 1 2 1076 6313
0 1135 5 1 1 1134
0 1136 7 1 2 6318 1135
0 1137 5 1 1 1136
0 1138 7 1 2 6339 1137
0 1139 5 1 1 1138
0 1140 7 1 2 6324 6330
0 1141 5 1 1 1140
0 1142 7 2 2 1139 1141
0 1143 5 1 1 6345
0 1144 7 2 2 6316 6343
0 1145 5 2 1 6347
0 1146 7 1 2 1143 6349
0 1147 5 2 1 1146
0 1148 7 1 2 6326 6331
0 1149 5 1 1 1148
0 1150 7 1 2 6320 1149
0 1151 5 1 1 1150
0 1152 7 3 2 6328 1151
0 1153 5 1 1 6353
0 1154 7 2 2 6351 1153
0 1155 5 2 1 6356
0 1156 7 1 2 6344 6358
0 1157 5 2 1 1156
0 1158 7 1 2 1128 6360
0 1159 5 1 1 1158
0 1160 7 1 2 6348 6354
0 1161 5 1 1 1160
0 1162 7 2 2 1159 1161
0 1163 5 1 1 6362
0 1164 7 1 2 5257 6359
0 1165 5 2 1 1164
0 1166 7 1 2 4875 6357
0 1167 5 1 1 1166
0 1168 7 3 2 6364 1167
0 1169 5 1 1 6366
0 1170 7 2 2 5249 6367
0 1171 7 2 2 6342 6369
0 1172 5 2 1 6371
0 1173 7 1 2 1163 6373
0 1174 5 2 1 1173
0 1175 7 1 2 6350 6355
0 1176 5 1 1 1175
0 1177 7 1 2 6346 1176
0 1178 5 1 1 1177
0 1179 7 3 2 6352 1178
0 1180 5 1 1 6377
0 1181 7 2 2 6375 1180
0 1182 5 2 1 6380
0 1183 7 1 2 5250 6382
0 1184 5 2 1 1183
0 1185 7 1 2 4867 6381
0 1186 5 1 1 1185
0 1187 7 3 2 6384 1186
0 1188 5 1 1 6386
0 1189 7 1 2 1132 6365
0 1190 5 1 1 1189
0 1191 7 1 2 6361 1190
0 1192 5 1 1 1191
0 1193 7 1 2 6370 6383
0 1194 5 2 1 1193
0 1195 7 1 2 1192 6389
0 1196 5 1 1 1195
0 1197 7 1 2 6372 6378
0 1198 5 1 1 1197
0 1199 7 2 2 1196 1198
0 1200 5 1 1 6391
0 1201 7 2 2 5242 6387
0 1202 7 2 2 6368 6393
0 1203 5 2 1 6395
0 1204 7 1 2 1200 6397
0 1205 5 2 1 1204
0 1206 7 1 2 6374 6379
0 1207 5 1 1 1206
0 1208 7 1 2 6363 1207
0 1209 5 1 1 1208
0 1210 7 3 2 6376 1209
0 1211 5 1 1 6401
0 1212 7 2 2 6399 1211
0 1213 5 2 1 6404
0 1214 7 1 2 5243 6406
0 1215 5 2 1 1214
0 1216 7 1 2 1188 6408
0 1217 5 1 1 1216
0 1218 7 1 2 6394 6407
0 1219 5 2 1 1218
0 1220 7 1 2 1217 6410
0 1221 5 1 1 1220
0 1222 7 1 2 4859 6405
0 1223 5 1 1 1222
0 1224 7 3 2 6409 1223
0 1225 5 1 1 6412
0 1226 7 2 2 5235 6413
0 1227 7 1 2 1169 6385
0 1228 5 1 1 1227
0 1229 7 1 2 6390 1228
0 1230 5 1 1 1229
0 1231 7 1 2 6411 1230
0 1232 5 1 1 1231
0 1233 7 1 2 6396 6402
0 1234 5 1 1 1233
0 1235 7 2 2 1232 1234
0 1236 5 1 1 6417
0 1237 7 2 2 6388 6415
0 1238 5 2 1 6419
0 1239 7 1 2 1236 6421
0 1240 5 2 1 1239
0 1241 7 1 2 6398 6403
0 1242 5 1 1 1241
0 1243 7 1 2 6392 1242
0 1244 5 1 1 1243
0 1245 7 3 2 6400 1244
0 1246 5 1 1 6425
0 1247 7 2 2 6423 1246
0 1248 5 2 1 6428
0 1249 7 1 2 6416 6430
0 1250 5 2 1 1249
0 1251 7 1 2 1221 6432
0 1252 5 1 1 1251
0 1253 7 1 2 6420 6426
0 1254 5 1 1 1253
0 1255 7 2 2 1252 1254
0 1256 5 1 1 6434
0 1257 7 1 2 5236 6431
0 1258 5 2 1 1257
0 1259 7 1 2 4851 6429
0 1260 5 1 1 1259
0 1261 7 3 2 6436 1260
0 1262 5 1 1 6438
0 1263 7 2 2 5228 6439
0 1264 7 2 2 6414 6441
0 1265 5 2 1 6443
0 1266 7 1 2 1256 6445
0 1267 5 2 1 1266
0 1268 7 1 2 6422 6427
0 1269 5 1 1 1268
0 1270 7 1 2 6418 1269
0 1271 5 1 1 1270
0 1272 7 3 2 6424 1271
0 1273 5 1 1 6449
0 1274 7 2 2 6447 1273
0 1275 5 2 1 6452
0 1276 7 1 2 5229 6454
0 1277 5 2 1 1276
0 1278 7 1 2 4843 6453
0 1279 5 1 1 1278
0 1280 7 3 2 6456 1279
0 1281 5 1 1 6458
0 1282 7 1 2 1225 6437
0 1283 5 1 1 1282
0 1284 7 1 2 6433 1283
0 1285 5 1 1 1284
0 1286 7 1 2 6442 6455
0 1287 5 2 1 1286
0 1288 7 1 2 1285 6461
0 1289 5 1 1 1288
0 1290 7 1 2 6444 6450
0 1291 5 1 1 1290
0 1292 7 2 2 1289 1291
0 1293 5 1 1 6463
0 1294 7 2 2 5221 6459
0 1295 7 2 2 6440 6465
0 1296 5 2 1 6467
0 1297 7 1 2 1293 6469
0 1298 5 2 1 1297
0 1299 7 1 2 6446 6451
0 1300 5 1 1 1299
0 1301 7 1 2 6435 1300
0 1302 5 1 1 1301
0 1303 7 3 2 6448 1302
0 1304 5 1 1 6473
0 1305 7 2 2 6471 1304
0 1306 5 2 1 6476
0 1307 7 1 2 5222 6478
0 1308 5 2 1 1307
0 1309 7 1 2 1281 6480
0 1310 5 1 1 1309
0 1311 7 1 2 6466 6479
0 1312 5 2 1 1311
0 1313 7 1 2 1310 6482
0 1314 5 1 1 1313
0 1315 7 1 2 4835 6477
0 1316 5 1 1 1315
0 1317 7 3 2 6481 1316
0 1318 5 1 1 6484
0 1319 7 2 2 5214 6485
0 1320 7 1 2 1262 6457
0 1321 5 1 1 1320
0 1322 7 1 2 6462 1321
0 1323 5 1 1 1322
0 1324 7 1 2 6483 1323
0 1325 5 1 1 1324
0 1326 7 1 2 6468 6474
0 1327 5 1 1 1326
0 1328 7 2 2 1325 1327
0 1329 5 1 1 6489
0 1330 7 2 2 6460 6487
0 1331 5 2 1 6491
0 1332 7 1 2 1329 6493
0 1333 5 2 1 1332
0 1334 7 1 2 6470 6475
0 1335 5 1 1 1334
0 1336 7 1 2 6464 1335
0 1337 5 1 1 1336
0 1338 7 3 2 6472 1337
0 1339 5 1 1 6497
0 1340 7 2 2 6495 1339
0 1341 5 2 1 6500
0 1342 7 1 2 6488 6502
0 1343 5 2 1 1342
0 1344 7 1 2 1314 6504
0 1345 5 1 1 1344
0 1346 7 1 2 6492 6498
0 1347 5 1 1 1346
0 1348 7 2 2 1345 1347
0 1349 5 1 1 6506
0 1350 7 1 2 5215 6503
0 1351 5 2 1 1350
0 1352 7 1 2 4827 6501
0 1353 5 1 1 1352
0 1354 7 3 2 6508 1353
0 1355 5 1 1 6510
0 1356 7 2 2 5207 6511
0 1357 7 2 2 6486 6513
0 1358 5 2 1 6515
0 1359 7 1 2 1349 6517
0 1360 5 2 1 1359
0 1361 7 1 2 6494 6499
0 1362 5 1 1 1361
0 1363 7 1 2 6490 1362
0 1364 5 1 1 1363
0 1365 7 3 2 6496 1364
0 1366 5 1 1 6521
0 1367 7 2 2 6519 1366
0 1368 5 2 1 6524
0 1369 7 1 2 5208 6526
0 1370 5 2 1 1369
0 1371 7 1 2 4819 6525
0 1372 5 1 1 1371
0 1373 7 3 2 6528 1372
0 1374 5 1 1 6530
0 1375 7 1 2 1318 6509
0 1376 5 1 1 1375
0 1377 7 1 2 6505 1376
0 1378 5 1 1 1377
0 1379 7 1 2 6514 6527
0 1380 5 2 1 1379
0 1381 7 1 2 1378 6533
0 1382 5 1 1 1381
0 1383 7 1 2 6516 6522
0 1384 5 1 1 1383
0 1385 7 2 2 1382 1384
0 1386 5 1 1 6535
0 1387 7 2 2 5200 6531
0 1388 7 2 2 6512 6537
0 1389 5 2 1 6539
0 1390 7 1 2 1386 6541
0 1391 5 2 1 1390
0 1392 7 1 2 6518 6523
0 1393 5 1 1 1392
0 1394 7 1 2 6507 1393
0 1395 5 1 1 1394
0 1396 7 3 2 6520 1395
0 1397 5 1 1 6545
0 1398 7 2 2 6543 1397
0 1399 5 2 1 6548
0 1400 7 1 2 5201 6550
0 1401 5 2 1 1400
0 1402 7 1 2 4811 6549
0 1403 5 1 1 1402
0 1404 7 3 2 6552 1403
0 1405 5 1 1 6554
0 1406 7 2 2 5193 6555
0 1407 7 1 2 6532 6557
0 1408 5 2 1 1407
0 1409 7 1 2 1355 6529
0 1410 5 1 1 1409
0 1411 7 1 2 6534 1410
0 1412 5 1 1 1411
0 1413 7 1 2 6538 6551
0 1414 5 2 1 1413
0 1415 7 1 2 1412 6561
0 1416 5 1 1 1415
0 1417 7 1 2 6540 6546
0 1418 5 1 1 1417
0 1419 7 2 2 1416 1418
0 1420 5 1 1 6563
0 1421 7 1 2 6559 1420
0 1422 5 2 1 1421
0 1423 7 1 2 6542 6547
0 1424 5 1 1 1423
0 1425 7 1 2 6536 1424
0 1426 5 1 1 1425
0 1427 7 2 2 6544 1426
0 1428 5 1 1 6567
0 1429 7 1 2 6560 6568
0 1430 5 1 1 1429
0 1431 7 1 2 6564 1430
0 1432 5 1 1 1431
0 1433 7 2 2 6565 1432
0 1434 5 2 1 6569
0 1435 7 1 2 1374 6553
0 1436 5 1 1 1435
0 1437 7 2 2 6562 1436
0 1438 5 1 1 6573
0 1439 7 2 2 6566 1428
0 1440 5 2 1 6575
0 1441 7 2 2 6558 6577
0 1442 5 1 1 6579
0 1443 7 1 2 1438 6580
0 1444 5 1 1 1443
0 1445 7 1 2 6574 1442
0 1446 5 1 1 1445
0 1447 7 1 2 1444 1446
0 1448 5 2 1 1447
0 1449 7 1 2 6571 6581
0 1450 5 1 1 1449
0 1451 7 1 2 5187 1450
0 1452 5 1 1 1451
0 1453 7 1 2 4788 6570
0 1454 5 1 1 1453
0 1455 7 1 2 5188 6572
0 1456 5 1 1 1455
0 1457 7 1 2 1454 1456
0 1458 7 1 2 6582 1457
0 1459 5 1 1 1458
0 1460 7 1 2 5180 6556
0 1461 5 1 1 1460
0 1462 7 1 2 4789 1405
0 1463 5 1 1 1462
0 1464 7 1 2 1461 1463
0 1465 5 1 1 1464
0 1466 7 1 2 4802 6578
0 1467 5 1 1 1466
0 1468 7 1 2 5194 6576
0 1469 5 1 1 1468
0 1470 7 1 2 1467 1469
0 1471 5 1 1 1470
0 1472 7 1 2 1465 1471
0 1473 7 1 2 1459 1472
0 1474 7 1 2 1452 1473
0 1475 5 1 1 1474
0 1476 7 3 2 5158 5168
0 1477 5 1 1 6583
0 1478 7 1 2 5177 1477
0 1479 5 2 1 1478
0 1480 7 1 2 5510 6586
0 1481 5 1 1 1480
0 1482 7 2 2 5525 6584
0 1483 5 1 1 6588
0 1484 7 1 2 1483 6587
0 1485 5 1 1 1484
0 1486 7 2 2 5148 1485
0 1487 5 2 1 6590
0 1488 7 4 2 1481 6592
0 1489 5 1 1 6594
0 1490 7 1 2 5178 6585
0 1491 5 2 1 1490
0 1492 7 1 2 5159 6598
0 1493 5 1 1 1492
0 1494 7 1 2 6593 1493
0 1495 5 1 1 1494
0 1496 7 1 2 5160 6591
0 1497 5 1 1 1496
0 1498 7 2 2 1495 1497
0 1499 5 1 1 6600
0 1500 7 1 2 5140 6595
0 1501 7 1 2 6601 1500
0 1502 5 2 1 1501
0 1503 7 2 2 5149 5161
0 1504 5 1 1 6604
0 1505 7 1 2 5526 6605
0 1506 5 1 1 1505
0 1507 7 1 2 5522 1504
0 1508 5 1 1 1507
0 1509 7 1 2 6599 1508
0 1510 7 1 2 1506 1509
0 1511 5 2 1 1510
0 1512 7 1 2 6602 6606
0 1513 5 1 1 1512
0 1514 7 2 2 5141 1513
0 1515 5 2 1 6608
0 1516 7 1 2 5503 6607
0 1517 5 1 1 1516
0 1518 7 3 2 6610 1517
0 1519 5 1 1 6612
0 1520 7 2 2 5132 6613
0 1521 7 1 2 6596 6615
0 1522 5 2 1 1521
0 1523 7 1 2 6597 6609
0 1524 5 2 1 1523
0 1525 7 1 2 1489 6611
0 1526 5 1 1 1525
0 1527 7 1 2 6619 1526
0 1528 5 1 1 1527
0 1529 7 1 2 1499 6620
0 1530 5 1 1 1529
0 1531 7 2 2 6603 1530
0 1532 5 2 1 6621
0 1533 7 1 2 6616 6622
0 1534 5 1 1 1533
0 1535 7 1 2 1528 1534
0 1536 5 1 1 1535
0 1537 7 1 2 6617 1536
0 1538 5 2 1 1537
0 1539 7 1 2 6618 6623
0 1540 5 1 1 1539
0 1541 7 2 2 5133 1540
0 1542 5 2 1 6627
0 1543 7 1 2 6614 6629
0 1544 5 1 1 1543
0 1545 7 1 2 1519 6628
0 1546 5 1 1 1545
0 1547 7 2 2 1544 1546
0 1548 5 1 1 6631
0 1549 7 1 2 5495 6624
0 1550 5 1 1 1549
0 1551 7 4 2 6630 1550
0 1552 5 1 1 6633
0 1553 7 1 2 5124 6634
0 1554 7 1 2 1548 1553
0 1555 5 2 1 1554
0 1556 7 1 2 6625 6637
0 1557 5 1 1 1556
0 1558 7 2 2 5125 1557
0 1559 5 2 1 6639
0 1560 7 1 2 5488 6626
0 1561 5 1 1 1560
0 1562 7 3 2 6641 1561
0 1563 5 1 1 6643
0 1564 7 1 2 6635 6640
0 1565 5 2 1 1564
0 1566 7 1 2 6632 6646
0 1567 5 1 1 1566
0 1568 7 1 2 6638 1567
0 1569 5 2 1 1568
0 1570 7 2 2 5116 6644
0 1571 7 1 2 6636 6650
0 1572 5 2 1 1571
0 1573 7 1 2 6648 6652
0 1574 5 2 1 1573
0 1575 7 1 2 5117 6654
0 1576 5 2 1 1575
0 1577 7 1 2 5481 6649
0 1578 5 1 1 1577
0 1579 7 4 2 6656 1578
0 1580 5 1 1 6658
0 1581 7 2 2 5108 6659
0 1582 7 1 2 6645 6662
0 1583 5 2 1 1582
0 1584 7 1 2 1563 6657
0 1585 5 1 1 1584
0 1586 7 1 2 6651 6655
0 1587 5 2 1 1586
0 1588 7 1 2 1585 6666
0 1589 5 1 1 1588
0 1590 7 1 2 1552 6642
0 1591 5 1 1 1590
0 1592 7 1 2 6647 1591
0 1593 5 1 1 1592
0 1594 7 1 2 6667 1593
0 1595 5 1 1 1594
0 1596 7 2 2 6653 1595
0 1597 5 2 1 6668
0 1598 7 1 2 6663 6669
0 1599 5 1 1 1598
0 1600 7 1 2 1589 1599
0 1601 5 1 1 1600
0 1602 7 1 2 6664 1601
0 1603 5 2 1 1602
0 1604 7 1 2 6665 6670
0 1605 5 1 1 1604
0 1606 7 2 2 5109 1605
0 1607 5 2 1 6674
0 1608 7 1 2 5474 6671
0 1609 5 1 1 1608
0 1610 7 2 2 6676 1609
0 1611 5 1 1 6678
0 1612 7 2 2 5100 6679
0 1613 7 1 2 6660 6680
0 1614 5 2 1 1613
0 1615 7 1 2 6672 6682
0 1616 5 2 1 1615
0 1617 7 1 2 5101 6684
0 1618 5 2 1 1617
0 1619 7 1 2 5467 6673
0 1620 5 1 1 1619
0 1621 7 4 2 6686 1620
0 1622 5 1 1 6688
0 1623 7 1 2 1611 6687
0 1624 5 1 1 1623
0 1625 7 1 2 6681 6685
0 1626 5 2 1 1625
0 1627 7 2 2 1624 6692
0 1628 5 1 1 6694
0 1629 7 1 2 5092 6689
0 1630 7 1 2 6695 1629
0 1631 5 2 1 1630
0 1632 7 1 2 6661 6677
0 1633 5 1 1 1632
0 1634 7 1 2 1580 6675
0 1635 5 1 1 1634
0 1636 7 1 2 1633 1635
0 1637 7 1 2 6693 1636
0 1638 5 1 1 1637
0 1639 7 1 2 6683 1638
0 1640 5 2 1 1639
0 1641 7 1 2 6696 6698
0 1642 5 1 1 1641
0 1643 7 2 2 5093 1642
0 1644 5 2 1 6700
0 1645 7 1 2 5460 6699
0 1646 5 1 1 1645
0 1647 7 3 2 6702 1646
0 1648 5 1 1 6704
0 1649 7 2 2 5084 6705
0 1650 7 1 2 6690 6707
0 1651 5 2 1 1650
0 1652 7 1 2 6691 6701
0 1653 5 2 1 1652
0 1654 7 1 2 1622 6703
0 1655 5 1 1 1654
0 1656 7 1 2 6711 1655
0 1657 5 1 1 1656
0 1658 7 1 2 1628 6712
0 1659 5 1 1 1658
0 1660 7 2 2 6697 1659
0 1661 5 2 1 6713
0 1662 7 1 2 6708 6714
0 1663 5 1 1 1662
0 1664 7 1 2 1657 1663
0 1665 5 1 1 1664
0 1666 7 1 2 6709 1665
0 1667 5 2 1 1666
0 1668 7 1 2 6710 6715
0 1669 5 1 1 1668
0 1670 7 2 2 5085 1669
0 1671 5 2 1 6719
0 1672 7 1 2 6706 6721
0 1673 5 1 1 1672
0 1674 7 1 2 1648 6720
0 1675 5 1 1 1674
0 1676 7 2 2 1673 1675
0 1677 5 1 1 6723
0 1678 7 1 2 5453 6716
0 1679 5 1 1 1678
0 1680 7 4 2 6722 1679
0 1681 5 1 1 6725
0 1682 7 1 2 5076 6726
0 1683 7 1 2 1677 1682
0 1684 5 2 1 1683
0 1685 7 1 2 6717 6729
0 1686 5 1 1 1685
0 1687 7 2 2 5077 1686
0 1688 5 2 1 6731
0 1689 7 1 2 5446 6718
0 1690 5 1 1 1689
0 1691 7 3 2 6733 1690
0 1692 5 1 1 6735
0 1693 7 1 2 6727 6732
0 1694 5 2 1 1693
0 1695 7 1 2 6724 6738
0 1696 5 1 1 1695
0 1697 7 1 2 6730 1696
0 1698 5 2 1 1697
0 1699 7 2 2 5068 6736
0 1700 7 1 2 6728 6742
0 1701 5 2 1 1700
0 1702 7 1 2 6740 6744
0 1703 5 2 1 1702
0 1704 7 1 2 5069 6746
0 1705 5 2 1 1704
0 1706 7 1 2 5439 6741
0 1707 5 1 1 1706
0 1708 7 4 2 6748 1707
0 1709 5 1 1 6750
0 1710 7 2 2 5060 6751
0 1711 7 1 2 6737 6754
0 1712 5 2 1 1711
0 1713 7 1 2 1692 6749
0 1714 5 1 1 1713
0 1715 7 1 2 6743 6747
0 1716 5 2 1 1715
0 1717 7 1 2 1714 6758
0 1718 5 1 1 1717
0 1719 7 1 2 1681 6734
0 1720 5 1 1 1719
0 1721 7 1 2 6739 1720
0 1722 5 1 1 1721
0 1723 7 1 2 6759 1722
0 1724 5 1 1 1723
0 1725 7 2 2 6745 1724
0 1726 5 2 1 6760
0 1727 7 1 2 6755 6761
0 1728 5 1 1 1727
0 1729 7 1 2 1718 1728
0 1730 5 1 1 1729
0 1731 7 1 2 6756 1730
0 1732 5 2 1 1731
0 1733 7 1 2 6757 6762
0 1734 5 1 1 1733
0 1735 7 2 2 5061 1734
0 1736 5 2 1 6766
0 1737 7 1 2 5432 6763
0 1738 5 1 1 1737
0 1739 7 2 2 6768 1738
0 1740 5 1 1 6770
0 1741 7 2 2 5052 6771
0 1742 7 1 2 6752 6772
0 1743 5 2 1 1742
0 1744 7 1 2 6764 6774
0 1745 5 2 1 1744
0 1746 7 1 2 5053 6776
0 1747 5 2 1 1746
0 1748 7 1 2 5425 6765
0 1749 5 1 1 1748
0 1750 7 4 2 6778 1749
0 1751 5 1 1 6780
0 1752 7 1 2 1740 6779
0 1753 5 1 1 1752
0 1754 7 1 2 6773 6777
0 1755 5 2 1 1754
0 1756 7 2 2 1753 6784
0 1757 5 1 1 6786
0 1758 7 1 2 5044 6781
0 1759 7 1 2 6787 1758
0 1760 5 2 1 1759
0 1761 7 1 2 6753 6769
0 1762 5 1 1 1761
0 1763 7 1 2 1709 6767
0 1764 5 1 1 1763
0 1765 7 1 2 1762 1764
0 1766 7 1 2 6785 1765
0 1767 5 1 1 1766
0 1768 7 1 2 6775 1767
0 1769 5 2 1 1768
0 1770 7 1 2 6788 6790
0 1771 5 1 1 1770
0 1772 7 2 2 5045 1771
0 1773 5 2 1 6792
0 1774 7 1 2 5418 6791
0 1775 5 1 1 1774
0 1776 7 3 2 6794 1775
0 1777 5 1 1 6796
0 1778 7 2 2 5036 6797
0 1779 7 1 2 6782 6799
0 1780 5 2 1 1779
0 1781 7 1 2 6783 6793
0 1782 5 2 1 1781
0 1783 7 1 2 1751 6795
0 1784 5 1 1 1783
0 1785 7 1 2 6803 1784
0 1786 5 1 1 1785
0 1787 7 1 2 1757 6804
0 1788 5 1 1 1787
0 1789 7 2 2 6789 1788
0 1790 5 2 1 6805
0 1791 7 1 2 6800 6806
0 1792 5 1 1 1791
0 1793 7 1 2 1786 1792
0 1794 5 1 1 1793
0 1795 7 1 2 6801 1794
0 1796 5 2 1 1795
0 1797 7 1 2 6802 6807
0 1798 5 1 1 1797
0 1799 7 2 2 5037 1798
0 1800 5 2 1 6811
0 1801 7 1 2 6798 6813
0 1802 5 1 1 1801
0 1803 7 1 2 1777 6812
0 1804 5 1 1 1803
0 1805 7 2 2 1802 1804
0 1806 5 1 1 6815
0 1807 7 1 2 5410 6808
0 1808 5 1 1 1807
0 1809 7 4 2 6814 1808
0 1810 5 1 1 6817
0 1811 7 1 2 5028 6818
0 1812 7 1 2 1806 1811
0 1813 5 2 1 1812
0 1814 7 1 2 6809 6821
0 1815 5 1 1 1814
0 1816 7 2 2 5029 1815
0 1817 5 2 1 6823
0 1818 7 1 2 5402 6810
0 1819 5 1 1 1818
0 1820 7 3 2 6825 1819
0 1821 5 1 1 6827
0 1822 7 1 2 6819 6824
0 1823 5 2 1 1822
0 1824 7 1 2 6816 6830
0 1825 5 1 1 1824
0 1826 7 1 2 6822 1825
0 1827 5 2 1 1826
0 1828 7 2 2 5020 6828
0 1829 7 1 2 6820 6834
0 1830 5 2 1 1829
0 1831 7 1 2 6832 6836
0 1832 5 2 1 1831
0 1833 7 1 2 5021 6838
0 1834 5 2 1 1833
0 1835 7 1 2 5394 6833
0 1836 5 1 1 1835
0 1837 7 4 2 6840 1836
0 1838 5 1 1 6842
0 1839 7 2 2 5012 6843
0 1840 7 1 2 6829 6846
0 1841 5 2 1 1840
0 1842 7 1 2 1821 6841
0 1843 5 1 1 1842
0 1844 7 1 2 6835 6839
0 1845 5 2 1 1844
0 1846 7 1 2 1843 6850
0 1847 5 1 1 1846
0 1848 7 1 2 1810 6826
0 1849 5 1 1 1848
0 1850 7 1 2 6831 1849
0 1851 5 1 1 1850
0 1852 7 1 2 6851 1851
0 1853 5 1 1 1852
0 1854 7 2 2 6837 1853
0 1855 5 2 1 6852
0 1856 7 1 2 6847 6853
0 1857 5 1 1 1856
0 1858 7 1 2 1847 1857
0 1859 5 1 1 1858
0 1860 7 1 2 6848 1859
0 1861 5 2 1 1860
0 1862 7 1 2 6849 6854
0 1863 5 1 1 1862
0 1864 7 2 2 5013 1863
0 1865 5 2 1 6858
0 1866 7 1 2 5386 6855
0 1867 5 1 1 1866
0 1868 7 2 2 6860 1867
0 1869 5 1 1 6862
0 1870 7 2 2 5004 6863
0 1871 7 1 2 6844 6864
0 1872 5 2 1 1871
0 1873 7 1 2 6856 6866
0 1874 5 2 1 1873
0 1875 7 1 2 5005 6868
0 1876 5 2 1 1875
0 1877 7 1 2 5378 6857
0 1878 5 1 1 1877
0 1879 7 4 2 6870 1878
0 1880 5 1 1 6872
0 1881 7 1 2 1869 6871
0 1882 5 1 1 1881
0 1883 7 1 2 6865 6869
0 1884 5 2 1 1883
0 1885 7 2 2 1882 6876
0 1886 5 1 1 6878
0 1887 7 1 2 4996 6873
0 1888 7 1 2 6879 1887
0 1889 5 2 1 1888
0 1890 7 1 2 6845 6861
0 1891 5 1 1 1890
0 1892 7 1 2 1838 6859
0 1893 5 1 1 1892
0 1894 7 1 2 1891 1893
0 1895 7 1 2 6877 1894
0 1896 5 1 1 1895
0 1897 7 1 2 6867 1896
0 1898 5 2 1 1897
0 1899 7 1 2 6880 6882
0 1900 5 1 1 1899
0 1901 7 2 2 4997 1900
0 1902 5 2 1 6884
0 1903 7 1 2 5370 6883
0 1904 5 1 1 1903
0 1905 7 3 2 6886 1904
0 1906 5 1 1 6888
0 1907 7 2 2 4988 6889
0 1908 7 1 2 6874 6891
0 1909 5 2 1 1908
0 1910 7 1 2 6875 6885
0 1911 5 2 1 1910
0 1912 7 1 2 1880 6887
0 1913 5 1 1 1912
0 1914 7 1 2 6895 1913
0 1915 5 1 1 1914
0 1916 7 1 2 1886 6896
0 1917 5 1 1 1916
0 1918 7 2 2 6881 1917
0 1919 5 2 1 6897
0 1920 7 1 2 6892 6898
0 1921 5 1 1 1920
0 1922 7 1 2 1915 1921
0 1923 5 1 1 1922
0 1924 7 1 2 6893 1923
0 1925 5 2 1 1924
0 1926 7 1 2 6894 6899
0 1927 5 1 1 1926
0 1928 7 2 2 4989 1927
0 1929 5 2 1 6903
0 1930 7 1 2 6890 6905
0 1931 5 1 1 1930
0 1932 7 1 2 1906 6904
0 1933 5 1 1 1932
0 1934 7 2 2 1931 1933
0 1935 5 1 1 6907
0 1936 7 1 2 5362 6900
0 1937 5 1 1 1936
0 1938 7 4 2 6906 1937
0 1939 5 1 1 6909
0 1940 7 1 2 4980 6910
0 1941 7 1 2 1935 1940
0 1942 5 2 1 1941
0 1943 7 1 2 6901 6913
0 1944 5 1 1 1943
0 1945 7 2 2 4981 1944
0 1946 5 2 1 6915
0 1947 7 1 2 5354 6902
0 1948 5 1 1 1947
0 1949 7 3 2 6917 1948
0 1950 5 1 1 6919
0 1951 7 1 2 6911 6916
0 1952 5 2 1 1951
0 1953 7 1 2 6908 6922
0 1954 5 1 1 1953
0 1955 7 1 2 6914 1954
0 1956 5 2 1 1955
0 1957 7 2 2 4972 6920
0 1958 7 1 2 6912 6926
0 1959 5 2 1 1958
0 1960 7 1 2 6924 6928
0 1961 5 2 1 1960
0 1962 7 1 2 4973 6930
0 1963 5 2 1 1962
0 1964 7 1 2 5346 6925
0 1965 5 1 1 1964
0 1966 7 4 2 6932 1965
0 1967 5 1 1 6934
0 1968 7 2 2 4964 6935
0 1969 7 1 2 6921 6938
0 1970 5 2 1 1969
0 1971 7 1 2 1950 6933
0 1972 5 1 1 1971
0 1973 7 1 2 6927 6931
0 1974 5 2 1 1973
0 1975 7 1 2 1972 6942
0 1976 5 1 1 1975
0 1977 7 1 2 1939 6918
0 1978 5 1 1 1977
0 1979 7 1 2 6923 1978
0 1980 5 1 1 1979
0 1981 7 1 2 6943 1980
0 1982 5 1 1 1981
0 1983 7 2 2 6929 1982
0 1984 5 2 1 6944
0 1985 7 1 2 6939 6945
0 1986 5 1 1 1985
0 1987 7 1 2 1976 1986
0 1988 5 1 1 1987
0 1989 7 1 2 6940 1988
0 1990 5 2 1 1989
0 1991 7 1 2 6941 6946
0 1992 5 1 1 1991
0 1993 7 2 2 4965 1992
0 1994 5 2 1 6950
0 1995 7 1 2 5338 6947
0 1996 5 1 1 1995
0 1997 7 2 2 6952 1996
0 1998 5 1 1 6954
0 1999 7 2 2 4956 6955
0 2000 7 1 2 6936 6956
0 2001 5 2 1 2000
0 2002 7 1 2 6948 6958
0 2003 5 2 1 2002
0 2004 7 1 2 4957 6960
0 2005 5 2 1 2004
0 2006 7 1 2 5330 6949
0 2007 5 1 1 2006
0 2008 7 4 2 6962 2007
0 2009 5 1 1 6964
0 2010 7 1 2 1998 6963
0 2011 5 1 1 2010
0 2012 7 1 2 6957 6961
0 2013 5 2 1 2012
0 2014 7 2 2 2011 6968
0 2015 5 1 1 6970
0 2016 7 1 2 4948 6965
0 2017 7 1 2 6971 2016
0 2018 5 2 1 2017
0 2019 7 1 2 6937 6953
0 2020 5 1 1 2019
0 2021 7 1 2 1967 6951
0 2022 5 1 1 2021
0 2023 7 1 2 2020 2022
0 2024 7 1 2 6969 2023
0 2025 5 1 1 2024
0 2026 7 1 2 6959 2025
0 2027 5 2 1 2026
0 2028 7 1 2 6972 6974
0 2029 5 1 1 2028
0 2030 7 2 2 4949 2029
0 2031 5 2 1 6976
0 2032 7 1 2 5322 6975
0 2033 5 1 1 2032
0 2034 7 3 2 6978 2033
0 2035 5 1 1 6980
0 2036 7 2 2 4940 6981
0 2037 7 1 2 6966 6983
0 2038 5 2 1 2037
0 2039 7 1 2 6967 6977
0 2040 5 2 1 2039
0 2041 7 1 2 2009 6979
0 2042 5 1 1 2041
0 2043 7 1 2 6987 2042
0 2044 5 1 1 2043
0 2045 7 1 2 2015 6988
0 2046 5 1 1 2045
0 2047 7 2 2 6973 2046
0 2048 5 2 1 6989
0 2049 7 1 2 6984 6990
0 2050 5 1 1 2049
0 2051 7 1 2 2044 2050
0 2052 5 1 1 2051
0 2053 7 1 2 6985 2052
0 2054 5 2 1 2053
0 2055 7 1 2 6986 6991
0 2056 5 1 1 2055
0 2057 7 2 2 4941 2056
0 2058 5 2 1 6995
0 2059 7 1 2 6982 6997
0 2060 5 1 1 2059
0 2061 7 1 2 2035 6996
0 2062 5 1 1 2061
0 2063 7 2 2 2060 2062
0 2064 5 1 1 6999
0 2065 7 1 2 5314 6992
0 2066 5 1 1 2065
0 2067 7 4 2 6998 2066
0 2068 5 1 1 7001
0 2069 7 1 2 4932 7002
0 2070 7 1 2 2064 2069
0 2071 5 2 1 2070
0 2072 7 1 2 6993 7005
0 2073 5 1 1 2072
0 2074 7 2 2 4933 2073
0 2075 5 2 1 7007
0 2076 7 1 2 5307 6994
0 2077 5 1 1 2076
0 2078 7 3 2 7009 2077
0 2079 5 1 1 7011
0 2080 7 1 2 7003 7008
0 2081 5 2 1 2080
0 2082 7 1 2 7000 7014
0 2083 5 1 1 2082
0 2084 7 1 2 7006 2083
0 2085 5 2 1 2084
0 2086 7 2 2 4924 7012
0 2087 7 1 2 7004 7018
0 2088 5 2 1 2087
0 2089 7 1 2 7016 7020
0 2090 5 2 1 2089
0 2091 7 1 2 4925 7022
0 2092 5 2 1 2091
0 2093 7 1 2 5300 7017
0 2094 5 1 1 2093
0 2095 7 4 2 7024 2094
0 2096 5 1 1 7026
0 2097 7 2 2 4916 7027
0 2098 7 1 2 7013 7030
0 2099 5 2 1 2098
0 2100 7 1 2 2079 7025
0 2101 5 1 1 2100
0 2102 7 1 2 7019 7023
0 2103 5 2 1 2102
0 2104 7 1 2 2101 7034
0 2105 5 1 1 2104
0 2106 7 1 2 2068 7010
0 2107 5 1 1 2106
0 2108 7 1 2 7015 2107
0 2109 5 1 1 2108
0 2110 7 1 2 7035 2109
0 2111 5 1 1 2110
0 2112 7 2 2 7021 2111
0 2113 5 2 1 7036
0 2114 7 1 2 7031 7037
0 2115 5 1 1 2114
0 2116 7 1 2 2105 2115
0 2117 5 1 1 2116
0 2118 7 1 2 7032 2117
0 2119 5 2 1 2118
0 2120 7 1 2 7033 7038
0 2121 5 1 1 2120
0 2122 7 2 2 4917 2121
0 2123 5 2 1 7042
0 2124 7 1 2 5293 7039
0 2125 5 1 1 2124
0 2126 7 2 2 7044 2125
0 2127 5 1 1 7046
0 2128 7 2 2 4908 7047
0 2129 7 1 2 7028 7048
0 2130 5 2 1 2129
0 2131 7 1 2 7040 7050
0 2132 5 2 1 2131
0 2133 7 1 2 4909 7052
0 2134 5 2 1 2133
0 2135 7 1 2 5286 7041
0 2136 5 1 1 2135
0 2137 7 4 2 7054 2136
0 2138 5 1 1 7056
0 2139 7 1 2 2127 7055
0 2140 5 1 1 2139
0 2141 7 1 2 7049 7053
0 2142 5 2 1 2141
0 2143 7 2 2 2140 7060
0 2144 5 1 1 7062
0 2145 7 1 2 4900 7057
0 2146 7 1 2 7063 2145
0 2147 5 2 1 2146
0 2148 7 1 2 7029 7045
0 2149 5 1 1 2148
0 2150 7 1 2 2096 7043
0 2151 5 1 1 2150
0 2152 7 1 2 2149 2151
0 2153 7 1 2 7061 2152
0 2154 5 1 1 2153
0 2155 7 1 2 7051 2154
0 2156 5 2 1 2155
0 2157 7 1 2 7064 7066
0 2158 5 1 1 2157
0 2159 7 2 2 4901 2158
0 2160 5 2 1 7068
0 2161 7 1 2 5279 7067
0 2162 5 1 1 2161
0 2163 7 3 2 7070 2162
0 2164 5 1 1 7072
0 2165 7 2 2 4892 7073
0 2166 7 1 2 7058 7075
0 2167 5 2 1 2166
0 2168 7 1 2 7059 7069
0 2169 5 2 1 2168
0 2170 7 1 2 2138 7071
0 2171 5 1 1 2170
0 2172 7 1 2 7079 2171
0 2173 5 1 1 2172
0 2174 7 1 2 2144 7080
0 2175 5 1 1 2174
0 2176 7 2 2 7065 2175
0 2177 5 2 1 7081
0 2178 7 1 2 7076 7082
0 2179 5 1 1 2178
0 2180 7 1 2 2173 2179
0 2181 5 1 1 2180
0 2182 7 1 2 7077 2181
0 2183 5 2 1 2182
0 2184 7 1 2 7078 7083
0 2185 5 1 1 2184
0 2186 7 2 2 4893 2185
0 2187 5 2 1 7087
0 2188 7 1 2 7074 7089
0 2189 5 1 1 2188
0 2190 7 1 2 2164 7088
0 2191 5 1 1 2190
0 2192 7 2 2 2189 2191
0 2193 5 1 1 7091
0 2194 7 1 2 5272 7084
0 2195 5 1 1 2194
0 2196 7 4 2 7090 2195
0 2197 5 1 1 7093
0 2198 7 1 2 4884 7094
0 2199 7 1 2 2193 2198
0 2200 5 2 1 2199
0 2201 7 1 2 7085 7097
0 2202 5 1 1 2201
0 2203 7 2 2 4885 2202
0 2204 5 2 1 7099
0 2205 7 1 2 5265 7086
0 2206 5 1 1 2205
0 2207 7 3 2 7101 2206
0 2208 5 1 1 7103
0 2209 7 1 2 7095 7100
0 2210 5 2 1 2209
0 2211 7 1 2 7092 7106
0 2212 5 1 1 2211
0 2213 7 1 2 7098 2212
0 2214 5 2 1 2213
0 2215 7 2 2 4876 7104
0 2216 7 1 2 7096 7110
0 2217 5 2 1 2216
0 2218 7 1 2 7108 7112
0 2219 5 2 1 2218
0 2220 7 1 2 4877 7114
0 2221 5 2 1 2220
0 2222 7 1 2 5258 7109
0 2223 5 1 1 2222
0 2224 7 4 2 7116 2223
0 2225 5 1 1 7118
0 2226 7 2 2 4868 7119
0 2227 7 1 2 7105 7122
0 2228 5 2 1 2227
0 2229 7 1 2 2208 7117
0 2230 5 1 1 2229
0 2231 7 1 2 7111 7115
0 2232 5 2 1 2231
0 2233 7 1 2 2230 7126
0 2234 5 1 1 2233
0 2235 7 1 2 2197 7102
0 2236 5 1 1 2235
0 2237 7 1 2 7107 2236
0 2238 5 1 1 2237
0 2239 7 1 2 7127 2238
0 2240 5 1 1 2239
0 2241 7 2 2 7113 2240
0 2242 5 2 1 7128
0 2243 7 1 2 7123 7129
0 2244 5 1 1 2243
0 2245 7 1 2 2234 2244
0 2246 5 1 1 2245
0 2247 7 1 2 7124 2246
0 2248 5 2 1 2247
0 2249 7 1 2 7125 7130
0 2250 5 1 1 2249
0 2251 7 2 2 4869 2250
0 2252 5 2 1 7134
0 2253 7 1 2 5251 7131
0 2254 5 1 1 2253
0 2255 7 2 2 7136 2254
0 2256 5 1 1 7138
0 2257 7 2 2 4860 7139
0 2258 7 1 2 7120 7140
0 2259 5 2 1 2258
0 2260 7 1 2 7132 7142
0 2261 5 2 1 2260
0 2262 7 1 2 4861 7144
0 2263 5 2 1 2262
0 2264 7 1 2 5244 7133
0 2265 5 1 1 2264
0 2266 7 4 2 7146 2265
0 2267 5 1 1 7148
0 2268 7 1 2 2256 7147
0 2269 5 1 1 2268
0 2270 7 1 2 7141 7145
0 2271 5 2 1 2270
0 2272 7 2 2 2269 7152
0 2273 5 1 1 7154
0 2274 7 1 2 4852 7149
0 2275 7 1 2 7155 2274
0 2276 5 2 1 2275
0 2277 7 1 2 7121 7137
0 2278 5 1 1 2277
0 2279 7 1 2 2225 7135
0 2280 5 1 1 2279
0 2281 7 1 2 2278 2280
0 2282 7 1 2 7153 2281
0 2283 5 1 1 2282
0 2284 7 1 2 7143 2283
0 2285 5 2 1 2284
0 2286 7 1 2 7156 7158
0 2287 5 1 1 2286
0 2288 7 2 2 4853 2287
0 2289 5 2 1 7160
0 2290 7 1 2 5237 7159
0 2291 5 1 1 2290
0 2292 7 3 2 7162 2291
0 2293 5 1 1 7164
0 2294 7 2 2 4844 7165
0 2295 7 1 2 7150 7167
0 2296 5 2 1 2295
0 2297 7 1 2 7151 7161
0 2298 5 2 1 2297
0 2299 7 1 2 2267 7163
0 2300 5 1 1 2299
0 2301 7 1 2 7171 2300
0 2302 5 1 1 2301
0 2303 7 1 2 2273 7172
0 2304 5 1 1 2303
0 2305 7 2 2 7157 2304
0 2306 5 2 1 7173
0 2307 7 1 2 7168 7174
0 2308 5 1 1 2307
0 2309 7 1 2 2302 2308
0 2310 5 1 1 2309
0 2311 7 1 2 7169 2310
0 2312 5 2 1 2311
0 2313 7 1 2 7170 7175
0 2314 5 1 1 2313
0 2315 7 2 2 4845 2314
0 2316 5 2 1 7179
0 2317 7 1 2 7166 7181
0 2318 5 1 1 2317
0 2319 7 1 2 2293 7180
0 2320 5 1 1 2319
0 2321 7 2 2 2318 2320
0 2322 5 1 1 7183
0 2323 7 1 2 5230 7176
0 2324 5 1 1 2323
0 2325 7 4 2 7182 2324
0 2326 5 1 1 7185
0 2327 7 1 2 4836 7186
0 2328 7 1 2 2322 2327
0 2329 5 2 1 2328
0 2330 7 1 2 7177 7189
0 2331 5 1 1 2330
0 2332 7 2 2 4837 2331
0 2333 5 2 1 7191
0 2334 7 1 2 5223 7178
0 2335 5 1 1 2334
0 2336 7 3 2 7193 2335
0 2337 5 1 1 7195
0 2338 7 1 2 7187 7192
0 2339 5 2 1 2338
0 2340 7 1 2 7184 7198
0 2341 5 1 1 2340
0 2342 7 1 2 7190 2341
0 2343 5 2 1 2342
0 2344 7 2 2 4828 7196
0 2345 7 1 2 7188 7202
0 2346 5 2 1 2345
0 2347 7 1 2 7200 7204
0 2348 5 2 1 2347
0 2349 7 1 2 4829 7206
0 2350 5 2 1 2349
0 2351 7 1 2 5216 7201
0 2352 5 1 1 2351
0 2353 7 4 2 7208 2352
0 2354 5 1 1 7210
0 2355 7 2 2 4820 7211
0 2356 7 1 2 7197 7214
0 2357 5 2 1 2356
0 2358 7 1 2 7203 7207
0 2359 5 2 1 2358
0 2360 7 1 2 2326 7194
0 2361 5 1 1 2360
0 2362 7 1 2 7199 2361
0 2363 5 1 1 2362
0 2364 7 1 2 7218 2363
0 2365 5 1 1 2364
0 2366 7 2 2 7205 2365
0 2367 5 2 1 7220
0 2368 7 1 2 7216 7222
0 2369 5 1 1 2368
0 2370 7 2 2 4821 2369
0 2371 5 2 1 7224
0 2372 7 1 2 5209 7223
0 2373 5 1 1 2372
0 2374 7 2 2 7226 2373
0 2375 5 1 1 7228
0 2376 7 1 2 2337 7209
0 2377 5 1 1 2376
0 2378 7 1 2 7219 2377
0 2379 5 1 1 2378
0 2380 7 1 2 7215 7221
0 2381 5 1 1 2380
0 2382 7 1 2 2379 2381
0 2383 5 1 1 2382
0 2384 7 1 2 7217 2383
0 2385 5 2 1 2384
0 2386 7 2 2 4812 7229
0 2387 7 1 2 7212 7232
0 2388 5 2 1 2387
0 2389 7 1 2 7230 7234
0 2390 5 2 1 2389
0 2391 7 1 2 4813 7236
0 2392 5 2 1 2391
0 2393 7 1 2 2375 7238
0 2394 5 1 1 2393
0 2395 7 1 2 7233 7237
0 2396 5 2 1 2395
0 2397 7 2 2 2394 7240
0 2398 5 1 1 7242
0 2399 7 1 2 5202 7231
0 2400 5 1 1 2399
0 2401 7 4 2 7239 2400
0 2402 5 1 1 7244
0 2403 7 1 2 4803 7245
0 2404 7 1 2 7243 2403
0 2405 5 2 1 2404
0 2406 7 1 2 7213 7227
0 2407 5 1 1 2406
0 2408 7 1 2 2354 7225
0 2409 5 1 1 2408
0 2410 7 1 2 2407 2409
0 2411 7 1 2 7241 2410
0 2412 5 1 1 2411
0 2413 7 1 2 7235 2412
0 2414 5 2 1 2413
0 2415 7 1 2 7248 7250
0 2416 5 1 1 2415
0 2417 7 2 2 4804 2416
0 2418 5 2 1 7252
0 2419 7 1 2 5195 7251
0 2420 5 1 1 2419
0 2421 7 3 2 7254 2420
0 2422 5 1 1 7256
0 2423 7 1 2 7246 7253
0 2424 5 2 1 2423
0 2425 7 1 2 2398 7259
0 2426 5 1 1 2425
0 2427 7 2 2 7249 2426
0 2428 5 2 1 7261
0 2429 7 2 2 4794 7257
0 2430 7 1 2 7247 7265
0 2431 5 2 1 2430
0 2432 7 1 2 7263 7267
0 2433 5 1 1 2432
0 2434 7 2 2 4795 2433
0 2435 5 2 1 7269
0 2436 7 1 2 7258 7271
0 2437 5 1 1 2436
0 2438 7 1 2 2422 7270
0 2439 5 1 1 2438
0 2440 7 2 2 2437 2439
0 2441 5 1 1 7273
0 2442 7 1 2 2402 7255
0 2443 5 1 1 2442
0 2444 7 1 2 7260 2443
0 2445 5 1 1 2444
0 2446 7 1 2 7262 7266
0 2447 5 1 1 2446
0 2448 7 1 2 2445 2447
0 2449 5 1 1 2448
0 2450 7 1 2 7268 2449
0 2451 5 1 1 2450
0 2452 7 1 2 5181 2451
0 2453 5 1 1 2452
0 2454 7 1 2 7274 2453
0 2455 5 1 1 2454
0 2456 7 1 2 5189 7264
0 2457 5 1 1 2456
0 2458 7 2 2 7272 2457
0 2459 5 1 1 7275
0 2460 7 1 2 5182 7276
0 2461 5 1 1 2460
0 2462 7 1 2 2459 2441
0 2463 5 1 1 2462
0 2464 7 1 2 2461 2463
0 2465 7 1 2 2455 2464
0 2466 5 1 1 2465
0 2467 7 1 2 5162 5527
0 2468 5 1 1 2467
0 2469 7 2 2 5536 2468
0 2470 7 2 2 5511 7277
0 2471 5 1 1 7279
0 2472 7 1 2 5169 5537
0 2473 7 1 2 2471 2472
0 2474 5 1 1 2473
0 2475 7 2 2 5545 2474
0 2476 5 1 1 7281
0 2477 7 1 2 5512 2476
0 2478 5 2 1 2477
0 2479 7 1 2 5150 7282
0 2480 5 1 1 2479
0 2481 7 2 2 7283 2480
0 2482 5 1 1 7285
0 2483 7 2 2 5504 7286
0 2484 5 2 1 7287
0 2485 7 1 2 7278 7284
0 2486 5 1 1 2485
0 2487 7 1 2 5513 6589
0 2488 5 1 1 2487
0 2489 7 2 2 2486 2488
0 2490 5 1 1 7291
0 2491 7 1 2 7289 7292
0 2492 5 2 1 2491
0 2493 7 1 2 5151 5543
0 2494 5 1 1 2493
0 2495 7 1 2 5170 7280
0 2496 5 1 1 2495
0 2497 7 2 2 2494 2496
0 2498 5 2 1 7295
0 2499 7 2 2 7293 7296
0 2500 5 1 1 7299
0 2501 7 1 2 5505 2500
0 2502 5 2 1 2501
0 2503 7 1 2 5142 7300
0 2504 5 1 1 2503
0 2505 7 2 2 7301 2504
0 2506 5 1 1 7303
0 2507 7 2 2 5496 7304
0 2508 5 2 1 7305
0 2509 7 1 2 2482 7302
0 2510 5 1 1 2509
0 2511 7 1 2 7288 7297
0 2512 5 1 1 2511
0 2513 7 2 2 2510 2512
0 2514 5 1 1 7309
0 2515 7 1 2 7307 2514
0 2516 5 2 1 2515
0 2517 7 1 2 7290 7298
0 2518 5 1 1 2517
0 2519 7 1 2 2490 2518
0 2520 5 1 1 2519
0 2521 7 3 2 7294 2520
0 2522 5 1 1 7313
0 2523 7 1 2 7308 7314
0 2524 5 1 1 2523
0 2525 7 1 2 7310 2524
0 2526 5 1 1 2525
0 2527 7 3 2 7311 2526
0 2528 5 1 1 7316
0 2529 7 2 2 7312 2522
0 2530 5 1 1 7319
0 2531 7 1 2 5497 2530
0 2532 5 2 1 2531
0 2533 7 1 2 5134 7320
0 2534 5 1 1 2533
0 2535 7 2 2 7321 2534
0 2536 5 1 1 7323
0 2537 7 2 2 5489 7324
0 2538 5 2 1 7325
0 2539 7 1 2 2506 7322
0 2540 5 1 1 2539
0 2541 7 1 2 7306 7315
0 2542 5 1 1 2541
0 2543 7 2 2 2540 2542
0 2544 5 1 1 7329
0 2545 7 1 2 7327 2544
0 2546 5 2 1 2545
0 2547 7 2 2 2528 7331
0 2548 5 1 1 7333
0 2549 7 1 2 5490 2548
0 2550 5 2 1 2549
0 2551 7 1 2 5126 7334
0 2552 5 1 1 2551
0 2553 7 2 2 7335 2552
0 2554 5 1 1 7337
0 2555 7 2 2 5482 7338
0 2556 5 2 1 7339
0 2557 7 1 2 2536 7336
0 2558 5 1 1 2557
0 2559 7 1 2 7317 7326
0 2560 5 1 1 2559
0 2561 7 2 2 2558 2560
0 2562 5 1 1 7343
0 2563 7 1 2 7341 2562
0 2564 5 2 1 2563
0 2565 7 1 2 7318 7328
0 2566 5 1 1 2565
0 2567 7 1 2 7330 2566
0 2568 5 1 1 2567
0 2569 7 3 2 7332 2568
0 2570 5 1 1 7347
0 2571 7 1 2 7342 7348
0 2572 5 1 1 2571
0 2573 7 1 2 7344 2572
0 2574 5 1 1 2573
0 2575 7 3 2 7345 2574
0 2576 5 1 1 7350
0 2577 7 2 2 7346 2570
0 2578 5 1 1 7353
0 2579 7 1 2 5483 2578
0 2580 5 2 1 2579
0 2581 7 1 2 5118 7354
0 2582 5 1 1 2581
0 2583 7 2 2 7355 2582
0 2584 5 1 1 7357
0 2585 7 2 2 5475 7358
0 2586 5 2 1 7359
0 2587 7 1 2 2554 7356
0 2588 5 1 1 2587
0 2589 7 1 2 7340 7349
0 2590 5 1 1 2589
0 2591 7 2 2 2588 2590
0 2592 5 1 1 7363
0 2593 7 1 2 7361 2592
0 2594 5 2 1 2593
0 2595 7 2 2 2576 7365
0 2596 5 1 1 7367
0 2597 7 1 2 5476 2596
0 2598 5 2 1 2597
0 2599 7 1 2 5110 7368
0 2600 5 1 1 2599
0 2601 7 2 2 7369 2600
0 2602 5 1 1 7371
0 2603 7 2 2 5468 7372
0 2604 5 2 1 7373
0 2605 7 1 2 2584 7370
0 2606 5 1 1 2605
0 2607 7 1 2 7351 7360
0 2608 5 1 1 2607
0 2609 7 2 2 2606 2608
0 2610 5 1 1 7377
0 2611 7 1 2 7375 2610
0 2612 5 2 1 2611
0 2613 7 1 2 7352 7362
0 2614 5 1 1 2613
0 2615 7 1 2 7364 2614
0 2616 5 1 1 2615
0 2617 7 3 2 7366 2616
0 2618 5 1 1 7381
0 2619 7 1 2 7376 7382
0 2620 5 1 1 2619
0 2621 7 1 2 7378 2620
0 2622 5 1 1 2621
0 2623 7 3 2 7379 2622
0 2624 5 1 1 7384
0 2625 7 2 2 7380 2618
0 2626 5 1 1 7387
0 2627 7 1 2 5469 2626
0 2628 5 2 1 2627
0 2629 7 1 2 5102 7388
0 2630 5 1 1 2629
0 2631 7 2 2 7389 2630
0 2632 5 1 1 7391
0 2633 7 2 2 5461 7392
0 2634 5 2 1 7393
0 2635 7 1 2 2602 7390
0 2636 5 1 1 2635
0 2637 7 1 2 7374 7383
0 2638 5 1 1 2637
0 2639 7 2 2 2636 2638
0 2640 5 1 1 7397
0 2641 7 1 2 7395 2640
0 2642 5 2 1 2641
0 2643 7 2 2 2624 7399
0 2644 5 1 1 7401
0 2645 7 1 2 5462 2644
0 2646 5 2 1 2645
0 2647 7 1 2 5094 7402
0 2648 5 1 1 2647
0 2649 7 2 2 7403 2648
0 2650 5 1 1 7405
0 2651 7 2 2 5454 7406
0 2652 5 2 1 7407
0 2653 7 1 2 2632 7404
0 2654 5 1 1 2653
0 2655 7 1 2 7385 7394
0 2656 5 1 1 2655
0 2657 7 2 2 2654 2656
0 2658 5 1 1 7411
0 2659 7 1 2 7409 2658
0 2660 5 2 1 2659
0 2661 7 1 2 7386 7396
0 2662 5 1 1 2661
0 2663 7 1 2 7398 2662
0 2664 5 1 1 2663
0 2665 7 3 2 7400 2664
0 2666 5 1 1 7415
0 2667 7 1 2 7410 7416
0 2668 5 1 1 2667
0 2669 7 1 2 7412 2668
0 2670 5 1 1 2669
0 2671 7 3 2 7413 2670
0 2672 5 1 1 7418
0 2673 7 2 2 7414 2666
0 2674 5 1 1 7421
0 2675 7 1 2 5455 2674
0 2676 5 2 1 2675
0 2677 7 1 2 5086 7422
0 2678 5 1 1 2677
0 2679 7 2 2 7423 2678
0 2680 5 1 1 7425
0 2681 7 2 2 5447 7426
0 2682 5 2 1 7427
0 2683 7 1 2 2650 7424
0 2684 5 1 1 2683
0 2685 7 1 2 7408 7417
0 2686 5 1 1 2685
0 2687 7 2 2 2684 2686
0 2688 5 1 1 7431
0 2689 7 1 2 7429 2688
0 2690 5 2 1 2689
0 2691 7 2 2 2672 7433
0 2692 5 1 1 7435
0 2693 7 1 2 5448 2692
0 2694 5 2 1 2693
0 2695 7 1 2 5078 7436
0 2696 5 1 1 2695
0 2697 7 2 2 7437 2696
0 2698 5 1 1 7439
0 2699 7 2 2 5440 7440
0 2700 5 2 1 7441
0 2701 7 1 2 2680 7438
0 2702 5 1 1 2701
0 2703 7 1 2 7419 7428
0 2704 5 1 1 2703
0 2705 7 2 2 2702 2704
0 2706 5 1 1 7445
0 2707 7 1 2 7443 2706
0 2708 5 2 1 2707
0 2709 7 1 2 7420 7430
0 2710 5 1 1 2709
0 2711 7 1 2 7432 2710
0 2712 5 1 1 2711
0 2713 7 3 2 7434 2712
0 2714 5 1 1 7449
0 2715 7 1 2 7444 7450
0 2716 5 1 1 2715
0 2717 7 1 2 7446 2716
0 2718 5 1 1 2717
0 2719 7 3 2 7447 2718
0 2720 5 1 1 7452
0 2721 7 2 2 7448 2714
0 2722 5 1 1 7455
0 2723 7 1 2 5441 2722
0 2724 5 2 1 2723
0 2725 7 1 2 5070 7456
0 2726 5 1 1 2725
0 2727 7 2 2 7457 2726
0 2728 5 1 1 7459
0 2729 7 2 2 5433 7460
0 2730 5 2 1 7461
0 2731 7 1 2 2698 7458
0 2732 5 1 1 2731
0 2733 7 1 2 7442 7451
0 2734 5 1 1 2733
0 2735 7 2 2 2732 2734
0 2736 5 1 1 7465
0 2737 7 1 2 7463 2736
0 2738 5 2 1 2737
0 2739 7 2 2 2720 7467
0 2740 5 1 1 7469
0 2741 7 1 2 5434 2740
0 2742 5 2 1 2741
0 2743 7 1 2 5062 7470
0 2744 5 1 1 2743
0 2745 7 2 2 7471 2744
0 2746 5 1 1 7473
0 2747 7 2 2 5426 7474
0 2748 5 2 1 7475
0 2749 7 1 2 2728 7472
0 2750 5 1 1 2749
0 2751 7 1 2 7453 7462
0 2752 5 1 1 2751
0 2753 7 2 2 2750 2752
0 2754 5 1 1 7479
0 2755 7 1 2 7477 2754
0 2756 5 2 1 2755
0 2757 7 1 2 7454 7464
0 2758 5 1 1 2757
0 2759 7 1 2 7466 2758
0 2760 5 1 1 2759
0 2761 7 3 2 7468 2760
0 2762 5 1 1 7483
0 2763 7 1 2 7478 7484
0 2764 5 1 1 2763
0 2765 7 1 2 7480 2764
0 2766 5 1 1 2765
0 2767 7 3 2 7481 2766
0 2768 5 1 1 7486
0 2769 7 2 2 7482 2762
0 2770 5 1 1 7489
0 2771 7 1 2 5427 2770
0 2772 5 2 1 2771
0 2773 7 1 2 5054 7490
0 2774 5 1 1 2773
0 2775 7 2 2 7491 2774
0 2776 5 1 1 7493
0 2777 7 2 2 5419 7494
0 2778 5 2 1 7495
0 2779 7 1 2 2746 7492
0 2780 5 1 1 2779
0 2781 7 1 2 7476 7485
0 2782 5 1 1 2781
0 2783 7 2 2 2780 2782
0 2784 5 1 1 7499
0 2785 7 1 2 7497 2784
0 2786 5 2 1 2785
0 2787 7 2 2 2768 7501
0 2788 5 1 1 7503
0 2789 7 1 2 5420 2788
0 2790 5 2 1 2789
0 2791 7 1 2 5046 7504
0 2792 5 1 1 2791
0 2793 7 2 2 7505 2792
0 2794 5 1 1 7507
0 2795 7 2 2 5411 7508
0 2796 5 2 1 7509
0 2797 7 1 2 2776 7506
0 2798 5 1 1 2797
0 2799 7 1 2 7487 7496
0 2800 5 1 1 2799
0 2801 7 2 2 2798 2800
0 2802 5 1 1 7513
0 2803 7 1 2 7511 2802
0 2804 5 2 1 2803
0 2805 7 1 2 7488 7498
0 2806 5 1 1 2805
0 2807 7 1 2 7500 2806
0 2808 5 1 1 2807
0 2809 7 3 2 7502 2808
0 2810 5 1 1 7517
0 2811 7 1 2 7512 7518
0 2812 5 1 1 2811
0 2813 7 1 2 7514 2812
0 2814 5 1 1 2813
0 2815 7 3 2 7515 2814
0 2816 5 1 1 7520
0 2817 7 2 2 7516 2810
0 2818 5 1 1 7523
0 2819 7 1 2 5412 2818
0 2820 5 2 1 2819
0 2821 7 1 2 5038 7524
0 2822 5 1 1 2821
0 2823 7 2 2 7525 2822
0 2824 5 1 1 7527
0 2825 7 2 2 5403 7528
0 2826 5 2 1 7529
0 2827 7 1 2 2794 7526
0 2828 5 1 1 2827
0 2829 7 1 2 7510 7519
0 2830 5 1 1 2829
0 2831 7 2 2 2828 2830
0 2832 5 1 1 7533
0 2833 7 1 2 7531 2832
0 2834 5 2 1 2833
0 2835 7 2 2 2816 7535
0 2836 5 1 1 7537
0 2837 7 1 2 5404 2836
0 2838 5 2 1 2837
0 2839 7 1 2 5030 7538
0 2840 5 1 1 2839
0 2841 7 2 2 7539 2840
0 2842 5 1 1 7541
0 2843 7 2 2 5395 7542
0 2844 5 2 1 7543
0 2845 7 1 2 2824 7540
0 2846 5 1 1 2845
0 2847 7 1 2 7521 7530
0 2848 5 1 1 2847
0 2849 7 2 2 2846 2848
0 2850 5 1 1 7547
0 2851 7 1 2 7545 2850
0 2852 5 2 1 2851
0 2853 7 1 2 7522 7532
0 2854 5 1 1 2853
0 2855 7 1 2 7534 2854
0 2856 5 1 1 2855
0 2857 7 3 2 7536 2856
0 2858 5 1 1 7551
0 2859 7 1 2 7546 7552
0 2860 5 1 1 2859
0 2861 7 1 2 7548 2860
0 2862 5 1 1 2861
0 2863 7 3 2 7549 2862
0 2864 5 1 1 7554
0 2865 7 2 2 7550 2858
0 2866 5 1 1 7557
0 2867 7 1 2 5396 2866
0 2868 5 2 1 2867
0 2869 7 1 2 5022 7558
0 2870 5 1 1 2869
0 2871 7 2 2 7559 2870
0 2872 5 1 1 7561
0 2873 7 2 2 5387 7562
0 2874 5 2 1 7563
0 2875 7 1 2 2842 7560
0 2876 5 1 1 2875
0 2877 7 1 2 7544 7553
0 2878 5 1 1 2877
0 2879 7 2 2 2876 2878
0 2880 5 1 1 7567
0 2881 7 1 2 7565 2880
0 2882 5 2 1 2881
0 2883 7 2 2 2864 7569
0 2884 5 1 1 7571
0 2885 7 1 2 5388 2884
0 2886 5 2 1 2885
0 2887 7 1 2 5014 7572
0 2888 5 1 1 2887
0 2889 7 2 2 7573 2888
0 2890 5 1 1 7575
0 2891 7 2 2 5379 7576
0 2892 5 2 1 7577
0 2893 7 1 2 2872 7574
0 2894 5 1 1 2893
0 2895 7 1 2 7555 7564
0 2896 5 1 1 2895
0 2897 7 2 2 2894 2896
0 2898 5 1 1 7581
0 2899 7 1 2 7579 2898
0 2900 5 2 1 2899
0 2901 7 1 2 7556 7566
0 2902 5 1 1 2901
0 2903 7 1 2 7568 2902
0 2904 5 1 1 2903
0 2905 7 3 2 7570 2904
0 2906 5 1 1 7585
0 2907 7 1 2 7580 7586
0 2908 5 1 1 2907
0 2909 7 1 2 7582 2908
0 2910 5 1 1 2909
0 2911 7 3 2 7583 2910
0 2912 5 1 1 7588
0 2913 7 2 2 7584 2906
0 2914 5 1 1 7591
0 2915 7 1 2 5380 2914
0 2916 5 2 1 2915
0 2917 7 1 2 5006 7592
0 2918 5 1 1 2917
0 2919 7 2 2 7593 2918
0 2920 5 1 1 7595
0 2921 7 2 2 5371 7596
0 2922 5 2 1 7597
0 2923 7 1 2 2890 7594
0 2924 5 1 1 2923
0 2925 7 1 2 7578 7587
0 2926 5 1 1 2925
0 2927 7 2 2 2924 2926
0 2928 5 1 1 7601
0 2929 7 1 2 7599 2928
0 2930 5 2 1 2929
0 2931 7 2 2 2912 7603
0 2932 5 1 1 7605
0 2933 7 1 2 5372 2932
0 2934 5 2 1 2933
0 2935 7 1 2 4998 7606
0 2936 5 1 1 2935
0 2937 7 2 2 7607 2936
0 2938 5 1 1 7609
0 2939 7 2 2 5363 7610
0 2940 5 2 1 7611
0 2941 7 1 2 2920 7608
0 2942 5 1 1 2941
0 2943 7 1 2 7589 7598
0 2944 5 1 1 2943
0 2945 7 2 2 2942 2944
0 2946 5 1 1 7615
0 2947 7 1 2 7613 2946
0 2948 5 2 1 2947
0 2949 7 1 2 7590 7600
0 2950 5 1 1 2949
0 2951 7 1 2 7602 2950
0 2952 5 1 1 2951
0 2953 7 3 2 7604 2952
0 2954 5 1 1 7619
0 2955 7 1 2 7614 7620
0 2956 5 1 1 2955
0 2957 7 1 2 7616 2956
0 2958 5 1 1 2957
0 2959 7 3 2 7617 2958
0 2960 5 1 1 7622
0 2961 7 2 2 7618 2954
0 2962 5 1 1 7625
0 2963 7 1 2 5364 2962
0 2964 5 2 1 2963
0 2965 7 1 2 4990 7626
0 2966 5 1 1 2965
0 2967 7 2 2 7627 2966
0 2968 5 1 1 7629
0 2969 7 2 2 5355 7630
0 2970 5 2 1 7631
0 2971 7 1 2 2938 7628
0 2972 5 1 1 2971
0 2973 7 1 2 7612 7621
0 2974 5 1 1 2973
0 2975 7 2 2 2972 2974
0 2976 5 1 1 7635
0 2977 7 1 2 7633 2976
0 2978 5 2 1 2977
0 2979 7 2 2 2960 7637
0 2980 5 1 1 7639
0 2981 7 1 2 5356 2980
0 2982 5 2 1 2981
0 2983 7 1 2 4982 7640
0 2984 5 1 1 2983
0 2985 7 2 2 7641 2984
0 2986 5 1 1 7643
0 2987 7 2 2 5347 7644
0 2988 5 2 1 7645
0 2989 7 1 2 2968 7642
0 2990 5 1 1 2989
0 2991 7 1 2 7623 7632
0 2992 5 1 1 2991
0 2993 7 2 2 2990 2992
0 2994 5 1 1 7649
0 2995 7 1 2 7647 2994
0 2996 5 2 1 2995
0 2997 7 1 2 7624 7634
0 2998 5 1 1 2997
0 2999 7 1 2 7636 2998
0 3000 5 1 1 2999
0 3001 7 3 2 7638 3000
0 3002 5 1 1 7653
0 3003 7 1 2 7648 7654
0 3004 5 1 1 3003
0 3005 7 1 2 7650 3004
0 3006 5 1 1 3005
0 3007 7 3 2 7651 3006
0 3008 5 1 1 7656
0 3009 7 2 2 7652 3002
0 3010 5 1 1 7659
0 3011 7 1 2 5348 3010
0 3012 5 2 1 3011
0 3013 7 1 2 4974 7660
0 3014 5 1 1 3013
0 3015 7 2 2 7661 3014
0 3016 5 1 1 7663
0 3017 7 2 2 5339 7664
0 3018 5 2 1 7665
0 3019 7 1 2 2986 7662
0 3020 5 1 1 3019
0 3021 7 1 2 7646 7655
0 3022 5 1 1 3021
0 3023 7 2 2 3020 3022
0 3024 5 1 1 7669
0 3025 7 1 2 7667 3024
0 3026 5 2 1 3025
0 3027 7 2 2 3008 7671
0 3028 5 1 1 7673
0 3029 7 1 2 5340 3028
0 3030 5 2 1 3029
0 3031 7 1 2 4966 7674
0 3032 5 1 1 3031
0 3033 7 2 2 7675 3032
0 3034 5 1 1 7677
0 3035 7 2 2 5331 7678
0 3036 5 2 1 7679
0 3037 7 1 2 3016 7676
0 3038 5 1 1 3037
0 3039 7 1 2 7657 7666
0 3040 5 1 1 3039
0 3041 7 2 2 3038 3040
0 3042 5 1 1 7683
0 3043 7 1 2 7681 3042
0 3044 5 2 1 3043
0 3045 7 1 2 7658 7668
0 3046 5 1 1 3045
0 3047 7 1 2 7670 3046
0 3048 5 1 1 3047
0 3049 7 3 2 7672 3048
0 3050 5 1 1 7687
0 3051 7 1 2 7682 7688
0 3052 5 1 1 3051
0 3053 7 1 2 7684 3052
0 3054 5 1 1 3053
0 3055 7 3 2 7685 3054
0 3056 5 1 1 7690
0 3057 7 2 2 7686 3050
0 3058 5 1 1 7693
0 3059 7 1 2 5332 3058
0 3060 5 2 1 3059
0 3061 7 1 2 4958 7694
0 3062 5 1 1 3061
0 3063 7 2 2 7695 3062
0 3064 5 1 1 7697
0 3065 7 2 2 5323 7698
0 3066 5 2 1 7699
0 3067 7 1 2 3034 7696
0 3068 5 1 1 3067
0 3069 7 1 2 7680 7689
0 3070 5 1 1 3069
0 3071 7 2 2 3068 3070
0 3072 5 1 1 7703
0 3073 7 1 2 7701 3072
0 3074 5 2 1 3073
0 3075 7 2 2 3056 7705
0 3076 5 1 1 7707
0 3077 7 1 2 5324 3076
0 3078 5 2 1 3077
0 3079 7 1 2 4950 7708
0 3080 5 1 1 3079
0 3081 7 2 2 7709 3080
0 3082 5 1 1 7711
0 3083 7 2 2 5315 7712
0 3084 5 2 1 7713
0 3085 7 1 2 3064 7710
0 3086 5 1 1 3085
0 3087 7 1 2 7691 7700
0 3088 5 1 1 3087
0 3089 7 2 2 3086 3088
0 3090 5 1 1 7717
0 3091 7 1 2 7715 3090
0 3092 5 2 1 3091
0 3093 7 1 2 7692 7702
0 3094 5 1 1 3093
0 3095 7 1 2 7704 3094
0 3096 5 1 1 3095
0 3097 7 3 2 7706 3096
0 3098 5 1 1 7721
0 3099 7 1 2 7716 7722
0 3100 5 1 1 3099
0 3101 7 1 2 7718 3100
0 3102 5 1 1 3101
0 3103 7 3 2 7719 3102
0 3104 5 1 1 7724
0 3105 7 2 2 7720 3098
0 3106 5 1 1 7727
0 3107 7 1 2 5316 3106
0 3108 5 2 1 3107
0 3109 7 1 2 4942 7728
0 3110 5 1 1 3109
0 3111 7 2 2 7729 3110
0 3112 5 1 1 7731
0 3113 7 2 2 5308 7732
0 3114 5 2 1 7733
0 3115 7 1 2 3082 7730
0 3116 5 1 1 3115
0 3117 7 1 2 7714 7723
0 3118 5 1 1 3117
0 3119 7 2 2 3116 3118
0 3120 5 1 1 7737
0 3121 7 1 2 7735 3120
0 3122 5 2 1 3121
0 3123 7 2 2 3104 7739
0 3124 5 1 1 7741
0 3125 7 1 2 5309 3124
0 3126 5 2 1 3125
0 3127 7 1 2 4934 7742
0 3128 5 1 1 3127
0 3129 7 2 2 7743 3128
0 3130 5 1 1 7745
0 3131 7 2 2 5301 7746
0 3132 5 2 1 7747
0 3133 7 1 2 3112 7744
0 3134 5 1 1 3133
0 3135 7 1 2 7725 7734
0 3136 5 1 1 3135
0 3137 7 2 2 3134 3136
0 3138 5 1 1 7751
0 3139 7 1 2 7749 3138
0 3140 5 2 1 3139
0 3141 7 1 2 7726 7736
0 3142 5 1 1 3141
0 3143 7 1 2 7738 3142
0 3144 5 1 1 3143
0 3145 7 3 2 7740 3144
0 3146 5 1 1 7755
0 3147 7 1 2 7750 7756
0 3148 5 1 1 3147
0 3149 7 1 2 7752 3148
0 3150 5 1 1 3149
0 3151 7 3 2 7753 3150
0 3152 5 1 1 7758
0 3153 7 2 2 7754 3146
0 3154 5 1 1 7761
0 3155 7 1 2 5302 3154
0 3156 5 2 1 3155
0 3157 7 1 2 4926 7762
0 3158 5 1 1 3157
0 3159 7 2 2 7763 3158
0 3160 5 1 1 7765
0 3161 7 2 2 5294 7766
0 3162 5 2 1 7767
0 3163 7 1 2 3130 7764
0 3164 5 1 1 3163
0 3165 7 1 2 7748 7757
0 3166 5 1 1 3165
0 3167 7 2 2 3164 3166
0 3168 5 1 1 7771
0 3169 7 1 2 7769 3168
0 3170 5 2 1 3169
0 3171 7 2 2 3152 7773
0 3172 5 1 1 7775
0 3173 7 1 2 5295 3172
0 3174 5 2 1 3173
0 3175 7 1 2 4918 7776
0 3176 5 1 1 3175
0 3177 7 2 2 7777 3176
0 3178 5 1 1 7779
0 3179 7 2 2 5287 7780
0 3180 5 2 1 7781
0 3181 7 1 2 3160 7778
0 3182 5 1 1 3181
0 3183 7 1 2 7759 7768
0 3184 5 1 1 3183
0 3185 7 2 2 3182 3184
0 3186 5 1 1 7785
0 3187 7 1 2 7783 3186
0 3188 5 2 1 3187
0 3189 7 1 2 7760 7770
0 3190 5 1 1 3189
0 3191 7 1 2 7772 3190
0 3192 5 1 1 3191
0 3193 7 3 2 7774 3192
0 3194 5 1 1 7789
0 3195 7 1 2 7784 7790
0 3196 5 1 1 3195
0 3197 7 1 2 7786 3196
0 3198 5 1 1 3197
0 3199 7 3 2 7787 3198
0 3200 5 1 1 7792
0 3201 7 2 2 7788 3194
0 3202 5 1 1 7795
0 3203 7 1 2 5288 3202
0 3204 5 2 1 3203
0 3205 7 1 2 4910 7796
0 3206 5 1 1 3205
0 3207 7 2 2 7797 3206
0 3208 5 1 1 7799
0 3209 7 2 2 5280 7800
0 3210 5 2 1 7801
0 3211 7 1 2 3178 7798
0 3212 5 1 1 3211
0 3213 7 1 2 7782 7791
0 3214 5 1 1 3213
0 3215 7 2 2 3212 3214
0 3216 5 1 1 7805
0 3217 7 1 2 7803 3216
0 3218 5 2 1 3217
0 3219 7 2 2 3200 7807
0 3220 5 1 1 7809
0 3221 7 1 2 5281 3220
0 3222 5 2 1 3221
0 3223 7 1 2 4902 7810
0 3224 5 1 1 3223
0 3225 7 2 2 7811 3224
0 3226 5 1 1 7813
0 3227 7 2 2 5273 7814
0 3228 5 2 1 7815
0 3229 7 1 2 3208 7812
0 3230 5 1 1 3229
0 3231 7 1 2 7793 7802
0 3232 5 1 1 3231
0 3233 7 2 2 3230 3232
0 3234 5 1 1 7819
0 3235 7 1 2 7817 3234
0 3236 5 2 1 3235
0 3237 7 1 2 7794 7804
0 3238 5 1 1 3237
0 3239 7 1 2 7806 3238
0 3240 5 1 1 3239
0 3241 7 3 2 7808 3240
0 3242 5 1 1 7823
0 3243 7 1 2 7818 7824
0 3244 5 1 1 3243
0 3245 7 1 2 7820 3244
0 3246 5 1 1 3245
0 3247 7 3 2 7821 3246
0 3248 5 1 1 7826
0 3249 7 2 2 7822 3242
0 3250 5 1 1 7829
0 3251 7 1 2 5274 3250
0 3252 5 2 1 3251
0 3253 7 1 2 4894 7830
0 3254 5 1 1 3253
0 3255 7 2 2 7831 3254
0 3256 5 1 1 7833
0 3257 7 2 2 5266 7834
0 3258 5 2 1 7835
0 3259 7 1 2 3226 7832
0 3260 5 1 1 3259
0 3261 7 1 2 7816 7825
0 3262 5 1 1 3261
0 3263 7 2 2 3260 3262
0 3264 5 1 1 7839
0 3265 7 1 2 7837 3264
0 3266 5 2 1 3265
0 3267 7 2 2 3248 7841
0 3268 5 1 1 7843
0 3269 7 1 2 5267 3268
0 3270 5 2 1 3269
0 3271 7 1 2 4886 7844
0 3272 5 1 1 3271
0 3273 7 2 2 7845 3272
0 3274 5 1 1 7847
0 3275 7 2 2 5259 7848
0 3276 5 2 1 7849
0 3277 7 1 2 3256 7846
0 3278 5 1 1 3277
0 3279 7 1 2 7827 7836
0 3280 5 1 1 3279
0 3281 7 2 2 3278 3280
0 3282 5 1 1 7853
0 3283 7 1 2 7851 3282
0 3284 5 2 1 3283
0 3285 7 1 2 7828 7838
0 3286 5 1 1 3285
0 3287 7 1 2 7840 3286
0 3288 5 1 1 3287
0 3289 7 3 2 7842 3288
0 3290 5 1 1 7857
0 3291 7 1 2 7852 7858
0 3292 5 1 1 3291
0 3293 7 1 2 7854 3292
0 3294 5 1 1 3293
0 3295 7 3 2 7855 3294
0 3296 5 1 1 7860
0 3297 7 2 2 7856 3290
0 3298 5 1 1 7863
0 3299 7 1 2 5260 3298
0 3300 5 2 1 3299
0 3301 7 1 2 4878 7864
0 3302 5 1 1 3301
0 3303 7 2 2 7865 3302
0 3304 5 1 1 7867
0 3305 7 2 2 5252 7868
0 3306 5 2 1 7869
0 3307 7 1 2 3274 7866
0 3308 5 1 1 3307
0 3309 7 1 2 7850 7859
0 3310 5 1 1 3309
0 3311 7 2 2 3308 3310
0 3312 5 1 1 7873
0 3313 7 1 2 7871 3312
0 3314 5 2 1 3313
0 3315 7 2 2 3296 7875
0 3316 5 1 1 7877
0 3317 7 1 2 5253 3316
0 3318 5 2 1 3317
0 3319 7 1 2 4870 7878
0 3320 5 1 1 3319
0 3321 7 2 2 7879 3320
0 3322 5 1 1 7881
0 3323 7 2 2 5245 7882
0 3324 5 2 1 7883
0 3325 7 1 2 3304 7880
0 3326 5 1 1 3325
0 3327 7 1 2 7861 7870
0 3328 5 1 1 3327
0 3329 7 2 2 3326 3328
0 3330 5 1 1 7887
0 3331 7 1 2 7885 3330
0 3332 5 2 1 3331
0 3333 7 1 2 7862 7872
0 3334 5 1 1 3333
0 3335 7 1 2 7874 3334
0 3336 5 1 1 3335
0 3337 7 3 2 7876 3336
0 3338 5 1 1 7891
0 3339 7 1 2 7886 7892
0 3340 5 1 1 3339
0 3341 7 1 2 7888 3340
0 3342 5 1 1 3341
0 3343 7 3 2 7889 3342
0 3344 5 1 1 7894
0 3345 7 2 2 7890 3338
0 3346 5 1 1 7897
0 3347 7 1 2 5246 3346
0 3348 5 2 1 3347
0 3349 7 1 2 4862 7898
0 3350 5 1 1 3349
0 3351 7 2 2 7899 3350
0 3352 5 1 1 7901
0 3353 7 2 2 5238 7902
0 3354 5 2 1 7903
0 3355 7 1 2 3322 7900
0 3356 5 1 1 3355
0 3357 7 1 2 7884 7893
0 3358 5 1 1 3357
0 3359 7 2 2 3356 3358
0 3360 5 1 1 7907
0 3361 7 1 2 7905 3360
0 3362 5 2 1 3361
0 3363 7 2 2 3344 7909
0 3364 5 1 1 7911
0 3365 7 1 2 5239 3364
0 3366 5 2 1 3365
0 3367 7 1 2 4854 7912
0 3368 5 1 1 3367
0 3369 7 2 2 7913 3368
0 3370 5 1 1 7915
0 3371 7 2 2 5231 7916
0 3372 5 2 1 7917
0 3373 7 1 2 3352 7914
0 3374 5 1 1 3373
0 3375 7 1 2 7895 7904
0 3376 5 1 1 3375
0 3377 7 2 2 3374 3376
0 3378 5 1 1 7921
0 3379 7 1 2 7919 3378
0 3380 5 2 1 3379
0 3381 7 1 2 7896 7906
0 3382 5 1 1 3381
0 3383 7 1 2 7908 3382
0 3384 5 1 1 3383
0 3385 7 3 2 7910 3384
0 3386 5 1 1 7925
0 3387 7 1 2 7920 7926
0 3388 5 1 1 3387
0 3389 7 1 2 7922 3388
0 3390 5 1 1 3389
0 3391 7 3 2 7923 3390
0 3392 5 1 1 7928
0 3393 7 2 2 7924 3386
0 3394 5 1 1 7931
0 3395 7 1 2 5232 3394
0 3396 5 2 1 3395
0 3397 7 1 2 4846 7932
0 3398 5 1 1 3397
0 3399 7 2 2 7933 3398
0 3400 5 1 1 7935
0 3401 7 2 2 5224 7936
0 3402 5 2 1 7937
0 3403 7 1 2 3370 7934
0 3404 5 1 1 3403
0 3405 7 1 2 7918 7927
0 3406 5 1 1 3405
0 3407 7 2 2 3404 3406
0 3408 5 1 1 7941
0 3409 7 1 2 7939 3408
0 3410 5 2 1 3409
0 3411 7 2 2 3392 7943
0 3412 5 1 1 7945
0 3413 7 1 2 5225 3412
0 3414 5 2 1 3413
0 3415 7 1 2 4838 7946
0 3416 5 1 1 3415
0 3417 7 2 2 7947 3416
0 3418 5 1 1 7949
0 3419 7 2 2 5217 7950
0 3420 5 2 1 7951
0 3421 7 1 2 3400 7948
0 3422 5 1 1 3421
0 3423 7 1 2 7929 7938
0 3424 5 1 1 3423
0 3425 7 2 2 3422 3424
0 3426 5 1 1 7955
0 3427 7 1 2 7953 3426
0 3428 5 2 1 3427
0 3429 7 1 2 7930 7940
0 3430 5 1 1 3429
0 3431 7 1 2 7942 3430
0 3432 5 1 1 3431
0 3433 7 3 2 7944 3432
0 3434 5 1 1 7959
0 3435 7 1 2 7954 7960
0 3436 5 1 1 3435
0 3437 7 1 2 7956 3436
0 3438 5 1 1 3437
0 3439 7 3 2 7957 3438
0 3440 5 1 1 7962
0 3441 7 2 2 7958 3434
0 3442 5 1 1 7965
0 3443 7 1 2 5218 3442
0 3444 5 2 1 3443
0 3445 7 1 2 4830 7966
0 3446 5 1 1 3445
0 3447 7 2 2 7967 3446
0 3448 5 1 1 7969
0 3449 7 2 2 5210 7970
0 3450 5 2 1 7971
0 3451 7 1 2 3418 7968
0 3452 5 1 1 3451
0 3453 7 1 2 7952 7961
0 3454 5 1 1 3453
0 3455 7 2 2 3452 3454
0 3456 5 1 1 7975
0 3457 7 1 2 7973 3456
0 3458 5 2 1 3457
0 3459 7 2 2 3440 7977
0 3460 5 1 1 7979
0 3461 7 1 2 5211 3460
0 3462 5 2 1 3461
0 3463 7 1 2 4822 7980
0 3464 5 1 1 3463
0 3465 7 2 2 7981 3464
0 3466 5 1 1 7983
0 3467 7 2 2 5203 7984
0 3468 5 2 1 7985
0 3469 7 1 2 3448 7982
0 3470 5 1 1 3469
0 3471 7 1 2 7963 7972
0 3472 5 1 1 3471
0 3473 7 2 2 3470 3472
0 3474 5 1 1 7989
0 3475 7 1 2 7987 3474
0 3476 5 2 1 3475
0 3477 7 1 2 7964 7974
0 3478 5 1 1 3477
0 3479 7 1 2 7976 3478
0 3480 5 1 1 3479
0 3481 7 3 2 7978 3480
0 3482 5 1 1 7993
0 3483 7 2 2 7991 3482
0 3484 5 1 1 7996
0 3485 7 1 2 5204 3484
0 3486 5 2 1 3485
0 3487 7 1 2 4814 7997
0 3488 5 1 1 3487
0 3489 7 3 2 7998 3488
0 3490 5 1 1 8000
0 3491 7 2 2 5196 8001
0 3492 5 2 1 8003
0 3493 7 1 2 3466 7999
0 3494 5 1 1 3493
0 3495 7 1 2 7986 7994
0 3496 5 1 1 3495
0 3497 7 2 2 3494 3496
0 3498 5 1 1 8007
0 3499 7 1 2 8005 3498
0 3500 5 2 1 3499
0 3501 7 1 2 7988 7995
0 3502 5 1 1 3501
0 3503 7 1 2 7990 3502
0 3504 5 1 1 3503
0 3505 7 3 2 7992 3504
0 3506 5 1 1 8011
0 3507 7 1 2 8006 8012
0 3508 5 1 1 3507
0 3509 7 1 2 8008 3508
0 3510 5 1 1 3509
0 3511 7 2 2 8009 3510
0 3512 5 1 1 8014
0 3513 7 1 2 5190 8015
0 3514 5 2 1 3513
0 3515 7 1 2 8004 8013
0 3516 5 2 1 3515
0 3517 7 2 2 8002 8018
0 3518 5 1 1 8020
0 3519 7 1 2 5191 3518
0 3520 5 1 1 3519
0 3521 7 1 2 4796 8021
0 3522 5 1 1 3521
0 3523 7 1 2 3520 3522
0 3524 7 1 2 8016 3523
0 3525 5 1 1 3524
0 3526 7 1 2 4790 3525
0 3527 5 1 1 3526
0 3528 7 1 2 5183 8017
0 3529 5 1 1 3528
0 3530 7 2 2 8010 3506
0 3531 5 1 1 8022
0 3532 7 1 2 5197 3531
0 3533 5 1 1 3532
0 3534 7 1 2 4805 8023
0 3535 5 1 1 3534
0 3536 7 2 2 3533 3535
0 3537 5 1 1 8024
0 3538 7 1 2 3529 8025
0 3539 7 1 2 3527 3538
0 3540 5 1 1 3539
0 3541 7 2 2 5163 111
0 3542 5 1 1 8026
0 3543 7 1 2 5171 5528
0 3544 5 2 1 3543
0 3545 7 1 2 5518 8028
0 3546 5 1 1 3545
0 3547 7 2 2 3542 3546
0 3548 5 1 1 8030
0 3549 7 1 2 5152 8031
0 3550 5 2 1 3549
0 3551 7 1 2 8027 8029
0 3552 5 1 1 3551
0 3553 7 3 2 5546 3552
0 3554 5 1 1 8034
0 3555 7 1 2 8032 8035
0 3556 5 1 1 3555
0 3557 7 1 2 5153 3554
0 3558 5 1 1 3557
0 3559 7 2 2 3556 3558
0 3560 5 1 1 8037
0 3561 7 2 2 5143 8038
0 3562 5 1 1 8039
0 3563 7 1 2 5154 8036
0 3564 5 1 1 3563
0 3565 7 1 2 3548 3564
0 3566 5 1 1 3565
0 3567 7 2 2 8033 3566
0 3568 5 2 1 8041
0 3569 7 1 2 5144 8043
0 3570 5 1 1 3569
0 3571 7 1 2 3560 3570
0 3572 5 1 1 3571
0 3573 7 2 2 3562 3572
0 3574 5 1 1 8045
0 3575 7 1 2 5135 8046
0 3576 5 2 1 3575
0 3577 7 1 2 8040 8044
0 3578 5 1 1 3577
0 3579 7 1 2 5506 8042
0 3580 5 1 1 3579
0 3581 7 2 2 3578 3580
0 3582 5 1 1 8049
0 3583 7 1 2 5136 3582
0 3584 5 2 1 3583
0 3585 7 1 2 3574 8051
0 3586 5 1 1 3585
0 3587 7 2 2 8047 3586
0 3588 5 1 1 8053
0 3589 7 1 2 5491 3588
0 3590 5 1 1 3589
0 3591 7 1 2 5498 8050
0 3592 5 1 1 3591
0 3593 7 1 2 3592 8052
0 3594 7 2 2 8048 3593
0 3595 5 1 1 8055
0 3596 7 1 2 5127 8056
0 3597 5 2 1 3596
0 3598 7 1 2 5128 8054
0 3599 5 2 1 3598
0 3600 7 1 2 8057 8059
0 3601 7 2 2 3590 3600
0 3602 5 1 1 8061
0 3603 7 1 2 5119 8062
0 3604 5 2 1 3603
0 3605 7 1 2 3595 8060
0 3606 5 1 1 3605
0 3607 7 2 2 8058 3606
0 3608 5 1 1 8065
0 3609 7 1 2 5120 8066
0 3610 5 2 1 3609
0 3611 7 1 2 3602 8067
0 3612 5 1 1 3611
0 3613 7 2 2 8063 3612
0 3614 5 1 1 8069
0 3615 7 1 2 5477 3614
0 3616 5 1 1 3615
0 3617 7 1 2 5484 3608
0 3618 5 1 1 3617
0 3619 7 1 2 8064 8068
0 3620 7 2 2 3618 3619
0 3621 5 1 1 8071
0 3622 7 1 2 5111 8072
0 3623 5 2 1 3622
0 3624 7 1 2 5112 8070
0 3625 5 2 1 3624
0 3626 7 1 2 8073 8075
0 3627 7 2 2 3616 3626
0 3628 5 1 1 8077
0 3629 7 1 2 5103 8078
0 3630 5 2 1 3629
0 3631 7 1 2 3621 8076
0 3632 5 1 1 3631
0 3633 7 2 2 8074 3632
0 3634 5 1 1 8081
0 3635 7 1 2 5104 8082
0 3636 5 2 1 3635
0 3637 7 1 2 3628 8083
0 3638 5 1 1 3637
0 3639 7 2 2 8079 3638
0 3640 5 1 1 8085
0 3641 7 1 2 5463 3640
0 3642 5 1 1 3641
0 3643 7 1 2 5470 3634
0 3644 5 1 1 3643
0 3645 7 1 2 8080 8084
0 3646 7 2 2 3644 3645
0 3647 5 1 1 8087
0 3648 7 1 2 5095 8088
0 3649 5 2 1 3648
0 3650 7 1 2 5096 8086
0 3651 5 2 1 3650
0 3652 7 1 2 8089 8091
0 3653 7 2 2 3642 3652
0 3654 5 1 1 8093
0 3655 7 1 2 5087 8094
0 3656 5 2 1 3655
0 3657 7 1 2 3647 8092
0 3658 5 1 1 3657
0 3659 7 2 2 8090 3658
0 3660 5 1 1 8097
0 3661 7 1 2 5088 8098
0 3662 5 2 1 3661
0 3663 7 1 2 3654 8099
0 3664 5 1 1 3663
0 3665 7 2 2 8095 3664
0 3666 5 1 1 8101
0 3667 7 1 2 5449 3666
0 3668 5 1 1 3667
0 3669 7 1 2 5456 3660
0 3670 5 1 1 3669
0 3671 7 1 2 8096 8100
0 3672 7 2 2 3670 3671
0 3673 5 1 1 8103
0 3674 7 1 2 5079 8104
0 3675 5 2 1 3674
0 3676 7 1 2 5080 8102
0 3677 5 2 1 3676
0 3678 7 1 2 8105 8107
0 3679 7 2 2 3668 3678
0 3680 5 1 1 8109
0 3681 7 1 2 5071 8110
0 3682 5 2 1 3681
0 3683 7 1 2 3673 8108
0 3684 5 1 1 3683
0 3685 7 2 2 8106 3684
0 3686 5 1 1 8113
0 3687 7 1 2 5072 8114
0 3688 5 2 1 3687
0 3689 7 1 2 3680 8115
0 3690 5 1 1 3689
0 3691 7 2 2 8111 3690
0 3692 5 1 1 8117
0 3693 7 1 2 5435 3692
0 3694 5 1 1 3693
0 3695 7 1 2 5442 3686
0 3696 5 1 1 3695
0 3697 7 1 2 8112 8116
0 3698 7 2 2 3696 3697
0 3699 5 1 1 8119
0 3700 7 1 2 5063 8120
0 3701 5 2 1 3700
0 3702 7 1 2 5064 8118
0 3703 5 2 1 3702
0 3704 7 1 2 8121 8123
0 3705 7 2 2 3694 3704
0 3706 5 1 1 8125
0 3707 7 1 2 5055 8126
0 3708 5 2 1 3707
0 3709 7 1 2 3699 8124
0 3710 5 1 1 3709
0 3711 7 2 2 8122 3710
0 3712 5 1 1 8129
0 3713 7 1 2 5056 8130
0 3714 5 2 1 3713
0 3715 7 1 2 3706 8131
0 3716 5 1 1 3715
0 3717 7 2 2 8127 3716
0 3718 5 1 1 8133
0 3719 7 1 2 5421 3718
0 3720 5 1 1 3719
0 3721 7 1 2 5428 3712
0 3722 5 1 1 3721
0 3723 7 1 2 8128 8132
0 3724 7 2 2 3722 3723
0 3725 5 1 1 8135
0 3726 7 1 2 5047 8136
0 3727 5 2 1 3726
0 3728 7 1 2 5048 8134
0 3729 5 2 1 3728
0 3730 7 1 2 8137 8139
0 3731 7 2 2 3720 3730
0 3732 5 1 1 8141
0 3733 7 1 2 5039 8142
0 3734 5 2 1 3733
0 3735 7 1 2 3725 8140
0 3736 5 1 1 3735
0 3737 7 2 2 8138 3736
0 3738 5 1 1 8145
0 3739 7 1 2 5040 8146
0 3740 5 2 1 3739
0 3741 7 1 2 3732 8147
0 3742 5 1 1 3741
0 3743 7 2 2 8143 3742
0 3744 5 1 1 8149
0 3745 7 1 2 5405 3744
0 3746 5 1 1 3745
0 3747 7 1 2 5413 3738
0 3748 5 1 1 3747
0 3749 7 1 2 8144 8148
0 3750 7 2 2 3748 3749
0 3751 5 1 1 8151
0 3752 7 1 2 5031 8152
0 3753 5 2 1 3752
0 3754 7 1 2 5032 8150
0 3755 5 2 1 3754
0 3756 7 1 2 8153 8155
0 3757 7 2 2 3746 3756
0 3758 5 1 1 8157
0 3759 7 1 2 5023 8158
0 3760 5 2 1 3759
0 3761 7 1 2 3751 8156
0 3762 5 1 1 3761
0 3763 7 2 2 8154 3762
0 3764 5 1 1 8161
0 3765 7 1 2 5024 8162
0 3766 5 2 1 3765
0 3767 7 1 2 3758 8163
0 3768 5 1 1 3767
0 3769 7 2 2 8159 3768
0 3770 5 1 1 8165
0 3771 7 1 2 5389 3770
0 3772 5 1 1 3771
0 3773 7 1 2 5397 3764
0 3774 5 1 1 3773
0 3775 7 1 2 8160 8164
0 3776 7 2 2 3774 3775
0 3777 5 1 1 8167
0 3778 7 1 2 5015 8168
0 3779 5 2 1 3778
0 3780 7 1 2 5016 8166
0 3781 5 2 1 3780
0 3782 7 1 2 8169 8171
0 3783 7 2 2 3772 3782
0 3784 5 1 1 8173
0 3785 7 1 2 5007 8174
0 3786 5 2 1 3785
0 3787 7 1 2 3777 8172
0 3788 5 1 1 3787
0 3789 7 2 2 8170 3788
0 3790 5 1 1 8177
0 3791 7 1 2 5008 8178
0 3792 5 2 1 3791
0 3793 7 1 2 3784 8179
0 3794 5 1 1 3793
0 3795 7 2 2 8175 3794
0 3796 5 1 1 8181
0 3797 7 1 2 5373 3796
0 3798 5 1 1 3797
0 3799 7 1 2 5381 3790
0 3800 5 1 1 3799
0 3801 7 1 2 8176 8180
0 3802 7 2 2 3800 3801
0 3803 5 1 1 8183
0 3804 7 1 2 4999 8184
0 3805 5 2 1 3804
0 3806 7 1 2 5000 8182
0 3807 5 2 1 3806
0 3808 7 1 2 8185 8187
0 3809 7 2 2 3798 3808
0 3810 5 1 1 8189
0 3811 7 1 2 4991 8190
0 3812 5 2 1 3811
0 3813 7 1 2 3803 8188
0 3814 5 1 1 3813
0 3815 7 2 2 8186 3814
0 3816 5 1 1 8193
0 3817 7 1 2 4992 8194
0 3818 5 2 1 3817
0 3819 7 1 2 3810 8195
0 3820 5 1 1 3819
0 3821 7 2 2 8191 3820
0 3822 5 1 1 8197
0 3823 7 1 2 5357 3822
0 3824 5 1 1 3823
0 3825 7 1 2 5365 3816
0 3826 5 1 1 3825
0 3827 7 1 2 8192 8196
0 3828 7 2 2 3826 3827
0 3829 5 1 1 8199
0 3830 7 1 2 4983 8200
0 3831 5 2 1 3830
0 3832 7 1 2 4984 8198
0 3833 5 2 1 3832
0 3834 7 1 2 8201 8203
0 3835 7 2 2 3824 3834
0 3836 5 1 1 8205
0 3837 7 1 2 4975 8206
0 3838 5 2 1 3837
0 3839 7 1 2 3829 8204
0 3840 5 1 1 3839
0 3841 7 2 2 8202 3840
0 3842 5 1 1 8209
0 3843 7 1 2 4976 8210
0 3844 5 2 1 3843
0 3845 7 1 2 3836 8211
0 3846 5 1 1 3845
0 3847 7 2 2 8207 3846
0 3848 5 1 1 8213
0 3849 7 1 2 5341 3848
0 3850 5 1 1 3849
0 3851 7 1 2 5349 3842
0 3852 5 1 1 3851
0 3853 7 1 2 8208 8212
0 3854 7 2 2 3852 3853
0 3855 5 1 1 8215
0 3856 7 1 2 4967 8216
0 3857 5 2 1 3856
0 3858 7 1 2 4968 8214
0 3859 5 2 1 3858
0 3860 7 1 2 8217 8219
0 3861 7 2 2 3850 3860
0 3862 5 1 1 8221
0 3863 7 1 2 4959 8222
0 3864 5 2 1 3863
0 3865 7 1 2 3855 8220
0 3866 5 1 1 3865
0 3867 7 2 2 8218 3866
0 3868 5 1 1 8225
0 3869 7 1 2 4960 8226
0 3870 5 2 1 3869
0 3871 7 1 2 3862 8227
0 3872 5 1 1 3871
0 3873 7 2 2 8223 3872
0 3874 5 1 1 8229
0 3875 7 1 2 5325 3874
0 3876 5 1 1 3875
0 3877 7 1 2 5333 3868
0 3878 5 1 1 3877
0 3879 7 1 2 8224 8228
0 3880 7 2 2 3878 3879
0 3881 5 1 1 8231
0 3882 7 1 2 4951 8232
0 3883 5 2 1 3882
0 3884 7 1 2 4952 8230
0 3885 5 2 1 3884
0 3886 7 1 2 8233 8235
0 3887 7 2 2 3876 3886
0 3888 5 1 1 8237
0 3889 7 1 2 4943 8238
0 3890 5 2 1 3889
0 3891 7 1 2 3881 8236
0 3892 5 1 1 3891
0 3893 7 2 2 8234 3892
0 3894 5 1 1 8241
0 3895 7 1 2 4944 8242
0 3896 5 2 1 3895
0 3897 7 1 2 3888 8243
0 3898 5 1 1 3897
0 3899 7 2 2 8239 3898
0 3900 5 1 1 8245
0 3901 7 1 2 5310 3900
0 3902 5 1 1 3901
0 3903 7 1 2 5317 3894
0 3904 5 1 1 3903
0 3905 7 1 2 8240 8244
0 3906 7 2 2 3904 3905
0 3907 5 1 1 8247
0 3908 7 1 2 4935 8248
0 3909 5 2 1 3908
0 3910 7 1 2 4936 8246
0 3911 5 2 1 3910
0 3912 7 1 2 8249 8251
0 3913 7 2 2 3902 3912
0 3914 5 1 1 8253
0 3915 7 1 2 4927 8254
0 3916 5 2 1 3915
0 3917 7 1 2 3907 8252
0 3918 5 1 1 3917
0 3919 7 2 2 8250 3918
0 3920 5 1 1 8257
0 3921 7 1 2 4928 8258
0 3922 5 2 1 3921
0 3923 7 1 2 3914 8259
0 3924 5 1 1 3923
0 3925 7 2 2 8255 3924
0 3926 5 1 1 8261
0 3927 7 1 2 5296 3926
0 3928 5 1 1 3927
0 3929 7 1 2 5303 3920
0 3930 5 1 1 3929
0 3931 7 1 2 8256 8260
0 3932 7 2 2 3930 3931
0 3933 5 1 1 8263
0 3934 7 1 2 4919 8264
0 3935 5 2 1 3934
0 3936 7 1 2 4920 8262
0 3937 5 2 1 3936
0 3938 7 1 2 8265 8267
0 3939 7 2 2 3928 3938
0 3940 5 1 1 8269
0 3941 7 1 2 4911 8270
0 3942 5 2 1 3941
0 3943 7 1 2 3933 8268
0 3944 5 1 1 3943
0 3945 7 2 2 8266 3944
0 3946 5 1 1 8273
0 3947 7 1 2 4912 8274
0 3948 5 2 1 3947
0 3949 7 1 2 3940 8275
0 3950 5 1 1 3949
0 3951 7 2 2 8271 3950
0 3952 5 1 1 8277
0 3953 7 1 2 5282 3952
0 3954 5 1 1 3953
0 3955 7 1 2 5289 3946
0 3956 5 1 1 3955
0 3957 7 1 2 8272 8276
0 3958 7 2 2 3956 3957
0 3959 5 1 1 8279
0 3960 7 1 2 4903 8280
0 3961 5 2 1 3960
0 3962 7 1 2 4904 8278
0 3963 5 2 1 3962
0 3964 7 1 2 8281 8283
0 3965 7 2 2 3954 3964
0 3966 5 1 1 8285
0 3967 7 1 2 4895 8286
0 3968 5 2 1 3967
0 3969 7 1 2 3959 8284
0 3970 5 1 1 3969
0 3971 7 2 2 8282 3970
0 3972 5 1 1 8289
0 3973 7 1 2 4896 8290
0 3974 5 2 1 3973
0 3975 7 1 2 3966 8291
0 3976 5 1 1 3975
0 3977 7 2 2 8287 3976
0 3978 5 1 1 8293
0 3979 7 1 2 5268 3978
0 3980 5 1 1 3979
0 3981 7 1 2 5275 3972
0 3982 5 1 1 3981
0 3983 7 1 2 8288 8292
0 3984 7 2 2 3982 3983
0 3985 5 1 1 8295
0 3986 7 1 2 4887 8296
0 3987 5 2 1 3986
0 3988 7 1 2 4888 8294
0 3989 5 2 1 3988
0 3990 7 1 2 8297 8299
0 3991 7 2 2 3980 3990
0 3992 5 1 1 8301
0 3993 7 1 2 4879 8302
0 3994 5 2 1 3993
0 3995 7 1 2 3985 8300
0 3996 5 1 1 3995
0 3997 7 2 2 8298 3996
0 3998 5 1 1 8305
0 3999 7 1 2 4880 8306
0 4000 5 2 1 3999
0 4001 7 1 2 3992 8307
0 4002 5 1 1 4001
0 4003 7 2 2 8303 4002
0 4004 5 1 1 8309
0 4005 7 1 2 5254 4004
0 4006 5 1 1 4005
0 4007 7 1 2 5261 3998
0 4008 5 1 1 4007
0 4009 7 1 2 8304 8308
0 4010 7 2 2 4008 4009
0 4011 5 1 1 8311
0 4012 7 1 2 4871 8312
0 4013 5 2 1 4012
0 4014 7 1 2 4872 8310
0 4015 5 2 1 4014
0 4016 7 1 2 8313 8315
0 4017 7 2 2 4006 4016
0 4018 5 1 1 8317
0 4019 7 1 2 4863 8318
0 4020 5 2 1 4019
0 4021 7 1 2 4011 8316
0 4022 5 1 1 4021
0 4023 7 2 2 8314 4022
0 4024 5 1 1 8321
0 4025 7 1 2 4864 8322
0 4026 5 2 1 4025
0 4027 7 1 2 4018 8323
0 4028 5 1 1 4027
0 4029 7 2 2 8319 4028
0 4030 5 1 1 8325
0 4031 7 1 2 5240 4030
0 4032 5 1 1 4031
0 4033 7 1 2 5247 4024
0 4034 5 1 1 4033
0 4035 7 1 2 8320 8324
0 4036 7 2 2 4034 4035
0 4037 5 1 1 8327
0 4038 7 1 2 4855 8328
0 4039 5 2 1 4038
0 4040 7 1 2 4856 8326
0 4041 5 2 1 4040
0 4042 7 1 2 8329 8331
0 4043 7 2 2 4032 4042
0 4044 5 1 1 8333
0 4045 7 1 2 4847 8334
0 4046 5 2 1 4045
0 4047 7 1 2 4037 8332
0 4048 5 1 1 4047
0 4049 7 2 2 8330 4048
0 4050 5 1 1 8337
0 4051 7 1 2 4848 8338
0 4052 5 2 1 4051
0 4053 7 1 2 4044 8339
0 4054 5 1 1 4053
0 4055 7 2 2 8335 4054
0 4056 5 1 1 8341
0 4057 7 1 2 5226 4056
0 4058 5 1 1 4057
0 4059 7 1 2 5233 4050
0 4060 5 1 1 4059
0 4061 7 1 2 8336 8340
0 4062 7 2 2 4060 4061
0 4063 5 1 1 8343
0 4064 7 1 2 4839 8344
0 4065 5 2 1 4064
0 4066 7 1 2 4840 8342
0 4067 5 2 1 4066
0 4068 7 1 2 8345 8347
0 4069 7 2 2 4058 4068
0 4070 5 1 1 8349
0 4071 7 1 2 4831 8350
0 4072 5 2 1 4071
0 4073 7 1 2 4063 8348
0 4074 5 1 1 4073
0 4075 7 2 2 8346 4074
0 4076 5 1 1 8353
0 4077 7 1 2 4832 8354
0 4078 5 2 1 4077
0 4079 7 1 2 4070 8355
0 4080 5 1 1 4079
0 4081 7 2 2 8351 4080
0 4082 5 1 1 8357
0 4083 7 1 2 5212 4082
0 4084 5 1 1 4083
0 4085 7 1 2 5219 4076
0 4086 5 1 1 4085
0 4087 7 1 2 8352 8356
0 4088 7 2 2 4086 4087
0 4089 5 1 1 8359
0 4090 7 1 2 4823 8360
0 4091 5 2 1 4090
0 4092 7 1 2 4824 8358
0 4093 5 2 1 4092
0 4094 7 1 2 8361 8363
0 4095 7 2 2 4084 4094
0 4096 5 1 1 8365
0 4097 7 1 2 4815 8366
0 4098 5 2 1 4097
0 4099 7 1 2 4089 8364
0 4100 5 1 1 4099
0 4101 7 2 2 8362 4100
0 4102 5 1 1 8369
0 4103 7 1 2 4816 8370
0 4104 5 2 1 4103
0 4105 7 1 2 4096 8371
0 4106 5 1 1 4105
0 4107 7 2 2 8367 4106
0 4108 5 1 1 8373
0 4109 7 1 2 5198 4108
0 4110 5 1 1 4109
0 4111 7 1 2 5205 4102
0 4112 5 1 1 4111
0 4113 7 1 2 8368 8372
0 4114 7 2 2 4112 4113
0 4115 5 1 1 8375
0 4116 7 1 2 4806 8376
0 4117 5 2 1 4116
0 4118 7 1 2 4807 8374
0 4119 5 2 1 4118
0 4120 7 1 2 8377 8379
0 4121 7 2 2 4110 4120
0 4122 5 1 1 8381
0 4123 7 1 2 4797 4122
0 4124 5 1 1 4123
0 4125 7 1 2 4115 8380
0 4126 5 1 1 4125
0 4127 7 1 2 8378 4126
0 4128 5 1 1 4127
0 4129 7 2 2 4791 4128
0 4130 5 1 1 8383
0 4131 7 1 2 4124 8384
0 4132 5 1 1 4131
0 4133 7 1 2 5184 8382
0 4134 5 1 1 4133
0 4135 7 1 2 4798 4130
0 4136 7 1 2 4134 4135
0 4137 5 1 1 4136
0 4138 7 1 2 4132 4137
0 4139 5 1 1 4138
0 4140 7 1 2 4808 3490
0 4141 5 1 1 4140
0 4142 7 1 2 5185 4799
0 4143 7 1 2 4141 4142
0 4144 7 1 2 8019 4143
0 4145 7 1 2 3512 4144
0 4146 7 1 2 3537 4145
0 4147 5 1 1 4146
0 4148 7 1 2 4139 4147
0 4149 7 1 2 3540 4148
0 4150 7 1 2 2466 4149
0 4151 7 2 2 1475 4150
0 4152 5 1 1 8385
0 4153 7 1 2 5199 5311
0 4154 5 2 1 4153
0 4155 7 1 2 4809 4937
0 4156 5 2 1 4155
0 4157 7 1 2 5192 5304
0 4158 5 2 1 4157
0 4159 7 1 2 4800 4929
0 4160 5 2 1 4159
0 4161 7 2 2 4792 4921
0 4162 5 3 1 8395
0 4163 7 1 2 8393 8397
0 4164 5 1 1 4163
0 4165 7 2 2 8391 4164
0 4166 5 2 1 8400
0 4167 7 1 2 8389 8402
0 4168 5 1 1 4167
0 4169 7 2 2 8387 4168
0 4170 5 1 1 8404
0 4171 7 1 2 5206 4170
0 4172 5 2 1 4171
0 4173 7 1 2 4817 8405
0 4174 5 2 1 4173
0 4175 7 1 2 5318 8408
0 4176 5 1 1 4175
0 4177 7 2 2 8406 4176
0 4178 5 1 1 8410
0 4179 7 1 2 5213 4178
0 4180 5 2 1 4179
0 4181 7 1 2 4825 8411
0 4182 5 2 1 4181
0 4183 7 1 2 5326 8414
0 4184 5 1 1 4183
0 4185 7 2 2 8412 4184
0 4186 5 1 1 8416
0 4187 7 1 2 5220 4186
0 4188 5 2 1 4187
0 4189 7 1 2 4833 8417
0 4190 5 2 1 4189
0 4191 7 1 2 5334 8420
0 4192 5 1 1 4191
0 4193 7 2 2 8418 4192
0 4194 5 1 1 8422
0 4195 7 1 2 5227 4194
0 4196 5 2 1 4195
0 4197 7 1 2 4841 8423
0 4198 5 2 1 4197
0 4199 7 1 2 5342 8426
0 4200 5 1 1 4199
0 4201 7 2 2 8424 4200
0 4202 5 1 1 8428
0 4203 7 1 2 5234 4202
0 4204 5 2 1 4203
0 4205 7 1 2 4849 8429
0 4206 5 2 1 4205
0 4207 7 1 2 5350 8432
0 4208 5 1 1 4207
0 4209 7 2 2 8430 4208
0 4210 5 1 1 8434
0 4211 7 1 2 5241 4210
0 4212 5 2 1 4211
0 4213 7 1 2 4857 8435
0 4214 5 2 1 4213
0 4215 7 1 2 5358 8438
0 4216 5 1 1 4215
0 4217 7 2 2 8436 4216
0 4218 5 1 1 8440
0 4219 7 1 2 5248 4218
0 4220 5 2 1 4219
0 4221 7 1 2 4865 8441
0 4222 5 2 1 4221
0 4223 7 1 2 5366 8444
0 4224 5 1 1 4223
0 4225 7 2 2 8442 4224
0 4226 5 1 1 8446
0 4227 7 1 2 5255 4226
0 4228 5 2 1 4227
0 4229 7 1 2 4873 8447
0 4230 5 2 1 4229
0 4231 7 1 2 5374 8450
0 4232 5 1 1 4231
0 4233 7 2 2 8448 4232
0 4234 5 1 1 8452
0 4235 7 1 2 5262 4234
0 4236 5 2 1 4235
0 4237 7 1 2 4881 8453
0 4238 5 2 1 4237
0 4239 7 1 2 5382 8456
0 4240 5 1 1 4239
0 4241 7 2 2 8454 4240
0 4242 5 1 1 8458
0 4243 7 1 2 5269 4242
0 4244 5 2 1 4243
0 4245 7 1 2 4889 8459
0 4246 5 2 1 4245
0 4247 7 1 2 5390 8462
0 4248 5 1 1 4247
0 4249 7 2 2 8460 4248
0 4250 5 1 1 8464
0 4251 7 1 2 5276 4250
0 4252 5 2 1 4251
0 4253 7 1 2 4897 8465
0 4254 5 2 1 4253
0 4255 7 1 2 5398 8468
0 4256 5 1 1 4255
0 4257 7 2 2 8466 4256
0 4258 5 1 1 8470
0 4259 7 1 2 5283 4258
0 4260 5 2 1 4259
0 4261 7 1 2 4905 8471
0 4262 5 2 1 4261
0 4263 7 2 2 8472 8474
0 4264 5 1 1 8476
0 4265 7 1 2 5033 8477
0 4266 5 1 1 4265
0 4267 7 1 2 5406 4264
0 4268 5 1 1 4267
0 4269 7 2 2 4266 4268
0 4270 5 1 1 8478
0 4271 7 1 2 5164 4270
0 4272 5 3 1 4271
0 4273 7 2 2 8467 8469
0 4274 5 1 1 8483
0 4275 7 1 2 5025 8484
0 4276 5 1 1 4275
0 4277 7 1 2 5399 4274
0 4278 5 1 1 4277
0 4279 7 2 2 4276 4278
0 4280 5 1 1 8485
0 4281 7 1 2 5155 4280
0 4282 5 3 1 4281
0 4283 7 1 2 5514 8486
0 4284 5 4 1 4283
0 4285 7 2 2 8461 8463
0 4286 5 1 1 8494
0 4287 7 1 2 5017 8495
0 4288 5 1 1 4287
0 4289 7 1 2 5391 4286
0 4290 5 1 1 4289
0 4291 7 2 2 4288 4290
0 4292 5 1 1 8496
0 4293 7 1 2 5145 4292
0 4294 5 3 1 4293
0 4295 7 1 2 5507 8497
0 4296 5 4 1 4295
0 4297 7 2 2 8455 8457
0 4298 5 1 1 8505
0 4299 7 1 2 5009 8506
0 4300 5 1 1 4299
0 4301 7 1 2 5383 4298
0 4302 5 1 1 4301
0 4303 7 2 2 4300 4302
0 4304 5 1 1 8507
0 4305 7 1 2 5137 4304
0 4306 5 4 1 4305
0 4307 7 2 2 8449 8451
0 4308 5 1 1 8513
0 4309 7 1 2 5001 8514
0 4310 5 1 1 4309
0 4311 7 1 2 5375 4308
0 4312 5 1 1 4311
0 4313 7 2 2 4310 4312
0 4314 5 1 1 8515
0 4315 7 3 2 5492 8516
0 4316 5 2 1 8517
0 4317 7 1 2 5499 8508
0 4318 5 4 1 4317
0 4319 7 2 2 8520 8522
0 4320 7 2 2 8443 8445
0 4321 5 1 1 8528
0 4322 7 1 2 4993 8529
0 4323 5 1 1 4322
0 4324 7 1 2 5367 4321
0 4325 5 1 1 4324
0 4326 7 2 2 4323 4325
0 4327 5 1 1 8530
0 4328 7 1 2 5121 4327
0 4329 5 3 1 4328
0 4330 7 1 2 5485 8531
0 4331 5 4 1 4330
0 4332 7 2 2 8437 8439
0 4333 5 1 1 8539
0 4334 7 1 2 4985 8540
0 4335 5 1 1 4334
0 4336 7 1 2 5359 4333
0 4337 5 1 1 4336
0 4338 7 2 2 4335 4337
0 4339 5 1 1 8541
0 4340 7 1 2 5113 4339
0 4341 5 3 1 4340
0 4342 7 1 2 5478 8542
0 4343 5 4 1 4342
0 4344 7 2 2 8431 8433
0 4345 5 1 1 8550
0 4346 7 1 2 4977 8551
0 4347 5 1 1 4346
0 4348 7 1 2 5351 4345
0 4349 5 1 1 4348
0 4350 7 2 2 4347 4349
0 4351 5 1 1 8552
0 4352 7 1 2 5105 4351
0 4353 5 4 1 4352
0 4354 7 1 2 5471 8553
0 4355 5 4 1 4354
0 4356 7 2 2 8425 8427
0 4357 5 1 1 8562
0 4358 7 1 2 4969 8563
0 4359 5 1 1 4358
0 4360 7 1 2 5343 4357
0 4361 5 1 1 4360
0 4362 7 2 2 4359 4361
0 4363 5 1 1 8564
0 4364 7 1 2 5097 4363
0 4365 5 4 1 4364
0 4366 7 2 2 8419 8421
0 4367 5 1 1 8570
0 4368 7 1 2 4961 8571
0 4369 5 1 1 4368
0 4370 7 1 2 5335 4367
0 4371 5 1 1 4370
0 4372 7 2 2 4369 4371
0 4373 5 1 1 8572
0 4374 7 1 2 5089 4373
0 4375 5 4 1 4374
0 4376 7 2 2 8413 8415
0 4377 5 1 1 8578
0 4378 7 1 2 4953 8579
0 4379 5 1 1 4378
0 4380 7 1 2 5327 4377
0 4381 5 1 1 4380
0 4382 7 2 2 4379 4381
0 4383 5 1 1 8580
0 4384 7 1 2 5450 8581
0 4385 5 4 1 4384
0 4386 7 1 2 5081 4383
0 4387 5 3 1 4386
0 4388 7 2 2 8407 8409
0 4389 5 1 1 8589
0 4390 7 1 2 4945 8590
0 4391 5 1 1 4390
0 4392 7 1 2 5319 4389
0 4393 5 1 1 4392
0 4394 7 2 2 4391 4393
0 4395 5 1 1 8591
0 4396 7 1 2 5443 8592
0 4397 5 4 1 4396
0 4398 7 1 2 5073 4395
0 4399 5 3 1 4398
0 4400 7 1 2 5186 5297
0 4401 5 1 1 4400
0 4402 7 2 2 8398 4401
0 4403 5 1 1 8600
0 4404 7 1 2 5049 4403
0 4405 5 1 1 4404
0 4406 7 2 2 8388 8390
0 4407 5 1 1 8602
0 4408 7 1 2 8401 4407
0 4409 5 1 1 4408
0 4410 7 1 2 8403 8603
0 4411 5 1 1 4410
0 4412 7 2 2 4409 4411
0 4413 5 1 1 8604
0 4414 7 1 2 5065 8605
0 4415 5 2 1 4414
0 4416 7 2 2 8392 8394
0 4417 5 1 1 8608
0 4418 7 1 2 8396 4417
0 4419 5 1 1 4418
0 4420 7 1 2 8399 8609
0 4421 5 1 1 4420
0 4422 7 2 2 4419 4421
0 4423 5 1 1 8610
0 4424 7 1 2 5057 8611
0 4425 5 1 1 4424
0 4426 7 2 2 8606 4425
0 4427 5 1 1 8612
0 4428 7 2 2 4405 8613
0 4429 5 1 1 8614
0 4430 7 2 2 5429 4423
0 4431 5 1 1 8616
0 4432 7 1 2 8607 8617
0 4433 5 1 1 4432
0 4434 7 1 2 5436 4413
0 4435 5 3 1 4434
0 4436 7 1 2 4433 8618
0 4437 7 2 2 4429 4436
0 4438 5 2 1 8621
0 4439 7 1 2 8597 8623
0 4440 5 1 1 4439
0 4441 7 2 2 8593 4440
0 4442 5 2 1 8625
0 4443 7 1 2 8586 8627
0 4444 5 1 1 4443
0 4445 7 2 2 8582 4444
0 4446 5 1 1 8629
0 4447 7 1 2 8574 4446
0 4448 5 2 1 4447
0 4449 7 1 2 5464 8565
0 4450 5 4 1 4449
0 4451 7 1 2 5457 8573
0 4452 5 4 1 4451
0 4453 7 2 2 8633 8637
0 4454 7 1 2 8631 8641
0 4455 5 1 1 4454
0 4456 7 2 2 8566 4455
0 4457 5 1 1 8643
0 4458 7 1 2 8558 4457
0 4459 5 1 1 4458
0 4460 7 2 2 8554 4459
0 4461 5 2 1 8645
0 4462 7 1 2 8546 8647
0 4463 5 1 1 4462
0 4464 7 2 2 8543 4463
0 4465 5 2 1 8649
0 4466 7 1 2 8535 8651
0 4467 5 1 1 4466
0 4468 7 3 2 8532 4467
0 4469 5 1 1 8653
0 4470 7 3 2 5129 4314
0 4471 5 2 1 8656
0 4472 7 1 2 8654 8659
0 4473 5 1 1 4472
0 4474 7 1 2 8526 4473
0 4475 5 1 1 4474
0 4476 7 1 2 8509 4475
0 4477 5 2 1 4476
0 4478 7 1 2 8501 8661
0 4479 5 1 1 4478
0 4480 7 2 2 8498 4479
0 4481 5 2 1 8663
0 4482 7 1 2 8490 8665
0 4483 5 1 1 4482
0 4484 7 2 2 8487 4483
0 4485 5 2 1 8667
0 4486 7 1 2 5519 8479
0 4487 5 4 1 4486
0 4488 7 1 2 8669 8671
0 4489 5 1 1 4488
0 4490 7 2 2 8480 4489
0 4491 5 2 1 8675
0 4492 7 1 2 5407 8475
0 4493 5 1 1 4492
0 4494 7 2 2 8473 4493
0 4495 5 1 1 8679
0 4496 7 1 2 5290 4495
0 4497 5 2 1 4496
0 4498 7 1 2 4913 8680
0 4499 5 2 1 4498
0 4500 7 2 2 8681 8683
0 4501 5 1 1 8685
0 4502 7 1 2 5041 8686
0 4503 5 1 1 4502
0 4504 7 1 2 5414 4501
0 4505 5 1 1 4504
0 4506 7 2 2 4503 4505
0 4507 5 1 1 8687
0 4508 7 1 2 5172 4507
0 4509 5 3 1 4508
0 4510 7 2 2 5523 8688
0 4511 5 3 1 8692
0 4512 7 2 2 8689 8694
0 4513 5 1 1 8697
0 4514 7 1 2 8676 4513
0 4515 5 1 1 4514
0 4516 7 1 2 8677 8698
0 4517 5 2 1 4516
0 4518 7 3 2 8481 8672
0 4519 5 2 1 8701
0 4520 7 1 2 8670 8704
0 4521 5 1 1 4520
0 4522 7 1 2 8668 8702
0 4523 5 1 1 4522
0 4524 7 1 2 4521 4523
0 4525 5 1 1 4524
0 4526 7 1 2 5415 8684
0 4527 5 1 1 4526
0 4528 7 2 2 8682 4527
0 4529 5 1 1 8706
0 4530 7 2 2 5179 4529
0 4531 5 2 1 8708
0 4532 7 3 2 8488 8491
0 4533 5 2 1 8712
0 4534 7 1 2 8664 8715
0 4535 5 1 1 4534
0 4536 7 1 2 8666 8713
0 4537 5 1 1 4536
0 4538 7 3 2 8499 8502
0 4539 5 2 1 8717
0 4540 7 1 2 8510 8720
0 4541 5 1 1 4540
0 4542 7 1 2 8662 8718
0 4543 5 1 1 4542
0 4544 7 1 2 8511 8523
0 4545 5 2 1 4544
0 4546 7 1 2 4469 8657
0 4547 5 1 1 4546
0 4548 7 1 2 8722 4547
0 4549 5 1 1 4548
0 4550 7 1 2 8518 8655
0 4551 5 1 1 4550
0 4552 7 3 2 8533 8536
0 4553 5 2 1 8724
0 4554 7 1 2 8650 8727
0 4555 5 1 1 4554
0 4556 7 1 2 8652 8725
0 4557 5 1 1 4556
0 4558 7 1 2 4555 4557
0 4559 5 1 1 4558
0 4560 7 3 2 8544 8547
0 4561 5 2 1 8729
0 4562 7 1 2 8648 8732
0 4563 5 1 1 4562
0 4564 7 1 2 8646 8730
0 4565 5 1 1 4564
0 4566 7 2 2 8555 8559
0 4567 5 2 1 8734
0 4568 7 1 2 8634 8736
0 4569 5 1 1 4568
0 4570 7 1 2 8644 8735
0 4571 5 1 1 4570
0 4572 7 2 2 8567 8635
0 4573 7 1 2 8632 8738
0 4574 5 1 1 4573
0 4575 7 1 2 8638 4574
0 4576 5 1 1 4575
0 4577 7 1 2 8575 8639
0 4578 5 2 1 4577
0 4579 7 1 2 8630 8740
0 4580 5 1 1 4579
0 4581 7 3 2 8583 8587
0 4582 5 2 1 8742
0 4583 7 1 2 8626 8743
0 4584 5 1 1 4583
0 4585 7 3 2 8594 8598
0 4586 5 2 1 8747
0 4587 7 1 2 8624 8748
0 4588 5 1 1 4587
0 4589 7 1 2 5422 8601
0 4590 5 1 1 4589
0 4591 7 1 2 4431 4590
0 4592 7 3 2 8619 4591
0 4593 5 1 1 8752
0 4594 7 1 2 8615 8753
0 4595 5 2 1 4594
0 4596 7 1 2 8622 8750
0 4597 5 1 1 4596
0 4598 7 1 2 8755 4597
0 4599 7 1 2 4588 4598
0 4600 5 1 1 4599
0 4601 7 1 2 8628 8745
0 4602 5 1 1 4601
0 4603 7 1 2 4600 4602
0 4604 7 1 2 4584 4603
0 4605 5 1 1 4604
0 4606 7 1 2 4580 4605
0 4607 7 1 2 4576 4606
0 4608 7 1 2 4571 4607
0 4609 7 1 2 4569 4608
0 4610 7 1 2 4565 4609
0 4611 7 1 2 4563 4610
0 4612 7 1 2 4559 4611
0 4613 5 1 1 4612
0 4614 7 1 2 4551 4613
0 4615 7 1 2 4549 4614
0 4616 7 1 2 4543 4615
0 4617 7 1 2 4541 4616
0 4618 7 1 2 4537 4617
0 4619 7 1 2 4535 4618
0 4620 7 1 2 8710 4619
0 4621 7 1 2 4525 4620
0 4622 7 1 2 8699 4621
0 4623 7 1 2 4515 4622
0 4624 7 2 2 5529 8707
0 4625 5 3 1 8757
0 4626 7 1 2 8678 8695
0 4627 5 1 1 4626
0 4628 7 2 2 8690 4627
0 4629 5 1 1 8762
0 4630 7 1 2 8759 4629
0 4631 5 2 1 4630
0 4632 7 1 2 8758 8763
0 4633 5 1 1 4632
0 4634 7 1 2 8764 4633
0 4635 7 1 2 4623 4634
0 4636 5 1 1 4635
0 4637 7 1 2 4427 8620
0 4638 5 1 1 4637
0 4639 7 2 2 4593 4638
0 4640 5 2 1 8766
0 4641 7 1 2 8595 8768
0 4642 5 1 1 4641
0 4643 7 2 2 8599 4642
0 4644 5 2 1 8770
0 4645 7 1 2 8584 8772
0 4646 5 1 1 4645
0 4647 7 2 2 8588 4646
0 4648 5 1 1 8774
0 4649 7 1 2 8640 4648
0 4650 5 2 1 4649
0 4651 7 1 2 8576 8776
0 4652 7 1 2 8568 4651
0 4653 5 1 1 4652
0 4654 7 1 2 8636 4653
0 4655 7 2 2 8560 4654
0 4656 5 1 1 8778
0 4657 7 2 2 8556 4656
0 4658 5 2 1 8780
0 4659 7 1 2 8548 8782
0 4660 5 1 1 4659
0 4661 7 2 2 8545 4660
0 4662 5 2 1 8784
0 4663 7 1 2 8537 8786
0 4664 5 1 1 4663
0 4665 7 2 2 8534 4664
0 4666 5 2 1 8788
0 4667 7 1 2 8521 8790
0 4668 5 1 1 4667
0 4669 7 1 2 8660 4668
0 4670 7 1 2 8512 4669
0 4671 5 1 1 4670
0 4672 7 2 2 8524 4671
0 4673 5 1 1 8792
0 4674 7 1 2 8503 8793
0 4675 5 1 1 4674
0 4676 7 2 2 8500 4675
0 4677 5 2 1 8794
0 4678 7 1 2 8492 8796
0 4679 5 1 1 4678
0 4680 7 2 2 8489 4679
0 4681 5 2 1 8798
0 4682 7 1 2 8673 8800
0 4683 5 1 1 4682
0 4684 7 3 2 8482 4683
0 4685 5 1 1 8802
0 4686 7 1 2 8700 4685
0 4687 5 1 1 4686
0 4688 7 1 2 8691 8803
0 4689 5 1 1 4688
0 4690 7 2 2 8696 8711
0 4691 7 1 2 4689 8805
0 4692 7 1 2 4687 4691
0 4693 5 1 1 4692
0 4694 7 1 2 8709 8804
0 4695 7 1 2 8693 4694
0 4696 5 1 1 4695
0 4697 7 1 2 4693 4696
0 4698 5 1 1 4697
0 4699 7 1 2 8716 8797
0 4700 5 1 1 4699
0 4701 7 1 2 8714 8795
0 4702 5 1 1 4701
0 4703 7 1 2 8719 4673
0 4704 5 1 1 4703
0 4705 7 1 2 8525 8721
0 4706 5 1 1 4705
0 4707 7 1 2 8519 8789
0 4708 5 1 1 4707
0 4709 7 1 2 8723 4708
0 4710 5 1 1 4709
0 4711 7 1 2 8658 8791
0 4712 5 1 1 4711
0 4713 7 1 2 8728 8785
0 4714 5 1 1 4713
0 4715 7 1 2 8726 8787
0 4716 5 1 1 4715
0 4717 7 1 2 8733 8781
0 4718 5 1 1 4717
0 4719 7 1 2 8731 8783
0 4720 5 1 1 4719
0 4721 7 1 2 8569 8737
0 4722 5 1 1 4721
0 4723 7 1 2 8557 8779
0 4724 5 1 1 4723
0 4725 7 1 2 8739 8777
0 4726 5 1 1 4725
0 4727 7 1 2 8577 4726
0 4728 5 1 1 4727
0 4729 7 1 2 8741 8775
0 4730 5 1 1 4729
0 4731 7 1 2 8744 8771
0 4732 5 1 1 4731
0 4733 7 1 2 8749 8769
0 4734 5 1 1 4733
0 4735 7 1 2 8751 8767
0 4736 5 1 1 4735
0 4737 7 1 2 8756 4736
0 4738 7 1 2 4734 4737
0 4739 5 1 1 4738
0 4740 7 1 2 8746 8773
0 4741 5 1 1 4740
0 4742 7 1 2 4739 4741
0 4743 7 1 2 4732 4742
0 4744 5 1 1 4743
0 4745 7 1 2 4730 4744
0 4746 7 1 2 4728 4745
0 4747 7 1 2 4724 4746
0 4748 7 1 2 4722 4747
0 4749 7 1 2 4720 4748
0 4750 7 1 2 4718 4749
0 4751 7 1 2 4716 4750
0 4752 7 1 2 4714 4751
0 4753 5 1 1 4752
0 4754 7 1 2 4712 4753
0 4755 7 1 2 4710 4754
0 4756 7 1 2 4706 4755
0 4757 7 1 2 4704 4756
0 4758 7 1 2 4702 4757
0 4759 7 1 2 4700 4758
0 4760 7 1 2 8760 4759
0 4761 7 1 2 8705 8801
0 4762 5 1 1 4761
0 4763 7 1 2 8703 8799
0 4764 5 1 1 4763
0 4765 7 1 2 4762 4764
0 4766 7 1 2 4760 4765
0 4767 7 1 2 4698 4766
0 4768 5 1 1 4767
0 4769 7 1 2 4636 4768
0 4770 7 1 2 4152 4769
0 4771 5 1 1 4770
0 4772 7 1 2 8596 8754
0 4773 7 1 2 8585 4772
0 4774 7 1 2 8642 4773
0 4775 7 1 2 8561 4774
0 4776 7 1 2 8549 4775
0 4777 7 1 2 8538 4776
0 4778 7 1 2 8527 4777
0 4779 7 1 2 8504 4778
0 4780 7 1 2 8493 4779
0 4781 7 1 2 8674 4780
0 4782 7 1 2 8761 4781
0 4783 7 1 2 8806 4782
0 4784 7 1 2 8765 4783
0 4785 5 1 1 4784
0 4786 7 1 2 8386 4785
0 4787 5 1 1 4786
3 9999 7 0 2 4771 4787
