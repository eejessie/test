1 0 0 3 0
2 11 1 0
2 12 1 0
2 13 1 0
1 1 0 2 0
2 14 1 1
2 15 1 1
1 2 0 2 0
2 16 1 2
2 39 1 2
1 3 0 2 0
2 59 1 3
2 78 1 3
1 4 0 2 0
2 101 1 4
2 121 1 4
1 5 0 2 0
2 124 1 5
2 125 1 5
1 6 0 2 0
2 126 1 6
2 127 1 6
1 7 0 2 0
2 128 1 7
2 129 1 7
1 8 0 2 0
2 130 1 8
2 131 1 8
1 9 0 2 0
2 132 1 9
2 133 1 9
1 10 0 2 0
2 134 1 10
2 135 1 10
2 136 1 17
2 137 1 17
2 138 1 29
2 139 1 29
2 140 1 29
2 141 1 31
2 142 1 31
2 143 1 31
2 144 1 32
2 145 1 32
2 146 1 43
2 147 1 43
2 148 1 43
2 149 1 45
2 150 1 45
2 151 1 45
2 152 1 45
2 153 1 47
2 154 1 47
2 155 1 47
2 156 1 48
2 157 1 48
2 158 1 55
2 159 1 55
2 160 1 55
2 161 1 63
2 162 1 63
2 163 1 63
2 164 1 63
2 165 1 65
2 166 1 65
2 167 1 65
2 168 1 73
2 169 1 73
2 170 1 73
2 171 1 80
2 172 1 80
2 173 1 82
2 174 1 82
2 175 1 82
2 176 1 84
2 177 1 84
2 178 1 84
2 179 1 85
2 180 1 85
2 181 1 87
2 182 1 87
2 183 1 90
2 184 1 90
2 185 1 98
2 186 1 98
2 187 1 105
2 188 1 105
2 189 1 107
2 190 1 107
2 191 1 108
2 192 1 108
2 193 1 116
2 194 1 116
0 17 5 2 1 11
0 18 5 1 1 14
0 19 5 1 1 16
0 20 5 1 1 59
0 21 5 1 1 101
0 22 5 1 1 124
0 23 5 1 1 126
0 24 5 1 1 128
0 25 5 1 1 130
0 26 5 1 1 132
0 27 5 1 1 134
0 28 7 1 2 125 135
0 29 5 3 1 28
0 30 7 1 2 22 27
0 31 5 3 1 30
0 32 7 2 2 138 141
0 33 5 1 1 144
0 34 7 1 2 12 33
0 35 5 1 1 34
0 36 7 1 2 136 145
0 37 5 1 1 36
0 38 7 1 2 35 37
3 594 5 0 1 38
0 40 7 1 2 13 142
0 41 5 1 1 40
0 42 7 1 2 139 41
0 43 5 3 1 42
0 44 7 1 2 15 127
0 45 5 4 1 44
0 46 7 1 2 18 23
0 47 5 3 1 46
0 48 7 2 2 149 153
0 49 5 1 1 156
0 50 7 1 2 146 49
0 51 5 1 1 50
0 52 7 1 2 137 140
0 53 5 1 1 52
0 54 7 1 2 143 53
0 55 5 3 1 54
0 56 7 1 2 157 158
0 57 5 1 1 56
0 58 7 1 2 51 57
3 595 5 0 1 58
0 60 7 1 2 147 154
0 61 5 1 1 60
0 62 7 1 2 39 129
0 63 5 4 1 62
0 64 7 1 2 19 24
0 65 5 3 1 64
0 66 7 1 2 161 165
0 67 5 1 1 66
0 68 7 1 2 150 67
0 69 7 1 2 61 68
0 70 5 1 1 69
0 71 7 1 2 151 159
0 72 5 1 1 71
0 73 7 3 2 155 166
0 74 5 1 1 168
0 75 7 1 2 162 169
0 76 7 1 2 72 75
0 77 5 1 1 76
3 596 7 0 2 70 77
0 79 7 1 2 148 170
0 80 5 2 1 79
0 81 7 1 2 78 131
0 82 5 3 1 81
0 83 7 1 2 20 25
0 84 5 3 1 83
0 85 7 2 2 173 176
0 86 5 1 1 179
0 87 7 2 2 152 163
0 88 5 1 1 181
0 89 7 1 2 167 88
0 90 5 2 1 89
0 91 7 1 2 86 183
0 92 7 1 2 171 91
0 93 5 1 1 92
0 94 7 1 2 164 74
0 95 5 1 1 94
0 96 7 1 2 160 182
0 97 5 1 1 96
0 98 7 2 2 95 97
0 99 7 1 2 180 185
0 100 5 1 1 99
3 597 7 0 2 93 100
0 102 7 1 2 177 186
0 103 5 1 1 102
0 104 7 1 2 121 133
0 105 5 2 1 104
0 106 7 1 2 21 26
0 107 5 2 1 106
0 108 7 2 2 187 189
0 109 5 1 1 191
0 110 7 1 2 174 192
0 111 7 1 2 103 110
0 112 5 1 1 111
0 113 7 1 2 175 184
0 114 7 1 2 172 113
0 115 5 1 1 114
0 116 7 2 2 178 115
0 117 5 1 1 193
0 118 7 1 2 109 194
0 119 5 1 1 118
0 120 7 1 2 112 119
3 598 5 0 1 120
0 122 7 1 2 188 117
0 123 5 1 1 122
3 599 7 0 2 190 123
