1 0 0 3 0
2 25 1 0
2 26 1 0
2 715 1 0
1 1 0 4 0
2 716 1 1
2 717 1 1
2 718 1 1
2 719 1 1
1 2 0 9 0
2 720 1 2
2 721 1 2
2 722 1 2
2 723 1 2
2 724 1 2
2 725 1 2
2 726 1 2
2 727 1 2
2 728 1 2
1 3 0 7 0
2 729 1 3
2 730 1 3
2 731 1 3
2 732 1 3
2 733 1 3
2 734 1 3
2 735 1 3
1 4 0 7 0
2 736 1 4
2 737 1 4
2 738 1 4
2 739 1 4
2 740 1 4
2 741 1 4
2 742 1 4
1 5 0 9 0
2 743 1 5
2 744 1 5
2 745 1 5
2 746 1 5
2 747 1 5
2 748 1 5
2 749 1 5
2 750 1 5
2 751 1 5
1 6 0 9 0
2 752 1 6
2 753 1 6
2 754 1 6
2 755 1 6
2 756 1 6
2 757 1 6
2 758 1 6
2 759 1 6
2 760 1 6
1 7 0 6 0
2 761 1 7
2 762 1 7
2 763 1 7
2 764 1 7
2 765 1 7
2 766 1 7
1 8 0 2 0
2 767 1 8
2 768 1 8
1 9 0 2 0
2 769 1 9
2 770 1 9
1 10 0 7 0
2 771 1 10
2 772 1 10
2 773 1 10
2 774 1 10
2 775 1 10
2 776 1 10
2 777 1 10
1 11 0 2 0
2 778 1 11
2 779 1 11
1 12 0 2 0
2 780 1 12
2 781 1 12
1 13 0 2 0
2 782 1 13
2 783 1 13
1 14 0 3 0
2 784 1 14
2 785 1 14
2 786 1 14
1 15 0 2 0
2 787 1 15
2 788 1 15
1 16 0 2 0
2 789 1 16
2 790 1 16
1 17 0 3 0
2 791 1 17
2 792 1 17
2 793 1 17
1 18 0 2 0
2 794 1 18
2 795 1 18
1 19 0 2 0
2 796 1 19
2 797 1 19
1 20 0 2 0
2 798 1 20
2 799 1 20
1 21 0 2 0
2 800 1 21
2 801 1 21
1 22 0 3 0
2 802 1 22
2 803 1 22
2 804 1 22
1 23 0 2 0
2 805 1 23
2 806 1 23
1 24 0 5 0
2 807 1 24
2 808 1 24
2 809 1 24
2 810 1 24
2 811 1 24
2 812 1 27
2 813 1 27
2 814 1 28
2 815 1 28
2 816 1 28
2 817 1 28
2 818 1 29
2 819 1 29
2 820 1 29
2 821 1 29
2 822 1 29
2 823 1 29
2 824 1 29
2 825 1 29
2 826 1 30
2 827 1 30
2 828 1 30
2 829 1 30
2 830 1 30
2 831 1 30
2 832 1 31
2 833 1 31
2 834 1 31
2 835 1 31
2 836 1 31
2 837 1 31
2 838 1 32
2 839 1 32
2 840 1 32
2 841 1 32
2 842 1 32
2 843 1 32
2 844 1 32
2 845 1 32
2 846 1 33
2 847 1 33
2 848 1 33
2 849 1 33
2 850 1 33
2 851 1 33
2 852 1 33
2 853 1 33
2 854 1 34
2 855 1 34
2 856 1 34
2 857 1 34
2 858 1 34
2 859 1 34
2 860 1 36
2 861 1 36
2 862 1 37
2 863 1 37
2 864 1 41
2 865 1 41
2 866 1 45
2 867 1 45
2 868 1 45
2 869 1 45
2 870 1 49
2 871 1 49
2 872 1 51
2 873 1 51
2 874 1 51
2 875 1 51
2 876 1 52
2 877 1 52
2 878 1 52
2 879 1 52
2 880 1 52
2 881 1 53
2 882 1 53
2 883 1 54
2 884 1 54
2 885 1 54
2 886 1 54
2 887 1 55
2 888 1 55
2 889 1 56
2 890 1 56
2 891 1 56
2 892 1 57
2 893 1 57
2 894 1 57
2 895 1 57
2 896 1 58
2 897 1 58
2 898 1 58
2 899 1 59
2 900 1 59
2 901 1 59
2 902 1 59
2 903 1 60
2 904 1 60
2 905 1 60
2 906 1 61
2 907 1 61
2 908 1 61
2 909 1 62
2 910 1 62
2 911 1 62
2 912 1 63
2 913 1 63
2 914 1 64
2 915 1 64
2 916 1 64
2 917 1 65
2 918 1 65
2 919 1 66
2 920 1 66
2 921 1 66
2 922 1 66
2 923 1 66
2 924 1 66
2 925 1 67
2 926 1 67
2 927 1 67
2 928 1 68
2 929 1 68
2 930 1 68
2 931 1 68
2 932 1 69
2 933 1 69
2 934 1 69
2 935 1 70
2 936 1 70
2 937 1 71
2 938 1 71
2 939 1 71
2 940 1 72
2 941 1 72
2 942 1 74
2 943 1 74
2 944 1 75
2 945 1 75
2 946 1 76
2 947 1 76
2 948 1 77
2 949 1 77
2 950 1 78
2 951 1 78
2 952 1 81
2 953 1 81
2 954 1 88
2 955 1 88
2 956 1 89
2 957 1 89
2 958 1 90
2 959 1 90
2 960 1 90
2 961 1 90
2 962 1 90
2 963 1 91
2 964 1 91
2 965 1 91
2 966 1 91
2 967 1 92
2 968 1 92
2 969 1 92
2 970 1 92
2 971 1 92
2 972 1 93
2 973 1 93
2 974 1 93
2 975 1 94
2 976 1 94
2 977 1 94
2 978 1 94
2 979 1 95
2 980 1 95
2 981 1 104
2 982 1 104
2 983 1 105
2 984 1 105
2 985 1 106
2 986 1 106
2 987 1 111
2 988 1 111
2 989 1 119
2 990 1 119
2 991 1 120
2 992 1 120
2 993 1 120
2 994 1 120
2 995 1 120
2 996 1 120
2 997 1 120
2 998 1 124
2 999 1 124
2 1000 1 125
2 1001 1 125
2 1002 1 134
2 1003 1 134
2 1004 1 140
2 1005 1 140
2 1006 1 141
2 1007 1 141
2 1008 1 141
2 1009 1 142
2 1010 1 142
2 1011 1 143
2 1012 1 143
2 1013 1 146
2 1014 1 146
2 1015 1 147
2 1016 1 147
2 1017 1 150
2 1018 1 150
2 1019 1 150
2 1020 1 150
2 1021 1 150
2 1022 1 150
2 1023 1 150
2 1024 1 150
2 1025 1 150
2 1026 1 150
2 1027 1 151
2 1028 1 151
2 1029 1 151
2 1030 1 151
2 1031 1 152
2 1032 1 152
2 1033 1 152
2 1034 1 152
2 1035 1 152
2 1036 1 154
2 1037 1 154
2 1038 1 157
2 1039 1 157
2 1040 1 157
2 1041 1 157
2 1042 1 157
2 1043 1 157
2 1044 1 157
2 1045 1 157
2 1046 1 157
2 1047 1 157
2 1048 1 158
2 1049 1 158
2 1050 1 159
2 1051 1 159
2 1052 1 159
2 1053 1 160
2 1054 1 160
2 1055 1 167
2 1056 1 167
2 1057 1 167
2 1058 1 167
2 1059 1 167
2 1060 1 167
2 1061 1 167
2 1062 1 172
2 1063 1 172
2 1064 1 172
2 1065 1 172
2 1066 1 177
2 1067 1 177
2 1068 1 177
2 1069 1 178
2 1070 1 178
2 1071 1 183
2 1072 1 183
2 1073 1 184
2 1074 1 184
2 1075 1 184
2 1076 1 186
2 1077 1 186
2 1078 1 189
2 1079 1 189
2 1080 1 194
2 1081 1 194
2 1082 1 194
2 1083 1 194
2 1084 1 204
2 1085 1 204
2 1086 1 206
2 1087 1 206
2 1088 1 207
2 1089 1 207
2 1090 1 207
2 1091 1 208
2 1092 1 208
2 1093 1 216
2 1094 1 216
2 1095 1 218
2 1096 1 218
2 1097 1 221
2 1098 1 221
2 1099 1 232
2 1100 1 232
2 1101 1 233
2 1102 1 233
2 1103 1 234
2 1104 1 234
2 1105 1 243
2 1106 1 243
2 1107 1 255
2 1108 1 255
2 1109 1 258
2 1110 1 258
2 1111 1 262
2 1112 1 262
2 1113 1 262
2 1114 1 270
2 1115 1 270
2 1116 1 270
2 1117 1 270
2 1118 1 270
2 1119 1 270
2 1120 1 277
2 1121 1 277
2 1122 1 279
2 1123 1 279
2 1124 1 300
2 1125 1 300
2 1126 1 304
2 1127 1 304
2 1128 1 304
2 1129 1 305
2 1130 1 305
2 1131 1 309
2 1132 1 309
2 1133 1 327
2 1134 1 327
2 1135 1 327
2 1136 1 330
2 1137 1 330
2 1138 1 330
2 1139 1 330
2 1140 1 334
2 1141 1 334
2 1142 1 334
2 1143 1 334
2 1144 1 362
2 1145 1 362
2 1146 1 374
2 1147 1 374
2 1148 1 374
2 1149 1 374
2 1150 1 375
2 1151 1 375
2 1152 1 375
2 1153 1 376
2 1154 1 376
2 1155 1 376
2 1156 1 376
2 1157 1 376
2 1158 1 376
2 1159 1 376
2 1160 1 377
2 1161 1 377
2 1162 1 377
2 1163 1 381
2 1164 1 381
2 1165 1 381
2 1166 1 381
2 1167 1 381
2 1168 1 427
2 1169 1 427
2 1170 1 427
2 1171 1 453
2 1172 1 453
2 1173 1 453
2 1174 1 453
2 1175 1 456
2 1176 1 456
2 1177 1 458
2 1178 1 458
2 1179 1 466
2 1180 1 466
2 1181 1 467
2 1182 1 467
2 1183 1 468
2 1184 1 468
2 1185 1 469
2 1186 1 469
2 1187 1 477
2 1188 1 477
2 1189 1 477
2 1190 1 477
2 1191 1 477
2 1192 1 477
2 1193 1 479
2 1194 1 479
2 1195 1 483
2 1196 1 483
2 1197 1 483
2 1198 1 483
2 1199 1 485
2 1200 1 485
2 1201 1 485
2 1202 1 485
2 1203 1 485
2 1204 1 500
2 1205 1 500
2 1206 1 500
2 1207 1 500
2 1208 1 507
2 1209 1 507
2 1210 1 509
2 1211 1 509
2 1212 1 515
2 1213 1 515
2 1214 1 519
2 1215 1 519
2 1216 1 534
2 1217 1 534
2 1218 1 534
2 1219 1 534
2 1220 1 537
2 1221 1 537
2 1222 1 537
2 1223 1 542
2 1224 1 542
2 1225 1 545
2 1226 1 545
2 1227 1 545
2 1228 1 548
2 1229 1 548
2 1230 1 549
2 1231 1 549
2 1232 1 550
2 1233 1 550
2 1234 1 552
2 1235 1 552
2 1236 1 561
2 1237 1 561
2 1238 1 623
2 1239 1 623
2 1240 1 623
2 1241 1 624
2 1242 1 624
2 1243 1 628
2 1244 1 628
2 1245 1 629
2 1246 1 629
2 1247 1 631
2 1248 1 631
2 1249 1 656
2 1250 1 656
2 1251 1 661
2 1252 1 661
0 27 5 2 1 25
0 28 5 4 1 716
0 29 5 8 1 720
0 30 5 6 1 729
0 31 5 6 1 736
0 32 5 8 1 743
0 33 5 8 1 752
0 34 5 6 1 761
0 35 5 1 1 767
0 36 5 2 1 769
0 37 5 2 1 771
0 38 5 1 1 778
0 39 5 1 1 780
0 40 5 1 1 782
0 41 5 2 1 784
0 42 5 1 1 787
0 43 5 1 1 789
0 44 5 1 1 791
0 45 5 4 1 794
0 46 5 1 1 796
0 47 5 1 1 798
0 48 5 1 1 800
0 49 5 2 1 802
0 50 5 1 1 805
0 51 5 4 1 807
0 52 7 5 2 781 47
0 53 5 2 1 876
0 54 7 4 2 39 799
0 55 5 2 1 883
0 56 7 3 2 881 887
0 57 7 4 2 783 48
0 58 5 3 1 892
0 59 7 4 2 40 801
0 60 5 3 1 899
0 61 7 3 2 896 903
0 62 7 3 2 785 870
0 63 5 2 1 909
0 64 7 3 2 864 803
0 65 5 2 1 914
0 66 7 6 2 912 917
0 67 7 3 2 770 44
0 68 5 4 1 925
0 69 7 3 2 860 792
0 70 5 2 1 932
0 71 7 3 2 768 43
0 72 5 2 1 937
0 73 7 1 2 26 938
0 74 5 2 1 73
0 75 7 2 2 35 790
0 76 5 2 1 944
0 77 7 2 2 812 945
0 78 5 2 1 948
0 79 7 1 2 717 950
0 80 5 1 1 79
0 81 7 2 2 942 80
0 82 7 1 2 933 952
0 83 5 1 1 82
0 84 7 1 2 814 949
0 85 5 1 1 84
0 86 7 1 2 83 85
0 87 5 1 1 86
0 88 7 2 2 928 87
0 89 5 2 1 954
0 90 7 5 2 772 866
0 91 5 4 1 958
0 92 7 5 2 862 795
0 93 5 3 1 967
0 94 7 4 2 963 972
0 95 5 2 1 975
0 96 7 1 2 721 979
0 97 5 1 1 96
0 98 7 1 2 818 964
0 99 5 1 1 98
0 100 7 1 2 730 99
0 101 7 1 2 97 100
0 102 7 1 2 956 101
0 103 5 1 1 102
0 104 7 2 2 718 926
0 105 5 2 1 981
0 106 7 2 2 946 982
0 107 5 1 1 985
0 108 7 1 2 927 939
0 109 5 1 1 108
0 110 7 1 2 719 935
0 111 5 2 1 110
0 112 7 1 2 109 987
0 113 5 1 1 112
0 114 7 1 2 929 940
0 115 5 1 1 114
0 116 7 1 2 715 115
0 117 7 1 2 113 116
0 118 5 1 1 117
0 119 7 2 2 107 118
0 120 5 7 1 989
0 121 7 1 2 965 990
0 122 5 1 1 121
0 123 7 1 2 813 941
0 124 5 2 1 123
0 125 7 2 2 986 998
0 126 7 1 2 959 1000
0 127 5 1 1 126
0 128 7 1 2 819 980
0 129 5 1 1 128
0 130 7 1 2 731 129
0 131 7 1 2 127 130
0 132 7 1 2 122 131
0 133 5 1 1 132
0 134 7 2 2 826 960
0 135 5 1 1 1002
0 136 7 1 2 722 1003
0 137 7 1 2 991 136
0 138 5 1 1 137
0 139 7 1 2 133 138
0 140 7 2 2 103 139
0 141 5 3 1 1004
0 142 7 2 2 42 806
0 143 5 2 1 1009
0 144 7 1 2 872 1011
0 145 5 1 1 144
0 146 7 2 2 788 50
0 147 5 2 1 1013
0 148 7 1 2 808 1015
0 149 5 1 1 148
0 150 7 10 2 145 149
0 151 7 4 2 737 744
0 152 7 5 2 753 854
0 153 5 1 1 1031
0 154 7 2 2 1027 1032
0 155 7 1 2 1017 1036
0 156 5 1 1 155
0 157 7 10 2 1012 1016
0 158 7 2 2 754 762
0 159 7 3 2 809 1048
0 160 7 2 2 1028 1050
0 161 7 1 2 1038 1053
0 162 5 1 1 161
0 163 7 1 2 156 162
0 164 5 1 1 163
0 165 7 1 2 1006 164
0 166 5 1 1 165
0 167 7 7 2 846 763
0 168 5 1 1 1055
0 169 7 1 2 1018 1056
0 170 5 1 1 169
0 171 7 1 2 847 855
0 172 7 4 2 873 171
0 173 7 1 2 1039 1062
0 174 5 1 1 173
0 175 7 1 2 170 174
0 176 5 1 1 175
0 177 7 3 2 832 838
0 178 7 2 2 820 968
0 179 5 1 1 1069
0 180 7 1 2 827 1070
0 181 7 1 2 957 180
0 182 5 1 1 181
0 183 7 2 2 947 999
0 184 5 3 1 1071
0 185 7 1 2 821 976
0 186 5 2 1 185
0 187 7 1 2 723 969
0 188 5 1 1 187
0 189 7 2 2 1076 188
0 190 5 1 1 1078
0 191 7 1 2 815 930
0 192 5 1 1 191
0 193 7 1 2 936 192
0 194 5 4 1 193
0 195 7 1 2 977 1080
0 196 5 1 1 195
0 197 7 1 2 1079 196
0 198 5 1 1 197
0 199 7 1 2 1073 198
0 200 5 1 1 199
0 201 7 1 2 983 190
0 202 5 1 1 201
0 203 7 1 2 724 773
0 204 7 2 2 867 203
0 205 5 1 1 1084
0 206 7 2 2 973 205
0 207 7 3 2 816 934
0 208 5 2 1 1088
0 209 7 1 2 1086 1089
0 210 5 1 1 209
0 211 7 1 2 202 210
0 212 7 1 2 200 211
0 213 5 1 1 212
0 214 7 1 2 828 213
0 215 5 1 1 214
0 216 7 2 2 732 970
0 217 5 1 1 1093
0 218 7 2 2 822 1090
0 219 5 1 1 1095
0 220 7 1 2 823 1074
0 221 7 2 2 1081 220
0 222 5 1 1 1097
0 223 7 1 2 219 222
0 224 5 1 1 223
0 225 7 1 2 1094 224
0 226 5 1 1 225
0 227 7 1 2 829 774
0 228 7 1 2 1098 227
0 229 5 1 1 228
0 230 7 1 2 226 229
0 231 7 1 2 215 230
0 232 7 2 2 182 231
0 233 5 2 1 1099
0 234 7 2 2 1066 1101
0 235 7 1 2 176 1103
0 236 5 1 1 235
0 237 7 1 2 166 236
0 238 5 1 1 237
0 239 7 1 2 919 238
0 240 5 1 1 239
0 241 7 1 2 755 1104
0 242 5 1 1 241
0 243 7 2 2 848 1029
0 244 7 1 2 1007 1105
0 245 5 1 1 244
0 246 7 1 2 242 245
0 247 5 1 1 246
0 248 7 1 2 764 865
0 249 7 1 2 804 248
0 250 5 1 1 249
0 251 7 1 2 856 786
0 252 7 1 2 871 251
0 253 5 1 1 252
0 254 7 1 2 250 253
0 255 5 2 1 254
0 256 7 1 2 1019 1107
0 257 5 1 1 256
0 258 7 2 2 765 810
0 259 5 1 1 1109
0 260 7 1 2 918 259
0 261 5 1 1 260
0 262 7 3 2 857 874
0 263 5 1 1 1111
0 264 7 1 2 913 263
0 265 5 1 1 264
0 266 7 1 2 1040 265
0 267 7 1 2 261 266
0 268 5 1 1 267
0 269 7 1 2 257 268
0 270 5 6 1 269
0 271 7 1 2 247 1114
0 272 5 1 1 271
0 273 7 1 2 240 272
0 274 5 1 1 273
0 275 7 1 2 906 274
0 276 5 1 1 275
0 277 7 2 2 893 1051
0 278 5 1 1 1120
0 279 7 2 2 900 1063
0 280 5 1 1 1122
0 281 7 1 2 278 280
0 282 5 1 1 281
0 283 7 1 2 1041 282
0 284 5 1 1 283
0 285 7 1 2 904 153
0 286 5 1 1 285
0 287 7 1 2 897 168
0 288 5 1 1 287
0 289 7 1 2 286 288
0 290 7 1 2 1020 289
0 291 5 1 1 290
0 292 7 1 2 284 291
0 293 5 1 1 292
0 294 7 1 2 920 293
0 295 5 1 1 294
0 296 7 1 2 849 898
0 297 5 1 1 296
0 298 7 1 2 756 905
0 299 5 1 1 298
0 300 7 2 2 297 299
0 301 7 1 2 1115 1124
0 302 5 1 1 301
0 303 7 1 2 295 302
0 304 5 3 1 303
0 305 7 2 2 833 745
0 306 5 1 1 1129
0 307 7 1 2 1102 1130
0 308 5 1 1 307
0 309 7 2 2 738 839
0 310 5 1 1 1131
0 311 7 1 2 1008 1132
0 312 5 1 1 311
0 313 7 1 2 308 312
0 314 5 1 1 313
0 315 7 1 2 1126 314
0 316 5 1 1 315
0 317 7 1 2 276 316
0 318 5 1 1 317
0 319 7 1 2 889 318
0 320 5 1 1 319
0 321 7 1 2 739 1100
0 322 5 1 1 321
0 323 7 1 2 840 882
0 324 5 1 1 323
0 325 7 1 2 746 888
0 326 5 1 1 325
0 327 7 3 2 324 326
0 328 7 1 2 1127 1133
0 329 5 1 1 328
0 330 7 4 2 841 884
0 331 5 1 1 1136
0 332 7 1 2 1064 1137
0 333 5 1 1 332
0 334 7 4 2 747 877
0 335 5 1 1 1140
0 336 7 1 2 1052 1141
0 337 5 1 1 336
0 338 7 1 2 333 337
0 339 5 1 1 338
0 340 7 1 2 1042 339
0 341 5 1 1 340
0 342 7 1 2 1057 1138
0 343 5 1 1 342
0 344 7 1 2 1033 1142
0 345 5 1 1 344
0 346 7 1 2 343 345
0 347 5 1 1 346
0 348 7 1 2 1021 347
0 349 5 1 1 348
0 350 7 1 2 341 349
0 351 5 1 1 350
0 352 7 1 2 921 351
0 353 5 1 1 352
0 354 7 1 2 757 331
0 355 5 1 1 354
0 356 7 1 2 850 335
0 357 5 1 1 356
0 358 7 1 2 355 357
0 359 7 1 2 1116 358
0 360 5 1 1 359
0 361 7 1 2 353 360
0 362 5 2 1 361
0 363 7 1 2 907 1144
0 364 5 1 1 363
0 365 7 1 2 329 364
0 366 5 1 1 365
0 367 7 1 2 834 1005
0 368 5 1 1 367
0 369 7 1 2 366 368
0 370 7 1 2 322 369
0 371 5 1 1 370
0 372 7 1 2 320 371
0 373 5 1 1 372
0 374 7 4 2 38 797
0 375 5 3 1 1146
0 376 7 7 2 779 46
0 377 5 3 1 1153
0 378 7 1 2 1150 1160
0 379 7 1 2 373 378
0 380 5 1 1 379
0 381 7 5 2 1067 1147
0 382 7 1 2 1065 1163
0 383 5 1 1 382
0 384 7 1 2 1054 1154
0 385 5 1 1 384
0 386 7 1 2 383 385
0 387 5 1 1 386
0 388 7 1 2 1043 387
0 389 5 1 1 388
0 390 7 1 2 1058 1164
0 391 5 1 1 390
0 392 7 1 2 1037 1155
0 393 5 1 1 392
0 394 7 1 2 391 393
0 395 5 1 1 394
0 396 7 1 2 1022 395
0 397 5 1 1 396
0 398 7 1 2 389 397
0 399 5 1 1 398
0 400 7 1 2 824 955
0 401 5 1 1 400
0 402 7 1 2 135 217
0 403 5 1 1 402
0 404 7 1 2 725 1001
0 405 5 1 1 404
0 406 7 1 2 403 405
0 407 7 1 2 401 406
0 408 5 1 1 407
0 409 7 1 2 1082 1087
0 410 5 1 1 409
0 411 7 1 2 1077 410
0 412 5 1 1 411
0 413 7 1 2 1075 412
0 414 5 1 1 413
0 415 7 1 2 775 1096
0 416 5 1 1 415
0 417 7 1 2 726 1091
0 418 5 1 1 417
0 419 7 1 2 978 984
0 420 7 1 2 418 419
0 421 5 1 1 420
0 422 7 1 2 416 421
0 423 7 1 2 414 422
0 424 5 1 1 423
0 425 7 1 2 733 424
0 426 5 1 1 425
0 427 7 3 2 727 974
0 428 5 1 1 1168
0 429 7 1 2 951 1169
0 430 5 1 1 429
0 431 7 1 2 988 430
0 432 5 1 1 431
0 433 7 1 2 817 861
0 434 7 1 2 793 433
0 435 5 1 1 434
0 436 7 1 2 1170 435
0 437 5 1 1 436
0 438 7 1 2 943 437
0 439 5 1 1 438
0 440 7 1 2 432 439
0 441 5 1 1 440
0 442 7 1 2 931 441
0 443 5 1 1 442
0 444 7 1 2 953 428
0 445 5 1 1 444
0 446 7 1 2 830 966
0 447 7 1 2 179 446
0 448 7 1 2 445 447
0 449 7 1 2 443 448
0 450 5 1 1 449
0 451 7 1 2 426 450
0 452 7 1 2 408 451
0 453 5 4 1 452
0 454 7 1 2 399 1171
0 455 5 1 1 454
0 456 7 2 2 811 992
0 457 7 1 2 748 758
0 458 7 2 2 1175 457
0 459 7 1 2 734 766
0 460 7 1 2 1085 459
0 461 7 1 2 1177 460
0 462 5 1 1 461
0 463 7 1 2 1072 1092
0 464 5 1 1 463
0 465 7 1 2 971 1083
0 466 7 2 2 464 465
0 467 7 2 2 1112 1179
0 468 7 2 2 825 831
0 469 7 2 2 851 1183
0 470 7 1 2 842 1185
0 471 7 1 2 1181 470
0 472 5 1 1 471
0 473 7 1 2 462 472
0 474 5 1 1 473
0 475 7 1 2 1044 474
0 476 5 1 1 475
0 477 7 6 2 1180 1184
0 478 5 1 1 1187
0 479 7 2 2 843 1188
0 480 5 1 1 1193
0 481 7 1 2 1059 1194
0 482 5 1 1 481
0 483 7 4 2 728 735
0 484 7 1 2 961 1195
0 485 7 5 2 993 484
0 486 5 1 1 1199
0 487 7 1 2 749 1034
0 488 7 1 2 1200 487
0 489 5 1 1 488
0 490 7 1 2 482 489
0 491 5 1 1 490
0 492 7 1 2 1023 491
0 493 5 1 1 492
0 494 7 1 2 476 493
0 495 5 1 1 494
0 496 7 1 2 835 1161
0 497 5 1 1 496
0 498 7 1 2 740 1151
0 499 5 1 1 498
0 500 7 4 2 497 499
0 501 7 1 2 495 1204
0 502 5 1 1 501
0 503 7 1 2 455 502
0 504 5 1 1 503
0 505 7 1 2 922 504
0 506 5 1 1 505
0 507 7 2 2 1106 1156
0 508 5 1 1 1208
0 509 7 2 2 759 1165
0 510 5 1 1 1210
0 511 7 1 2 508 510
0 512 5 1 1 511
0 513 7 1 2 1172 512
0 514 5 1 1 513
0 515 7 2 2 852 1201
0 516 5 1 1 1212
0 517 7 1 2 480 516
0 518 5 1 1 517
0 519 7 2 2 844 853
0 520 5 1 1 1214
0 521 7 1 2 1205 520
0 522 7 1 2 518 521
0 523 5 1 1 522
0 524 7 1 2 514 523
0 525 5 1 1 524
0 526 7 1 2 1117 525
0 527 5 1 1 526
0 528 7 1 2 506 527
0 529 5 1 1 528
0 530 7 1 2 890 529
0 531 5 1 1 530
0 532 7 1 2 1173 1206
0 533 5 1 1 532
0 534 7 4 2 741 1157
0 535 7 1 2 1189 1216
0 536 5 1 1 535
0 537 7 3 2 836 1148
0 538 7 1 2 1202 1220
0 539 5 1 1 538
0 540 7 1 2 536 539
0 541 7 1 2 533 540
0 542 5 2 1 541
0 543 7 1 2 1145 1223
0 544 5 1 1 543
0 545 7 3 2 1190 1221
0 546 7 1 2 1060 1225
0 547 5 1 1 546
0 548 7 2 2 962 1158
0 549 7 2 2 994 1228
0 550 7 2 2 742 1196
0 551 7 1 2 1035 1232
0 552 7 2 2 1230 551
0 553 5 1 1 1234
0 554 7 1 2 547 553
0 555 5 1 1 554
0 556 7 1 2 1024 555
0 557 5 1 1 556
0 558 7 1 2 1186 1222
0 559 7 1 2 1182 558
0 560 5 1 1 559
0 561 7 2 2 776 1197
0 562 7 1 2 868 1049
0 563 7 1 2 1217 562
0 564 7 1 2 1236 563
0 565 7 1 2 1176 564
0 566 5 1 1 565
0 567 7 1 2 560 566
0 568 5 1 1 567
0 569 7 1 2 1045 568
0 570 5 1 1 569
0 571 7 1 2 557 570
0 572 5 1 1 571
0 573 7 1 2 923 572
0 574 5 1 1 573
0 575 7 1 2 1213 1218
0 576 5 1 1 575
0 577 7 1 2 760 1226
0 578 5 1 1 577
0 579 7 1 2 576 578
0 580 5 1 1 579
0 581 7 1 2 1118 580
0 582 5 1 1 581
0 583 7 1 2 574 582
0 584 5 1 1 583
0 585 7 1 2 1134 584
0 586 5 1 1 585
0 587 7 1 2 544 586
0 588 7 1 2 531 587
0 589 5 1 1 588
0 590 7 1 2 908 589
0 591 5 1 1 590
0 592 7 1 2 306 1162
0 593 5 1 1 592
0 594 7 1 2 310 1152
0 595 5 1 1 594
0 596 7 1 2 593 595
0 597 7 1 2 1174 596
0 598 5 1 1 597
0 599 7 1 2 845 486
0 600 5 1 1 599
0 601 7 1 2 750 478
0 602 5 1 1 601
0 603 7 1 2 1207 602
0 604 7 1 2 600 603
0 605 5 1 1 604
0 606 7 1 2 598 605
0 607 5 1 1 606
0 608 7 1 2 891 607
0 609 5 1 1 608
0 610 7 1 2 1135 1224
0 611 5 1 1 610
0 612 7 1 2 1143 1227
0 613 5 1 1 612
0 614 7 1 2 1139 1219
0 615 7 1 2 1203 614
0 616 5 1 1 615
0 617 7 1 2 613 616
0 618 7 1 2 611 617
0 619 7 1 2 609 618
0 620 5 1 1 619
0 621 7 1 2 1128 620
0 622 5 1 1 621
0 623 7 3 2 885 1191
0 624 7 2 2 1166 1238
0 625 5 1 1 1241
0 626 7 1 2 1113 1242
0 627 5 1 1 626
0 628 7 2 2 869 878
0 629 7 2 2 1030 1198
0 630 7 1 2 1159 1245
0 631 7 2 2 1243 630
0 632 7 1 2 777 1110
0 633 7 1 2 1247 632
0 634 7 1 2 995 633
0 635 5 1 1 634
0 636 7 1 2 627 635
0 637 5 1 1 636
0 638 7 1 2 1046 637
0 639 5 1 1 638
0 640 7 1 2 858 1248
0 641 7 1 2 996 640
0 642 5 1 1 641
0 643 7 1 2 625 642
0 644 5 1 1 643
0 645 7 1 2 859 863
0 646 5 1 1 645
0 647 7 1 2 1025 646
0 648 7 1 2 644 647
0 649 5 1 1 648
0 650 7 1 2 639 649
0 651 5 1 1 650
0 652 7 1 2 924 1125
0 653 7 1 2 651 652
0 654 5 1 1 653
0 655 7 1 2 901 1149
0 656 7 2 2 1239 655
0 657 7 1 2 837 875
0 658 7 1 2 1215 657
0 659 7 1 2 1249 658
0 660 5 1 1 659
0 661 7 2 2 879 894
0 662 7 1 2 1233 1229
0 663 7 1 2 1251 662
0 664 7 1 2 1178 663
0 665 5 1 1 664
0 666 7 1 2 660 665
0 667 5 1 1 666
0 668 7 1 2 1047 1108
0 669 7 1 2 667 668
0 670 5 1 1 669
0 671 7 1 2 910 1061
0 672 7 1 2 1068 671
0 673 7 1 2 1250 672
0 674 5 1 1 673
0 675 7 1 2 751 915
0 676 7 1 2 1252 675
0 677 7 1 2 1235 676
0 678 5 1 1 677
0 679 7 1 2 674 678
0 680 5 1 1 679
0 681 7 1 2 1026 680
0 682 5 1 1 681
0 683 7 1 2 895 1211
0 684 7 1 2 1240 683
0 685 5 1 1 684
0 686 7 1 2 902 1237
0 687 7 1 2 1244 686
0 688 7 1 2 1209 687
0 689 7 1 2 997 688
0 690 5 1 1 689
0 691 7 1 2 685 690
0 692 5 1 1 691
0 693 7 1 2 1119 692
0 694 5 1 1 693
0 695 7 1 2 880 911
0 696 7 1 2 1010 695
0 697 7 1 2 1246 696
0 698 7 1 2 1121 697
0 699 7 1 2 1231 698
0 700 5 1 1 699
0 701 7 1 2 886 916
0 702 7 1 2 1014 701
0 703 7 1 2 1167 702
0 704 7 1 2 1123 703
0 705 7 1 2 1192 704
0 706 5 1 1 705
0 707 7 1 2 700 706
0 708 7 1 2 694 707
0 709 7 1 2 682 708
0 710 7 1 2 670 709
0 711 7 1 2 654 710
0 712 7 1 2 622 711
0 713 7 1 2 591 712
0 714 7 1 2 380 713
3 1999 5 0 1 714
