1 0 0 2 0
2 64 1 0
2 65 1 0
1 1 0 2 0
2 66 1 1
2 67 1 1
1 2 0 2 0
2 68 1 2
2 69 1 2
1 3 0 2 0
2 70 1 3
2 71 1 3
1 4 0 2 0
2 72 1 4
2 73 1 4
1 5 0 2 0
2 74 1 5
2 75 1 5
1 6 0 2 0
2 76 1 6
2 77 1 6
1 7 0 2 0
2 78 1 7
2 79 1 7
1 8 0 2 0
2 80 1 8
2 81 1 8
1 9 0 2 0
2 82 1 9
2 83 1 9
1 10 0 2 0
2 84 1 10
2 85 1 10
1 11 0 2 0
2 86 1 11
2 87 1 11
1 12 0 2 0
2 88 1 12
2 89 1 12
1 13 0 2 0
2 90 1 13
2 91 1 13
1 14 0 2 0
2 92 1 14
2 93 1 14
1 15 0 2 0
2 94 1 15
2 95 1 15
1 16 0 2 0
2 96 1 16
2 165 1 16
1 17 0 2 0
2 177 1 17
2 192 1 17
1 18 0 2 0
2 207 1 18
2 222 1 18
1 19 0 2 0
2 237 1 19
2 252 1 19
1 20 0 2 0
2 267 1 20
2 282 1 20
1 21 0 2 0
2 297 1 21
2 312 1 21
1 22 0 2 0
2 327 1 22
2 342 1 22
1 23 0 2 0
2 357 1 23
2 372 1 23
1 24 0 2 0
2 387 1 24
2 402 1 24
1 25 0 2 0
2 417 1 25
2 432 1 25
1 26 0 2 0
2 447 1 26
2 462 1 26
1 27 0 2 0
2 477 1 27
2 492 1 27
1 28 0 2 0
2 507 1 28
2 522 1 28
1 29 0 2 0
2 537 1 29
2 552 1 29
1 30 0 2 0
2 567 1 30
2 582 1 30
1 31 0 2 0
2 597 1 31
2 612 1 31
1 32 0 2 0
2 628 1 32
2 631 1 32
1 33 0 2 0
2 632 1 33
2 633 1 33
1 34 0 2 0
2 634 1 34
2 635 1 34
1 35 0 2 0
2 636 1 35
2 637 1 35
1 36 0 2 0
2 638 1 36
2 639 1 36
1 37 0 2 0
2 640 1 37
2 641 1 37
1 38 0 2 0
2 642 1 38
2 643 1 38
1 39 0 2 0
2 644 1 39
2 645 1 39
1 40 0 2 0
2 646 1 40
2 647 1 40
1 41 0 2 0
2 648 1 41
2 649 1 41
1 42 0 2 0
2 650 1 42
2 651 1 42
1 43 0 2 0
2 652 1 43
2 653 1 43
1 44 0 2 0
2 654 1 44
2 655 1 44
1 45 0 2 0
2 656 1 45
2 657 1 45
1 46 0 2 0
2 658 1 46
2 659 1 46
1 47 0 2 0
2 660 1 47
2 661 1 47
1 48 0 2 0
2 662 1 48
2 663 1 48
1 49 0 2 0
2 664 1 49
2 665 1 49
1 50 0 2 0
2 666 1 50
2 667 1 50
1 51 0 2 0
2 668 1 51
2 669 1 51
1 52 0 2 0
2 670 1 52
2 671 1 52
1 53 0 2 0
2 672 1 53
2 673 1 53
1 54 0 2 0
2 674 1 54
2 675 1 54
1 55 0 2 0
2 676 1 55
2 677 1 55
1 56 0 2 0
2 678 1 56
2 679 1 56
1 57 0 2 0
2 680 1 57
2 681 1 57
1 58 0 2 0
2 682 1 58
2 683 1 58
1 59 0 2 0
2 684 1 59
2 685 1 59
1 60 0 2 0
2 686 1 60
2 687 1 60
1 61 0 2 0
2 688 1 61
2 689 1 61
1 62 0 2 0
2 690 1 62
2 691 1 62
1 63 0 2 0
2 692 1 63
2 693 1 63
2 694 1 131
2 695 1 131
2 696 1 132
2 697 1 132
2 698 1 133
2 699 1 133
2 700 1 134
2 701 1 134
2 702 1 135
2 703 1 135
2 704 1 136
2 705 1 136
2 706 1 137
2 707 1 137
2 708 1 138
2 709 1 138
2 710 1 139
2 711 1 139
2 712 1 140
2 713 1 140
2 714 1 141
2 715 1 141
2 716 1 142
2 717 1 142
2 718 1 143
2 719 1 143
2 720 1 144
2 721 1 144
2 722 1 145
2 723 1 145
2 724 1 146
2 725 1 146
2 726 1 147
2 727 1 147
2 728 1 148
2 729 1 148
2 730 1 149
2 731 1 149
2 732 1 150
2 733 1 150
2 734 1 151
2 735 1 151
2 736 1 152
2 737 1 152
2 738 1 153
2 739 1 153
2 740 1 154
2 741 1 154
2 742 1 155
2 743 1 155
2 744 1 156
2 745 1 156
2 746 1 157
2 747 1 157
2 748 1 158
2 749 1 158
2 750 1 159
2 751 1 159
2 752 1 161
2 753 1 161
2 754 1 162
2 755 1 162
2 756 1 162
2 757 1 167
2 758 1 167
2 759 1 169
2 760 1 169
2 761 1 170
2 762 1 170
2 763 1 180
2 764 1 180
2 765 1 183
2 766 1 183
2 767 1 185
2 768 1 185
2 769 1 186
2 770 1 186
2 771 1 195
2 772 1 195
2 773 1 198
2 774 1 198
2 775 1 200
2 776 1 200
2 777 1 201
2 778 1 201
2 779 1 210
2 780 1 210
2 781 1 213
2 782 1 213
2 783 1 215
2 784 1 215
2 785 1 216
2 786 1 216
2 787 1 225
2 788 1 225
2 789 1 228
2 790 1 228
2 791 1 230
2 792 1 230
2 793 1 231
2 794 1 231
2 795 1 240
2 796 1 240
2 797 1 243
2 798 1 243
2 799 1 245
2 800 1 245
2 801 1 246
2 802 1 246
2 803 1 255
2 804 1 255
2 805 1 258
2 806 1 258
2 807 1 260
2 808 1 260
2 809 1 261
2 810 1 261
2 811 1 270
2 812 1 270
2 813 1 273
2 814 1 273
2 815 1 275
2 816 1 275
2 817 1 276
2 818 1 276
2 819 1 285
2 820 1 285
2 821 1 288
2 822 1 288
2 823 1 290
2 824 1 290
2 825 1 291
2 826 1 291
2 827 1 300
2 828 1 300
2 829 1 303
2 830 1 303
2 831 1 305
2 832 1 305
2 833 1 306
2 834 1 306
2 835 1 315
2 836 1 315
2 837 1 318
2 838 1 318
2 839 1 320
2 840 1 320
2 841 1 321
2 842 1 321
2 843 1 330
2 844 1 330
2 845 1 333
2 846 1 333
2 847 1 335
2 848 1 335
2 849 1 336
2 850 1 336
2 851 1 345
2 852 1 345
2 853 1 348
2 854 1 348
2 855 1 350
2 856 1 350
2 857 1 351
2 858 1 351
2 859 1 360
2 860 1 360
2 861 1 363
2 862 1 363
2 863 1 365
2 864 1 365
2 865 1 366
2 866 1 366
2 867 1 375
2 868 1 375
2 869 1 378
2 870 1 378
2 871 1 380
2 872 1 380
2 873 1 381
2 874 1 381
2 875 1 390
2 876 1 390
2 877 1 393
2 878 1 393
2 879 1 395
2 880 1 395
2 881 1 396
2 882 1 396
2 883 1 405
2 884 1 405
2 885 1 408
2 886 1 408
2 887 1 410
2 888 1 410
2 889 1 411
2 890 1 411
2 891 1 420
2 892 1 420
2 893 1 423
2 894 1 423
2 895 1 425
2 896 1 425
2 897 1 426
2 898 1 426
2 899 1 435
2 900 1 435
2 901 1 438
2 902 1 438
2 903 1 440
2 904 1 440
2 905 1 441
2 906 1 441
2 907 1 450
2 908 1 450
2 909 1 453
2 910 1 453
2 911 1 455
2 912 1 455
2 913 1 456
2 914 1 456
2 915 1 465
2 916 1 465
2 917 1 468
2 918 1 468
2 919 1 470
2 920 1 470
2 921 1 471
2 922 1 471
2 923 1 480
2 924 1 480
2 925 1 483
2 926 1 483
2 927 1 485
2 928 1 485
2 929 1 486
2 930 1 486
2 931 1 495
2 932 1 495
2 933 1 498
2 934 1 498
2 935 1 500
2 936 1 500
2 937 1 501
2 938 1 501
2 939 1 510
2 940 1 510
2 941 1 513
2 942 1 513
2 943 1 515
2 944 1 515
2 945 1 516
2 946 1 516
2 947 1 525
2 948 1 525
2 949 1 528
2 950 1 528
2 951 1 530
2 952 1 530
2 953 1 531
2 954 1 531
2 955 1 540
2 956 1 540
2 957 1 543
2 958 1 543
2 959 1 545
2 960 1 545
2 961 1 546
2 962 1 546
2 963 1 555
2 964 1 555
2 965 1 558
2 966 1 558
2 967 1 560
2 968 1 560
2 969 1 561
2 970 1 561
2 971 1 570
2 972 1 570
2 973 1 573
2 974 1 573
2 975 1 575
2 976 1 575
2 977 1 576
2 978 1 576
2 979 1 585
2 980 1 585
2 981 1 588
2 982 1 588
2 983 1 590
2 984 1 590
2 985 1 591
2 986 1 591
2 987 1 600
2 988 1 600
2 989 1 603
2 990 1 603
2 991 1 605
2 992 1 605
2 993 1 606
2 994 1 606
2 995 1 615
2 996 1 615
2 997 1 616
2 998 1 616
2 999 1 618
2 1000 1 618
2 1001 1 620
2 1002 1 620
2 1003 1 621
2 1004 1 621
0 97 5 1 1 64
0 98 5 1 1 66
0 99 5 1 1 68
0 100 5 1 1 70
0 101 5 1 1 72
0 102 5 1 1 74
0 103 5 1 1 76
0 104 5 1 1 78
0 105 5 1 1 80
0 106 5 1 1 82
0 107 5 1 1 84
0 108 5 1 1 86
0 109 5 1 1 88
0 110 5 1 1 90
0 111 5 1 1 92
0 112 5 1 1 94
0 113 5 1 1 96
0 114 5 1 1 177
0 115 5 1 1 207
0 116 5 1 1 237
0 117 5 1 1 267
0 118 5 1 1 297
0 119 5 1 1 327
0 120 5 1 1 357
0 121 5 1 1 387
0 122 5 1 1 417
0 123 5 1 1 447
0 124 5 1 1 477
0 125 5 1 1 507
0 126 5 1 1 537
0 127 5 1 1 567
0 128 5 1 1 597
0 129 5 1 1 628
0 130 5 1 1 632
0 131 5 2 1 634
0 132 5 2 1 636
0 133 5 2 1 638
0 134 5 2 1 640
0 135 5 2 1 642
0 136 5 2 1 644
0 137 5 2 1 646
0 138 5 2 1 648
0 139 5 2 1 650
0 140 5 2 1 652
0 141 5 2 1 654
0 142 5 2 1 656
0 143 5 2 1 658
0 144 5 2 1 660
0 145 5 2 1 662
0 146 5 2 1 664
0 147 5 2 1 666
0 148 5 2 1 668
0 149 5 2 1 670
0 150 5 2 1 672
0 151 5 2 1 674
0 152 5 2 1 676
0 153 5 2 1 678
0 154 5 2 1 680
0 155 5 2 1 682
0 156 5 2 1 684
0 157 5 2 1 686
0 158 5 2 1 688
0 159 5 2 1 690
0 160 5 1 1 692
0 161 7 2 2 65 631
0 162 5 3 1 752
0 163 7 1 2 97 129
0 164 5 1 1 163
3 1267 7 0 2 754 164
0 166 7 1 2 67 633
0 167 5 2 1 166
0 168 7 1 2 98 130
0 169 5 2 1 168
0 170 7 2 2 757 759
0 171 5 1 1 761
0 172 7 1 2 753 171
0 173 5 1 1 172
0 174 7 1 2 755 762
0 175 5 1 1 174
0 176 7 1 2 173 175
3 1268 5 0 1 176
0 178 7 1 2 756 758
0 179 5 1 1 178
0 180 7 2 2 760 179
0 181 5 1 1 763
0 182 7 1 2 99 181
0 183 5 2 1 182
0 184 7 1 2 69 764
0 185 5 2 1 184
0 186 7 2 2 765 767
0 187 5 1 1 769
0 188 7 1 2 635 770
0 189 5 1 1 188
0 190 7 1 2 694 187
0 191 5 1 1 190
3 1269 7 0 2 189 191
0 193 7 1 2 695 768
0 194 5 1 1 193
0 195 7 2 2 766 194
0 196 5 1 1 771
0 197 7 1 2 100 196
0 198 5 2 1 197
0 199 7 1 2 71 772
0 200 5 2 1 199
0 201 7 2 2 773 775
0 202 5 1 1 777
0 203 7 1 2 637 778
0 204 5 1 1 203
0 205 7 1 2 696 202
0 206 5 1 1 205
3 1270 7 0 2 204 206
0 208 7 1 2 697 776
0 209 5 1 1 208
0 210 7 2 2 774 209
0 211 5 1 1 779
0 212 7 1 2 101 211
0 213 5 2 1 212
0 214 7 1 2 73 780
0 215 5 2 1 214
0 216 7 2 2 781 783
0 217 5 1 1 785
0 218 7 1 2 639 786
0 219 5 1 1 218
0 220 7 1 2 698 217
0 221 5 1 1 220
3 1271 7 0 2 219 221
0 223 7 1 2 699 784
0 224 5 1 1 223
0 225 7 2 2 782 224
0 226 5 1 1 787
0 227 7 1 2 102 226
0 228 5 2 1 227
0 229 7 1 2 75 788
0 230 5 2 1 229
0 231 7 2 2 789 791
0 232 5 1 1 793
0 233 7 1 2 641 794
0 234 5 1 1 233
0 235 7 1 2 700 232
0 236 5 1 1 235
3 1272 7 0 2 234 236
0 238 7 1 2 701 792
0 239 5 1 1 238
0 240 7 2 2 790 239
0 241 5 1 1 795
0 242 7 1 2 103 241
0 243 5 2 1 242
0 244 7 1 2 77 796
0 245 5 2 1 244
0 246 7 2 2 797 799
0 247 5 1 1 801
0 248 7 1 2 643 802
0 249 5 1 1 248
0 250 7 1 2 702 247
0 251 5 1 1 250
3 1273 7 0 2 249 251
0 253 7 1 2 703 800
0 254 5 1 1 253
0 255 7 2 2 798 254
0 256 5 1 1 803
0 257 7 1 2 79 804
0 258 5 2 1 257
0 259 7 1 2 104 256
0 260 5 2 1 259
0 261 7 2 2 805 807
0 262 5 1 1 809
0 263 7 1 2 645 810
0 264 5 1 1 263
0 265 7 1 2 704 262
0 266 5 1 1 265
3 1274 7 0 2 264 266
0 268 7 1 2 705 806
0 269 5 1 1 268
0 270 7 2 2 808 269
0 271 5 1 1 811
0 272 7 1 2 105 271
0 273 5 2 1 272
0 274 7 1 2 81 812
0 275 5 2 1 274
0 276 7 2 2 813 815
0 277 5 1 1 817
0 278 7 1 2 647 818
0 279 5 1 1 278
0 280 7 1 2 706 277
0 281 5 1 1 280
3 1275 7 0 2 279 281
0 283 7 1 2 707 816
0 284 5 1 1 283
0 285 7 2 2 814 284
0 286 5 1 1 819
0 287 7 1 2 106 286
0 288 5 2 1 287
0 289 7 1 2 83 820
0 290 5 2 1 289
0 291 7 2 2 821 823
0 292 5 1 1 825
0 293 7 1 2 649 826
0 294 5 1 1 293
0 295 7 1 2 708 292
0 296 5 1 1 295
3 1276 7 0 2 294 296
0 298 7 1 2 709 824
0 299 5 1 1 298
0 300 7 2 2 822 299
0 301 5 1 1 827
0 302 7 1 2 107 301
0 303 5 2 1 302
0 304 7 1 2 85 828
0 305 5 2 1 304
0 306 7 2 2 829 831
0 307 5 1 1 833
0 308 7 1 2 651 834
0 309 5 1 1 308
0 310 7 1 2 710 307
0 311 5 1 1 310
3 1277 7 0 2 309 311
0 313 7 1 2 711 832
0 314 5 1 1 313
0 315 7 2 2 830 314
0 316 5 1 1 835
0 317 7 1 2 108 316
0 318 5 2 1 317
0 319 7 1 2 87 836
0 320 5 2 1 319
0 321 7 2 2 837 839
0 322 5 1 1 841
0 323 7 1 2 653 842
0 324 5 1 1 323
0 325 7 1 2 712 322
0 326 5 1 1 325
3 1278 7 0 2 324 326
0 328 7 1 2 713 840
0 329 5 1 1 328
0 330 7 2 2 838 329
0 331 5 1 1 843
0 332 7 1 2 109 331
0 333 5 2 1 332
0 334 7 1 2 89 844
0 335 5 2 1 334
0 336 7 2 2 845 847
0 337 5 1 1 849
0 338 7 1 2 655 850
0 339 5 1 1 338
0 340 7 1 2 714 337
0 341 5 1 1 340
3 1279 7 0 2 339 341
0 343 7 1 2 715 848
0 344 5 1 1 343
0 345 7 2 2 846 344
0 346 5 1 1 851
0 347 7 1 2 110 346
0 348 5 2 1 347
0 349 7 1 2 91 852
0 350 5 2 1 349
0 351 7 2 2 853 855
0 352 5 1 1 857
0 353 7 1 2 657 858
0 354 5 1 1 353
0 355 7 1 2 716 352
0 356 5 1 1 355
3 1280 7 0 2 354 356
0 358 7 1 2 717 856
0 359 5 1 1 358
0 360 7 2 2 854 359
0 361 5 1 1 859
0 362 7 1 2 93 860
0 363 5 2 1 362
0 364 7 1 2 111 361
0 365 5 2 1 364
0 366 7 2 2 861 863
0 367 5 1 1 865
0 368 7 1 2 659 866
0 369 5 1 1 368
0 370 7 1 2 718 367
0 371 5 1 1 370
3 1281 7 0 2 369 371
0 373 7 1 2 719 862
0 374 5 1 1 373
0 375 7 2 2 864 374
0 376 5 1 1 867
0 377 7 1 2 112 376
0 378 5 2 1 377
0 379 7 1 2 95 868
0 380 5 2 1 379
0 381 7 2 2 869 871
0 382 5 1 1 873
0 383 7 1 2 661 874
0 384 5 1 1 383
0 385 7 1 2 720 382
0 386 5 1 1 385
3 1282 7 0 2 384 386
0 388 7 1 2 721 872
0 389 5 1 1 388
0 390 7 2 2 870 389
0 391 5 1 1 875
0 392 7 1 2 113 391
0 393 5 2 1 392
0 394 7 1 2 165 876
0 395 5 2 1 394
0 396 7 2 2 877 879
0 397 5 1 1 881
0 398 7 1 2 663 882
0 399 5 1 1 398
0 400 7 1 2 722 397
0 401 5 1 1 400
3 1283 7 0 2 399 401
0 403 7 1 2 723 880
0 404 5 1 1 403
0 405 7 2 2 878 404
0 406 5 1 1 883
0 407 7 1 2 114 406
0 408 5 2 1 407
0 409 7 1 2 192 884
0 410 5 2 1 409
0 411 7 2 2 885 887
0 412 5 1 1 889
0 413 7 1 2 665 890
0 414 5 1 1 413
0 415 7 1 2 724 412
0 416 5 1 1 415
3 1284 7 0 2 414 416
0 418 7 1 2 725 888
0 419 5 1 1 418
0 420 7 2 2 886 419
0 421 5 1 1 891
0 422 7 1 2 115 421
0 423 5 2 1 422
0 424 7 1 2 222 892
0 425 5 2 1 424
0 426 7 2 2 893 895
0 427 5 1 1 897
0 428 7 1 2 667 898
0 429 5 1 1 428
0 430 7 1 2 726 427
0 431 5 1 1 430
3 1285 7 0 2 429 431
0 433 7 1 2 727 896
0 434 5 1 1 433
0 435 7 2 2 894 434
0 436 5 1 1 899
0 437 7 1 2 116 436
0 438 5 2 1 437
0 439 7 1 2 252 900
0 440 5 2 1 439
0 441 7 2 2 901 903
0 442 5 1 1 905
0 443 7 1 2 669 906
0 444 5 1 1 443
0 445 7 1 2 728 442
0 446 5 1 1 445
3 1286 7 0 2 444 446
0 448 7 1 2 729 904
0 449 5 1 1 448
0 450 7 2 2 902 449
0 451 5 1 1 907
0 452 7 1 2 117 451
0 453 5 2 1 452
0 454 7 1 2 282 908
0 455 5 2 1 454
0 456 7 2 2 909 911
0 457 5 1 1 913
0 458 7 1 2 671 914
0 459 5 1 1 458
0 460 7 1 2 730 457
0 461 5 1 1 460
3 1287 7 0 2 459 461
0 463 7 1 2 731 912
0 464 5 1 1 463
0 465 7 2 2 910 464
0 466 5 1 1 915
0 467 7 1 2 118 466
0 468 5 2 1 467
0 469 7 1 2 312 916
0 470 5 2 1 469
0 471 7 2 2 917 919
0 472 5 1 1 921
0 473 7 1 2 673 922
0 474 5 1 1 473
0 475 7 1 2 732 472
0 476 5 1 1 475
3 1288 7 0 2 474 476
0 478 7 1 2 733 920
0 479 5 1 1 478
0 480 7 2 2 918 479
0 481 5 1 1 923
0 482 7 1 2 119 481
0 483 5 2 1 482
0 484 7 1 2 342 924
0 485 5 2 1 484
0 486 7 2 2 925 927
0 487 5 1 1 929
0 488 7 1 2 675 930
0 489 5 1 1 488
0 490 7 1 2 734 487
0 491 5 1 1 490
3 1289 7 0 2 489 491
0 493 7 1 2 735 928
0 494 5 1 1 493
0 495 7 2 2 926 494
0 496 5 1 1 931
0 497 7 1 2 120 496
0 498 5 2 1 497
0 499 7 1 2 372 932
0 500 5 2 1 499
0 501 7 2 2 933 935
0 502 5 1 1 937
0 503 7 1 2 677 938
0 504 5 1 1 503
0 505 7 1 2 736 502
0 506 5 1 1 505
3 1290 7 0 2 504 506
0 508 7 1 2 737 936
0 509 5 1 1 508
0 510 7 2 2 934 509
0 511 5 1 1 939
0 512 7 1 2 121 511
0 513 5 2 1 512
0 514 7 1 2 402 940
0 515 5 2 1 514
0 516 7 2 2 941 943
0 517 5 1 1 945
0 518 7 1 2 679 946
0 519 5 1 1 518
0 520 7 1 2 738 517
0 521 5 1 1 520
3 1291 7 0 2 519 521
0 523 7 1 2 739 944
0 524 5 1 1 523
0 525 7 2 2 942 524
0 526 5 1 1 947
0 527 7 1 2 122 526
0 528 5 2 1 527
0 529 7 1 2 432 948
0 530 5 2 1 529
0 531 7 2 2 949 951
0 532 5 1 1 953
0 533 7 1 2 681 954
0 534 5 1 1 533
0 535 7 1 2 740 532
0 536 5 1 1 535
3 1292 7 0 2 534 536
0 538 7 1 2 741 952
0 539 5 1 1 538
0 540 7 2 2 950 539
0 541 5 1 1 955
0 542 7 1 2 123 541
0 543 5 2 1 542
0 544 7 1 2 462 956
0 545 5 2 1 544
0 546 7 2 2 957 959
0 547 5 1 1 961
0 548 7 1 2 683 962
0 549 5 1 1 548
0 550 7 1 2 742 547
0 551 5 1 1 550
3 1293 7 0 2 549 551
0 553 7 1 2 743 960
0 554 5 1 1 553
0 555 7 2 2 958 554
0 556 5 1 1 963
0 557 7 1 2 124 556
0 558 5 2 1 557
0 559 7 1 2 492 964
0 560 5 2 1 559
0 561 7 2 2 965 967
0 562 5 1 1 969
0 563 7 1 2 685 970
0 564 5 1 1 563
0 565 7 1 2 744 562
0 566 5 1 1 565
3 1294 7 0 2 564 566
0 568 7 1 2 745 968
0 569 5 1 1 568
0 570 7 2 2 966 569
0 571 5 1 1 971
0 572 7 1 2 125 571
0 573 5 2 1 572
0 574 7 1 2 522 972
0 575 5 2 1 574
0 576 7 2 2 973 975
0 577 5 1 1 977
0 578 7 1 2 687 978
0 579 5 1 1 578
0 580 7 1 2 746 577
0 581 5 1 1 580
3 1295 7 0 2 579 581
0 583 7 1 2 747 976
0 584 5 1 1 583
0 585 7 2 2 974 584
0 586 5 1 1 979
0 587 7 1 2 126 586
0 588 5 2 1 587
0 589 7 1 2 552 980
0 590 5 2 1 589
0 591 7 2 2 981 983
0 592 5 1 1 985
0 593 7 1 2 689 986
0 594 5 1 1 593
0 595 7 1 2 748 592
0 596 5 1 1 595
3 1296 7 0 2 594 596
0 598 7 1 2 749 984
0 599 5 1 1 598
0 600 7 2 2 982 599
0 601 5 1 1 987
0 602 7 1 2 127 601
0 603 5 2 1 602
0 604 7 1 2 582 988
0 605 5 2 1 604
0 606 7 2 2 989 991
0 607 5 1 1 993
0 608 7 1 2 691 994
0 609 5 1 1 608
0 610 7 1 2 750 607
0 611 5 1 1 610
3 1297 7 0 2 609 611
0 613 7 1 2 751 992
0 614 5 1 1 613
0 615 7 2 2 990 614
0 616 5 2 1 995
0 617 7 1 2 128 160
0 618 5 2 1 617
0 619 7 1 2 612 693
0 620 5 2 1 619
0 621 7 2 2 999 1001
0 622 5 1 1 1003
0 623 7 1 2 996 622
0 624 5 1 1 623
0 625 7 1 2 997 1004
0 626 5 1 1 625
0 627 7 1 2 624 626
3 1298 5 0 1 627
0 629 7 1 2 998 1002
0 630 5 1 1 629
3 1299 7 0 2 1000 630
