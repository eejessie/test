1 0 0 2 0
2 49 1 0
2 730 1 0
1 1 0 2 0
2 731 1 1
2 732 1 1
1 2 0 2 0
2 733 1 2
2 734 1 2
1 3 0 2 0
2 735 1 3
2 736 1 3
1 4 0 2 0
2 737 1 4
2 738 1 4
1 5 0 2 0
2 739 1 5
2 740 1 5
1 6 0 2 0
2 741 1 6
2 742 1 6
1 7 0 2 0
2 743 1 7
2 744 1 7
1 8 0 2 0
2 745 1 8
2 746 1 8
1 9 0 2 0
2 747 1 9
2 748 1 9
1 10 0 2 0
2 749 1 10
2 750 1 10
1 11 0 2 0
2 751 1 11
2 752 1 11
1 12 0 2 0
2 753 1 12
2 754 1 12
1 13 0 2 0
2 755 1 13
2 756 1 13
1 14 0 2 0
2 757 1 14
2 758 1 14
1 15 0 2 0
2 759 1 15
2 760 1 15
1 16 0 2 0
2 761 1 16
2 762 1 16
1 17 0 2 0
2 763 1 17
2 764 1 17
1 18 0 2 0
2 765 1 18
2 766 1 18
1 19 0 2 0
2 767 1 19
2 768 1 19
1 20 0 2 0
2 769 1 20
2 770 1 20
1 21 0 2 0
2 771 1 21
2 772 1 21
1 22 0 2 0
2 773 1 22
2 774 1 22
1 23 0 2 0
2 775 1 23
2 776 1 23
1 24 0 2 0
2 777 1 24
2 778 1 24
1 25 0 2 0
2 779 1 25
2 780 1 25
1 26 0 2 0
2 781 1 26
2 782 1 26
1 27 0 2 0
2 783 1 27
2 784 1 27
1 28 0 2 0
2 785 1 28
2 786 1 28
1 29 0 2 0
2 787 1 29
2 788 1 29
1 30 0 2 0
2 789 1 30
2 790 1 30
1 31 0 2 0
2 791 1 31
2 792 1 31
1 32 0 2 0
2 793 1 32
2 794 1 32
1 33 0 2 0
2 795 1 33
2 796 1 33
1 34 0 2 0
2 797 1 34
2 798 1 34
1 35 0 2 0
2 799 1 35
2 800 1 35
1 36 0 2 0
2 801 1 36
2 802 1 36
1 37 0 2 0
2 803 1 37
2 804 1 37
1 38 0 2 0
2 805 1 38
2 806 1 38
1 39 0 2 0
2 807 1 39
2 808 1 39
1 40 0 2 0
2 809 1 40
2 810 1 40
1 41 0 2 0
2 811 1 41
2 812 1 41
1 42 0 2 0
2 813 1 42
2 814 1 42
1 43 0 2 0
2 815 1 43
2 816 1 43
1 44 0 2 0
2 817 1 44
2 818 1 44
1 45 0 2 0
2 819 1 45
2 820 1 45
1 46 0 2 0
2 821 1 46
2 822 1 46
1 47 0 2 0
2 823 1 47
2 824 1 47
1 48 0 2 0
2 825 1 48
2 826 1 48
2 827 1 69
2 828 1 69
2 829 1 70
2 830 1 70
2 831 1 71
2 832 1 71
2 833 1 72
2 834 1 72
2 835 1 73
2 836 1 73
2 837 1 74
2 838 1 74
2 839 1 75
2 840 1 75
2 841 1 76
2 842 1 76
2 843 1 77
2 844 1 77
2 845 1 78
2 846 1 78
2 847 1 79
2 848 1 79
2 849 1 80
2 850 1 80
2 851 1 81
2 852 1 81
2 853 1 100
2 854 1 100
2 855 1 102
2 856 1 102
2 857 1 104
2 858 1 104
2 859 1 106
2 860 1 106
2 861 1 107
2 862 1 107
2 863 1 108
2 864 1 108
2 865 1 108
2 866 1 111
2 867 1 111
2 868 1 112
2 869 1 112
2 870 1 115
2 871 1 115
2 872 1 118
2 873 1 118
2 874 1 120
2 875 1 120
2 876 1 123
2 877 1 123
2 878 1 126
2 879 1 126
2 880 1 128
2 881 1 128
2 882 1 131
2 883 1 131
2 884 1 134
2 885 1 134
2 886 1 136
2 887 1 136
2 888 1 139
2 889 1 139
2 890 1 142
2 891 1 142
2 892 1 144
2 893 1 144
2 894 1 147
2 895 1 147
2 896 1 150
2 897 1 150
2 898 1 152
2 899 1 152
2 900 1 155
2 901 1 155
2 902 1 158
2 903 1 158
2 904 1 160
2 905 1 160
2 906 1 163
2 907 1 163
2 908 1 166
2 909 1 166
2 910 1 168
2 911 1 168
2 912 1 171
2 913 1 171
2 914 1 174
2 915 1 174
2 916 1 176
2 917 1 176
2 918 1 179
2 919 1 179
2 920 1 182
2 921 1 182
2 922 1 184
2 923 1 184
2 924 1 187
2 925 1 187
2 926 1 190
2 927 1 190
2 928 1 192
2 929 1 192
2 930 1 195
2 931 1 195
2 932 1 198
2 933 1 198
2 934 1 200
2 935 1 200
2 936 1 203
2 937 1 203
2 938 1 206
2 939 1 206
2 940 1 208
2 941 1 208
2 942 1 211
2 943 1 211
2 944 1 214
2 945 1 214
2 946 1 216
2 947 1 216
2 948 1 219
2 949 1 219
2 950 1 221
2 951 1 221
2 952 1 222
2 953 1 222
2 954 1 223
2 955 1 223
2 956 1 224
2 957 1 224
2 958 1 225
2 959 1 225
2 960 1 231
2 961 1 231
2 962 1 234
2 963 1 234
2 964 1 234
2 965 1 235
2 966 1 235
2 967 1 241
2 968 1 241
2 969 1 244
2 970 1 244
2 971 1 244
2 972 1 244
2 973 1 246
2 974 1 246
2 975 1 246
2 976 1 247
2 977 1 247
2 978 1 253
2 979 1 253
2 980 1 256
2 981 1 256
2 982 1 256
2 983 1 256
2 984 1 258
2 985 1 258
2 986 1 258
2 987 1 259
2 988 1 259
2 989 1 265
2 990 1 265
2 991 1 268
2 992 1 268
2 993 1 268
2 994 1 268
2 995 1 270
2 996 1 270
2 997 1 270
2 998 1 271
2 999 1 271
2 1000 1 277
2 1001 1 277
2 1002 1 280
2 1003 1 280
2 1004 1 280
2 1005 1 280
2 1006 1 281
2 1007 1 281
2 1008 1 287
2 1009 1 287
2 1010 1 290
2 1011 1 290
2 1012 1 290
2 1013 1 290
2 1014 1 292
2 1015 1 292
2 1016 1 292
2 1017 1 292
2 1018 1 293
2 1019 1 293
2 1020 1 299
2 1021 1 299
2 1022 1 302
2 1023 1 302
2 1024 1 302
2 1025 1 302
2 1026 1 304
2 1027 1 304
2 1028 1 304
2 1029 1 304
2 1030 1 305
2 1031 1 305
2 1032 1 311
2 1033 1 311
2 1034 1 314
2 1035 1 314
2 1036 1 314
2 1037 1 316
2 1038 1 316
2 1039 1 316
2 1040 1 317
2 1041 1 317
2 1042 1 323
2 1043 1 323
2 1044 1 326
2 1045 1 326
2 1046 1 326
2 1047 1 326
2 1048 1 328
2 1049 1 328
2 1050 1 328
2 1051 1 328
2 1052 1 329
2 1053 1 329
2 1054 1 335
2 1055 1 335
2 1056 1 338
2 1057 1 338
2 1058 1 338
2 1059 1 338
2 1060 1 340
2 1061 1 340
2 1062 1 340
2 1063 1 340
2 1064 1 341
2 1065 1 341
2 1066 1 347
2 1067 1 347
2 1068 1 350
2 1069 1 350
2 1070 1 350
2 1071 1 350
2 1072 1 352
2 1073 1 352
2 1074 1 352
2 1075 1 353
2 1076 1 353
2 1077 1 359
2 1078 1 359
2 1079 1 362
2 1080 1 362
2 1081 1 362
2 1082 1 364
2 1083 1 364
2 1084 1 364
2 1085 1 364
2 1086 1 365
2 1087 1 365
2 1088 1 371
2 1089 1 371
2 1090 1 374
2 1091 1 374
2 1092 1 374
2 1093 1 374
2 1094 1 376
2 1095 1 376
2 1096 1 376
2 1097 1 377
2 1098 1 377
2 1099 1 383
2 1100 1 383
2 1101 1 386
2 1102 1 386
2 1103 1 386
2 1104 1 386
2 1105 1 387
2 1106 1 387
2 1107 1 393
2 1108 1 393
2 1109 1 396
2 1110 1 396
2 1111 1 398
2 1112 1 398
2 1113 1 401
2 1114 1 401
2 1115 1 405
2 1116 1 405
2 1117 1 406
2 1118 1 406
2 1119 1 407
2 1120 1 407
2 1121 1 411
2 1122 1 411
2 1123 1 411
2 1124 1 413
2 1125 1 413
2 1126 1 415
2 1127 1 415
2 1128 1 415
2 1129 1 419
2 1130 1 419
2 1131 1 421
2 1132 1 421
2 1133 1 423
2 1134 1 423
2 1135 1 429
2 1136 1 429
2 1137 1 431
2 1138 1 431
2 1139 1 432
2 1140 1 432
2 1141 1 435
2 1142 1 435
2 1143 1 438
2 1144 1 438
2 1145 1 442
2 1146 1 442
2 1147 1 447
2 1148 1 447
2 1149 1 447
2 1150 1 447
2 1151 1 450
2 1152 1 450
2 1153 1 454
2 1154 1 454
2 1155 1 460
2 1156 1 460
2 1157 1 462
2 1158 1 462
2 1159 1 462
2 1160 1 465
2 1161 1 465
2 1162 1 469
2 1163 1 469
2 1164 1 473
2 1165 1 473
2 1166 1 473
2 1167 1 474
2 1168 1 474
2 1169 1 479
2 1170 1 479
2 1171 1 479
2 1172 1 485
2 1173 1 485
2 1174 1 485
2 1175 1 491
2 1176 1 491
2 1177 1 492
2 1178 1 492
2 1179 1 495
2 1180 1 495
2 1181 1 500
2 1182 1 500
2 1183 1 506
2 1184 1 506
2 1185 1 509
2 1186 1 509
2 1187 1 509
2 1188 1 510
2 1189 1 510
2 1190 1 514
2 1191 1 514
2 1192 1 520
2 1193 1 520
2 1194 1 525
2 1195 1 525
2 1196 1 526
2 1197 1 526
2 1198 1 529
2 1199 1 529
2 1200 1 530
2 1201 1 530
2 1202 1 535
2 1203 1 535
2 1204 1 536
2 1205 1 536
2 1206 1 540
2 1207 1 540
2 1208 1 540
2 1209 1 545
2 1210 1 545
2 1211 1 581
2 1212 1 581
2 1213 1 581
2 1214 1 585
2 1215 1 585
2 1216 1 585
2 1217 1 589
2 1218 1 589
2 1219 1 591
2 1220 1 591
2 1221 1 593
2 1222 1 593
2 1223 1 594
2 1224 1 594
2 1225 1 597
2 1226 1 597
2 1227 1 601
2 1228 1 601
2 1229 1 603
2 1230 1 603
2 1231 1 604
2 1232 1 604
2 1233 1 607
2 1234 1 607
2 1235 1 610
2 1236 1 610
2 1237 1 614
2 1238 1 614
2 1239 1 619
2 1240 1 619
2 1241 1 623
2 1242 1 623
2 1243 1 624
2 1244 1 624
2 1245 1 627
2 1246 1 627
2 1247 1 628
2 1248 1 628
2 1249 1 631
2 1250 1 631
2 1251 1 632
2 1252 1 632
2 1253 1 719
2 1254 1 719
0 50 5 1 1 49
0 51 5 1 1 731
0 52 5 1 1 733
0 53 5 1 1 735
0 54 5 1 1 737
0 55 5 1 1 739
0 56 5 1 1 741
0 57 5 1 1 743
0 58 5 1 1 745
0 59 5 1 1 747
0 60 5 1 1 749
0 61 5 1 1 751
0 62 5 1 1 753
0 63 5 1 1 755
0 64 5 1 1 757
0 65 5 1 1 759
0 66 5 1 1 761
0 67 5 1 1 763
0 68 5 1 1 765
0 69 5 2 1 767
0 70 5 2 1 769
0 71 5 2 1 771
0 72 5 2 1 773
0 73 5 2 1 775
0 74 5 2 1 777
0 75 5 2 1 779
0 76 5 2 1 781
0 77 5 2 1 783
0 78 5 2 1 785
0 79 5 2 1 787
0 80 5 2 1 789
0 81 5 2 1 791
0 82 5 1 1 793
0 83 5 1 1 795
0 84 5 1 1 797
0 85 5 1 1 799
0 86 5 1 1 801
0 87 5 1 1 803
0 88 5 1 1 805
0 89 5 1 1 807
0 90 5 1 1 809
0 91 5 1 1 811
0 92 5 1 1 813
0 93 5 1 1 815
0 94 5 1 1 817
0 95 5 1 1 819
0 96 5 1 1 821
0 97 5 1 1 823
0 98 5 1 1 825
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 734 766
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 732 764
0 106 5 2 1 105
0 107 7 2 2 730 762
0 108 5 3 1 861
0 109 7 1 2 859 863
0 110 5 1 1 109
0 111 7 2 2 857 110
0 112 5 2 1 866
0 113 7 1 2 855 868
0 114 5 1 1 113
0 115 7 2 2 853 114
0 116 5 1 1 870
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 736 871
0 120 5 2 1 119
0 121 7 1 2 827 874
0 122 5 1 1 121
0 123 7 2 2 872 122
0 124 5 1 1 876
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 738 877
0 128 5 2 1 127
0 129 7 1 2 829 880
0 130 5 1 1 129
0 131 7 2 2 878 130
0 132 5 1 1 882
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 740 883
0 136 5 2 1 135
0 137 7 1 2 831 886
0 138 5 1 1 137
0 139 7 2 2 884 138
0 140 5 1 1 888
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 742 889
0 144 5 2 1 143
0 145 7 1 2 833 892
0 146 5 1 1 145
0 147 7 2 2 890 146
0 148 5 1 1 894
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 744 895
0 152 5 2 1 151
0 153 7 1 2 835 898
0 154 5 1 1 153
0 155 7 2 2 896 154
0 156 5 1 1 900
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 746 901
0 160 5 2 1 159
0 161 7 1 2 837 904
0 162 5 1 1 161
0 163 7 2 2 902 162
0 164 5 1 1 906
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 748 907
0 168 5 2 1 167
0 169 7 1 2 839 910
0 170 5 1 1 169
0 171 7 2 2 908 170
0 172 5 1 1 912
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 750 913
0 176 5 2 1 175
0 177 7 1 2 841 916
0 178 5 1 1 177
0 179 7 2 2 914 178
0 180 5 1 1 918
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 752 919
0 184 5 2 1 183
0 185 7 1 2 843 922
0 186 5 1 1 185
0 187 7 2 2 920 186
0 188 5 1 1 924
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 754 925
0 192 5 2 1 191
0 193 7 1 2 845 928
0 194 5 1 1 193
0 195 7 2 2 926 194
0 196 5 1 1 930
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 756 931
0 200 5 2 1 199
0 201 7 1 2 847 934
0 202 5 1 1 201
0 203 7 2 2 932 202
0 204 5 1 1 936
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 758 937
0 208 5 2 1 207
0 209 7 1 2 849 940
0 210 5 1 1 209
0 211 7 2 2 938 210
0 212 5 1 1 942
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 760 943
0 216 5 2 1 215
0 217 7 1 2 851 946
0 218 5 1 1 217
0 219 7 2 2 944 218
0 220 5 1 1 948
0 221 7 2 2 826 220
0 222 5 2 1 950
0 223 7 2 2 98 949
0 224 5 2 1 954
0 225 7 2 2 945 947
0 226 5 1 1 958
0 227 7 1 2 792 226
0 228 5 1 1 227
0 229 7 1 2 852 959
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 960
0 233 7 1 2 824 961
0 234 5 3 1 233
0 235 7 2 2 939 941
0 236 5 1 1 965
0 237 7 1 2 790 966
0 238 5 1 1 237
0 239 7 1 2 850 236
0 240 5 1 1 239
0 241 7 2 2 238 240
0 242 5 1 1 967
0 243 7 1 2 822 242
0 244 5 4 1 243
0 245 7 1 2 96 968
0 246 5 3 1 245
0 247 7 2 2 933 935
0 248 5 1 1 976
0 249 7 1 2 788 977
0 250 5 1 1 249
0 251 7 1 2 848 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 978
0 255 7 1 2 820 254
0 256 5 4 1 255
0 257 7 1 2 95 979
0 258 5 3 1 257
0 259 7 2 2 927 929
0 260 5 1 1 987
0 261 7 1 2 786 988
0 262 5 1 1 261
0 263 7 1 2 846 260
0 264 5 1 1 263
0 265 7 2 2 262 264
0 266 5 1 1 989
0 267 7 1 2 818 266
0 268 5 4 1 267
0 269 7 1 2 94 990
0 270 5 3 1 269
0 271 7 2 2 921 923
0 272 5 1 1 998
0 273 7 1 2 784 999
0 274 5 1 1 273
0 275 7 1 2 844 272
0 276 5 1 1 275
0 277 7 2 2 274 276
0 278 5 1 1 1000
0 279 7 1 2 816 278
0 280 5 4 1 279
0 281 7 2 2 915 917
0 282 5 1 1 1006
0 283 7 1 2 782 1007
0 284 5 1 1 283
0 285 7 1 2 842 282
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 1008
0 289 7 1 2 814 288
0 290 5 4 1 289
0 291 7 1 2 92 1009
0 292 5 4 1 291
0 293 7 2 2 909 911
0 294 5 1 1 1018
0 295 7 1 2 780 1019
0 296 5 1 1 295
0 297 7 1 2 840 294
0 298 5 1 1 297
0 299 7 2 2 296 298
0 300 5 1 1 1020
0 301 7 1 2 812 300
0 302 5 4 1 301
0 303 7 1 2 91 1021
0 304 5 4 1 303
0 305 7 2 2 903 905
0 306 5 1 1 1030
0 307 7 1 2 778 1031
0 308 5 1 1 307
0 309 7 1 2 838 306
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 1032
0 313 7 1 2 810 312
0 314 5 3 1 313
0 315 7 1 2 90 1033
0 316 5 3 1 315
0 317 7 2 2 897 899
0 318 5 1 1 1040
0 319 7 1 2 776 1041
0 320 5 1 1 319
0 321 7 1 2 836 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1042
0 325 7 1 2 808 324
0 326 5 4 1 325
0 327 7 1 2 89 1043
0 328 5 4 1 327
0 329 7 2 2 891 893
0 330 5 1 1 1052
0 331 7 1 2 774 1053
0 332 5 1 1 331
0 333 7 1 2 834 330
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 1054
0 337 7 1 2 806 336
0 338 5 4 1 337
0 339 7 1 2 88 1055
0 340 5 4 1 339
0 341 7 2 2 885 887
0 342 5 1 1 1064
0 343 7 1 2 772 1065
0 344 5 1 1 343
0 345 7 1 2 832 342
0 346 5 1 1 345
0 347 7 2 2 344 346
0 348 5 1 1 1066
0 349 7 1 2 87 1067
0 350 5 4 1 349
0 351 7 1 2 804 348
0 352 5 3 1 351
0 353 7 2 2 879 881
0 354 5 1 1 1075
0 355 7 1 2 770 1076
0 356 5 1 1 355
0 357 7 1 2 830 354
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 1077
0 361 7 1 2 802 360
0 362 5 3 1 361
0 363 7 1 2 86 1078
0 364 5 4 1 363
0 365 7 2 2 873 875
0 366 5 1 1 1086
0 367 7 1 2 768 1087
0 368 5 1 1 367
0 369 7 1 2 828 366
0 370 5 1 1 369
0 371 7 2 2 368 370
0 372 5 1 1 1088
0 373 7 1 2 85 1089
0 374 5 4 1 373
0 375 7 1 2 800 372
0 376 5 3 1 375
0 377 7 2 2 854 856
0 378 5 1 1 1097
0 379 7 1 2 867 378
0 380 5 1 1 379
0 381 7 1 2 869 1098
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 1099
0 385 7 1 2 84 384
0 386 5 4 1 385
0 387 7 2 2 858 860
0 388 5 1 1 1105
0 389 7 1 2 862 388
0 390 5 1 1 389
0 391 7 1 2 864 1106
0 392 5 1 1 391
0 393 7 2 2 390 392
0 394 5 1 1 1107
0 395 7 1 2 83 394
0 396 5 2 1 395
0 397 7 1 2 796 1108
0 398 5 2 1 397
0 399 7 1 2 50 66
0 400 5 1 1 399
0 401 7 2 2 865 400
0 402 5 1 1 1113
0 403 7 1 2 794 402
0 404 5 1 1 403
0 405 7 2 2 1111 404
0 406 5 2 1 1115
0 407 7 2 2 1109 1117
0 408 7 1 2 1101 1119
0 409 5 1 1 408
0 410 7 1 2 798 1100
0 411 5 3 1 410
0 412 7 1 2 409 1121
0 413 7 2 2 1094 412
0 414 5 1 1 1124
0 415 7 3 2 1090 414
0 416 5 1 1 1126
0 417 7 1 2 1082 1127
0 418 5 1 1 417
0 419 7 2 2 1079 418
0 420 5 1 1 1129
0 421 7 2 2 1072 1130
0 422 5 1 1 1131
0 423 7 2 2 1068 422
0 424 5 1 1 1133
0 425 7 1 2 1060 1134
0 426 5 1 1 425
0 427 7 1 2 1056 426
0 428 5 1 1 427
0 429 7 2 2 1048 428
0 430 5 1 1 1135
0 431 7 2 2 1044 430
0 432 5 2 1 1137
0 433 7 1 2 1037 1139
0 434 5 1 1 433
0 435 7 2 2 1034 434
0 436 5 1 1 1141
0 437 7 1 2 1026 436
0 438 5 2 1 437
0 439 7 1 2 1022 1143
0 440 5 1 1 439
0 441 7 1 2 1014 440
0 442 5 2 1 441
0 443 7 1 2 1010 1145
0 444 7 1 2 1002 443
0 445 5 1 1 444
0 446 7 1 2 93 1001
0 447 5 4 1 446
0 448 7 1 2 445 1147
0 449 7 1 2 995 448
0 450 5 2 1 449
0 451 7 1 2 991 1151
0 452 5 1 1 451
0 453 7 1 2 984 452
0 454 5 2 1 453
0 455 7 1 2 980 1153
0 456 5 1 1 455
0 457 7 1 2 973 456
0 458 5 1 1 457
0 459 7 1 2 969 458
0 460 5 2 1 459
0 461 7 1 2 97 232
0 462 5 3 1 461
0 463 7 1 2 1155 1157
0 464 5 1 1 463
0 465 7 2 2 962 464
0 466 5 1 1 1160
0 467 7 1 2 956 466
0 468 5 1 1 467
0 469 7 2 2 952 468
0 470 5 1 1 1162
0 471 7 1 2 955 1161
0 472 5 1 1 471
0 473 7 3 2 1158 963
0 474 5 2 1 1164
0 475 7 1 2 970 1167
0 476 5 1 1 475
0 477 7 1 2 1156 1165
0 478 5 1 1 477
0 479 7 3 2 971 974
0 480 5 1 1 1169
0 481 7 1 2 1154 1170
0 482 5 1 1 481
0 483 7 1 2 981 482
0 484 5 1 1 483
0 485 7 3 2 982 985
0 486 5 1 1 1172
0 487 7 1 2 1152 1173
0 488 5 1 1 487
0 489 7 1 2 992 488
0 490 5 1 1 489
0 491 7 2 2 993 996
0 492 5 2 1 1175
0 493 7 1 2 1003 1177
0 494 5 1 1 493
0 495 7 2 2 1004 1148
0 496 7 1 2 1146 1179
0 497 5 1 1 496
0 498 7 1 2 1011 497
0 499 5 1 1 498
0 500 7 2 2 1012 1015
0 501 7 1 2 1144 1181
0 502 5 1 1 501
0 503 7 1 2 1023 502
0 504 5 1 1 503
0 505 7 1 2 1024 1027
0 506 5 2 1 505
0 507 7 1 2 1142 1183
0 508 5 1 1 507
0 509 7 3 2 1035 1038
0 510 5 2 1 1185
0 511 7 1 2 1138 1186
0 512 5 1 1 511
0 513 7 1 2 1045 1049
0 514 5 2 1 513
0 515 7 1 2 1057 1190
0 516 5 1 1 515
0 517 7 1 2 1046 1136
0 518 5 1 1 517
0 519 7 1 2 1058 1061
0 520 5 2 1 519
0 521 7 1 2 424 1192
0 522 5 1 1 521
0 523 7 1 2 1069 1132
0 524 5 1 1 523
0 525 7 2 2 1070 1073
0 526 5 2 1 1194
0 527 7 1 2 420 1196
0 528 5 1 1 527
0 529 7 2 2 1080 1083
0 530 5 2 1 1198
0 531 7 1 2 1128 1199
0 532 5 1 1 531
0 533 7 1 2 1091 1125
0 534 5 1 1 533
0 535 7 2 2 1092 1095
0 536 5 2 1 1202
0 537 7 1 2 1102 1204
0 538 5 1 1 537
0 539 7 1 2 1103 1122
0 540 5 3 1 539
0 541 7 1 2 1120 1206
0 542 5 1 1 541
0 543 7 1 2 82 1114
0 544 5 1 1 543
0 545 7 2 2 1110 544
0 546 5 1 1 1209
0 547 7 1 2 1116 1210
0 548 5 1 1 547
0 549 7 1 2 542 548
0 550 7 1 2 538 549
0 551 7 1 2 534 550
0 552 5 1 1 551
0 553 7 1 2 416 1200
0 554 5 1 1 553
0 555 7 1 2 552 554
0 556 7 1 2 532 555
0 557 5 1 1 556
0 558 7 1 2 528 557
0 559 7 1 2 524 558
0 560 5 1 1 559
0 561 7 1 2 522 560
0 562 7 1 2 518 561
0 563 7 1 2 516 562
0 564 5 1 1 563
0 565 7 1 2 1140 1188
0 566 5 1 1 565
0 567 7 1 2 564 566
0 568 7 1 2 512 567
0 569 5 1 1 568
0 570 7 1 2 508 569
0 571 7 1 2 504 570
0 572 7 1 2 499 571
0 573 7 1 2 494 572
0 574 7 1 2 490 573
0 575 7 1 2 484 574
0 576 7 1 2 478 575
0 577 7 1 2 476 576
0 578 7 1 2 472 577
0 579 7 1 2 1163 578
0 580 5 1 1 579
0 581 7 3 2 1112 546
0 582 5 1 1 1211
0 583 7 1 2 1123 1212
0 584 5 1 1 583
0 585 7 3 2 1104 584
0 586 5 1 1 1214
0 587 7 1 2 1093 1215
0 588 5 1 1 587
0 589 7 2 2 1096 588
0 590 5 1 1 1217
0 591 7 2 2 1081 1218
0 592 5 1 1 1219
0 593 7 2 2 1084 592
0 594 5 2 1 1221
0 595 7 1 2 1074 1223
0 596 5 1 1 595
0 597 7 2 2 1071 596
0 598 7 1 2 1062 1225
0 599 5 1 1 598
0 600 7 1 2 1059 599
0 601 7 2 2 1047 600
0 602 5 1 1 1227
0 603 7 2 2 1050 602
0 604 5 2 1 1229
0 605 7 1 2 1036 1231
0 606 5 1 1 605
0 607 7 2 2 1039 606
0 608 5 1 1 1233
0 609 7 1 2 1025 608
0 610 5 2 1 609
0 611 7 1 2 1028 1235
0 612 5 1 1 611
0 613 7 1 2 1013 612
0 614 5 2 1 613
0 615 7 1 2 1016 1237
0 616 5 1 1 615
0 617 7 1 2 1005 616
0 618 5 1 1 617
0 619 7 2 2 1149 618
0 620 5 1 1 1239
0 621 7 1 2 997 1240
0 622 5 1 1 621
0 623 7 2 2 994 622
0 624 5 2 1 1241
0 625 7 1 2 986 1243
0 626 5 1 1 625
0 627 7 2 2 983 626
0 628 5 2 1 1245
0 629 7 1 2 975 1247
0 630 5 1 1 629
0 631 7 2 2 972 630
0 632 5 2 1 1249
0 633 7 1 2 1166 1251
0 634 5 1 1 633
0 635 7 1 2 1168 1250
0 636 5 1 1 635
0 637 7 1 2 634 636
0 638 5 1 1 637
0 639 7 1 2 1174 1242
0 640 5 1 1 639
0 641 7 1 2 486 1244
0 642 5 1 1 641
0 643 7 1 2 1176 620
0 644 5 1 1 643
0 645 7 1 2 1150 1178
0 646 5 1 1 645
0 647 7 1 2 1180 1238
0 648 5 1 1 647
0 649 7 1 2 1017 648
0 650 5 1 1 649
0 651 7 1 2 1182 1236
0 652 5 1 1 651
0 653 7 1 2 1029 652
0 654 5 1 1 653
0 655 7 1 2 1184 1234
0 656 5 1 1 655
0 657 7 1 2 1187 1230
0 658 5 1 1 657
0 659 7 1 2 1051 1228
0 660 5 1 1 659
0 661 7 1 2 1063 1191
0 662 5 1 1 661
0 663 7 1 2 1193 1226
0 664 5 1 1 663
0 665 7 1 2 1195 1222
0 666 5 1 1 665
0 667 7 1 2 1085 1220
0 668 5 1 1 667
0 669 7 1 2 1201 590
0 670 5 1 1 669
0 671 7 1 2 1203 1216
0 672 5 1 1 671
0 673 7 1 2 1205 586
0 674 5 1 1 673
0 675 7 1 2 1207 1213
0 676 5 1 1 675
0 677 7 1 2 1118 1208
0 678 5 1 1 677
0 679 7 1 2 582 678
0 680 5 1 1 679
0 681 7 1 2 676 680
0 682 7 1 2 674 681
0 683 7 1 2 672 682
0 684 5 1 1 683
0 685 7 1 2 670 684
0 686 7 1 2 668 685
0 687 5 1 1 686
0 688 7 1 2 1197 1224
0 689 5 1 1 688
0 690 7 1 2 687 689
0 691 7 1 2 666 690
0 692 5 1 1 691
0 693 7 1 2 664 692
0 694 7 1 2 662 693
0 695 7 1 2 660 694
0 696 5 1 1 695
0 697 7 1 2 1189 1232
0 698 5 1 1 697
0 699 7 1 2 696 698
0 700 7 1 2 658 699
0 701 5 1 1 700
0 702 7 1 2 656 701
0 703 7 1 2 654 702
0 704 7 1 2 650 703
0 705 7 1 2 646 704
0 706 7 1 2 644 705
0 707 7 1 2 642 706
0 708 7 1 2 640 707
0 709 7 1 2 957 708
0 710 7 1 2 480 1248
0 711 5 1 1 710
0 712 7 1 2 1171 1246
0 713 5 1 1 712
0 714 7 1 2 711 713
0 715 7 1 2 709 714
0 716 7 1 2 638 715
0 717 7 1 2 1159 1252
0 718 5 1 1 717
0 719 7 2 2 964 718
0 720 5 1 1 1253
0 721 7 1 2 951 720
0 722 5 1 1 721
0 723 7 1 2 953 1254
0 724 5 1 1 723
0 725 7 1 2 722 724
0 726 7 1 2 716 725
0 727 7 1 2 470 726
0 728 5 1 1 727
0 729 7 1 2 580 728
3 4099 5 0 1 729
