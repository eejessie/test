1 0 0 2 0
2 49 1 0
2 1720 1 0
1 1 0 2 0
2 1721 1 1
2 1722 1 1
1 2 0 2 0
2 1723 1 2
2 1724 1 2
1 3 0 2 0
2 1725 1 3
2 1726 1 3
1 4 0 2 0
2 1727 1 4
2 1728 1 4
1 5 0 2 0
2 1729 1 5
2 1730 1 5
1 6 0 2 0
2 1731 1 6
2 1732 1 6
1 7 0 2 0
2 1733 1 7
2 1734 1 7
1 8 0 2 0
2 1735 1 8
2 1736 1 8
1 9 0 2 0
2 1737 1 9
2 1738 1 9
1 10 0 2 0
2 1739 1 10
2 1740 1 10
1 11 0 2 0
2 1741 1 11
2 1742 1 11
1 12 0 2 0
2 1743 1 12
2 1744 1 12
1 13 0 2 0
2 1745 1 13
2 1746 1 13
1 14 0 2 0
2 1747 1 14
2 1748 1 14
1 15 0 2 0
2 1749 1 15
2 1750 1 15
1 16 0 2 0
2 1751 1 16
2 1752 1 16
1 17 0 2 0
2 1753 1 17
2 1754 1 17
1 18 0 2 0
2 1755 1 18
2 1756 1 18
1 19 0 2 0
2 1757 1 19
2 1758 1 19
1 20 0 2 0
2 1759 1 20
2 1760 1 20
1 21 0 2 0
2 1761 1 21
2 1762 1 21
1 22 0 2 0
2 1763 1 22
2 1764 1 22
1 23 0 2 0
2 1765 1 23
2 1766 1 23
1 24 0 2 0
2 1767 1 24
2 1768 1 24
1 25 0 2 0
2 1769 1 25
2 1770 1 25
1 26 0 2 0
2 1771 1 26
2 1772 1 26
1 27 0 2 0
2 1773 1 27
2 1774 1 27
1 28 0 2 0
2 1775 1 28
2 1776 1 28
1 29 0 2 0
2 1777 1 29
2 1778 1 29
1 30 0 2 0
2 1779 1 30
2 1780 1 30
1 31 0 2 0
2 1781 1 31
2 1782 1 31
1 32 0 2 0
2 1783 1 32
2 1784 1 32
1 33 0 2 0
2 1785 1 33
2 1786 1 33
1 34 0 2 0
2 1787 1 34
2 1788 1 34
1 35 0 2 0
2 1789 1 35
2 1790 1 35
1 36 0 2 0
2 1791 1 36
2 1792 1 36
1 37 0 2 0
2 1793 1 37
2 1794 1 37
1 38 0 2 0
2 1795 1 38
2 1796 1 38
1 39 0 2 0
2 1797 1 39
2 1798 1 39
1 40 0 2 0
2 1799 1 40
2 1800 1 40
1 41 0 2 0
2 1801 1 41
2 1802 1 41
1 42 0 2 0
2 1803 1 42
2 1804 1 42
1 43 0 2 0
2 1805 1 43
2 1806 1 43
1 44 0 2 0
2 1807 1 44
2 1808 1 44
1 45 0 2 0
2 1809 1 45
2 1810 1 45
1 46 0 2 0
2 1811 1 46
2 1812 1 46
1 47 0 2 0
2 1813 1 47
2 1814 1 47
1 48 0 2 0
2 1815 1 48
2 1816 1 48
2 1817 1 69
2 1818 1 69
2 1819 1 70
2 1820 1 70
2 1821 1 71
2 1822 1 71
2 1823 1 72
2 1824 1 72
2 1825 1 73
2 1826 1 73
2 1827 1 74
2 1828 1 74
2 1829 1 75
2 1830 1 75
2 1831 1 76
2 1832 1 76
2 1833 1 77
2 1834 1 77
2 1835 1 78
2 1836 1 78
2 1837 1 79
2 1838 1 79
2 1839 1 80
2 1840 1 80
2 1841 1 99
2 1842 1 99
2 1843 1 100
2 1844 1 100
2 1845 1 101
2 1846 1 101
2 1847 1 102
2 1848 1 102
2 1849 1 104
2 1850 1 104
2 1851 1 106
2 1852 1 106
2 1853 1 108
2 1854 1 108
2 1855 1 110
2 1856 1 110
2 1857 1 111
2 1858 1 111
2 1859 1 112
2 1860 1 112
2 1861 1 112
2 1862 1 115
2 1863 1 115
2 1864 1 116
2 1865 1 116
2 1866 1 119
2 1867 1 119
2 1868 1 122
2 1869 1 122
2 1870 1 124
2 1871 1 124
2 1872 1 127
2 1873 1 127
2 1874 1 130
2 1875 1 130
2 1876 1 132
2 1877 1 132
2 1878 1 135
2 1879 1 135
2 1880 1 138
2 1881 1 138
2 1882 1 140
2 1883 1 140
2 1884 1 143
2 1885 1 143
2 1886 1 146
2 1887 1 146
2 1888 1 148
2 1889 1 148
2 1890 1 151
2 1891 1 151
2 1892 1 154
2 1893 1 154
2 1894 1 156
2 1895 1 156
2 1896 1 159
2 1897 1 159
2 1898 1 162
2 1899 1 162
2 1900 1 164
2 1901 1 164
2 1902 1 167
2 1903 1 167
2 1904 1 170
2 1905 1 170
2 1906 1 172
2 1907 1 172
2 1908 1 175
2 1909 1 175
2 1910 1 178
2 1911 1 178
2 1912 1 180
2 1913 1 180
2 1914 1 183
2 1915 1 183
2 1916 1 186
2 1917 1 186
2 1918 1 188
2 1919 1 188
2 1920 1 191
2 1921 1 191
2 1922 1 194
2 1923 1 194
2 1924 1 196
2 1925 1 196
2 1926 1 199
2 1927 1 199
2 1928 1 202
2 1929 1 202
2 1930 1 204
2 1931 1 204
2 1932 1 207
2 1933 1 207
2 1934 1 210
2 1935 1 210
2 1936 1 212
2 1937 1 212
2 1938 1 215
2 1939 1 215
2 1940 1 215
2 1941 1 216
2 1942 1 216
2 1943 1 216
2 1944 1 219
2 1945 1 219
2 1946 1 219
2 1947 1 220
2 1948 1 220
2 1949 1 221
2 1950 1 221
2 1951 1 222
2 1952 1 222
2 1953 1 222
2 1954 1 222
2 1955 1 223
2 1956 1 223
2 1957 1 224
2 1958 1 224
2 1959 1 224
2 1960 1 224
2 1961 1 225
2 1962 1 225
2 1963 1 231
2 1964 1 231
2 1965 1 231
2 1966 1 232
2 1967 1 232
2 1968 1 234
2 1969 1 234
2 1970 1 234
2 1971 1 236
2 1972 1 236
2 1973 1 236
2 1974 1 237
2 1975 1 237
2 1976 1 243
2 1977 1 243
2 1978 1 243
2 1979 1 243
2 1980 1 244
2 1981 1 244
2 1982 1 244
2 1983 1 246
2 1984 1 246
2 1985 1 246
2 1986 1 248
2 1987 1 248
2 1988 1 248
2 1989 1 249
2 1990 1 249
2 1991 1 255
2 1992 1 255
2 1993 1 255
2 1994 1 255
2 1995 1 256
2 1996 1 256
2 1997 1 256
2 1998 1 258
2 1999 1 258
2 2000 1 258
2 2001 1 260
2 2002 1 260
2 2003 1 260
2 2004 1 261
2 2005 1 261
2 2006 1 267
2 2007 1 267
2 2008 1 267
2 2009 1 267
2 2010 1 268
2 2011 1 268
2 2012 1 268
2 2013 1 270
2 2014 1 270
2 2015 1 270
2 2016 1 272
2 2017 1 272
2 2018 1 272
2 2019 1 273
2 2020 1 273
2 2021 1 279
2 2022 1 279
2 2023 1 279
2 2024 1 279
2 2025 1 280
2 2026 1 280
2 2027 1 280
2 2028 1 282
2 2029 1 282
2 2030 1 282
2 2031 1 284
2 2032 1 284
2 2033 1 284
2 2034 1 285
2 2035 1 285
2 2036 1 291
2 2037 1 291
2 2038 1 291
2 2039 1 291
2 2040 1 292
2 2041 1 292
2 2042 1 292
2 2043 1 294
2 2044 1 294
2 2045 1 294
2 2046 1 296
2 2047 1 296
2 2048 1 296
2 2049 1 297
2 2050 1 297
2 2051 1 303
2 2052 1 303
2 2053 1 303
2 2054 1 303
2 2055 1 304
2 2056 1 304
2 2057 1 304
2 2058 1 306
2 2059 1 306
2 2060 1 306
2 2061 1 308
2 2062 1 308
2 2063 1 308
2 2064 1 309
2 2065 1 309
2 2066 1 315
2 2067 1 315
2 2068 1 315
2 2069 1 315
2 2070 1 316
2 2071 1 316
2 2072 1 316
2 2073 1 318
2 2074 1 318
2 2075 1 318
2 2076 1 320
2 2077 1 320
2 2078 1 320
2 2079 1 321
2 2080 1 321
2 2081 1 327
2 2082 1 327
2 2083 1 327
2 2084 1 327
2 2085 1 328
2 2086 1 328
2 2087 1 328
2 2088 1 330
2 2089 1 330
2 2090 1 330
2 2091 1 332
2 2092 1 332
2 2093 1 332
2 2094 1 333
2 2095 1 333
2 2096 1 339
2 2097 1 339
2 2098 1 339
2 2099 1 339
2 2100 1 340
2 2101 1 340
2 2102 1 340
2 2103 1 342
2 2104 1 342
2 2105 1 342
2 2106 1 344
2 2107 1 344
2 2108 1 344
2 2109 1 345
2 2110 1 345
2 2111 1 351
2 2112 1 351
2 2113 1 351
2 2114 1 351
2 2115 1 352
2 2116 1 352
2 2117 1 352
2 2118 1 354
2 2119 1 354
2 2120 1 354
2 2121 1 356
2 2122 1 356
2 2123 1 356
2 2124 1 357
2 2125 1 357
2 2126 1 363
2 2127 1 363
2 2128 1 363
2 2129 1 363
2 2130 1 364
2 2131 1 364
2 2132 1 364
2 2133 1 366
2 2134 1 366
2 2135 1 366
2 2136 1 368
2 2137 1 368
2 2138 1 368
2 2139 1 369
2 2140 1 369
2 2141 1 375
2 2142 1 375
2 2143 1 375
2 2144 1 375
2 2145 1 376
2 2146 1 376
2 2147 1 376
2 2148 1 378
2 2149 1 378
2 2150 1 378
2 2151 1 380
2 2152 1 380
2 2153 1 380
2 2154 1 381
2 2155 1 381
2 2156 1 387
2 2157 1 387
2 2158 1 387
2 2159 1 387
2 2160 1 387
2 2161 1 388
2 2162 1 388
2 2163 1 388
2 2164 1 390
2 2165 1 390
2 2166 1 390
2 2167 1 392
2 2168 1 392
2 2169 1 392
2 2170 1 393
2 2171 1 393
2 2172 1 397
2 2173 1 397
2 2174 1 399
2 2175 1 399
2 2176 1 399
2 2177 1 400
2 2178 1 400
2 2179 1 400
2 2180 1 402
2 2181 1 402
2 2182 1 402
2 2183 1 404
2 2184 1 404
2 2185 1 404
2 2186 1 406
2 2187 1 406
2 2188 1 407
2 2189 1 407
2 2190 1 408
2 2191 1 408
2 2192 1 408
2 2193 1 409
2 2194 1 409
2 2195 1 409
2 2196 1 410
2 2197 1 410
2 2198 1 410
2 2199 1 412
2 2200 1 412
2 2201 1 413
2 2202 1 413
2 2203 1 413
2 2204 1 417
2 2205 1 417
2 2206 1 418
2 2207 1 418
2 2208 1 421
2 2209 1 421
2 2210 1 422
2 2211 1 422
2 2212 1 425
2 2213 1 425
2 2214 1 426
2 2215 1 426
2 2216 1 429
2 2217 1 429
2 2218 1 430
2 2219 1 430
2 2220 1 433
2 2221 1 433
2 2222 1 434
2 2223 1 434
2 2224 1 437
2 2225 1 437
2 2226 1 438
2 2227 1 438
2 2228 1 441
2 2229 1 441
2 2230 1 442
2 2231 1 442
2 2232 1 445
2 2233 1 445
2 2234 1 446
2 2235 1 446
2 2236 1 449
2 2237 1 449
2 2238 1 450
2 2239 1 450
2 2240 1 453
2 2241 1 453
2 2242 1 454
2 2243 1 454
2 2244 1 457
2 2245 1 457
2 2246 1 458
2 2247 1 458
2 2248 1 461
2 2249 1 461
2 2250 1 462
2 2251 1 462
2 2252 1 465
2 2253 1 465
2 2254 1 466
2 2255 1 466
2 2256 1 469
2 2257 1 469
2 2258 1 469
2 2259 1 470
2 2260 1 470
2 2261 1 470
2 2262 1 473
2 2263 1 473
2 2264 1 473
2 2265 1 474
2 2266 1 474
2 2267 1 475
2 2268 1 475
2 2269 1 475
2 2270 1 476
2 2271 1 476
2 2272 1 481
2 2273 1 481
2 2274 1 481
2 2275 1 482
2 2276 1 482
2 2277 1 483
2 2278 1 483
2 2279 1 483
2 2280 1 484
2 2281 1 484
2 2282 1 489
2 2283 1 489
2 2284 1 492
2 2285 1 492
2 2286 1 493
2 2287 1 493
2 2288 1 493
2 2289 1 494
2 2290 1 494
2 2291 1 499
2 2292 1 499
2 2293 1 499
2 2294 1 500
2 2295 1 500
2 2296 1 501
2 2297 1 501
2 2298 1 501
2 2299 1 502
2 2300 1 502
2 2301 1 507
2 2302 1 507
2 2303 1 507
2 2304 1 508
2 2305 1 508
2 2306 1 510
2 2307 1 510
2 2308 1 511
2 2309 1 511
2 2310 1 511
2 2311 1 512
2 2312 1 512
2 2313 1 517
2 2314 1 517
2 2315 1 517
2 2316 1 518
2 2317 1 518
2 2318 1 520
2 2319 1 520
2 2320 1 521
2 2321 1 521
2 2322 1 521
2 2323 1 522
2 2324 1 522
2 2325 1 527
2 2326 1 527
2 2327 1 527
2 2328 1 528
2 2329 1 528
2 2330 1 530
2 2331 1 530
2 2332 1 531
2 2333 1 531
2 2334 1 531
2 2335 1 532
2 2336 1 532
2 2337 1 537
2 2338 1 537
2 2339 1 537
2 2340 1 538
2 2341 1 538
2 2342 1 540
2 2343 1 540
2 2344 1 541
2 2345 1 541
2 2346 1 541
2 2347 1 542
2 2348 1 542
2 2349 1 547
2 2350 1 547
2 2351 1 547
2 2352 1 548
2 2353 1 548
2 2354 1 550
2 2355 1 550
2 2356 1 551
2 2357 1 551
2 2358 1 551
2 2359 1 552
2 2360 1 552
2 2361 1 557
2 2362 1 557
2 2363 1 557
2 2364 1 558
2 2365 1 558
2 2366 1 560
2 2367 1 560
2 2368 1 561
2 2369 1 561
2 2370 1 561
2 2371 1 562
2 2372 1 562
2 2373 1 567
2 2374 1 567
2 2375 1 567
2 2376 1 568
2 2377 1 568
2 2378 1 570
2 2379 1 570
2 2380 1 571
2 2381 1 571
2 2382 1 571
2 2383 1 572
2 2384 1 572
2 2385 1 577
2 2386 1 577
2 2387 1 577
2 2388 1 578
2 2389 1 578
2 2390 1 580
2 2391 1 580
2 2392 1 581
2 2393 1 581
2 2394 1 581
2 2395 1 582
2 2396 1 582
2 2397 1 587
2 2398 1 587
2 2399 1 587
2 2400 1 588
2 2401 1 588
2 2402 1 590
2 2403 1 590
2 2404 1 591
2 2405 1 591
2 2406 1 591
2 2407 1 592
2 2408 1 592
2 2409 1 597
2 2410 1 597
2 2411 1 597
2 2412 1 598
2 2413 1 598
2 2414 1 600
2 2415 1 600
2 2416 1 601
2 2417 1 601
2 2418 1 601
2 2419 1 602
2 2420 1 602
2 2421 1 607
2 2422 1 607
2 2423 1 607
2 2424 1 608
2 2425 1 608
2 2426 1 610
2 2427 1 610
2 2428 1 611
2 2429 1 611
2 2430 1 611
2 2431 1 612
2 2432 1 612
2 2433 1 617
2 2434 1 617
2 2435 1 617
2 2436 1 618
2 2437 1 618
2 2438 1 620
2 2439 1 620
2 2440 1 621
2 2441 1 621
2 2442 1 621
2 2443 1 622
2 2444 1 622
2 2445 1 624
2 2446 1 624
2 2447 1 627
2 2448 1 627
2 2449 1 627
2 2450 1 630
2 2451 1 630
2 2452 1 631
2 2453 1 631
2 2454 1 631
2 2455 1 632
2 2456 1 632
2 2457 1 633
2 2458 1 633
2 2459 1 633
2 2460 1 634
2 2461 1 634
2 2462 1 635
2 2463 1 635
2 2464 1 636
2 2465 1 636
2 2466 1 639
2 2467 1 639
2 2468 1 642
2 2469 1 642
2 2470 1 643
2 2471 1 643
2 2472 1 647
2 2473 1 647
2 2474 1 650
2 2475 1 650
2 2476 1 651
2 2477 1 651
2 2478 1 655
2 2479 1 655
2 2480 1 658
2 2481 1 658
2 2482 1 659
2 2483 1 659
2 2484 1 663
2 2485 1 663
2 2486 1 666
2 2487 1 666
2 2488 1 667
2 2489 1 667
2 2490 1 671
2 2491 1 671
2 2492 1 674
2 2493 1 674
2 2494 1 675
2 2495 1 675
2 2496 1 679
2 2497 1 679
2 2498 1 682
2 2499 1 682
2 2500 1 683
2 2501 1 683
2 2502 1 687
2 2503 1 687
2 2504 1 690
2 2505 1 690
2 2506 1 691
2 2507 1 691
2 2508 1 695
2 2509 1 695
2 2510 1 698
2 2511 1 698
2 2512 1 699
2 2513 1 699
2 2514 1 703
2 2515 1 703
2 2516 1 706
2 2517 1 706
2 2518 1 707
2 2519 1 707
2 2520 1 711
2 2521 1 711
2 2522 1 714
2 2523 1 714
2 2524 1 715
2 2525 1 715
2 2526 1 719
2 2527 1 719
2 2528 1 722
2 2529 1 722
2 2530 1 723
2 2531 1 723
2 2532 1 727
2 2533 1 727
2 2534 1 730
2 2535 1 730
2 2536 1 731
2 2537 1 731
2 2538 1 735
2 2539 1 735
2 2540 1 738
2 2541 1 738
2 2542 1 739
2 2543 1 739
2 2544 1 743
2 2545 1 743
2 2546 1 746
2 2547 1 746
2 2548 1 747
2 2549 1 747
2 2550 1 753
2 2551 1 753
2 2552 1 761
2 2553 1 761
2 2554 1 763
2 2555 1 763
2 2556 1 765
2 2557 1 765
2 2558 1 767
2 2559 1 767
2 2560 1 769
2 2561 1 769
2 2562 1 771
2 2563 1 771
2 2564 1 773
2 2565 1 773
2 2566 1 775
2 2567 1 775
2 2568 1 777
2 2569 1 777
2 2570 1 779
2 2571 1 779
2 2572 1 781
2 2573 1 781
2 2574 1 783
2 2575 1 783
2 2576 1 785
2 2577 1 785
2 2578 1 787
2 2579 1 787
2 2580 1 789
2 2581 1 789
2 2582 1 791
2 2583 1 791
2 2584 1 794
2 2585 1 794
2 2586 1 797
2 2587 1 797
2 2588 1 800
2 2589 1 800
2 2590 1 803
2 2591 1 803
2 2592 1 804
2 2593 1 804
2 2594 1 808
2 2595 1 808
2 2596 1 811
2 2597 1 811
2 2598 1 812
2 2599 1 812
2 2600 1 816
2 2601 1 816
2 2602 1 819
2 2603 1 819
2 2604 1 820
2 2605 1 820
2 2606 1 824
2 2607 1 824
2 2608 1 827
2 2609 1 827
2 2610 1 828
2 2611 1 828
2 2612 1 832
2 2613 1 832
2 2614 1 835
2 2615 1 835
2 2616 1 836
2 2617 1 836
2 2618 1 840
2 2619 1 840
2 2620 1 843
2 2621 1 843
2 2622 1 844
2 2623 1 844
2 2624 1 848
2 2625 1 848
2 2626 1 851
2 2627 1 851
2 2628 1 852
2 2629 1 852
2 2630 1 856
2 2631 1 856
2 2632 1 859
2 2633 1 859
2 2634 1 860
2 2635 1 860
2 2636 1 864
2 2637 1 864
2 2638 1 867
2 2639 1 867
2 2640 1 868
2 2641 1 868
2 2642 1 872
2 2643 1 872
2 2644 1 875
2 2645 1 875
2 2646 1 876
2 2647 1 876
2 2648 1 880
2 2649 1 880
2 2650 1 883
2 2651 1 883
2 2652 1 884
2 2653 1 884
2 2654 1 888
2 2655 1 888
2 2656 1 891
2 2657 1 891
2 2658 1 892
2 2659 1 892
2 2660 1 896
2 2661 1 896
2 2662 1 899
2 2663 1 899
2 2664 1 900
2 2665 1 900
2 2666 1 904
2 2667 1 904
2 2668 1 906
2 2669 1 906
2 2670 1 907
2 2671 1 907
2 2672 1 910
2 2673 1 910
2 2674 1 910
2 2675 1 910
2 2676 1 911
2 2677 1 911
2 2678 1 912
2 2679 1 912
2 2680 1 913
2 2681 1 913
2 2682 1 914
2 2683 1 914
2 2684 1 915
2 2685 1 915
2 2686 1 934
2 2687 1 934
2 2688 1 934
2 2689 1 935
2 2690 1 935
2 2691 1 938
2 2692 1 938
2 2693 1 938
2 2694 1 942
2 2695 1 942
2 2696 1 950
2 2697 1 950
2 2698 1 950
2 2699 1 951
2 2700 1 951
2 2701 1 954
2 2702 1 954
2 2703 1 962
2 2704 1 962
2 2705 1 966
2 2706 1 966
2 2707 1 966
2 2708 1 970
2 2709 1 970
2 2710 1 978
2 2711 1 978
2 2712 1 982
2 2713 1 982
2 2714 1 982
2 2715 1 983
2 2716 1 983
2 2717 1 986
2 2718 1 986
2 2719 1 994
2 2720 1 994
2 2721 1 998
2 2722 1 998
2 2723 1 998
2 2724 1 999
2 2725 1 999
2 2726 1 1002
2 2727 1 1002
2 2728 1 1010
2 2729 1 1010
2 2730 1 1014
2 2731 1 1014
2 2732 1 1014
2 2733 1 1015
2 2734 1 1015
2 2735 1 1018
2 2736 1 1018
2 2737 1 1026
2 2738 1 1026
2 2739 1 1030
2 2740 1 1030
2 2741 1 1030
2 2742 1 1034
2 2743 1 1034
2 2744 1 1044
2 2745 1 1044
2 2746 1 1044
2 2747 1 1045
2 2748 1 1045
2 2749 1 1048
2 2750 1 1048
2 2751 1 1052
2 2752 1 1052
2 2753 1 1056
2 2754 1 1056
2 2755 1 1062
2 2756 1 1062
2 2757 1 1068
2 2758 1 1068
2 2759 1 1072
2 2760 1 1072
2 2761 1 1085
2 2762 1 1085
2 2763 1 1091
2 2764 1 1091
2 2765 1 1092
2 2766 1 1092
2 2767 1 1101
2 2768 1 1101
2 2769 1 1107
2 2770 1 1107
2 2771 1 1117
2 2772 1 1117
2 2773 1 1123
2 2774 1 1123
2 2775 1 1133
2 2776 1 1133
2 2777 1 1139
2 2778 1 1139
2 2779 1 1140
2 2780 1 1140
2 2781 1 1149
2 2782 1 1149
2 2783 1 1155
2 2784 1 1155
2 2785 1 1169
2 2786 1 1169
2 2787 1 1189
2 2788 1 1189
2 2789 1 1190
2 2790 1 1190
2 2791 1 1193
2 2792 1 1193
2 2793 1 1194
2 2794 1 1194
2 2795 1 1197
2 2796 1 1197
2 2797 1 1198
2 2798 1 1198
2 2799 1 1201
2 2800 1 1201
2 2801 1 1202
2 2802 1 1202
2 2803 1 1205
2 2804 1 1205
2 2805 1 1206
2 2806 1 1206
2 2807 1 1209
2 2808 1 1209
2 2809 1 1210
2 2810 1 1210
2 2811 1 1213
2 2812 1 1213
2 2813 1 1214
2 2814 1 1214
2 2815 1 1217
2 2816 1 1217
2 2817 1 1218
2 2818 1 1218
2 2819 1 1221
2 2820 1 1221
2 2821 1 1222
2 2822 1 1222
2 2823 1 1225
2 2824 1 1225
2 2825 1 1226
2 2826 1 1226
2 2827 1 1229
2 2828 1 1229
2 2829 1 1230
2 2830 1 1230
2 2831 1 1233
2 2832 1 1233
2 2833 1 1234
2 2834 1 1234
2 2835 1 1237
2 2836 1 1237
2 2837 1 1238
2 2838 1 1238
2 2839 1 1243
2 2840 1 1243
2 2841 1 1243
2 2842 1 1244
2 2843 1 1244
2 2844 1 1249
2 2845 1 1249
2 2846 1 1249
2 2847 1 1250
2 2848 1 1250
2 2849 1 1252
2 2850 1 1252
2 2851 1 1257
2 2852 1 1257
2 2853 1 1257
2 2854 1 1258
2 2855 1 1258
2 2856 1 1263
2 2857 1 1263
2 2858 1 1263
2 2859 1 1264
2 2860 1 1264
2 2861 1 1266
2 2862 1 1266
2 2863 1 1271
2 2864 1 1271
2 2865 1 1271
2 2866 1 1272
2 2867 1 1272
2 2868 1 1274
2 2869 1 1274
2 2870 1 1279
2 2871 1 1279
2 2872 1 1279
2 2873 1 1280
2 2874 1 1280
2 2875 1 1282
2 2876 1 1282
2 2877 1 1287
2 2878 1 1287
2 2879 1 1287
2 2880 1 1288
2 2881 1 1288
2 2882 1 1290
2 2883 1 1290
2 2884 1 1295
2 2885 1 1295
2 2886 1 1295
2 2887 1 1296
2 2888 1 1296
2 2889 1 1298
2 2890 1 1298
2 2891 1 1303
2 2892 1 1303
2 2893 1 1303
2 2894 1 1304
2 2895 1 1304
2 2896 1 1306
2 2897 1 1306
2 2898 1 1311
2 2899 1 1311
2 2900 1 1311
2 2901 1 1312
2 2902 1 1312
2 2903 1 1314
2 2904 1 1314
2 2905 1 1319
2 2906 1 1319
2 2907 1 1319
2 2908 1 1320
2 2909 1 1320
2 2910 1 1322
2 2911 1 1322
2 2912 1 1327
2 2913 1 1327
2 2914 1 1327
2 2915 1 1328
2 2916 1 1328
2 2917 1 1330
2 2918 1 1330
2 2919 1 1335
2 2920 1 1335
2 2921 1 1335
2 2922 1 1336
2 2923 1 1336
2 2924 1 1338
2 2925 1 1338
2 2926 1 1343
2 2927 1 1343
2 2928 1 1344
2 2929 1 1344
2 2930 1 1346
2 2931 1 1346
2 2932 1 1347
2 2933 1 1347
2 2934 1 1348
2 2935 1 1348
2 2936 1 1351
2 2937 1 1351
2 2938 1 1354
2 2939 1 1354
2 2940 1 1355
2 2941 1 1355
2 2942 1 1359
2 2943 1 1359
2 2944 1 1362
2 2945 1 1362
2 2946 1 1363
2 2947 1 1363
2 2948 1 1367
2 2949 1 1367
2 2950 1 1370
2 2951 1 1370
2 2952 1 1371
2 2953 1 1371
2 2954 1 1375
2 2955 1 1375
2 2956 1 1378
2 2957 1 1378
2 2958 1 1379
2 2959 1 1379
2 2960 1 1383
2 2961 1 1383
2 2962 1 1386
2 2963 1 1386
2 2964 1 1387
2 2965 1 1387
2 2966 1 1391
2 2967 1 1391
2 2968 1 1394
2 2969 1 1394
2 2970 1 1395
2 2971 1 1395
2 2972 1 1399
2 2973 1 1399
2 2974 1 1402
2 2975 1 1402
2 2976 1 1403
2 2977 1 1403
2 2978 1 1407
2 2979 1 1407
2 2980 1 1410
2 2981 1 1410
2 2982 1 1411
2 2983 1 1411
2 2984 1 1415
2 2985 1 1415
2 2986 1 1418
2 2987 1 1418
2 2988 1 1419
2 2989 1 1419
2 2990 1 1423
2 2991 1 1423
2 2992 1 1426
2 2993 1 1426
2 2994 1 1427
2 2995 1 1427
2 2996 1 1431
2 2997 1 1431
2 2998 1 1434
2 2999 1 1434
2 3000 1 1435
2 3001 1 1435
2 3002 1 1439
2 3003 1 1439
2 3004 1 1442
2 3005 1 1442
2 3006 1 1443
2 3007 1 1443
2 3008 1 1447
2 3009 1 1447
2 3010 1 1448
2 3011 1 1448
2 3012 1 1453
2 3013 1 1453
2 3014 1 1453
2 3015 1 1454
2 3016 1 1454
2 3017 1 1456
2 3018 1 1456
2 3019 1 1459
2 3020 1 1459
2 3021 1 1462
2 3022 1 1462
2 3023 1 1465
2 3024 1 1465
2 3025 1 1469
2 3026 1 1469
2 3027 1 1473
2 3028 1 1473
2 3029 1 1477
2 3030 1 1477
2 3031 1 1485
2 3032 1 1485
2 3033 1 1489
2 3034 1 1489
2 3035 1 1497
2 3036 1 1497
2 3037 1 1501
2 3038 1 1501
2 3039 1 1509
2 3040 1 1509
2 3041 1 1517
2 3042 1 1517
2 3043 1 1525
2 3044 1 1525
2 3045 1 1531
2 3046 1 1531
2 3047 1 1543
2 3048 1 1543
2 3049 1 1547
2 3050 1 1547
2 3051 1 1563
2 3052 1 1563
2 3053 1 1575
2 3054 1 1575
2 3055 1 1587
2 3056 1 1587
2 3057 1 1599
2 3058 1 1599
2 3059 1 1607
2 3060 1 1607
2 3061 1 1619
2 3062 1 1619
2 3063 1 1627
2 3064 1 1627
2 3065 1 1635
2 3066 1 1635
2 3067 1 1639
2 3068 1 1639
2 3069 1 1643
2 3070 1 1643
2 3071 1 1643
2 3072 1 1644
2 3073 1 1644
2 3074 1 1644
2 3075 1 1649
2 3076 1 1649
2 3077 1 1652
2 3078 1 1652
2 3079 1 1655
2 3080 1 1655
2 3081 1 1658
2 3082 1 1658
2 3083 1 1664
2 3084 1 1664
2 3085 1 1667
2 3086 1 1667
2 3087 1 1668
2 3088 1 1668
2 3089 1 1671
2 3090 1 1671
2 3091 1 1674
2 3092 1 1674
2 3093 1 1677
2 3094 1 1677
2 3095 1 1680
2 3096 1 1680
2 3097 1 1682
2 3098 1 1682
2 3099 1 1693
2 3100 1 1693
2 3101 1 1699
2 3102 1 1699
2 3103 1 1702
2 3104 1 1702
2 3105 1 1704
2 3106 1 1704
0 50 5 1 1 49
0 51 5 1 1 1721
0 52 5 1 1 1723
0 53 5 1 1 1725
0 54 5 1 1 1727
0 55 5 1 1 1729
0 56 5 1 1 1731
0 57 5 1 1 1733
0 58 5 1 1 1735
0 59 5 1 1 1737
0 60 5 1 1 1739
0 61 5 1 1 1741
0 62 5 1 1 1743
0 63 5 1 1 1745
0 64 5 1 1 1747
0 65 5 1 1 1749
0 66 5 1 1 1751
0 67 5 1 1 1753
0 68 5 1 1 1755
0 69 5 2 1 1757
0 70 5 2 1 1759
0 71 5 2 1 1761
0 72 5 2 1 1763
0 73 5 2 1 1765
0 74 5 2 1 1767
0 75 5 2 1 1769
0 76 5 2 1 1771
0 77 5 2 1 1773
0 78 5 2 1 1775
0 79 5 2 1 1777
0 80 5 2 1 1779
0 81 5 1 1 1781
0 82 5 1 1 1783
0 83 5 1 1 1785
0 84 5 1 1 1787
0 85 5 1 1 1789
0 86 5 1 1 1791
0 87 5 1 1 1793
0 88 5 1 1 1795
0 89 5 1 1 1797
0 90 5 1 1 1799
0 91 5 1 1 1801
0 92 5 1 1 1803
0 93 5 1 1 1805
0 94 5 1 1 1807
0 95 5 1 1 1809
0 96 5 1 1 1811
0 97 5 1 1 1813
0 98 5 1 1 1815
0 99 7 2 2 65 81
0 100 5 2 1 1841
0 101 7 2 2 1750 1782
0 102 5 2 1 1845
0 103 7 1 2 52 68
0 104 5 2 1 103
0 105 7 1 2 1724 1756
0 106 5 2 1 105
0 107 7 1 2 51 67
0 108 5 2 1 107
0 109 7 1 2 1722 1754
0 110 5 2 1 109
0 111 7 2 2 1720 1752
0 112 5 3 1 1857
0 113 7 1 2 1855 1859
0 114 5 1 1 113
0 115 7 2 2 1853 114
0 116 5 2 1 1862
0 117 7 1 2 1851 1864
0 118 5 1 1 117
0 119 7 2 2 1849 118
0 120 5 1 1 1866
0 121 7 1 2 53 120
0 122 5 2 1 121
0 123 7 1 2 1726 1867
0 124 5 2 1 123
0 125 7 1 2 1817 1870
0 126 5 1 1 125
0 127 7 2 2 1868 126
0 128 5 1 1 1872
0 129 7 1 2 54 128
0 130 5 2 1 129
0 131 7 1 2 1728 1873
0 132 5 2 1 131
0 133 7 1 2 1819 1876
0 134 5 1 1 133
0 135 7 2 2 1874 134
0 136 5 1 1 1878
0 137 7 1 2 55 136
0 138 5 2 1 137
0 139 7 1 2 1730 1879
0 140 5 2 1 139
0 141 7 1 2 1821 1882
0 142 5 1 1 141
0 143 7 2 2 1880 142
0 144 5 1 1 1884
0 145 7 1 2 56 144
0 146 5 2 1 145
0 147 7 1 2 1732 1885
0 148 5 2 1 147
0 149 7 1 2 1823 1888
0 150 5 1 1 149
0 151 7 2 2 1886 150
0 152 5 1 1 1890
0 153 7 1 2 57 152
0 154 5 2 1 153
0 155 7 1 2 1734 1891
0 156 5 2 1 155
0 157 7 1 2 1825 1894
0 158 5 1 1 157
0 159 7 2 2 1892 158
0 160 5 1 1 1896
0 161 7 1 2 58 160
0 162 5 2 1 161
0 163 7 1 2 1736 1897
0 164 5 2 1 163
0 165 7 1 2 1827 1900
0 166 5 1 1 165
0 167 7 2 2 1898 166
0 168 5 1 1 1902
0 169 7 1 2 59 168
0 170 5 2 1 169
0 171 7 1 2 1738 1903
0 172 5 2 1 171
0 173 7 1 2 1829 1906
0 174 5 1 1 173
0 175 7 2 2 1904 174
0 176 5 1 1 1908
0 177 7 1 2 60 176
0 178 5 2 1 177
0 179 7 1 2 1740 1909
0 180 5 2 1 179
0 181 7 1 2 1831 1912
0 182 5 1 1 181
0 183 7 2 2 1910 182
0 184 5 1 1 1914
0 185 7 1 2 61 184
0 186 5 2 1 185
0 187 7 1 2 1742 1915
0 188 5 2 1 187
0 189 7 1 2 1833 1918
0 190 5 1 1 189
0 191 7 2 2 1916 190
0 192 5 1 1 1920
0 193 7 1 2 62 192
0 194 5 2 1 193
0 195 7 1 2 1744 1921
0 196 5 2 1 195
0 197 7 1 2 1835 1924
0 198 5 1 1 197
0 199 7 2 2 1922 198
0 200 5 1 1 1926
0 201 7 1 2 63 200
0 202 5 2 1 201
0 203 7 1 2 1746 1927
0 204 5 2 1 203
0 205 7 1 2 1837 1930
0 206 5 1 1 205
0 207 7 2 2 1928 206
0 208 5 1 1 1932
0 209 7 1 2 64 208
0 210 5 2 1 209
0 211 7 1 2 1748 1933
0 212 5 2 1 211
0 213 7 1 2 1839 1936
0 214 5 1 1 213
0 215 7 3 2 1934 214
0 216 5 3 1 1938
0 217 7 1 2 1847 1941
0 218 5 1 1 217
0 219 7 3 2 1843 218
0 220 5 2 1 1944
0 221 7 2 2 98 1945
0 222 5 4 1 1949
0 223 7 2 2 1816 1947
0 224 5 4 1 1955
0 225 7 2 2 1844 1848
0 226 5 1 1 1961
0 227 7 1 2 1939 226
0 228 5 1 1 227
0 229 7 1 2 1942 1962
0 230 5 1 1 229
0 231 7 3 2 228 230
0 232 5 2 1 1963
0 233 7 1 2 97 1966
0 234 5 3 1 233
0 235 7 1 2 1814 1964
0 236 5 3 1 235
0 237 7 2 2 1935 1937
0 238 5 1 1 1974
0 239 7 1 2 1780 1975
0 240 5 1 1 239
0 241 7 1 2 1840 238
0 242 5 1 1 241
0 243 7 4 2 240 242
0 244 5 3 1 1976
0 245 7 1 2 96 1977
0 246 5 3 1 245
0 247 7 1 2 1812 1980
0 248 5 3 1 247
0 249 7 2 2 1929 1931
0 250 5 1 1 1989
0 251 7 1 2 1778 1990
0 252 5 1 1 251
0 253 7 1 2 1838 250
0 254 5 1 1 253
0 255 7 4 2 252 254
0 256 5 3 1 1991
0 257 7 1 2 95 1992
0 258 5 3 1 257
0 259 7 1 2 1810 1995
0 260 5 3 1 259
0 261 7 2 2 1923 1925
0 262 5 1 1 2004
0 263 7 1 2 1776 2005
0 264 5 1 1 263
0 265 7 1 2 1836 262
0 266 5 1 1 265
0 267 7 4 2 264 266
0 268 5 3 1 2006
0 269 7 1 2 94 2007
0 270 5 3 1 269
0 271 7 1 2 1808 2010
0 272 5 3 1 271
0 273 7 2 2 1917 1919
0 274 5 1 1 2019
0 275 7 1 2 1774 2020
0 276 5 1 1 275
0 277 7 1 2 1834 274
0 278 5 1 1 277
0 279 7 4 2 276 278
0 280 5 3 1 2021
0 281 7 1 2 93 2022
0 282 5 3 1 281
0 283 7 1 2 1806 2025
0 284 5 3 1 283
0 285 7 2 2 1911 1913
0 286 5 1 1 2034
0 287 7 1 2 1772 2035
0 288 5 1 1 287
0 289 7 1 2 1832 286
0 290 5 1 1 289
0 291 7 4 2 288 290
0 292 5 3 1 2036
0 293 7 1 2 92 2037
0 294 5 3 1 293
0 295 7 1 2 1804 2040
0 296 5 3 1 295
0 297 7 2 2 1905 1907
0 298 5 1 1 2049
0 299 7 1 2 1770 2050
0 300 5 1 1 299
0 301 7 1 2 1830 298
0 302 5 1 1 301
0 303 7 4 2 300 302
0 304 5 3 1 2051
0 305 7 1 2 91 2052
0 306 5 3 1 305
0 307 7 1 2 1802 2055
0 308 5 3 1 307
0 309 7 2 2 1899 1901
0 310 5 1 1 2064
0 311 7 1 2 1768 2065
0 312 5 1 1 311
0 313 7 1 2 1828 310
0 314 5 1 1 313
0 315 7 4 2 312 314
0 316 5 3 1 2066
0 317 7 1 2 90 2067
0 318 5 3 1 317
0 319 7 1 2 1800 2070
0 320 5 3 1 319
0 321 7 2 2 1893 1895
0 322 5 1 1 2079
0 323 7 1 2 1766 2080
0 324 5 1 1 323
0 325 7 1 2 1826 322
0 326 5 1 1 325
0 327 7 4 2 324 326
0 328 5 3 1 2081
0 329 7 1 2 89 2082
0 330 5 3 1 329
0 331 7 1 2 1798 2085
0 332 5 3 1 331
0 333 7 2 2 1887 1889
0 334 5 1 1 2094
0 335 7 1 2 1764 2095
0 336 5 1 1 335
0 337 7 1 2 1824 334
0 338 5 1 1 337
0 339 7 4 2 336 338
0 340 5 3 1 2096
0 341 7 1 2 88 2097
0 342 5 3 1 341
0 343 7 1 2 1796 2100
0 344 5 3 1 343
0 345 7 2 2 1881 1883
0 346 5 1 1 2109
0 347 7 1 2 1762 2110
0 348 5 1 1 347
0 349 7 1 2 1822 346
0 350 5 1 1 349
0 351 7 4 2 348 350
0 352 5 3 1 2111
0 353 7 1 2 87 2112
0 354 5 3 1 353
0 355 7 1 2 1794 2115
0 356 5 3 1 355
0 357 7 2 2 1875 1877
0 358 5 1 1 2124
0 359 7 1 2 1760 2125
0 360 5 1 1 359
0 361 7 1 2 1820 358
0 362 5 1 1 361
0 363 7 4 2 360 362
0 364 5 3 1 2126
0 365 7 1 2 86 2127
0 366 5 3 1 365
0 367 7 1 2 1792 2130
0 368 5 3 1 367
0 369 7 2 2 1869 1871
0 370 5 1 1 2139
0 371 7 1 2 1758 2140
0 372 5 1 1 371
0 373 7 1 2 1818 370
0 374 5 1 1 373
0 375 7 4 2 372 374
0 376 5 3 1 2141
0 377 7 1 2 85 2142
0 378 5 3 1 377
0 379 7 1 2 1790 2145
0 380 5 3 1 379
0 381 7 2 2 1850 1852
0 382 5 1 1 2154
0 383 7 1 2 1863 382
0 384 5 1 1 383
0 385 7 1 2 1865 2155
0 386 5 1 1 385
0 387 7 5 2 384 386
0 388 5 3 1 2156
0 389 7 1 2 84 2161
0 390 5 3 1 389
0 391 7 1 2 1788 2157
0 392 5 3 1 391
0 393 7 2 2 1854 1856
0 394 5 1 1 2170
0 395 7 1 2 1858 394
0 396 5 1 1 395
0 397 7 2 2 1860 2171
0 398 5 1 1 2172
0 399 7 3 2 396 398
0 400 5 3 1 2174
0 401 7 1 2 1786 2175
0 402 5 3 1 401
0 403 7 1 2 83 2177
0 404 5 3 1 403
0 405 7 1 2 50 66
0 406 5 2 1 405
0 407 7 2 2 1861 2186
0 408 5 3 1 2188
0 409 7 3 2 1784 2190
0 410 5 3 1 2193
0 411 7 1 2 2183 2194
0 412 5 2 1 411
0 413 7 3 2 2180 2199
0 414 5 1 1 2201
0 415 7 1 2 2167 2202
0 416 5 1 1 415
0 417 7 2 2 2164 416
0 418 5 2 1 2204
0 419 7 1 2 2151 2206
0 420 5 1 1 419
0 421 7 2 2 2148 420
0 422 5 2 1 2208
0 423 7 1 2 2136 2210
0 424 5 1 1 423
0 425 7 2 2 2133 424
0 426 5 2 1 2212
0 427 7 1 2 2121 2214
0 428 5 1 1 427
0 429 7 2 2 2118 428
0 430 5 2 1 2216
0 431 7 1 2 2106 2218
0 432 5 1 1 431
0 433 7 2 2 2103 432
0 434 5 2 1 2220
0 435 7 1 2 2091 2222
0 436 5 1 1 435
0 437 7 2 2 2088 436
0 438 5 2 1 2224
0 439 7 1 2 2076 2226
0 440 5 1 1 439
0 441 7 2 2 2073 440
0 442 5 2 1 2228
0 443 7 1 2 2061 2230
0 444 5 1 1 443
0 445 7 2 2 2058 444
0 446 5 2 1 2232
0 447 7 1 2 2046 2234
0 448 5 1 1 447
0 449 7 2 2 2043 448
0 450 5 2 1 2236
0 451 7 1 2 2031 2238
0 452 5 1 1 451
0 453 7 2 2 2028 452
0 454 5 2 1 2240
0 455 7 1 2 2016 2242
0 456 5 1 1 455
0 457 7 2 2 2013 456
0 458 5 2 1 2244
0 459 7 1 2 2001 2246
0 460 5 1 1 459
0 461 7 2 2 1998 460
0 462 5 2 1 2248
0 463 7 1 2 1986 2250
0 464 5 1 1 463
0 465 7 2 2 1983 464
0 466 5 2 1 2252
0 467 7 1 2 1971 2254
0 468 5 1 1 467
0 469 7 3 2 1968 468
0 470 5 3 1 2256
0 471 7 1 2 1957 2259
0 472 5 1 1 471
0 473 7 3 2 1951 472
0 474 5 2 1 2262
0 475 7 3 2 1984 1987
0 476 5 2 1 2267
0 477 7 1 2 2249 2270
0 478 5 1 1 477
0 479 7 1 2 2251 2268
0 480 5 1 1 479
0 481 7 3 2 478 480
0 482 5 2 1 2272
0 483 7 3 2 1952 1958
0 484 5 2 1 2277
0 485 7 1 2 2257 2280
0 486 5 1 1 485
0 487 7 1 2 2260 2278
0 488 5 1 1 487
0 489 7 2 2 486 488
0 490 5 1 1 2282
0 491 7 1 2 2273 2283
0 492 5 2 1 491
0 493 7 3 2 1969 1972
0 494 5 2 1 2286
0 495 7 1 2 2253 2289
0 496 5 1 1 495
0 497 7 1 2 2255 2287
0 498 5 1 1 497
0 499 7 3 2 496 498
0 500 5 2 1 2291
0 501 7 3 2 1999 2002
0 502 5 2 1 2296
0 503 7 1 2 2245 2299
0 504 5 1 1 503
0 505 7 1 2 2247 2297
0 506 5 1 1 505
0 507 7 3 2 504 506
0 508 5 2 1 2301
0 509 7 1 2 2292 2302
0 510 5 2 1 509
0 511 7 3 2 2014 2017
0 512 5 2 1 2308
0 513 7 1 2 2241 2311
0 514 5 1 1 513
0 515 7 1 2 2243 2309
0 516 5 1 1 515
0 517 7 3 2 514 516
0 518 5 2 1 2313
0 519 7 1 2 2274 2314
0 520 5 2 1 519
0 521 7 3 2 2029 2032
0 522 5 2 1 2320
0 523 7 1 2 2237 2323
0 524 5 1 1 523
0 525 7 1 2 2239 2321
0 526 5 1 1 525
0 527 7 3 2 524 526
0 528 5 2 1 2325
0 529 7 1 2 2303 2326
0 530 5 2 1 529
0 531 7 3 2 2044 2047
0 532 5 2 1 2332
0 533 7 1 2 2233 2335
0 534 5 1 1 533
0 535 7 1 2 2235 2333
0 536 5 1 1 535
0 537 7 3 2 534 536
0 538 5 2 1 2337
0 539 7 1 2 2315 2338
0 540 5 2 1 539
0 541 7 3 2 2059 2062
0 542 5 2 1 2344
0 543 7 1 2 2229 2347
0 544 5 1 1 543
0 545 7 1 2 2231 2345
0 546 5 1 1 545
0 547 7 3 2 544 546
0 548 5 2 1 2349
0 549 7 1 2 2327 2350
0 550 5 2 1 549
0 551 7 3 2 2074 2077
0 552 5 2 1 2356
0 553 7 1 2 2225 2359
0 554 5 1 1 553
0 555 7 1 2 2227 2357
0 556 5 1 1 555
0 557 7 3 2 554 556
0 558 5 2 1 2361
0 559 7 1 2 2339 2362
0 560 5 2 1 559
0 561 7 3 2 2089 2092
0 562 5 2 1 2368
0 563 7 1 2 2221 2371
0 564 5 1 1 563
0 565 7 1 2 2223 2369
0 566 5 1 1 565
0 567 7 3 2 564 566
0 568 5 2 1 2373
0 569 7 1 2 2351 2374
0 570 5 2 1 569
0 571 7 3 2 2104 2107
0 572 5 2 1 2380
0 573 7 1 2 2217 2383
0 574 5 1 1 573
0 575 7 1 2 2219 2381
0 576 5 1 1 575
0 577 7 3 2 574 576
0 578 5 2 1 2385
0 579 7 1 2 2363 2386
0 580 5 2 1 579
0 581 7 3 2 2119 2122
0 582 5 2 1 2392
0 583 7 1 2 2213 2395
0 584 5 1 1 583
0 585 7 1 2 2215 2393
0 586 5 1 1 585
0 587 7 3 2 584 586
0 588 5 2 1 2397
0 589 7 1 2 2375 2398
0 590 5 2 1 589
0 591 7 3 2 2134 2137
0 592 5 2 1 2404
0 593 7 1 2 2209 2407
0 594 5 1 1 593
0 595 7 1 2 2211 2405
0 596 5 1 1 595
0 597 7 3 2 594 596
0 598 5 2 1 2409
0 599 7 1 2 2387 2410
0 600 5 2 1 599
0 601 7 3 2 2149 2152
0 602 5 2 1 2416
0 603 7 1 2 2205 2419
0 604 5 1 1 603
0 605 7 1 2 2207 2417
0 606 5 1 1 605
0 607 7 3 2 604 606
0 608 5 2 1 2421
0 609 7 1 2 2399 2422
0 610 5 2 1 609
0 611 7 3 2 2165 2168
0 612 5 2 1 2428
0 613 7 1 2 414 2429
0 614 5 1 1 613
0 615 7 1 2 2203 2431
0 616 5 1 1 615
0 617 7 3 2 614 616
0 618 5 2 1 2433
0 619 7 1 2 2411 2436
0 620 5 2 1 619
0 621 7 3 2 2181 2184
0 622 5 2 1 2440
0 623 7 1 2 2195 2443
0 624 5 2 1 623
0 625 7 1 2 2196 2441
0 626 5 1 1 625
0 627 7 3 2 2445 626
0 628 5 1 1 2447
0 629 7 1 2 2423 2448
0 630 5 2 1 629
0 631 7 3 2 82 2189
0 632 5 2 1 2452
0 633 7 3 2 2197 2455
0 634 5 2 1 2457
0 635 7 2 2 2437 2460
0 636 5 2 1 2462
0 637 7 1 2 2424 628
0 638 5 1 1 637
0 639 7 2 2 2450 638
0 640 5 1 1 2466
0 641 7 1 2 2463 2467
0 642 5 2 1 641
0 643 7 2 2 2451 2468
0 644 5 1 1 2470
0 645 7 1 2 2412 2434
0 646 5 1 1 645
0 647 7 2 2 2438 646
0 648 5 1 1 2472
0 649 7 1 2 644 2473
0 650 5 2 1 649
0 651 7 2 2 2439 2474
0 652 5 1 1 2476
0 653 7 1 2 2400 2425
0 654 5 1 1 653
0 655 7 2 2 2426 654
0 656 5 1 1 2478
0 657 7 1 2 652 2479
0 658 5 2 1 657
0 659 7 2 2 2427 2480
0 660 5 1 1 2482
0 661 7 1 2 2388 2413
0 662 5 1 1 661
0 663 7 2 2 2414 662
0 664 5 1 1 2484
0 665 7 1 2 660 2485
0 666 5 2 1 665
0 667 7 2 2 2415 2486
0 668 5 1 1 2488
0 669 7 1 2 2376 2401
0 670 5 1 1 669
0 671 7 2 2 2402 670
0 672 5 1 1 2490
0 673 7 1 2 668 2491
0 674 5 2 1 673
0 675 7 2 2 2403 2492
0 676 5 1 1 2494
0 677 7 1 2 2364 2389
0 678 5 1 1 677
0 679 7 2 2 2390 678
0 680 5 1 1 2496
0 681 7 1 2 676 2497
0 682 5 2 1 681
0 683 7 2 2 2391 2498
0 684 5 1 1 2500
0 685 7 1 2 2352 2377
0 686 5 1 1 685
0 687 7 2 2 2378 686
0 688 5 1 1 2502
0 689 7 1 2 684 2503
0 690 5 2 1 689
0 691 7 2 2 2379 2504
0 692 5 1 1 2506
0 693 7 1 2 2340 2365
0 694 5 1 1 693
0 695 7 2 2 2366 694
0 696 5 1 1 2508
0 697 7 1 2 692 2509
0 698 5 2 1 697
0 699 7 2 2 2367 2510
0 700 5 1 1 2512
0 701 7 1 2 2328 2353
0 702 5 1 1 701
0 703 7 2 2 2354 702
0 704 5 1 1 2514
0 705 7 1 2 700 2515
0 706 5 2 1 705
0 707 7 2 2 2355 2516
0 708 5 1 1 2518
0 709 7 1 2 2316 2341
0 710 5 1 1 709
0 711 7 2 2 2342 710
0 712 5 1 1 2520
0 713 7 1 2 708 2521
0 714 5 2 1 713
0 715 7 2 2 2343 2522
0 716 5 1 1 2524
0 717 7 1 2 2304 2329
0 718 5 1 1 717
0 719 7 2 2 2330 718
0 720 5 1 1 2526
0 721 7 1 2 716 2527
0 722 5 2 1 721
0 723 7 2 2 2331 2528
0 724 5 1 1 2530
0 725 7 1 2 2275 2317
0 726 5 1 1 725
0 727 7 2 2 2318 726
0 728 5 1 1 2532
0 729 7 1 2 724 2533
0 730 5 2 1 729
0 731 7 2 2 2319 2534
0 732 5 1 1 2536
0 733 7 1 2 2294 2305
0 734 5 1 1 733
0 735 7 2 2 2306 734
0 736 5 1 1 2538
0 737 7 1 2 732 2539
0 738 5 2 1 737
0 739 7 2 2 2307 2540
0 740 5 1 1 2542
0 741 7 1 2 2276 490
0 742 5 1 1 741
0 743 7 2 2 2284 742
0 744 5 1 1 2544
0 745 7 1 2 740 2545
0 746 5 2 1 745
0 747 7 2 2 2285 2546
0 748 5 1 1 2548
0 749 7 1 2 2263 2293
0 750 5 1 1 749
0 751 7 1 2 2265 2295
0 752 5 1 1 751
0 753 7 2 2 750 752
0 754 5 1 1 2550
0 755 7 1 2 748 2551
0 756 5 1 1 755
0 757 7 1 2 1950 2261
0 758 5 1 1 757
0 759 7 1 2 1956 2258
0 760 5 1 1 759
0 761 7 2 2 758 760
0 762 5 1 1 2552
0 763 7 2 2 756 2553
0 764 7 1 2 1846 1940
0 765 5 2 1 764
0 766 7 1 2 1967 1978
0 767 5 2 1 766
0 768 7 1 2 1979 1993
0 769 5 2 1 768
0 770 7 1 2 1994 2008
0 771 5 2 1 770
0 772 7 1 2 2009 2023
0 773 5 2 1 772
0 774 7 1 2 2024 2038
0 775 5 2 1 774
0 776 7 1 2 2039 2053
0 777 5 2 1 776
0 778 7 1 2 2054 2068
0 779 5 2 1 778
0 780 7 1 2 2069 2083
0 781 5 2 1 780
0 782 7 1 2 2084 2098
0 783 5 2 1 782
0 784 7 1 2 2099 2113
0 785 5 2 1 784
0 786 7 1 2 2114 2128
0 787 5 2 1 786
0 788 7 1 2 2129 2143
0 789 5 2 1 788
0 790 7 1 2 2144 2162
0 791 5 2 1 790
0 792 7 1 2 2146 2158
0 793 5 1 1 792
0 794 7 2 2 2582 793
0 795 5 1 1 2584
0 796 7 1 2 2173 2187
0 797 5 2 1 796
0 798 7 1 2 2159 2586
0 799 5 1 1 798
0 800 7 2 2 2178 799
0 801 5 1 1 2588
0 802 7 1 2 2585 2589
0 803 5 2 1 802
0 804 7 2 2 2583 2590
0 805 5 1 1 2592
0 806 7 1 2 2131 2147
0 807 5 1 1 806
0 808 7 2 2 2580 807
0 809 5 1 1 2594
0 810 7 1 2 805 2595
0 811 5 2 1 810
0 812 7 2 2 2581 2596
0 813 5 1 1 2598
0 814 7 1 2 2116 2132
0 815 5 1 1 814
0 816 7 2 2 2578 815
0 817 5 1 1 2600
0 818 7 1 2 813 2601
0 819 5 2 1 818
0 820 7 2 2 2579 2602
0 821 5 1 1 2604
0 822 7 1 2 2101 2117
0 823 5 1 1 822
0 824 7 2 2 2576 823
0 825 5 1 1 2606
0 826 7 1 2 821 2607
0 827 5 2 1 826
0 828 7 2 2 2577 2608
0 829 5 1 1 2610
0 830 7 1 2 2086 2102
0 831 5 1 1 830
0 832 7 2 2 2574 831
0 833 5 1 1 2612
0 834 7 1 2 829 2613
0 835 5 2 1 834
0 836 7 2 2 2575 2614
0 837 5 1 1 2616
0 838 7 1 2 2071 2087
0 839 5 1 1 838
0 840 7 2 2 2572 839
0 841 5 1 1 2618
0 842 7 1 2 837 2619
0 843 5 2 1 842
0 844 7 2 2 2573 2620
0 845 5 1 1 2622
0 846 7 1 2 2056 2072
0 847 5 1 1 846
0 848 7 2 2 2570 847
0 849 5 1 1 2624
0 850 7 1 2 845 2625
0 851 5 2 1 850
0 852 7 2 2 2571 2626
0 853 5 1 1 2628
0 854 7 1 2 2041 2057
0 855 5 1 1 854
0 856 7 2 2 2568 855
0 857 5 1 1 2630
0 858 7 1 2 853 2631
0 859 5 2 1 858
0 860 7 2 2 2569 2632
0 861 5 1 1 2634
0 862 7 1 2 2026 2042
0 863 5 1 1 862
0 864 7 2 2 2566 863
0 865 5 1 1 2636
0 866 7 1 2 861 2637
0 867 5 2 1 866
0 868 7 2 2 2567 2638
0 869 5 1 1 2640
0 870 7 1 2 2011 2027
0 871 5 1 1 870
0 872 7 2 2 2564 871
0 873 5 1 1 2642
0 874 7 1 2 869 2643
0 875 5 2 1 874
0 876 7 2 2 2565 2644
0 877 5 1 1 2646
0 878 7 1 2 1996 2012
0 879 5 1 1 878
0 880 7 2 2 2562 879
0 881 5 1 1 2648
0 882 7 1 2 877 2649
0 883 5 2 1 882
0 884 7 2 2 2563 2650
0 885 5 1 1 2652
0 886 7 1 2 1981 1997
0 887 5 1 1 886
0 888 7 2 2 2560 887
0 889 5 1 1 2654
0 890 7 1 2 885 2655
0 891 5 2 1 890
0 892 7 2 2 2561 2656
0 893 5 1 1 2658
0 894 7 1 2 1965 1982
0 895 5 1 1 894
0 896 7 2 2 2558 895
0 897 5 1 1 2660
0 898 7 1 2 893 2661
0 899 5 2 1 898
0 900 7 2 2 2559 2662
0 901 5 1 1 2664
0 902 7 1 2 1842 1943
0 903 5 1 1 902
0 904 7 2 2 2556 903
0 905 5 1 1 2666
0 906 7 2 2 901 2667
0 907 5 2 1 2668
0 908 7 1 2 1946 2669
0 909 5 1 1 908
0 910 7 4 2 2557 909
0 911 5 2 1 2672
0 912 7 2 2 2549 754
0 913 5 2 1 2678
0 914 7 2 2 1948 2670
0 915 5 2 1 2682
0 916 7 1 2 2679 2684
0 917 5 1 1 916
0 918 7 1 2 2673 917
0 919 5 1 1 918
0 920 7 1 2 2554 919
0 921 5 1 1 920
0 922 7 1 2 762 2680
0 923 5 1 1 922
0 924 7 1 2 2676 923
0 925 5 1 1 924
0 926 7 1 2 2681 2683
0 927 5 1 1 926
0 928 7 1 2 2555 927
0 929 5 1 1 928
0 930 7 1 2 925 929
0 931 5 1 1 930
0 932 7 1 2 2665 905
0 933 5 1 1 932
0 934 7 3 2 2671 933
0 935 5 2 1 2686
0 936 7 1 2 2659 897
0 937 5 1 1 936
0 938 7 3 2 2663 937
0 939 5 1 1 2691
0 940 7 1 2 2537 736
0 941 5 1 1 940
0 942 7 2 2 2541 941
0 943 5 1 1 2694
0 944 7 1 2 939 2695
0 945 5 1 1 944
0 946 7 1 2 2692 943
0 947 5 1 1 946
0 948 7 1 2 2653 889
0 949 5 1 1 948
0 950 7 3 2 2657 949
0 951 5 2 1 2696
0 952 7 1 2 2531 728
0 953 5 1 1 952
0 954 7 2 2 2535 953
0 955 5 1 1 2701
0 956 7 1 2 2699 2702
0 957 5 1 1 956
0 958 7 1 2 2697 955
0 959 5 1 1 958
0 960 7 1 2 2525 720
0 961 5 1 1 960
0 962 7 2 2 2529 961
0 963 5 1 1 2703
0 964 7 1 2 2641 873
0 965 5 1 1 964
0 966 7 3 2 2645 965
0 967 5 1 1 2705
0 968 7 1 2 2519 712
0 969 5 1 1 968
0 970 7 2 2 2523 969
0 971 5 1 1 2708
0 972 7 1 2 967 2709
0 973 5 1 1 972
0 974 7 1 2 2706 971
0 975 5 1 1 974
0 976 7 1 2 2513 704
0 977 5 1 1 976
0 978 7 2 2 2517 977
0 979 5 1 1 2710
0 980 7 1 2 2629 857
0 981 5 1 1 980
0 982 7 3 2 2633 981
0 983 5 2 1 2712
0 984 7 1 2 2507 696
0 985 5 1 1 984
0 986 7 2 2 2511 985
0 987 5 1 1 2717
0 988 7 1 2 2715 2718
0 989 5 1 1 988
0 990 7 1 2 2713 987
0 991 5 1 1 990
0 992 7 1 2 2501 688
0 993 5 1 1 992
0 994 7 2 2 2505 993
0 995 5 1 1 2719
0 996 7 1 2 2617 841
0 997 5 1 1 996
0 998 7 3 2 2621 997
0 999 5 2 1 2721
0 1000 7 1 2 2495 680
0 1001 5 1 1 1000
0 1002 7 2 2 2499 1001
0 1003 5 1 1 2726
0 1004 7 1 2 2724 2727
0 1005 5 1 1 1004
0 1006 7 1 2 2722 1003
0 1007 5 1 1 1006
0 1008 7 1 2 2489 672
0 1009 5 1 1 1008
0 1010 7 2 2 2493 1009
0 1011 5 1 1 2728
0 1012 7 1 2 2605 825
0 1013 5 1 1 1012
0 1014 7 3 2 2609 1013
0 1015 5 2 1 2730
0 1016 7 1 2 2483 664
0 1017 5 1 1 1016
0 1018 7 2 2 2487 1017
0 1019 5 1 1 2735
0 1020 7 1 2 2733 2736
0 1021 5 1 1 1020
0 1022 7 1 2 2731 1019
0 1023 5 1 1 1022
0 1024 7 1 2 2477 656
0 1025 5 1 1 1024
0 1026 7 2 2 2481 1025
0 1027 5 1 1 2737
0 1028 7 1 2 2593 809
0 1029 5 1 1 1028
0 1030 7 3 2 2597 1029
0 1031 5 1 1 2739
0 1032 7 1 2 2471 648
0 1033 5 1 1 1032
0 1034 7 2 2 2475 1033
0 1035 5 1 1 2742
0 1036 7 1 2 1031 2743
0 1037 5 1 1 1036
0 1038 7 1 2 2740 1035
0 1039 5 1 1 1038
0 1040 7 1 2 2464 640
0 1041 5 1 1 1040
0 1042 7 1 2 795 801
0 1043 5 1 1 1042
0 1044 7 3 2 2591 1043
0 1045 5 2 1 2744
0 1046 7 1 2 2435 2458
0 1047 5 1 1 1046
0 1048 7 2 2 2465 1047
0 1049 5 1 1 2749
0 1050 7 1 2 2176 2191
0 1051 5 1 1 1050
0 1052 7 2 2 2587 1051
0 1053 5 1 1 2751
0 1054 7 1 2 2449 1053
0 1055 5 1 1 1054
0 1056 7 2 2 2200 1055
0 1057 5 1 1 2753
0 1058 7 1 2 2750 1057
0 1059 5 1 1 1058
0 1060 7 1 2 1049 2754
0 1061 5 1 1 1060
0 1062 7 2 2 2179 2192
0 1063 5 1 1 2755
0 1064 7 1 2 2163 2756
0 1065 5 1 1 1064
0 1066 7 1 2 2160 1063
0 1067 5 1 1 1066
0 1068 7 2 2 1065 1067
0 1069 5 1 1 2757
0 1070 7 1 2 1061 1069
0 1071 5 1 1 1070
0 1072 7 2 2 1059 1071
0 1073 5 1 1 2759
0 1074 7 1 2 2745 2760
0 1075 5 1 1 1074
0 1076 7 1 2 2469 1075
0 1077 7 1 2 1041 1076
0 1078 5 1 1 1077
0 1079 7 1 2 2747 1073
0 1080 5 1 1 1079
0 1081 7 1 2 1078 1080
0 1082 5 1 1 1081
0 1083 7 1 2 1039 1082
0 1084 5 1 1 1083
0 1085 7 2 2 1037 1084
0 1086 5 1 1 2761
0 1087 7 1 2 2738 1086
0 1088 5 1 1 1087
0 1089 7 1 2 2599 817
0 1090 5 1 1 1089
0 1091 7 2 2 2603 1090
0 1092 5 2 1 2763
0 1093 7 1 2 1027 2762
0 1094 5 1 1 1093
0 1095 7 1 2 2765 1094
0 1096 5 1 1 1095
0 1097 7 1 2 1088 1096
0 1098 5 1 1 1097
0 1099 7 1 2 1023 1098
0 1100 5 1 1 1099
0 1101 7 2 2 1021 1100
0 1102 5 1 1 2767
0 1103 7 1 2 2729 1102
0 1104 5 1 1 1103
0 1105 7 1 2 2611 833
0 1106 5 1 1 1105
0 1107 7 2 2 2615 1106
0 1108 5 1 1 2769
0 1109 7 1 2 1011 2768
0 1110 5 1 1 1109
0 1111 7 1 2 1108 1110
0 1112 5 1 1 1111
0 1113 7 1 2 1104 1112
0 1114 5 1 1 1113
0 1115 7 1 2 1007 1114
0 1116 5 1 1 1115
0 1117 7 2 2 1005 1116
0 1118 5 1 1 2771
0 1119 7 1 2 2720 1118
0 1120 5 1 1 1119
0 1121 7 1 2 2623 849
0 1122 5 1 1 1121
0 1123 7 2 2 2627 1122
0 1124 5 1 1 2773
0 1125 7 1 2 995 2772
0 1126 5 1 1 1125
0 1127 7 1 2 1124 1126
0 1128 5 1 1 1127
0 1129 7 1 2 1120 1128
0 1130 5 1 1 1129
0 1131 7 1 2 991 1130
0 1132 5 1 1 1131
0 1133 7 2 2 989 1132
0 1134 5 1 1 2775
0 1135 7 1 2 2711 1134
0 1136 5 1 1 1135
0 1137 7 1 2 2635 865
0 1138 5 1 1 1137
0 1139 7 2 2 2639 1138
0 1140 5 2 1 2777
0 1141 7 1 2 979 2776
0 1142 5 1 1 1141
0 1143 7 1 2 2779 1142
0 1144 5 1 1 1143
0 1145 7 1 2 1136 1144
0 1146 5 1 1 1145
0 1147 7 1 2 975 1146
0 1148 5 1 1 1147
0 1149 7 2 2 973 1148
0 1150 5 1 1 2781
0 1151 7 1 2 2704 1150
0 1152 5 1 1 1151
0 1153 7 1 2 2647 881
0 1154 5 1 1 1153
0 1155 7 2 2 2651 1154
0 1156 5 1 1 2783
0 1157 7 1 2 963 2782
0 1158 5 1 1 1157
0 1159 7 1 2 1156 1158
0 1160 5 1 1 1159
0 1161 7 1 2 1152 1160
0 1162 5 1 1 1161
0 1163 7 1 2 959 1162
0 1164 5 1 1 1163
0 1165 7 1 2 957 1164
0 1166 5 1 1 1165
0 1167 7 1 2 947 1166
0 1168 5 1 1 1167
0 1169 7 2 2 945 1168
0 1170 5 1 1 2785
0 1171 7 1 2 2689 1170
0 1172 5 1 1 1171
0 1173 7 1 2 2687 2786
0 1174 5 1 1 1173
0 1175 7 1 2 2543 744
0 1176 5 1 1 1175
0 1177 7 1 2 2547 1176
0 1178 7 1 2 1174 1177
0 1179 5 1 1 1178
0 1180 7 1 2 1172 1179
0 1181 7 1 2 931 1180
0 1182 5 1 1 1181
0 1183 7 1 2 921 1182
0 1184 5 1 1 1183
0 1185 7 1 2 2266 1184
0 1186 5 1 1 1185
0 1187 7 1 2 2182 2453
0 1188 5 1 1 1187
0 1189 7 2 2 2185 1188
0 1190 5 2 1 2787
0 1191 7 1 2 2169 2789
0 1192 5 1 1 1191
0 1193 7 2 2 2166 1192
0 1194 5 2 1 2791
0 1195 7 1 2 2153 2793
0 1196 5 1 1 1195
0 1197 7 2 2 2150 1196
0 1198 5 2 1 2795
0 1199 7 1 2 2138 2797
0 1200 5 1 1 1199
0 1201 7 2 2 2135 1200
0 1202 5 2 1 2799
0 1203 7 1 2 2123 2801
0 1204 5 1 1 1203
0 1205 7 2 2 2120 1204
0 1206 5 2 1 2803
0 1207 7 1 2 2108 2805
0 1208 5 1 1 1207
0 1209 7 2 2 2105 1208
0 1210 5 2 1 2807
0 1211 7 1 2 2093 2809
0 1212 5 1 1 1211
0 1213 7 2 2 2090 1212
0 1214 5 2 1 2811
0 1215 7 1 2 2078 2813
0 1216 5 1 1 1215
0 1217 7 2 2 2075 1216
0 1218 5 2 1 2815
0 1219 7 1 2 2063 2817
0 1220 5 1 1 1219
0 1221 7 2 2 2060 1220
0 1222 5 2 1 2819
0 1223 7 1 2 2048 2821
0 1224 5 1 1 1223
0 1225 7 2 2 2045 1224
0 1226 5 2 1 2823
0 1227 7 1 2 2033 2825
0 1228 5 1 1 1227
0 1229 7 2 2 2030 1228
0 1230 5 2 1 2827
0 1231 7 1 2 2018 2829
0 1232 5 1 1 1231
0 1233 7 2 2 2015 1232
0 1234 5 2 1 2831
0 1235 7 1 2 2003 2833
0 1236 5 1 1 1235
0 1237 7 2 2 2000 1236
0 1238 5 2 1 2835
0 1239 7 1 2 2269 2836
0 1240 5 1 1 1239
0 1241 7 1 2 2271 2837
0 1242 5 1 1 1241
0 1243 7 3 2 1240 1242
0 1244 5 2 1 2839
0 1245 7 1 2 2312 2828
0 1246 5 1 1 1245
0 1247 7 1 2 2310 2830
0 1248 5 1 1 1247
0 1249 7 3 2 1246 1248
0 1250 5 2 1 2844
0 1251 7 1 2 2840 2847
0 1252 5 2 1 1251
0 1253 7 1 2 2298 2832
0 1254 5 1 1 1253
0 1255 7 1 2 2300 2834
0 1256 5 1 1 1255
0 1257 7 3 2 1254 1256
0 1258 5 2 1 2851
0 1259 7 1 2 2324 2824
0 1260 5 1 1 1259
0 1261 7 1 2 2322 2826
0 1262 5 1 1 1261
0 1263 7 3 2 1260 1262
0 1264 5 2 1 2856
0 1265 7 1 2 2852 2859
0 1266 5 2 1 1265
0 1267 7 1 2 2336 2820
0 1268 5 1 1 1267
0 1269 7 1 2 2334 2822
0 1270 5 1 1 1269
0 1271 7 3 2 1268 1270
0 1272 5 2 1 2863
0 1273 7 1 2 2848 2866
0 1274 5 2 1 1273
0 1275 7 1 2 2348 2816
0 1276 5 1 1 1275
0 1277 7 1 2 2346 2818
0 1278 5 1 1 1277
0 1279 7 3 2 1276 1278
0 1280 5 2 1 2870
0 1281 7 1 2 2860 2873
0 1282 5 2 1 1281
0 1283 7 1 2 2360 2812
0 1284 5 1 1 1283
0 1285 7 1 2 2358 2814
0 1286 5 1 1 1285
0 1287 7 3 2 1284 1286
0 1288 5 2 1 2877
0 1289 7 1 2 2867 2880
0 1290 5 2 1 1289
0 1291 7 1 2 2372 2808
0 1292 5 1 1 1291
0 1293 7 1 2 2370 2810
0 1294 5 1 1 1293
0 1295 7 3 2 1292 1294
0 1296 5 2 1 2884
0 1297 7 1 2 2874 2887
0 1298 5 2 1 1297
0 1299 7 1 2 2384 2804
0 1300 5 1 1 1299
0 1301 7 1 2 2382 2806
0 1302 5 1 1 1301
0 1303 7 3 2 1300 1302
0 1304 5 2 1 2891
0 1305 7 1 2 2881 2894
0 1306 5 2 1 1305
0 1307 7 1 2 2396 2800
0 1308 5 1 1 1307
0 1309 7 1 2 2394 2802
0 1310 5 1 1 1309
0 1311 7 3 2 1308 1310
0 1312 5 2 1 2898
0 1313 7 1 2 2888 2901
0 1314 5 2 1 1313
0 1315 7 1 2 2408 2796
0 1316 5 1 1 1315
0 1317 7 1 2 2406 2798
0 1318 5 1 1 1317
0 1319 7 3 2 1316 1318
0 1320 5 2 1 2905
0 1321 7 1 2 2895 2908
0 1322 5 2 1 1321
0 1323 7 1 2 2420 2792
0 1324 5 1 1 1323
0 1325 7 1 2 2418 2794
0 1326 5 1 1 1325
0 1327 7 3 2 1324 1326
0 1328 5 2 1 2912
0 1329 7 1 2 2902 2915
0 1330 5 2 1 1329
0 1331 7 1 2 2432 2788
0 1332 5 1 1 1331
0 1333 7 1 2 2430 2790
0 1334 5 1 1 1333
0 1335 7 3 2 1332 1334
0 1336 5 2 1 2919
0 1337 7 1 2 2909 2922
0 1338 5 2 1 1337
0 1339 7 1 2 2442 2456
0 1340 5 1 1 1339
0 1341 7 1 2 2444 2454
0 1342 5 1 1 1341
0 1343 7 2 2 1340 1342
0 1344 5 2 1 2926
0 1345 7 1 2 2916 2927
0 1346 5 2 1 1345
0 1347 7 2 2 2461 2923
0 1348 5 2 1 2932
0 1349 7 1 2 2913 2928
0 1350 5 1 1 1349
0 1351 7 2 2 2930 1350
0 1352 5 1 1 2936
0 1353 7 1 2 2933 2937
0 1354 5 2 1 1353
0 1355 7 2 2 2931 2938
0 1356 5 1 1 2940
0 1357 7 1 2 2906 2920
0 1358 5 1 1 1357
0 1359 7 2 2 2924 1358
0 1360 5 1 1 2942
0 1361 7 1 2 1356 2943
0 1362 5 2 1 1361
0 1363 7 2 2 2925 2944
0 1364 5 1 1 2946
0 1365 7 1 2 2899 2914
0 1366 5 1 1 1365
0 1367 7 2 2 2917 1366
0 1368 5 1 1 2948
0 1369 7 1 2 1364 2949
0 1370 5 2 1 1369
0 1371 7 2 2 2918 2950
0 1372 5 1 1 2952
0 1373 7 1 2 2892 2907
0 1374 5 1 1 1373
0 1375 7 2 2 2910 1374
0 1376 5 1 1 2954
0 1377 7 1 2 1372 2955
0 1378 5 2 1 1377
0 1379 7 2 2 2911 2956
0 1380 5 1 1 2958
0 1381 7 1 2 2885 2900
0 1382 5 1 1 1381
0 1383 7 2 2 2903 1382
0 1384 5 1 1 2960
0 1385 7 1 2 1380 2961
0 1386 5 2 1 1385
0 1387 7 2 2 2904 2962
0 1388 5 1 1 2964
0 1389 7 1 2 2878 2893
0 1390 5 1 1 1389
0 1391 7 2 2 2896 1390
0 1392 5 1 1 2966
0 1393 7 1 2 1388 2967
0 1394 5 2 1 1393
0 1395 7 2 2 2897 2968
0 1396 5 1 1 2970
0 1397 7 1 2 2871 2886
0 1398 5 1 1 1397
0 1399 7 2 2 2889 1398
0 1400 5 1 1 2972
0 1401 7 1 2 1396 2973
0 1402 5 2 1 1401
0 1403 7 2 2 2890 2974
0 1404 5 1 1 2976
0 1405 7 1 2 2864 2879
0 1406 5 1 1 1405
0 1407 7 2 2 2882 1406
0 1408 5 1 1 2978
0 1409 7 1 2 1404 2979
0 1410 5 2 1 1409
0 1411 7 2 2 2883 2980
0 1412 5 1 1 2982
0 1413 7 1 2 2857 2872
0 1414 5 1 1 1413
0 1415 7 2 2 2875 1414
0 1416 5 1 1 2984
0 1417 7 1 2 1412 2985
0 1418 5 2 1 1417
0 1419 7 2 2 2876 2986
0 1420 5 1 1 2988
0 1421 7 1 2 2845 2865
0 1422 5 1 1 1421
0 1423 7 2 2 2868 1422
0 1424 5 1 1 2990
0 1425 7 1 2 1420 2991
0 1426 5 2 1 1425
0 1427 7 2 2 2869 2992
0 1428 5 1 1 2994
0 1429 7 1 2 2854 2858
0 1430 5 1 1 1429
0 1431 7 2 2 2861 1430
0 1432 5 1 1 2996
0 1433 7 1 2 1428 2997
0 1434 5 2 1 1433
0 1435 7 2 2 2862 2998
0 1436 5 1 1 3000
0 1437 7 1 2 2842 2846
0 1438 5 1 1 1437
0 1439 7 2 2 2849 1438
0 1440 5 1 1 3002
0 1441 7 1 2 1436 3003
0 1442 5 2 1 1441
0 1443 7 2 2 2850 3004
0 1444 5 1 1 3006
0 1445 7 1 2 1988 2838
0 1446 5 1 1 1445
0 1447 7 2 2 1985 1446
0 1448 5 2 1 3008
0 1449 7 1 2 2288 3009
0 1450 5 1 1 1449
0 1451 7 1 2 2290 3010
0 1452 5 1 1 1451
0 1453 7 3 2 1450 1452
0 1454 5 2 1 3012
0 1455 7 1 2 2853 3013
0 1456 5 2 1 1455
0 1457 7 1 2 2855 3015
0 1458 5 1 1 1457
0 1459 7 2 2 3017 1458
0 1460 5 1 1 3019
0 1461 7 1 2 1444 3020
0 1462 5 2 1 1461
0 1463 7 1 2 3007 1460
0 1464 5 1 1 1463
0 1465 7 2 2 3021 1464
0 1466 5 1 1 3023
0 1467 7 1 2 2995 1432
0 1468 5 1 1 1467
0 1469 7 2 2 2999 1468
0 1470 5 1 1 3025
0 1471 7 1 2 2989 1424
0 1472 5 1 1 1471
0 1473 7 2 2 2993 1472
0 1474 5 1 1 3027
0 1475 7 1 2 2983 1416
0 1476 5 1 1 1475
0 1477 7 2 2 2987 1476
0 1478 5 1 1 3029
0 1479 7 1 2 2778 1478
0 1480 5 1 1 1479
0 1481 7 1 2 2780 3030
0 1482 5 1 1 1481
0 1483 7 1 2 2971 1400
0 1484 5 1 1 1483
0 1485 7 2 2 2975 1484
0 1486 5 1 1 3031
0 1487 7 1 2 2965 1392
0 1488 5 1 1 1487
0 1489 7 2 2 2969 1488
0 1490 5 1 1 3033
0 1491 7 1 2 2723 1490
0 1492 5 1 1 1491
0 1493 7 1 2 2725 3034
0 1494 5 1 1 1493
0 1495 7 1 2 2959 1384
0 1496 5 1 1 1495
0 1497 7 2 2 2963 1496
0 1498 5 1 1 3035
0 1499 7 1 2 2953 1376
0 1500 5 1 1 1499
0 1501 7 2 2 2957 1500
0 1502 5 1 1 3037
0 1503 7 1 2 2732 1502
0 1504 5 1 1 1503
0 1505 7 1 2 2734 3038
0 1506 5 1 1 1505
0 1507 7 1 2 2947 1368
0 1508 5 1 1 1507
0 1509 7 2 2 2951 1508
0 1510 5 1 1 3039
0 1511 7 1 2 2764 1510
0 1512 5 1 1 1511
0 1513 7 1 2 2766 3040
0 1514 5 1 1 1513
0 1515 7 1 2 2934 1352
0 1516 5 1 1 1515
0 1517 7 2 2 2939 1516
0 1518 5 1 1 3041
0 1519 7 1 2 2746 1518
0 1520 5 1 1 1519
0 1521 7 1 2 2748 3042
0 1522 5 1 1 1521
0 1523 7 1 2 2459 2921
0 1524 5 1 1 1523
0 1525 7 2 2 2935 1524
0 1526 5 1 1 3043
0 1527 7 1 2 2198 2929
0 1528 5 1 1 1527
0 1529 7 1 2 2446 2752
0 1530 5 1 1 1529
0 1531 7 2 2 1528 1530
0 1532 5 1 1 3045
0 1533 7 1 2 3044 3046
0 1534 5 1 1 1533
0 1535 7 1 2 2758 1534
0 1536 5 1 1 1535
0 1537 7 1 2 1526 1532
0 1538 5 1 1 1537
0 1539 7 1 2 1536 1538
0 1540 5 1 1 1539
0 1541 7 1 2 1522 1540
0 1542 5 1 1 1541
0 1543 7 2 2 1520 1542
0 1544 5 1 1 3047
0 1545 7 1 2 2941 1360
0 1546 5 1 1 1545
0 1547 7 2 2 2945 1546
0 1548 5 1 1 3049
0 1549 7 1 2 3048 3050
0 1550 5 1 1 1549
0 1551 7 1 2 2741 1550
0 1552 5 1 1 1551
0 1553 7 1 2 1544 1548
0 1554 5 1 1 1553
0 1555 7 1 2 1552 1554
0 1556 5 1 1 1555
0 1557 7 1 2 1514 1556
0 1558 5 1 1 1557
0 1559 7 1 2 1512 1558
0 1560 5 1 1 1559
0 1561 7 1 2 1506 1560
0 1562 5 1 1 1561
0 1563 7 2 2 1504 1562
0 1564 5 1 1 3051
0 1565 7 1 2 3036 3052
0 1566 5 1 1 1565
0 1567 7 1 2 2770 1566
0 1568 5 1 1 1567
0 1569 7 1 2 1498 1564
0 1570 5 1 1 1569
0 1571 7 1 2 1568 1570
0 1572 5 1 1 1571
0 1573 7 1 2 1494 1572
0 1574 5 1 1 1573
0 1575 7 2 2 1492 1574
0 1576 5 1 1 3053
0 1577 7 1 2 3032 3054
0 1578 5 1 1 1577
0 1579 7 1 2 2774 1578
0 1580 5 1 1 1579
0 1581 7 1 2 1486 1576
0 1582 5 1 1 1581
0 1583 7 1 2 1580 1582
0 1584 5 1 1 1583
0 1585 7 1 2 2977 1408
0 1586 5 1 1 1585
0 1587 7 2 2 2981 1586
0 1588 5 1 1 3055
0 1589 7 1 2 2716 3056
0 1590 5 1 1 1589
0 1591 7 1 2 1584 1590
0 1592 5 1 1 1591
0 1593 7 1 2 2714 1588
0 1594 5 1 1 1593
0 1595 7 1 2 1592 1594
0 1596 5 1 1 1595
0 1597 7 1 2 1482 1596
0 1598 5 1 1 1597
0 1599 7 2 2 1480 1598
0 1600 5 1 1 3057
0 1601 7 1 2 3028 3058
0 1602 5 1 1 1601
0 1603 7 1 2 2707 1602
0 1604 5 1 1 1603
0 1605 7 1 2 1474 1600
0 1606 5 1 1 1605
0 1607 7 2 2 1604 1606
0 1608 5 1 1 3059
0 1609 7 1 2 3026 3060
0 1610 5 1 1 1609
0 1611 7 1 2 2784 1610
0 1612 5 1 1 1611
0 1613 7 1 2 1470 1608
0 1614 5 1 1 1613
0 1615 7 1 2 1612 1614
0 1616 5 1 1 1615
0 1617 7 1 2 3001 1440
0 1618 5 1 1 1617
0 1619 7 2 2 3005 1618
0 1620 5 1 1 3061
0 1621 7 1 2 2700 3062
0 1622 5 1 1 1621
0 1623 7 1 2 1616 1622
0 1624 5 1 1 1623
0 1625 7 1 2 2698 1620
0 1626 5 1 1 1625
0 1627 7 2 2 1624 1626
0 1628 5 1 1 3063
0 1629 7 1 2 3024 3064
0 1630 5 1 1 1629
0 1631 7 1 2 2693 1630
0 1632 5 1 1 1631
0 1633 7 1 2 1466 1628
0 1634 5 1 1 1633
0 1635 7 2 2 1632 1634
0 1636 5 1 1 3065
0 1637 7 1 2 2688 1636
0 1638 5 1 1 1637
0 1639 7 2 2 3018 3022
0 1640 5 1 1 3067
0 1641 7 1 2 1973 3011
0 1642 5 1 1 1641
0 1643 7 3 2 1970 1642
0 1644 5 3 1 3069
0 1645 7 1 2 2279 3070
0 1646 5 1 1 1645
0 1647 7 1 2 2281 3072
0 1648 5 1 1 1647
0 1649 7 2 2 1646 1648
0 1650 5 1 1 3075
0 1651 7 1 2 2841 3076
0 1652 5 2 1 1651
0 1653 7 1 2 2843 1650
0 1654 5 1 1 1653
0 1655 7 2 2 3077 1654
0 1656 5 1 1 3079
0 1657 7 1 2 1640 3080
0 1658 5 2 1 1657
0 1659 7 1 2 3068 1656
0 1660 5 1 1 1659
0 1661 7 1 2 3081 1660
0 1662 7 1 2 1638 1661
0 1663 5 1 1 1662
0 1664 7 2 2 3078 3082
0 1665 5 1 1 3083
0 1666 7 1 2 1959 3073
0 1667 5 2 1 1666
0 1668 7 2 2 1953 3085
0 1669 5 1 1 3087
0 1670 7 1 2 3014 1669
0 1671 5 2 1 1670
0 1672 7 1 2 3016 3088
0 1673 5 1 1 1672
0 1674 7 2 2 3089 1673
0 1675 5 1 1 3091
0 1676 7 1 2 1665 3092
0 1677 5 2 1 1676
0 1678 7 1 2 3084 1675
0 1679 5 1 1 1678
0 1680 7 2 2 3093 1679
0 1681 5 1 1 3095
0 1682 7 2 2 2674 2685
0 1683 5 1 1 3097
0 1684 7 1 2 3096 1683
0 1685 5 1 1 1684
0 1686 7 1 2 2690 3066
0 1687 5 1 1 1686
0 1688 7 1 2 1685 1687
0 1689 7 1 2 1663 1688
0 1690 5 1 1 1689
0 1691 7 1 2 1681 3098
0 1692 5 1 1 1691
0 1693 7 2 2 3090 3094
0 1694 5 1 1 3099
0 1695 7 1 2 1960 3071
0 1696 5 1 1 1695
0 1697 7 1 2 1954 3074
0 1698 5 1 1 1697
0 1699 7 2 2 1696 1698
0 1700 5 1 1 3101
0 1701 7 1 2 1694 3102
0 1702 5 2 1 1701
0 1703 7 1 2 3100 1700
0 1704 5 2 1 1703
0 1705 7 1 2 3103 3105
0 1706 5 1 1 1705
0 1707 7 1 2 2677 1706
0 1708 5 1 1 1707
0 1709 7 1 2 1692 1708
0 1710 7 1 2 1690 1709
0 1711 5 1 1 1710
0 1712 7 1 2 2675 3106
0 1713 5 1 1 1712
0 1714 7 1 2 2264 3086
0 1715 7 1 2 3104 1714
0 1716 7 1 2 1713 1715
0 1717 7 1 2 1711 1716
0 1718 5 1 1 1717
0 1719 7 1 2 1186 1718
3 3499 5 0 1 1719
