1 0 0 2 0
2 49 1 0
2 704 1 0
1 1 0 2 0
2 705 1 1
2 706 1 1
1 2 0 2 0
2 707 1 2
2 708 1 2
1 3 0 2 0
2 709 1 3
2 710 1 3
1 4 0 2 0
2 711 1 4
2 712 1 4
1 5 0 2 0
2 713 1 5
2 714 1 5
1 6 0 2 0
2 715 1 6
2 716 1 6
1 7 0 2 0
2 717 1 7
2 718 1 7
1 8 0 2 0
2 719 1 8
2 720 1 8
1 9 0 2 0
2 721 1 9
2 722 1 9
1 10 0 2 0
2 723 1 10
2 724 1 10
1 11 0 2 0
2 725 1 11
2 726 1 11
1 12 0 2 0
2 727 1 12
2 728 1 12
1 13 0 2 0
2 729 1 13
2 730 1 13
1 14 0 2 0
2 731 1 14
2 732 1 14
1 15 0 2 0
2 733 1 15
2 734 1 15
1 16 0 2 0
2 735 1 16
2 736 1 16
1 17 0 2 0
2 737 1 17
2 738 1 17
1 18 0 2 0
2 739 1 18
2 740 1 18
1 19 0 2 0
2 741 1 19
2 742 1 19
1 20 0 2 0
2 743 1 20
2 744 1 20
1 21 0 2 0
2 745 1 21
2 746 1 21
1 22 0 2 0
2 747 1 22
2 748 1 22
1 23 0 2 0
2 749 1 23
2 750 1 23
1 24 0 2 0
2 751 1 24
2 752 1 24
1 25 0 2 0
2 753 1 25
2 754 1 25
1 26 0 2 0
2 755 1 26
2 756 1 26
1 27 0 2 0
2 757 1 27
2 758 1 27
1 28 0 2 0
2 759 1 28
2 760 1 28
1 29 0 2 0
2 761 1 29
2 762 1 29
1 30 0 2 0
2 763 1 30
2 764 1 30
1 31 0 2 0
2 765 1 31
2 766 1 31
1 32 0 2 0
2 767 1 32
2 768 1 32
1 33 0 3 0
2 769 1 33
2 770 1 33
2 771 1 33
1 34 0 3 0
2 772 1 34
2 773 1 34
2 774 1 34
1 35 0 3 0
2 775 1 35
2 776 1 35
2 777 1 35
1 36 0 3 0
2 778 1 36
2 779 1 36
2 780 1 36
1 37 0 3 0
2 781 1 37
2 782 1 37
2 783 1 37
1 38 0 3 0
2 784 1 38
2 785 1 38
2 786 1 38
1 39 0 3 0
2 787 1 39
2 788 1 39
2 789 1 39
1 40 0 3 0
2 790 1 40
2 791 1 40
2 792 1 40
1 41 0 3 0
2 793 1 41
2 794 1 41
2 795 1 41
1 42 0 3 0
2 796 1 42
2 797 1 42
2 798 1 42
1 43 0 3 0
2 799 1 43
2 800 1 43
2 801 1 43
1 44 0 3 0
2 802 1 44
2 803 1 44
2 804 1 44
1 45 0 2 0
2 805 1 45
2 806 1 45
1 46 0 3 0
2 807 1 46
2 808 1 46
2 809 1 46
1 47 0 3 0
2 810 1 47
2 811 1 47
2 812 1 47
1 48 0 2 0
2 813 1 48
2 814 1 48
2 815 1 69
2 816 1 69
2 817 1 70
2 818 1 70
2 819 1 71
2 820 1 71
2 821 1 72
2 822 1 72
2 823 1 73
2 824 1 73
2 825 1 74
2 826 1 74
2 827 1 75
2 828 1 75
2 829 1 76
2 830 1 76
2 831 1 77
2 832 1 77
2 833 1 78
2 834 1 78
2 835 1 79
2 836 1 79
2 837 1 80
2 838 1 80
2 839 1 83
2 840 1 83
2 841 1 84
2 842 1 84
2 843 1 85
2 844 1 85
2 845 1 86
2 846 1 86
2 847 1 87
2 848 1 87
2 849 1 88
2 850 1 88
2 851 1 89
2 852 1 89
2 853 1 90
2 854 1 90
2 855 1 91
2 856 1 91
2 857 1 92
2 858 1 92
2 859 1 93
2 860 1 93
2 861 1 94
2 862 1 94
2 863 1 95
2 864 1 95
2 865 1 96
2 866 1 96
2 867 1 97
2 868 1 97
2 869 1 98
2 870 1 98
2 871 1 98
2 872 1 100
2 873 1 100
2 874 1 102
2 875 1 102
2 876 1 104
2 877 1 104
2 878 1 106
2 879 1 106
2 880 1 107
2 881 1 107
2 882 1 108
2 883 1 108
2 884 1 108
2 885 1 111
2 886 1 111
2 887 1 112
2 888 1 112
2 889 1 115
2 890 1 115
2 891 1 118
2 892 1 118
2 893 1 120
2 894 1 120
2 895 1 123
2 896 1 123
2 897 1 126
2 898 1 126
2 899 1 128
2 900 1 128
2 901 1 131
2 902 1 131
2 903 1 134
2 904 1 134
2 905 1 136
2 906 1 136
2 907 1 139
2 908 1 139
2 909 1 142
2 910 1 142
2 911 1 144
2 912 1 144
2 913 1 147
2 914 1 147
2 915 1 150
2 916 1 150
2 917 1 152
2 918 1 152
2 919 1 155
2 920 1 155
2 921 1 158
2 922 1 158
2 923 1 160
2 924 1 160
2 925 1 163
2 926 1 163
2 927 1 166
2 928 1 166
2 929 1 168
2 930 1 168
2 931 1 171
2 932 1 171
2 933 1 174
2 934 1 174
2 935 1 176
2 936 1 176
2 937 1 179
2 938 1 179
2 939 1 182
2 940 1 182
2 941 1 184
2 942 1 184
2 943 1 187
2 944 1 187
2 945 1 190
2 946 1 190
2 947 1 192
2 948 1 192
2 949 1 195
2 950 1 195
2 951 1 198
2 952 1 198
2 953 1 200
2 954 1 200
2 955 1 203
2 956 1 203
2 957 1 206
2 958 1 206
2 959 1 208
2 960 1 208
2 961 1 209
2 962 1 209
2 963 1 215
2 964 1 215
2 965 1 216
2 966 1 216
2 967 1 218
2 968 1 218
2 969 1 220
2 970 1 220
2 971 1 221
2 972 1 221
2 973 1 227
2 974 1 227
2 975 1 228
2 976 1 228
2 977 1 230
2 978 1 230
2 979 1 232
2 980 1 232
2 981 1 233
2 982 1 233
2 983 1 239
2 984 1 239
2 985 1 239
2 986 1 242
2 987 1 242
2 988 1 244
2 989 1 244
2 990 1 245
2 991 1 245
2 992 1 246
2 993 1 246
2 994 1 251
2 995 1 251
2 996 1 251
2 997 1 254
2 998 1 254
2 999 1 256
2 1000 1 256
2 1001 1 259
2 1002 1 259
2 1003 1 261
2 1004 1 261
2 1005 1 261
2 1006 1 265
2 1007 1 265
2 1008 1 266
2 1009 1 266
2 1010 1 269
2 1011 1 269
2 1012 1 272
2 1013 1 272
2 1014 1 274
2 1015 1 274
2 1016 1 275
2 1017 1 275
2 1018 1 281
2 1019 1 281
2 1020 1 281
2 1021 1 285
2 1022 1 285
2 1023 1 286
2 1024 1 286
2 1025 1 289
2 1026 1 289
2 1027 1 292
2 1028 1 292
2 1029 1 293
2 1030 1 293
2 1031 1 299
2 1032 1 299
2 1033 1 299
2 1034 1 302
2 1035 1 302
2 1036 1 305
2 1037 1 305
2 1038 1 308
2 1039 1 308
2 1040 1 309
2 1041 1 309
2 1042 1 315
2 1043 1 315
2 1044 1 316
2 1045 1 316
2 1046 1 316
2 1047 1 318
2 1048 1 318
2 1049 1 321
2 1050 1 321
2 1051 1 324
2 1052 1 324
2 1053 1 325
2 1054 1 325
2 1055 1 331
2 1056 1 331
2 1057 1 331
2 1058 1 334
2 1059 1 334
2 1060 1 337
2 1061 1 337
2 1062 1 340
2 1063 1 340
2 1064 1 341
2 1065 1 341
2 1066 1 347
2 1067 1 347
2 1068 1 347
2 1069 1 348
2 1070 1 348
2 1071 1 350
2 1072 1 350
2 1073 1 353
2 1074 1 353
2 1075 1 356
2 1076 1 356
2 1077 1 357
2 1078 1 357
2 1079 1 363
2 1080 1 363
2 1081 1 363
2 1082 1 366
2 1083 1 366
2 1084 1 369
2 1085 1 369
2 1086 1 372
2 1087 1 372
2 1088 1 373
2 1089 1 373
2 1090 1 379
2 1091 1 379
2 1092 1 380
2 1093 1 380
2 1094 1 380
2 1095 1 382
2 1096 1 382
2 1097 1 385
2 1098 1 385
2 1099 1 388
2 1100 1 388
2 1101 1 389
2 1102 1 389
2 1103 1 395
2 1104 1 395
2 1105 1 395
2 1106 1 398
2 1107 1 398
2 1108 1 401
2 1109 1 401
2 1110 1 404
2 1111 1 404
2 1112 1 405
2 1113 1 405
2 1114 1 411
2 1115 1 411
2 1116 1 412
2 1117 1 412
2 1118 1 412
2 1119 1 414
2 1120 1 414
2 1121 1 417
2 1122 1 417
2 1123 1 420
2 1124 1 420
2 1125 1 421
2 1126 1 421
2 1127 1 427
2 1128 1 427
2 1129 1 427
2 1130 1 428
2 1131 1 428
2 1132 1 430
2 1133 1 430
2 1134 1 433
2 1135 1 433
2 1136 1 433
2 1137 1 435
2 1138 1 435
2 1139 1 438
2 1140 1 438
2 1141 1 438
2 1142 1 445
2 1143 1 445
2 1144 1 446
2 1145 1 446
2 1146 1 448
2 1147 1 448
2 1148 1 450
2 1149 1 450
2 1150 1 451
2 1151 1 451
2 1152 1 457
2 1153 1 457
2 1154 1 457
2 1155 1 458
2 1156 1 458
2 1157 1 462
2 1158 1 462
2 1159 1 471
2 1160 1 471
2 1161 1 473
2 1162 1 473
2 1163 1 477
2 1164 1 477
2 1165 1 481
2 1166 1 481
2 1167 1 485
2 1168 1 485
2 1169 1 489
2 1170 1 489
2 1171 1 491
2 1172 1 491
2 1173 1 493
2 1174 1 493
2 1175 1 497
2 1176 1 497
2 1177 1 501
2 1178 1 501
2 1179 1 509
2 1180 1 509
2 1181 1 513
2 1182 1 513
2 1183 1 521
2 1184 1 521
2 1185 1 530
2 1186 1 530
2 1187 1 608
2 1188 1 608
2 1189 1 619
2 1190 1 619
2 1191 1 630
2 1192 1 630
2 1193 1 641
2 1194 1 641
2 1195 1 652
2 1196 1 652
2 1197 1 663
2 1198 1 663
2 1199 1 675
2 1200 1 675
2 1201 1 687
2 1202 1 687
0 50 5 1 1 49
0 51 5 1 1 705
0 52 5 1 1 707
0 53 5 1 1 709
0 54 5 1 1 711
0 55 5 1 1 713
0 56 5 1 1 715
0 57 5 1 1 717
0 58 5 1 1 719
0 59 5 1 1 721
0 60 5 1 1 723
0 61 5 1 1 725
0 62 5 1 1 727
0 63 5 1 1 729
0 64 5 1 1 731
0 65 5 1 1 733
0 66 5 1 1 735
0 67 5 1 1 737
0 68 5 1 1 739
0 69 5 2 1 741
0 70 5 2 1 743
0 71 5 2 1 745
0 72 5 2 1 747
0 73 5 2 1 749
0 74 5 2 1 751
0 75 5 2 1 753
0 76 5 2 1 755
0 77 5 2 1 757
0 78 5 2 1 759
0 79 5 2 1 761
0 80 5 2 1 763
0 81 5 1 1 765
0 82 5 1 1 767
0 83 5 2 1 769
0 84 5 2 1 772
0 85 5 2 1 775
0 86 5 2 1 778
0 87 5 2 1 781
0 88 5 2 1 784
0 89 5 2 1 787
0 90 5 2 1 790
0 91 5 2 1 793
0 92 5 2 1 796
0 93 5 2 1 799
0 94 5 2 1 802
0 95 5 2 1 805
0 96 5 2 1 807
0 97 5 2 1 810
0 98 5 3 1 813
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 708 740
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 706 738
0 106 5 2 1 105
0 107 7 2 2 704 736
0 108 5 3 1 880
0 109 7 1 2 878 882
0 110 5 1 1 109
0 111 7 2 2 876 110
0 112 5 2 1 885
0 113 7 1 2 874 887
0 114 5 1 1 113
0 115 7 2 2 872 114
0 116 5 1 1 889
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 710 890
0 120 5 2 1 119
0 121 7 1 2 815 893
0 122 5 1 1 121
0 123 7 2 2 891 122
0 124 5 1 1 895
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 712 896
0 128 5 2 1 127
0 129 7 1 2 817 899
0 130 5 1 1 129
0 131 7 2 2 897 130
0 132 5 1 1 901
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 714 902
0 136 5 2 1 135
0 137 7 1 2 819 905
0 138 5 1 1 137
0 139 7 2 2 903 138
0 140 5 1 1 907
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 716 908
0 144 5 2 1 143
0 145 7 1 2 821 911
0 146 5 1 1 145
0 147 7 2 2 909 146
0 148 5 1 1 913
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 718 914
0 152 5 2 1 151
0 153 7 1 2 823 917
0 154 5 1 1 153
0 155 7 2 2 915 154
0 156 5 1 1 919
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 720 920
0 160 5 2 1 159
0 161 7 1 2 825 923
0 162 5 1 1 161
0 163 7 2 2 921 162
0 164 5 1 1 925
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 722 926
0 168 5 2 1 167
0 169 7 1 2 827 929
0 170 5 1 1 169
0 171 7 2 2 927 170
0 172 5 1 1 931
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 724 932
0 176 5 2 1 175
0 177 7 1 2 829 935
0 178 5 1 1 177
0 179 7 2 2 933 178
0 180 5 1 1 937
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 726 938
0 184 5 2 1 183
0 185 7 1 2 831 941
0 186 5 1 1 185
0 187 7 2 2 939 186
0 188 5 1 1 943
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 728 944
0 192 5 2 1 191
0 193 7 1 2 833 947
0 194 5 1 1 193
0 195 7 2 2 945 194
0 196 5 1 1 949
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 730 950
0 200 5 2 1 199
0 201 7 1 2 835 953
0 202 5 1 1 201
0 203 7 2 2 951 202
0 204 5 1 1 955
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 732 956
0 208 5 2 1 207
0 209 7 2 2 957 959
0 210 5 1 1 961
0 211 7 1 2 764 962
0 212 5 1 1 211
0 213 7 1 2 837 210
0 214 5 1 1 213
0 215 7 2 2 212 214
0 216 5 2 1 963
0 217 7 1 2 865 964
0 218 5 2 1 217
0 219 7 1 2 808 965
0 220 5 2 1 219
0 221 7 2 2 898 900
0 222 5 1 1 971
0 223 7 1 2 744 972
0 224 5 1 1 223
0 225 7 1 2 818 222
0 226 5 1 1 225
0 227 7 2 2 224 226
0 228 5 2 1 973
0 229 7 1 2 779 975
0 230 5 2 1 229
0 231 7 1 2 845 974
0 232 5 2 1 231
0 233 7 2 2 873 875
0 234 5 1 1 981
0 235 7 1 2 886 234
0 236 5 1 1 235
0 237 7 1 2 888 982
0 238 5 1 1 237
0 239 7 3 2 236 238
0 240 5 1 1 983
0 241 7 1 2 841 240
0 242 5 2 1 241
0 243 7 1 2 773 984
0 244 5 2 1 243
0 245 7 2 2 877 879
0 246 5 2 1 990
0 247 7 1 2 881 992
0 248 5 1 1 247
0 249 7 1 2 883 991
0 250 5 1 1 249
0 251 7 3 2 248 250
0 252 5 1 1 994
0 253 7 1 2 839 252
0 254 5 2 1 253
0 255 7 1 2 770 995
0 256 5 2 1 255
0 257 7 1 2 50 66
0 258 5 1 1 257
0 259 7 2 2 884 258
0 260 5 1 1 1001
0 261 7 3 2 82 1002
0 262 5 1 1 1003
0 263 7 1 2 999 1004
0 264 5 1 1 263
0 265 7 2 2 997 264
0 266 5 2 1 1006
0 267 7 1 2 988 1008
0 268 5 1 1 267
0 269 7 2 2 986 268
0 270 5 1 1 1010
0 271 7 1 2 776 1011
0 272 5 2 1 271
0 273 7 1 2 843 270
0 274 5 2 1 273
0 275 7 2 2 892 894
0 276 5 1 1 1016
0 277 7 1 2 742 1017
0 278 5 1 1 277
0 279 7 1 2 816 276
0 280 5 1 1 279
0 281 7 3 2 278 280
0 282 5 1 1 1018
0 283 7 1 2 1014 282
0 284 5 1 1 283
0 285 7 2 2 1012 284
0 286 5 2 1 1021
0 287 7 1 2 979 1023
0 288 5 1 1 287
0 289 7 2 2 977 288
0 290 5 1 1 1025
0 291 7 1 2 782 290
0 292 5 2 1 291
0 293 7 2 2 904 906
0 294 5 1 1 1029
0 295 7 1 2 746 1030
0 296 5 1 1 295
0 297 7 1 2 820 294
0 298 5 1 1 297
0 299 7 3 2 296 298
0 300 5 1 1 1031
0 301 7 1 2 847 1026
0 302 5 2 1 301
0 303 7 1 2 300 1034
0 304 5 1 1 303
0 305 7 2 2 1027 304
0 306 5 1 1 1036
0 307 7 1 2 785 306
0 308 5 2 1 307
0 309 7 2 2 910 912
0 310 5 1 1 1040
0 311 7 1 2 748 1041
0 312 5 1 1 311
0 313 7 1 2 822 310
0 314 5 1 1 313
0 315 7 2 2 312 314
0 316 5 3 1 1042
0 317 7 1 2 849 1037
0 318 5 2 1 317
0 319 7 1 2 1044 1047
0 320 5 1 1 319
0 321 7 2 2 1038 320
0 322 5 1 1 1049
0 323 7 1 2 788 322
0 324 5 2 1 323
0 325 7 2 2 916 918
0 326 5 1 1 1053
0 327 7 1 2 750 1054
0 328 5 1 1 327
0 329 7 1 2 824 326
0 330 5 1 1 329
0 331 7 3 2 328 330
0 332 5 1 1 1055
0 333 7 1 2 851 1050
0 334 5 2 1 333
0 335 7 1 2 332 1058
0 336 5 1 1 335
0 337 7 2 2 1051 336
0 338 5 1 1 1060
0 339 7 1 2 791 338
0 340 5 2 1 339
0 341 7 2 2 922 924
0 342 5 1 1 1064
0 343 7 1 2 752 1065
0 344 5 1 1 343
0 345 7 1 2 826 342
0 346 5 1 1 345
0 347 7 3 2 344 346
0 348 5 2 1 1066
0 349 7 1 2 853 1061
0 350 5 2 1 349
0 351 7 1 2 1069 1071
0 352 5 1 1 351
0 353 7 2 2 1062 352
0 354 5 1 1 1073
0 355 7 1 2 794 354
0 356 5 2 1 355
0 357 7 2 2 928 930
0 358 5 1 1 1077
0 359 7 1 2 754 1078
0 360 5 1 1 359
0 361 7 1 2 828 358
0 362 5 1 1 361
0 363 7 3 2 360 362
0 364 5 1 1 1079
0 365 7 1 2 855 1074
0 366 5 2 1 365
0 367 7 1 2 364 1082
0 368 5 1 1 367
0 369 7 2 2 1075 368
0 370 5 1 1 1084
0 371 7 1 2 797 370
0 372 5 2 1 371
0 373 7 2 2 934 936
0 374 5 1 1 1088
0 375 7 1 2 756 1089
0 376 5 1 1 375
0 377 7 1 2 830 374
0 378 5 1 1 377
0 379 7 2 2 376 378
0 380 5 3 1 1090
0 381 7 1 2 857 1085
0 382 5 2 1 381
0 383 7 1 2 1092 1095
0 384 5 1 1 383
0 385 7 2 2 1086 384
0 386 5 1 1 1097
0 387 7 1 2 800 386
0 388 5 2 1 387
0 389 7 2 2 940 942
0 390 5 1 1 1101
0 391 7 1 2 758 1102
0 392 5 1 1 391
0 393 7 1 2 832 390
0 394 5 1 1 393
0 395 7 3 2 392 394
0 396 5 1 1 1103
0 397 7 1 2 859 1098
0 398 5 2 1 397
0 399 7 1 2 396 1106
0 400 5 1 1 399
0 401 7 2 2 1099 400
0 402 5 1 1 1108
0 403 7 1 2 803 402
0 404 5 2 1 403
0 405 7 2 2 946 948
0 406 5 1 1 1112
0 407 7 1 2 760 1113
0 408 5 1 1 407
0 409 7 1 2 834 406
0 410 5 1 1 409
0 411 7 2 2 408 410
0 412 5 3 1 1114
0 413 7 1 2 861 1109
0 414 5 2 1 413
0 415 7 1 2 1116 1119
0 416 5 1 1 415
0 417 7 2 2 1110 416
0 418 5 1 1 1121
0 419 7 1 2 806 418
0 420 5 2 1 419
0 421 7 2 2 952 954
0 422 5 1 1 1125
0 423 7 1 2 762 1126
0 424 5 1 1 423
0 425 7 1 2 836 422
0 426 5 1 1 425
0 427 7 3 2 424 426
0 428 5 2 1 1127
0 429 7 1 2 863 1122
0 430 5 2 1 429
0 431 7 1 2 1130 1132
0 432 5 1 1 431
0 433 7 3 2 1123 432
0 434 5 1 1 1134
0 435 7 2 2 969 1135
0 436 5 1 1 1137
0 437 7 1 2 967 436
0 438 5 3 1 437
0 439 7 1 2 867 1139
0 440 5 1 1 439
0 441 7 1 2 869 440
0 442 5 1 1 441
0 443 7 1 2 838 960
0 444 5 1 1 443
0 445 7 2 2 958 444
0 446 5 2 1 1142
0 447 7 1 2 65 81
0 448 5 2 1 447
0 449 7 1 2 734 766
0 450 5 2 1 449
0 451 7 2 2 1146 1148
0 452 5 1 1 1150
0 453 7 1 2 1143 452
0 454 5 1 1 453
0 455 7 1 2 1144 1151
0 456 5 1 1 455
0 457 7 3 2 454 456
0 458 5 2 1 1152
0 459 7 1 2 442 1153
0 460 5 1 1 459
0 461 7 1 2 870 1155
0 462 5 2 1 461
0 463 7 1 2 1140 1157
0 464 5 1 1 463
0 465 7 1 2 811 464
0 466 5 1 1 465
0 467 7 1 2 809 434
0 468 5 1 1 467
0 469 7 1 2 866 1136
0 470 5 1 1 469
0 471 7 2 2 468 470
0 472 5 1 1 1159
0 473 7 2 2 1124 1133
0 474 5 1 1 1161
0 475 7 1 2 1128 474
0 476 5 1 1 475
0 477 7 2 2 1111 1120
0 478 5 1 1 1163
0 479 7 1 2 1117 478
0 480 5 1 1 479
0 481 7 2 2 1100 1107
0 482 5 1 1 1165
0 483 7 1 2 1104 482
0 484 5 1 1 483
0 485 7 2 2 1087 1096
0 486 5 1 1 1167
0 487 7 1 2 1093 486
0 488 5 1 1 487
0 489 7 2 2 1076 1083
0 490 5 1 1 1169
0 491 7 2 2 1063 1072
0 492 5 1 1 1171
0 493 7 2 2 1052 1059
0 494 5 1 1 1173
0 495 7 1 2 1056 494
0 496 5 1 1 495
0 497 7 2 2 1039 1048
0 498 5 1 1 1175
0 499 7 1 2 1045 498
0 500 5 1 1 499
0 501 7 2 2 1028 1035
0 502 5 1 1 1177
0 503 7 1 2 1032 502
0 504 5 1 1 503
0 505 7 1 2 780 1022
0 506 5 1 1 505
0 507 7 1 2 846 1024
0 508 5 1 1 507
0 509 7 2 2 506 508
0 510 5 1 1 1179
0 511 7 1 2 976 1180
0 512 5 1 1 511
0 513 7 2 2 1013 1015
0 514 5 1 1 1181
0 515 7 1 2 1019 514
0 516 5 1 1 515
0 517 7 1 2 842 1007
0 518 5 1 1 517
0 519 7 1 2 774 1009
0 520 5 1 1 519
0 521 7 2 2 518 520
0 522 5 1 1 1183
0 523 7 1 2 996 262
0 524 5 1 1 523
0 525 7 1 2 771 524
0 526 5 1 1 525
0 527 7 1 2 993 1005
0 528 5 1 1 527
0 529 7 1 2 768 260
0 530 5 2 1 529
0 531 7 1 2 840 1185
0 532 7 1 2 528 531
0 533 5 1 1 532
0 534 7 1 2 526 533
0 535 7 1 2 522 534
0 536 5 1 1 535
0 537 7 1 2 985 1184
0 538 5 1 1 537
0 539 7 1 2 536 538
0 540 7 1 2 1182 539
0 541 5 1 1 540
0 542 7 1 2 516 541
0 543 7 1 2 510 542
0 544 5 1 1 543
0 545 7 1 2 512 544
0 546 7 1 2 1178 545
0 547 5 1 1 546
0 548 7 1 2 504 547
0 549 7 1 2 1176 548
0 550 5 1 1 549
0 551 7 1 2 500 550
0 552 7 1 2 1174 551
0 553 5 1 1 552
0 554 7 1 2 496 553
0 555 5 1 1 554
0 556 7 1 2 1172 555
0 557 5 1 1 556
0 558 7 1 2 1067 492
0 559 5 1 1 558
0 560 7 1 2 557 559
0 561 5 1 1 560
0 562 7 1 2 1170 561
0 563 5 1 1 562
0 564 7 1 2 1080 490
0 565 5 1 1 564
0 566 7 1 2 563 565
0 567 7 1 2 1168 566
0 568 5 1 1 567
0 569 7 1 2 488 568
0 570 7 1 2 1166 569
0 571 5 1 1 570
0 572 7 1 2 484 571
0 573 7 1 2 1164 572
0 574 5 1 1 573
0 575 7 1 2 480 574
0 576 7 1 2 1162 575
0 577 5 1 1 576
0 578 7 1 2 476 577
0 579 7 1 2 1160 578
0 580 5 1 1 579
0 581 7 1 2 966 472
0 582 5 1 1 581
0 583 7 1 2 580 582
0 584 7 1 2 466 583
0 585 7 1 2 460 584
0 586 5 1 1 585
0 587 7 1 2 804 1118
0 588 5 1 1 587
0 589 7 1 2 862 1115
0 590 5 1 1 589
0 591 7 1 2 798 1094
0 592 5 1 1 591
0 593 7 1 2 858 1091
0 594 5 1 1 593
0 595 7 1 2 792 1070
0 596 5 1 1 595
0 597 7 1 2 854 1068
0 598 5 1 1 597
0 599 7 1 2 786 1046
0 600 5 1 1 599
0 601 7 1 2 850 1043
0 602 5 1 1 601
0 603 7 1 2 1000 1186
0 604 5 1 1 603
0 605 7 1 2 987 998
0 606 7 1 2 604 605
0 607 5 1 1 606
0 608 7 2 2 989 607
0 609 5 1 1 1187
0 610 7 1 2 844 1188
0 611 5 1 1 610
0 612 7 1 2 777 609
0 613 5 1 1 612
0 614 7 1 2 1020 613
0 615 5 1 1 614
0 616 7 1 2 611 615
0 617 7 1 2 980 616
0 618 5 1 1 617
0 619 7 2 2 978 618
0 620 5 1 1 1189
0 621 7 1 2 783 620
0 622 5 1 1 621
0 623 7 1 2 1033 622
0 624 5 1 1 623
0 625 7 1 2 848 1190
0 626 5 1 1 625
0 627 7 1 2 624 626
0 628 7 1 2 602 627
0 629 5 1 1 628
0 630 7 2 2 600 629
0 631 5 1 1 1191
0 632 7 1 2 789 631
0 633 5 1 1 632
0 634 7 1 2 1057 633
0 635 5 1 1 634
0 636 7 1 2 852 1192
0 637 5 1 1 636
0 638 7 1 2 635 637
0 639 7 1 2 598 638
0 640 5 1 1 639
0 641 7 2 2 596 640
0 642 5 1 1 1193
0 643 7 1 2 795 642
0 644 5 1 1 643
0 645 7 1 2 1081 644
0 646 5 1 1 645
0 647 7 1 2 856 1194
0 648 5 1 1 647
0 649 7 1 2 646 648
0 650 7 1 2 594 649
0 651 5 1 1 650
0 652 7 2 2 592 651
0 653 5 1 1 1195
0 654 7 1 2 801 653
0 655 5 1 1 654
0 656 7 1 2 1105 655
0 657 5 1 1 656
0 658 7 1 2 860 1196
0 659 5 1 1 658
0 660 7 1 2 657 659
0 661 7 1 2 590 660
0 662 5 1 1 661
0 663 7 2 2 588 662
0 664 5 1 1 1197
0 665 7 1 2 1131 664
0 666 5 1 1 665
0 667 7 1 2 864 666
0 668 5 1 1 667
0 669 7 1 2 1129 1198
0 670 5 1 1 669
0 671 7 1 2 668 670
0 672 5 1 1 671
0 673 7 1 2 970 672
0 674 5 1 1 673
0 675 7 2 2 968 674
0 676 5 1 1 1199
0 677 7 1 2 871 676
0 678 5 1 1 677
0 679 7 1 2 1141 1156
0 680 5 1 1 679
0 681 7 1 2 678 680
0 682 5 1 1 681
0 683 7 1 2 868 682
0 684 5 1 1 683
0 685 7 1 2 1145 1149
0 686 5 1 1 685
0 687 7 2 2 1147 686
0 688 5 1 1 1201
0 689 7 1 2 1158 688
0 690 5 1 1 689
0 691 7 1 2 812 1154
0 692 5 1 1 691
0 693 7 1 2 814 692
0 694 5 1 1 693
0 695 7 1 2 1202 694
0 696 5 1 1 695
0 697 7 1 2 1138 1200
0 698 7 1 2 696 697
0 699 5 1 1 698
0 700 7 1 2 690 699
0 701 5 1 1 700
0 702 7 1 2 684 701
0 703 7 1 2 586 702
3 3499 5 0 1 703
