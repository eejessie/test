1 0 0 273 0
2 25 1 0
2 26 1 0
2 57275 1 0
2 57276 1 0
2 57277 1 0
2 57278 1 0
2 57279 1 0
2 57280 1 0
2 57281 1 0
2 57282 1 0
2 57283 1 0
2 57284 1 0
2 57285 1 0
2 57286 1 0
2 57287 1 0
2 57288 1 0
2 57289 1 0
2 57290 1 0
2 57291 1 0
2 57292 1 0
2 57293 1 0
2 57294 1 0
2 57295 1 0
2 57296 1 0
2 57297 1 0
2 57298 1 0
2 57299 1 0
2 57300 1 0
2 57301 1 0
2 57302 1 0
2 57303 1 0
2 57304 1 0
2 57305 1 0
2 57306 1 0
2 57307 1 0
2 57308 1 0
2 57309 1 0
2 57310 1 0
2 57311 1 0
2 57312 1 0
2 57313 1 0
2 57314 1 0
2 57315 1 0
2 57316 1 0
2 57317 1 0
2 57318 1 0
2 57319 1 0
2 57320 1 0
2 57321 1 0
2 57322 1 0
2 57323 1 0
2 57324 1 0
2 57325 1 0
2 57326 1 0
2 57327 1 0
2 57328 1 0
2 57329 1 0
2 57330 1 0
2 57331 1 0
2 57332 1 0
2 57333 1 0
2 57334 1 0
2 57335 1 0
2 57336 1 0
2 57337 1 0
2 57338 1 0
2 57339 1 0
2 57340 1 0
2 57341 1 0
2 57342 1 0
2 57343 1 0
2 57344 1 0
2 57345 1 0
2 57346 1 0
2 57347 1 0
2 57348 1 0
2 57349 1 0
2 57350 1 0
2 57351 1 0
2 57352 1 0
2 57353 1 0
2 57354 1 0
2 57355 1 0
2 57356 1 0
2 57357 1 0
2 57358 1 0
2 57359 1 0
2 57360 1 0
2 57361 1 0
2 57362 1 0
2 57363 1 0
2 57364 1 0
2 57365 1 0
2 57366 1 0
2 57367 1 0
2 57368 1 0
2 57369 1 0
2 57370 1 0
2 57371 1 0
2 57372 1 0
2 57373 1 0
2 57374 1 0
2 57375 1 0
2 57376 1 0
2 57377 1 0
2 57378 1 0
2 57379 1 0
2 57380 1 0
2 57381 1 0
2 57382 1 0
2 57383 1 0
2 57384 1 0
2 57385 1 0
2 57386 1 0
2 57387 1 0
2 57388 1 0
2 57389 1 0
2 57390 1 0
2 57391 1 0
2 57392 1 0
2 57393 1 0
2 57394 1 0
2 57395 1 0
2 57396 1 0
2 57397 1 0
2 57398 1 0
2 57399 1 0
2 57400 1 0
2 57401 1 0
2 57402 1 0
2 57403 1 0
2 57404 1 0
2 57405 1 0
2 57406 1 0
2 57407 1 0
2 57408 1 0
2 57409 1 0
2 57410 1 0
2 57411 1 0
2 57412 1 0
2 57413 1 0
2 57414 1 0
2 57415 1 0
2 57416 1 0
2 57417 1 0
2 57418 1 0
2 57419 1 0
2 57420 1 0
2 57421 1 0
2 57422 1 0
2 57423 1 0
2 57424 1 0
2 57425 1 0
2 57426 1 0
2 57427 1 0
2 57428 1 0
2 57429 1 0
2 57430 1 0
2 57431 1 0
2 57432 1 0
2 57433 1 0
2 57434 1 0
2 57435 1 0
2 57436 1 0
2 57437 1 0
2 57438 1 0
2 57439 1 0
2 57440 1 0
2 57441 1 0
2 57442 1 0
2 57443 1 0
2 57444 1 0
2 57445 1 0
2 57446 1 0
2 57447 1 0
2 57448 1 0
2 57449 1 0
2 57450 1 0
2 57451 1 0
2 57452 1 0
2 57453 1 0
2 57454 1 0
2 57455 1 0
2 57456 1 0
2 57457 1 0
2 57458 1 0
2 57459 1 0
2 57460 1 0
2 57461 1 0
2 57462 1 0
2 57463 1 0
2 57464 1 0
2 57465 1 0
2 57466 1 0
2 57467 1 0
2 57468 1 0
2 57469 1 0
2 57470 1 0
2 57471 1 0
2 57472 1 0
2 57473 1 0
2 57474 1 0
2 57475 1 0
2 57476 1 0
2 57477 1 0
2 57478 1 0
2 57479 1 0
2 57480 1 0
2 57481 1 0
2 57482 1 0
2 57483 1 0
2 57484 1 0
2 57485 1 0
2 57486 1 0
2 57487 1 0
2 57488 1 0
2 57489 1 0
2 57490 1 0
2 57491 1 0
2 57492 1 0
2 57493 1 0
2 57494 1 0
2 57495 1 0
2 57496 1 0
2 57497 1 0
2 57498 1 0
2 57499 1 0
2 57500 1 0
2 57501 1 0
2 57502 1 0
2 57503 1 0
2 57504 1 0
2 57505 1 0
2 57506 1 0
2 57507 1 0
2 57508 1 0
2 57509 1 0
2 57510 1 0
2 57511 1 0
2 57512 1 0
2 57513 1 0
2 57514 1 0
2 57515 1 0
2 57516 1 0
2 57517 1 0
2 57518 1 0
2 57519 1 0
2 57520 1 0
2 57521 1 0
2 57522 1 0
2 57523 1 0
2 57524 1 0
2 57525 1 0
2 57526 1 0
2 57527 1 0
2 57528 1 0
2 57529 1 0
2 57530 1 0
2 57531 1 0
2 57532 1 0
2 57533 1 0
2 57534 1 0
2 57535 1 0
2 57536 1 0
2 57537 1 0
2 57538 1 0
2 57539 1 0
2 57540 1 0
2 57541 1 0
2 57542 1 0
2 57543 1 0
2 57544 1 0
2 57545 1 0
1 1 0 277 0
2 57546 1 1
2 57547 1 1
2 57548 1 1
2 57549 1 1
2 57550 1 1
2 57551 1 1
2 57552 1 1
2 57553 1 1
2 57554 1 1
2 57555 1 1
2 57556 1 1
2 57557 1 1
2 57558 1 1
2 57559 1 1
2 57560 1 1
2 57561 1 1
2 57562 1 1
2 57563 1 1
2 57564 1 1
2 57565 1 1
2 57566 1 1
2 57567 1 1
2 57568 1 1
2 57569 1 1
2 57570 1 1
2 57571 1 1
2 57572 1 1
2 57573 1 1
2 57574 1 1
2 57575 1 1
2 57576 1 1
2 57577 1 1
2 57578 1 1
2 57579 1 1
2 57580 1 1
2 57581 1 1
2 57582 1 1
2 57583 1 1
2 57584 1 1
2 57585 1 1
2 57586 1 1
2 57587 1 1
2 57588 1 1
2 57589 1 1
2 57590 1 1
2 57591 1 1
2 57592 1 1
2 57593 1 1
2 57594 1 1
2 57595 1 1
2 57596 1 1
2 57597 1 1
2 57598 1 1
2 57599 1 1
2 57600 1 1
2 57601 1 1
2 57602 1 1
2 57603 1 1
2 57604 1 1
2 57605 1 1
2 57606 1 1
2 57607 1 1
2 57608 1 1
2 57609 1 1
2 57610 1 1
2 57611 1 1
2 57612 1 1
2 57613 1 1
2 57614 1 1
2 57615 1 1
2 57616 1 1
2 57617 1 1
2 57618 1 1
2 57619 1 1
2 57620 1 1
2 57621 1 1
2 57622 1 1
2 57623 1 1
2 57624 1 1
2 57625 1 1
2 57626 1 1
2 57627 1 1
2 57628 1 1
2 57629 1 1
2 57630 1 1
2 57631 1 1
2 57632 1 1
2 57633 1 1
2 57634 1 1
2 57635 1 1
2 57636 1 1
2 57637 1 1
2 57638 1 1
2 57639 1 1
2 57640 1 1
2 57641 1 1
2 57642 1 1
2 57643 1 1
2 57644 1 1
2 57645 1 1
2 57646 1 1
2 57647 1 1
2 57648 1 1
2 57649 1 1
2 57650 1 1
2 57651 1 1
2 57652 1 1
2 57653 1 1
2 57654 1 1
2 57655 1 1
2 57656 1 1
2 57657 1 1
2 57658 1 1
2 57659 1 1
2 57660 1 1
2 57661 1 1
2 57662 1 1
2 57663 1 1
2 57664 1 1
2 57665 1 1
2 57666 1 1
2 57667 1 1
2 57668 1 1
2 57669 1 1
2 57670 1 1
2 57671 1 1
2 57672 1 1
2 57673 1 1
2 57674 1 1
2 57675 1 1
2 57676 1 1
2 57677 1 1
2 57678 1 1
2 57679 1 1
2 57680 1 1
2 57681 1 1
2 57682 1 1
2 57683 1 1
2 57684 1 1
2 57685 1 1
2 57686 1 1
2 57687 1 1
2 57688 1 1
2 57689 1 1
2 57690 1 1
2 57691 1 1
2 57692 1 1
2 57693 1 1
2 57694 1 1
2 57695 1 1
2 57696 1 1
2 57697 1 1
2 57698 1 1
2 57699 1 1
2 57700 1 1
2 57701 1 1
2 57702 1 1
2 57703 1 1
2 57704 1 1
2 57705 1 1
2 57706 1 1
2 57707 1 1
2 57708 1 1
2 57709 1 1
2 57710 1 1
2 57711 1 1
2 57712 1 1
2 57713 1 1
2 57714 1 1
2 57715 1 1
2 57716 1 1
2 57717 1 1
2 57718 1 1
2 57719 1 1
2 57720 1 1
2 57721 1 1
2 57722 1 1
2 57723 1 1
2 57724 1 1
2 57725 1 1
2 57726 1 1
2 57727 1 1
2 57728 1 1
2 57729 1 1
2 57730 1 1
2 57731 1 1
2 57732 1 1
2 57733 1 1
2 57734 1 1
2 57735 1 1
2 57736 1 1
2 57737 1 1
2 57738 1 1
2 57739 1 1
2 57740 1 1
2 57741 1 1
2 57742 1 1
2 57743 1 1
2 57744 1 1
2 57745 1 1
2 57746 1 1
2 57747 1 1
2 57748 1 1
2 57749 1 1
2 57750 1 1
2 57751 1 1
2 57752 1 1
2 57753 1 1
2 57754 1 1
2 57755 1 1
2 57756 1 1
2 57757 1 1
2 57758 1 1
2 57759 1 1
2 57760 1 1
2 57761 1 1
2 57762 1 1
2 57763 1 1
2 57764 1 1
2 57765 1 1
2 57766 1 1
2 57767 1 1
2 57768 1 1
2 57769 1 1
2 57770 1 1
2 57771 1 1
2 57772 1 1
2 57773 1 1
2 57774 1 1
2 57775 1 1
2 57776 1 1
2 57777 1 1
2 57778 1 1
2 57779 1 1
2 57780 1 1
2 57781 1 1
2 57782 1 1
2 57783 1 1
2 57784 1 1
2 57785 1 1
2 57786 1 1
2 57787 1 1
2 57788 1 1
2 57789 1 1
2 57790 1 1
2 57791 1 1
2 57792 1 1
2 57793 1 1
2 57794 1 1
2 57795 1 1
2 57796 1 1
2 57797 1 1
2 57798 1 1
2 57799 1 1
2 57800 1 1
2 57801 1 1
2 57802 1 1
2 57803 1 1
2 57804 1 1
2 57805 1 1
2 57806 1 1
2 57807 1 1
2 57808 1 1
2 57809 1 1
2 57810 1 1
2 57811 1 1
2 57812 1 1
2 57813 1 1
2 57814 1 1
2 57815 1 1
2 57816 1 1
2 57817 1 1
2 57818 1 1
2 57819 1 1
2 57820 1 1
2 57821 1 1
2 57822 1 1
1 2 0 278 0
2 57823 1 2
2 57824 1 2
2 57825 1 2
2 57826 1 2
2 57827 1 2
2 57828 1 2
2 57829 1 2
2 57830 1 2
2 57831 1 2
2 57832 1 2
2 57833 1 2
2 57834 1 2
2 57835 1 2
2 57836 1 2
2 57837 1 2
2 57838 1 2
2 57839 1 2
2 57840 1 2
2 57841 1 2
2 57842 1 2
2 57843 1 2
2 57844 1 2
2 57845 1 2
2 57846 1 2
2 57847 1 2
2 57848 1 2
2 57849 1 2
2 57850 1 2
2 57851 1 2
2 57852 1 2
2 57853 1 2
2 57854 1 2
2 57855 1 2
2 57856 1 2
2 57857 1 2
2 57858 1 2
2 57859 1 2
2 57860 1 2
2 57861 1 2
2 57862 1 2
2 57863 1 2
2 57864 1 2
2 57865 1 2
2 57866 1 2
2 57867 1 2
2 57868 1 2
2 57869 1 2
2 57870 1 2
2 57871 1 2
2 57872 1 2
2 57873 1 2
2 57874 1 2
2 57875 1 2
2 57876 1 2
2 57877 1 2
2 57878 1 2
2 57879 1 2
2 57880 1 2
2 57881 1 2
2 57882 1 2
2 57883 1 2
2 57884 1 2
2 57885 1 2
2 57886 1 2
2 57887 1 2
2 57888 1 2
2 57889 1 2
2 57890 1 2
2 57891 1 2
2 57892 1 2
2 57893 1 2
2 57894 1 2
2 57895 1 2
2 57896 1 2
2 57897 1 2
2 57898 1 2
2 57899 1 2
2 57900 1 2
2 57901 1 2
2 57902 1 2
2 57903 1 2
2 57904 1 2
2 57905 1 2
2 57906 1 2
2 57907 1 2
2 57908 1 2
2 57909 1 2
2 57910 1 2
2 57911 1 2
2 57912 1 2
2 57913 1 2
2 57914 1 2
2 57915 1 2
2 57916 1 2
2 57917 1 2
2 57918 1 2
2 57919 1 2
2 57920 1 2
2 57921 1 2
2 57922 1 2
2 57923 1 2
2 57924 1 2
2 57925 1 2
2 57926 1 2
2 57927 1 2
2 57928 1 2
2 57929 1 2
2 57930 1 2
2 57931 1 2
2 57932 1 2
2 57933 1 2
2 57934 1 2
2 57935 1 2
2 57936 1 2
2 57937 1 2
2 57938 1 2
2 57939 1 2
2 57940 1 2
2 57941 1 2
2 57942 1 2
2 57943 1 2
2 57944 1 2
2 57945 1 2
2 57946 1 2
2 57947 1 2
2 57948 1 2
2 57949 1 2
2 57950 1 2
2 57951 1 2
2 57952 1 2
2 57953 1 2
2 57954 1 2
2 57955 1 2
2 57956 1 2
2 57957 1 2
2 57958 1 2
2 57959 1 2
2 57960 1 2
2 57961 1 2
2 57962 1 2
2 57963 1 2
2 57964 1 2
2 57965 1 2
2 57966 1 2
2 57967 1 2
2 57968 1 2
2 57969 1 2
2 57970 1 2
2 57971 1 2
2 57972 1 2
2 57973 1 2
2 57974 1 2
2 57975 1 2
2 57976 1 2
2 57977 1 2
2 57978 1 2
2 57979 1 2
2 57980 1 2
2 57981 1 2
2 57982 1 2
2 57983 1 2
2 57984 1 2
2 57985 1 2
2 57986 1 2
2 57987 1 2
2 57988 1 2
2 57989 1 2
2 57990 1 2
2 57991 1 2
2 57992 1 2
2 57993 1 2
2 57994 1 2
2 57995 1 2
2 57996 1 2
2 57997 1 2
2 57998 1 2
2 57999 1 2
2 58000 1 2
2 58001 1 2
2 58002 1 2
2 58003 1 2
2 58004 1 2
2 58005 1 2
2 58006 1 2
2 58007 1 2
2 58008 1 2
2 58009 1 2
2 58010 1 2
2 58011 1 2
2 58012 1 2
2 58013 1 2
2 58014 1 2
2 58015 1 2
2 58016 1 2
2 58017 1 2
2 58018 1 2
2 58019 1 2
2 58020 1 2
2 58021 1 2
2 58022 1 2
2 58023 1 2
2 58024 1 2
2 58025 1 2
2 58026 1 2
2 58027 1 2
2 58028 1 2
2 58029 1 2
2 58030 1 2
2 58031 1 2
2 58032 1 2
2 58033 1 2
2 58034 1 2
2 58035 1 2
2 58036 1 2
2 58037 1 2
2 58038 1 2
2 58039 1 2
2 58040 1 2
2 58041 1 2
2 58042 1 2
2 58043 1 2
2 58044 1 2
2 58045 1 2
2 58046 1 2
2 58047 1 2
2 58048 1 2
2 58049 1 2
2 58050 1 2
2 58051 1 2
2 58052 1 2
2 58053 1 2
2 58054 1 2
2 58055 1 2
2 58056 1 2
2 58057 1 2
2 58058 1 2
2 58059 1 2
2 58060 1 2
2 58061 1 2
2 58062 1 2
2 58063 1 2
2 58064 1 2
2 58065 1 2
2 58066 1 2
2 58067 1 2
2 58068 1 2
2 58069 1 2
2 58070 1 2
2 58071 1 2
2 58072 1 2
2 58073 1 2
2 58074 1 2
2 58075 1 2
2 58076 1 2
2 58077 1 2
2 58078 1 2
2 58079 1 2
2 58080 1 2
2 58081 1 2
2 58082 1 2
2 58083 1 2
2 58084 1 2
2 58085 1 2
2 58086 1 2
2 58087 1 2
2 58088 1 2
2 58089 1 2
2 58090 1 2
2 58091 1 2
2 58092 1 2
2 58093 1 2
2 58094 1 2
2 58095 1 2
2 58096 1 2
2 58097 1 2
2 58098 1 2
2 58099 1 2
2 58100 1 2
1 3 0 275 0
2 58101 1 3
2 58102 1 3
2 58103 1 3
2 58104 1 3
2 58105 1 3
2 58106 1 3
2 58107 1 3
2 58108 1 3
2 58109 1 3
2 58110 1 3
2 58111 1 3
2 58112 1 3
2 58113 1 3
2 58114 1 3
2 58115 1 3
2 58116 1 3
2 58117 1 3
2 58118 1 3
2 58119 1 3
2 58120 1 3
2 58121 1 3
2 58122 1 3
2 58123 1 3
2 58124 1 3
2 58125 1 3
2 58126 1 3
2 58127 1 3
2 58128 1 3
2 58129 1 3
2 58130 1 3
2 58131 1 3
2 58132 1 3
2 58133 1 3
2 58134 1 3
2 58135 1 3
2 58136 1 3
2 58137 1 3
2 58138 1 3
2 58139 1 3
2 58140 1 3
2 58141 1 3
2 58142 1 3
2 58143 1 3
2 58144 1 3
2 58145 1 3
2 58146 1 3
2 58147 1 3
2 58148 1 3
2 58149 1 3
2 58150 1 3
2 58151 1 3
2 58152 1 3
2 58153 1 3
2 58154 1 3
2 58155 1 3
2 58156 1 3
2 58157 1 3
2 58158 1 3
2 58159 1 3
2 58160 1 3
2 58161 1 3
2 58162 1 3
2 58163 1 3
2 58164 1 3
2 58165 1 3
2 58166 1 3
2 58167 1 3
2 58168 1 3
2 58169 1 3
2 58170 1 3
2 58171 1 3
2 58172 1 3
2 58173 1 3
2 58174 1 3
2 58175 1 3
2 58176 1 3
2 58177 1 3
2 58178 1 3
2 58179 1 3
2 58180 1 3
2 58181 1 3
2 58182 1 3
2 58183 1 3
2 58184 1 3
2 58185 1 3
2 58186 1 3
2 58187 1 3
2 58188 1 3
2 58189 1 3
2 58190 1 3
2 58191 1 3
2 58192 1 3
2 58193 1 3
2 58194 1 3
2 58195 1 3
2 58196 1 3
2 58197 1 3
2 58198 1 3
2 58199 1 3
2 58200 1 3
2 58201 1 3
2 58202 1 3
2 58203 1 3
2 58204 1 3
2 58205 1 3
2 58206 1 3
2 58207 1 3
2 58208 1 3
2 58209 1 3
2 58210 1 3
2 58211 1 3
2 58212 1 3
2 58213 1 3
2 58214 1 3
2 58215 1 3
2 58216 1 3
2 58217 1 3
2 58218 1 3
2 58219 1 3
2 58220 1 3
2 58221 1 3
2 58222 1 3
2 58223 1 3
2 58224 1 3
2 58225 1 3
2 58226 1 3
2 58227 1 3
2 58228 1 3
2 58229 1 3
2 58230 1 3
2 58231 1 3
2 58232 1 3
2 58233 1 3
2 58234 1 3
2 58235 1 3
2 58236 1 3
2 58237 1 3
2 58238 1 3
2 58239 1 3
2 58240 1 3
2 58241 1 3
2 58242 1 3
2 58243 1 3
2 58244 1 3
2 58245 1 3
2 58246 1 3
2 58247 1 3
2 58248 1 3
2 58249 1 3
2 58250 1 3
2 58251 1 3
2 58252 1 3
2 58253 1 3
2 58254 1 3
2 58255 1 3
2 58256 1 3
2 58257 1 3
2 58258 1 3
2 58259 1 3
2 58260 1 3
2 58261 1 3
2 58262 1 3
2 58263 1 3
2 58264 1 3
2 58265 1 3
2 58266 1 3
2 58267 1 3
2 58268 1 3
2 58269 1 3
2 58270 1 3
2 58271 1 3
2 58272 1 3
2 58273 1 3
2 58274 1 3
2 58275 1 3
2 58276 1 3
2 58277 1 3
2 58278 1 3
2 58279 1 3
2 58280 1 3
2 58281 1 3
2 58282 1 3
2 58283 1 3
2 58284 1 3
2 58285 1 3
2 58286 1 3
2 58287 1 3
2 58288 1 3
2 58289 1 3
2 58290 1 3
2 58291 1 3
2 58292 1 3
2 58293 1 3
2 58294 1 3
2 58295 1 3
2 58296 1 3
2 58297 1 3
2 58298 1 3
2 58299 1 3
2 58300 1 3
2 58301 1 3
2 58302 1 3
2 58303 1 3
2 58304 1 3
2 58305 1 3
2 58306 1 3
2 58307 1 3
2 58308 1 3
2 58309 1 3
2 58310 1 3
2 58311 1 3
2 58312 1 3
2 58313 1 3
2 58314 1 3
2 58315 1 3
2 58316 1 3
2 58317 1 3
2 58318 1 3
2 58319 1 3
2 58320 1 3
2 58321 1 3
2 58322 1 3
2 58323 1 3
2 58324 1 3
2 58325 1 3
2 58326 1 3
2 58327 1 3
2 58328 1 3
2 58329 1 3
2 58330 1 3
2 58331 1 3
2 58332 1 3
2 58333 1 3
2 58334 1 3
2 58335 1 3
2 58336 1 3
2 58337 1 3
2 58338 1 3
2 58339 1 3
2 58340 1 3
2 58341 1 3
2 58342 1 3
2 58343 1 3
2 58344 1 3
2 58345 1 3
2 58346 1 3
2 58347 1 3
2 58348 1 3
2 58349 1 3
2 58350 1 3
2 58351 1 3
2 58352 1 3
2 58353 1 3
2 58354 1 3
2 58355 1 3
2 58356 1 3
2 58357 1 3
2 58358 1 3
2 58359 1 3
2 58360 1 3
2 58361 1 3
2 58362 1 3
2 58363 1 3
2 58364 1 3
2 58365 1 3
2 58366 1 3
2 58367 1 3
2 58368 1 3
2 58369 1 3
2 58370 1 3
2 58371 1 3
2 58372 1 3
2 58373 1 3
2 58374 1 3
2 58375 1 3
1 4 0 323 0
2 58376 1 4
2 58377 1 4
2 58378 1 4
2 58379 1 4
2 58380 1 4
2 58381 1 4
2 58382 1 4
2 58383 1 4
2 58384 1 4
2 58385 1 4
2 58386 1 4
2 58387 1 4
2 58388 1 4
2 58389 1 4
2 58390 1 4
2 58391 1 4
2 58392 1 4
2 58393 1 4
2 58394 1 4
2 58395 1 4
2 58396 1 4
2 58397 1 4
2 58398 1 4
2 58399 1 4
2 58400 1 4
2 58401 1 4
2 58402 1 4
2 58403 1 4
2 58404 1 4
2 58405 1 4
2 58406 1 4
2 58407 1 4
2 58408 1 4
2 58409 1 4
2 58410 1 4
2 58411 1 4
2 58412 1 4
2 58413 1 4
2 58414 1 4
2 58415 1 4
2 58416 1 4
2 58417 1 4
2 58418 1 4
2 58419 1 4
2 58420 1 4
2 58421 1 4
2 58422 1 4
2 58423 1 4
2 58424 1 4
2 58425 1 4
2 58426 1 4
2 58427 1 4
2 58428 1 4
2 58429 1 4
2 58430 1 4
2 58431 1 4
2 58432 1 4
2 58433 1 4
2 58434 1 4
2 58435 1 4
2 58436 1 4
2 58437 1 4
2 58438 1 4
2 58439 1 4
2 58440 1 4
2 58441 1 4
2 58442 1 4
2 58443 1 4
2 58444 1 4
2 58445 1 4
2 58446 1 4
2 58447 1 4
2 58448 1 4
2 58449 1 4
2 58450 1 4
2 58451 1 4
2 58452 1 4
2 58453 1 4
2 58454 1 4
2 58455 1 4
2 58456 1 4
2 58457 1 4
2 58458 1 4
2 58459 1 4
2 58460 1 4
2 58461 1 4
2 58462 1 4
2 58463 1 4
2 58464 1 4
2 58465 1 4
2 58466 1 4
2 58467 1 4
2 58468 1 4
2 58469 1 4
2 58470 1 4
2 58471 1 4
2 58472 1 4
2 58473 1 4
2 58474 1 4
2 58475 1 4
2 58476 1 4
2 58477 1 4
2 58478 1 4
2 58479 1 4
2 58480 1 4
2 58481 1 4
2 58482 1 4
2 58483 1 4
2 58484 1 4
2 58485 1 4
2 58486 1 4
2 58487 1 4
2 58488 1 4
2 58489 1 4
2 58490 1 4
2 58491 1 4
2 58492 1 4
2 58493 1 4
2 58494 1 4
2 58495 1 4
2 58496 1 4
2 58497 1 4
2 58498 1 4
2 58499 1 4
2 58500 1 4
2 58501 1 4
2 58502 1 4
2 58503 1 4
2 58504 1 4
2 58505 1 4
2 58506 1 4
2 58507 1 4
2 58508 1 4
2 58509 1 4
2 58510 1 4
2 58511 1 4
2 58512 1 4
2 58513 1 4
2 58514 1 4
2 58515 1 4
2 58516 1 4
2 58517 1 4
2 58518 1 4
2 58519 1 4
2 58520 1 4
2 58521 1 4
2 58522 1 4
2 58523 1 4
2 58524 1 4
2 58525 1 4
2 58526 1 4
2 58527 1 4
2 58528 1 4
2 58529 1 4
2 58530 1 4
2 58531 1 4
2 58532 1 4
2 58533 1 4
2 58534 1 4
2 58535 1 4
2 58536 1 4
2 58537 1 4
2 58538 1 4
2 58539 1 4
2 58540 1 4
2 58541 1 4
2 58542 1 4
2 58543 1 4
2 58544 1 4
2 58545 1 4
2 58546 1 4
2 58547 1 4
2 58548 1 4
2 58549 1 4
2 58550 1 4
2 58551 1 4
2 58552 1 4
2 58553 1 4
2 58554 1 4
2 58555 1 4
2 58556 1 4
2 58557 1 4
2 58558 1 4
2 58559 1 4
2 58560 1 4
2 58561 1 4
2 58562 1 4
2 58563 1 4
2 58564 1 4
2 58565 1 4
2 58566 1 4
2 58567 1 4
2 58568 1 4
2 58569 1 4
2 58570 1 4
2 58571 1 4
2 58572 1 4
2 58573 1 4
2 58574 1 4
2 58575 1 4
2 58576 1 4
2 58577 1 4
2 58578 1 4
2 58579 1 4
2 58580 1 4
2 58581 1 4
2 58582 1 4
2 58583 1 4
2 58584 1 4
2 58585 1 4
2 58586 1 4
2 58587 1 4
2 58588 1 4
2 58589 1 4
2 58590 1 4
2 58591 1 4
2 58592 1 4
2 58593 1 4
2 58594 1 4
2 58595 1 4
2 58596 1 4
2 58597 1 4
2 58598 1 4
2 58599 1 4
2 58600 1 4
2 58601 1 4
2 58602 1 4
2 58603 1 4
2 58604 1 4
2 58605 1 4
2 58606 1 4
2 58607 1 4
2 58608 1 4
2 58609 1 4
2 58610 1 4
2 58611 1 4
2 58612 1 4
2 58613 1 4
2 58614 1 4
2 58615 1 4
2 58616 1 4
2 58617 1 4
2 58618 1 4
2 58619 1 4
2 58620 1 4
2 58621 1 4
2 58622 1 4
2 58623 1 4
2 58624 1 4
2 58625 1 4
2 58626 1 4
2 58627 1 4
2 58628 1 4
2 58629 1 4
2 58630 1 4
2 58631 1 4
2 58632 1 4
2 58633 1 4
2 58634 1 4
2 58635 1 4
2 58636 1 4
2 58637 1 4
2 58638 1 4
2 58639 1 4
2 58640 1 4
2 58641 1 4
2 58642 1 4
2 58643 1 4
2 58644 1 4
2 58645 1 4
2 58646 1 4
2 58647 1 4
2 58648 1 4
2 58649 1 4
2 58650 1 4
2 58651 1 4
2 58652 1 4
2 58653 1 4
2 58654 1 4
2 58655 1 4
2 58656 1 4
2 58657 1 4
2 58658 1 4
2 58659 1 4
2 58660 1 4
2 58661 1 4
2 58662 1 4
2 58663 1 4
2 58664 1 4
2 58665 1 4
2 58666 1 4
2 58667 1 4
2 58668 1 4
2 58669 1 4
2 58670 1 4
2 58671 1 4
2 58672 1 4
2 58673 1 4
2 58674 1 4
2 58675 1 4
2 58676 1 4
2 58677 1 4
2 58678 1 4
2 58679 1 4
2 58680 1 4
2 58681 1 4
2 58682 1 4
2 58683 1 4
2 58684 1 4
2 58685 1 4
2 58686 1 4
2 58687 1 4
2 58688 1 4
2 58689 1 4
2 58690 1 4
2 58691 1 4
2 58692 1 4
2 58693 1 4
2 58694 1 4
2 58695 1 4
2 58696 1 4
2 58697 1 4
2 58698 1 4
1 5 0 122 0
2 58699 1 5
2 58700 1 5
2 58701 1 5
2 58702 1 5
2 58703 1 5
2 58704 1 5
2 58705 1 5
2 58706 1 5
2 58707 1 5
2 58708 1 5
2 58709 1 5
2 58710 1 5
2 58711 1 5
2 58712 1 5
2 58713 1 5
2 58714 1 5
2 58715 1 5
2 58716 1 5
2 58717 1 5
2 58718 1 5
2 58719 1 5
2 58720 1 5
2 58721 1 5
2 58722 1 5
2 58723 1 5
2 58724 1 5
2 58725 1 5
2 58726 1 5
2 58727 1 5
2 58728 1 5
2 58729 1 5
2 58730 1 5
2 58731 1 5
2 58732 1 5
2 58733 1 5
2 58734 1 5
2 58735 1 5
2 58736 1 5
2 58737 1 5
2 58738 1 5
2 58739 1 5
2 58740 1 5
2 58741 1 5
2 58742 1 5
2 58743 1 5
2 58744 1 5
2 58745 1 5
2 58746 1 5
2 58747 1 5
2 58748 1 5
2 58749 1 5
2 58750 1 5
2 58751 1 5
2 58752 1 5
2 58753 1 5
2 58754 1 5
2 58755 1 5
2 58756 1 5
2 58757 1 5
2 58758 1 5
2 58759 1 5
2 58760 1 5
2 58761 1 5
2 58762 1 5
2 58763 1 5
2 58764 1 5
2 58765 1 5
2 58766 1 5
2 58767 1 5
2 58768 1 5
2 58769 1 5
2 58770 1 5
2 58771 1 5
2 58772 1 5
2 58773 1 5
2 58774 1 5
2 58775 1 5
2 58776 1 5
2 58777 1 5
2 58778 1 5
2 58779 1 5
2 58780 1 5
2 58781 1 5
2 58782 1 5
2 58783 1 5
2 58784 1 5
2 58785 1 5
2 58786 1 5
2 58787 1 5
2 58788 1 5
2 58789 1 5
2 58790 1 5
2 58791 1 5
2 58792 1 5
2 58793 1 5
2 58794 1 5
2 58795 1 5
2 58796 1 5
2 58797 1 5
2 58798 1 5
2 58799 1 5
2 58800 1 5
2 58801 1 5
2 58802 1 5
2 58803 1 5
2 58804 1 5
2 58805 1 5
2 58806 1 5
2 58807 1 5
2 58808 1 5
2 58809 1 5
2 58810 1 5
2 58811 1 5
2 58812 1 5
2 58813 1 5
2 58814 1 5
2 58815 1 5
2 58816 1 5
2 58817 1 5
2 58818 1 5
2 58819 1 5
2 58820 1 5
1 6 0 84 0
2 58821 1 6
2 58822 1 6
2 58823 1 6
2 58824 1 6
2 58825 1 6
2 58826 1 6
2 58827 1 6
2 58828 1 6
2 58829 1 6
2 58830 1 6
2 58831 1 6
2 58832 1 6
2 58833 1 6
2 58834 1 6
2 58835 1 6
2 58836 1 6
2 58837 1 6
2 58838 1 6
2 58839 1 6
2 58840 1 6
2 58841 1 6
2 58842 1 6
2 58843 1 6
2 58844 1 6
2 58845 1 6
2 58846 1 6
2 58847 1 6
2 58848 1 6
2 58849 1 6
2 58850 1 6
2 58851 1 6
2 58852 1 6
2 58853 1 6
2 58854 1 6
2 58855 1 6
2 58856 1 6
2 58857 1 6
2 58858 1 6
2 58859 1 6
2 58860 1 6
2 58861 1 6
2 58862 1 6
2 58863 1 6
2 58864 1 6
2 58865 1 6
2 58866 1 6
2 58867 1 6
2 58868 1 6
2 58869 1 6
2 58870 1 6
2 58871 1 6
2 58872 1 6
2 58873 1 6
2 58874 1 6
2 58875 1 6
2 58876 1 6
2 58877 1 6
2 58878 1 6
2 58879 1 6
2 58880 1 6
2 58881 1 6
2 58882 1 6
2 58883 1 6
2 58884 1 6
2 58885 1 6
2 58886 1 6
2 58887 1 6
2 58888 1 6
2 58889 1 6
2 58890 1 6
2 58891 1 6
2 58892 1 6
2 58893 1 6
2 58894 1 6
2 58895 1 6
2 58896 1 6
2 58897 1 6
2 58898 1 6
2 58899 1 6
2 58900 1 6
2 58901 1 6
2 58902 1 6
2 58903 1 6
2 58904 1 6
1 7 0 13 0
2 58905 1 7
2 58906 1 7
2 58907 1 7
2 58908 1 7
2 58909 1 7
2 58910 1 7
2 58911 1 7
2 58912 1 7
2 58913 1 7
2 58914 1 7
2 58915 1 7
2 58916 1 7
2 58917 1 7
1 8 0 121 0
2 58918 1 8
2 58919 1 8
2 58920 1 8
2 58921 1 8
2 58922 1 8
2 58923 1 8
2 58924 1 8
2 58925 1 8
2 58926 1 8
2 58927 1 8
2 58928 1 8
2 58929 1 8
2 58930 1 8
2 58931 1 8
2 58932 1 8
2 58933 1 8
2 58934 1 8
2 58935 1 8
2 58936 1 8
2 58937 1 8
2 58938 1 8
2 58939 1 8
2 58940 1 8
2 58941 1 8
2 58942 1 8
2 58943 1 8
2 58944 1 8
2 58945 1 8
2 58946 1 8
2 58947 1 8
2 58948 1 8
2 58949 1 8
2 58950 1 8
2 58951 1 8
2 58952 1 8
2 58953 1 8
2 58954 1 8
2 58955 1 8
2 58956 1 8
2 58957 1 8
2 58958 1 8
2 58959 1 8
2 58960 1 8
2 58961 1 8
2 58962 1 8
2 58963 1 8
2 58964 1 8
2 58965 1 8
2 58966 1 8
2 58967 1 8
2 58968 1 8
2 58969 1 8
2 58970 1 8
2 58971 1 8
2 58972 1 8
2 58973 1 8
2 58974 1 8
2 58975 1 8
2 58976 1 8
2 58977 1 8
2 58978 1 8
2 58979 1 8
2 58980 1 8
2 58981 1 8
2 58982 1 8
2 58983 1 8
2 58984 1 8
2 58985 1 8
2 58986 1 8
2 58987 1 8
2 58988 1 8
2 58989 1 8
2 58990 1 8
2 58991 1 8
2 58992 1 8
2 58993 1 8
2 58994 1 8
2 58995 1 8
2 58996 1 8
2 58997 1 8
2 58998 1 8
2 58999 1 8
2 59000 1 8
2 59001 1 8
2 59002 1 8
2 59003 1 8
2 59004 1 8
2 59005 1 8
2 59006 1 8
2 59007 1 8
2 59008 1 8
2 59009 1 8
2 59010 1 8
2 59011 1 8
2 59012 1 8
2 59013 1 8
2 59014 1 8
2 59015 1 8
2 59016 1 8
2 59017 1 8
2 59018 1 8
2 59019 1 8
2 59020 1 8
2 59021 1 8
2 59022 1 8
2 59023 1 8
2 59024 1 8
2 59025 1 8
2 59026 1 8
2 59027 1 8
2 59028 1 8
2 59029 1 8
2 59030 1 8
2 59031 1 8
2 59032 1 8
2 59033 1 8
2 59034 1 8
2 59035 1 8
2 59036 1 8
2 59037 1 8
2 59038 1 8
1 9 0 140 0
2 59039 1 9
2 59040 1 9
2 59041 1 9
2 59042 1 9
2 59043 1 9
2 59044 1 9
2 59045 1 9
2 59046 1 9
2 59047 1 9
2 59048 1 9
2 59049 1 9
2 59050 1 9
2 59051 1 9
2 59052 1 9
2 59053 1 9
2 59054 1 9
2 59055 1 9
2 59056 1 9
2 59057 1 9
2 59058 1 9
2 59059 1 9
2 59060 1 9
2 59061 1 9
2 59062 1 9
2 59063 1 9
2 59064 1 9
2 59065 1 9
2 59066 1 9
2 59067 1 9
2 59068 1 9
2 59069 1 9
2 59070 1 9
2 59071 1 9
2 59072 1 9
2 59073 1 9
2 59074 1 9
2 59075 1 9
2 59076 1 9
2 59077 1 9
2 59078 1 9
2 59079 1 9
2 59080 1 9
2 59081 1 9
2 59082 1 9
2 59083 1 9
2 59084 1 9
2 59085 1 9
2 59086 1 9
2 59087 1 9
2 59088 1 9
2 59089 1 9
2 59090 1 9
2 59091 1 9
2 59092 1 9
2 59093 1 9
2 59094 1 9
2 59095 1 9
2 59096 1 9
2 59097 1 9
2 59098 1 9
2 59099 1 9
2 59100 1 9
2 59101 1 9
2 59102 1 9
2 59103 1 9
2 59104 1 9
2 59105 1 9
2 59106 1 9
2 59107 1 9
2 59108 1 9
2 59109 1 9
2 59110 1 9
2 59111 1 9
2 59112 1 9
2 59113 1 9
2 59114 1 9
2 59115 1 9
2 59116 1 9
2 59117 1 9
2 59118 1 9
2 59119 1 9
2 59120 1 9
2 59121 1 9
2 59122 1 9
2 59123 1 9
2 59124 1 9
2 59125 1 9
2 59126 1 9
2 59127 1 9
2 59128 1 9
2 59129 1 9
2 59130 1 9
2 59131 1 9
2 59132 1 9
2 59133 1 9
2 59134 1 9
2 59135 1 9
2 59136 1 9
2 59137 1 9
2 59138 1 9
2 59139 1 9
2 59140 1 9
2 59141 1 9
2 59142 1 9
2 59143 1 9
2 59144 1 9
2 59145 1 9
2 59146 1 9
2 59147 1 9
2 59148 1 9
2 59149 1 9
2 59150 1 9
2 59151 1 9
2 59152 1 9
2 59153 1 9
2 59154 1 9
2 59155 1 9
2 59156 1 9
2 59157 1 9
2 59158 1 9
2 59159 1 9
2 59160 1 9
2 59161 1 9
2 59162 1 9
2 59163 1 9
2 59164 1 9
2 59165 1 9
2 59166 1 9
2 59167 1 9
2 59168 1 9
2 59169 1 9
2 59170 1 9
2 59171 1 9
2 59172 1 9
2 59173 1 9
2 59174 1 9
2 59175 1 9
2 59176 1 9
2 59177 1 9
2 59178 1 9
1 10 0 217 0
2 59179 1 10
2 59180 1 10
2 59181 1 10
2 59182 1 10
2 59183 1 10
2 59184 1 10
2 59185 1 10
2 59186 1 10
2 59187 1 10
2 59188 1 10
2 59189 1 10
2 59190 1 10
2 59191 1 10
2 59192 1 10
2 59193 1 10
2 59194 1 10
2 59195 1 10
2 59196 1 10
2 59197 1 10
2 59198 1 10
2 59199 1 10
2 59200 1 10
2 59201 1 10
2 59202 1 10
2 59203 1 10
2 59204 1 10
2 59205 1 10
2 59206 1 10
2 59207 1 10
2 59208 1 10
2 59209 1 10
2 59210 1 10
2 59211 1 10
2 59212 1 10
2 59213 1 10
2 59214 1 10
2 59215 1 10
2 59216 1 10
2 59217 1 10
2 59218 1 10
2 59219 1 10
2 59220 1 10
2 59221 1 10
2 59222 1 10
2 59223 1 10
2 59224 1 10
2 59225 1 10
2 59226 1 10
2 59227 1 10
2 59228 1 10
2 59229 1 10
2 59230 1 10
2 59231 1 10
2 59232 1 10
2 59233 1 10
2 59234 1 10
2 59235 1 10
2 59236 1 10
2 59237 1 10
2 59238 1 10
2 59239 1 10
2 59240 1 10
2 59241 1 10
2 59242 1 10
2 59243 1 10
2 59244 1 10
2 59245 1 10
2 59246 1 10
2 59247 1 10
2 59248 1 10
2 59249 1 10
2 59250 1 10
2 59251 1 10
2 59252 1 10
2 59253 1 10
2 59254 1 10
2 59255 1 10
2 59256 1 10
2 59257 1 10
2 59258 1 10
2 59259 1 10
2 59260 1 10
2 59261 1 10
2 59262 1 10
2 59263 1 10
2 59264 1 10
2 59265 1 10
2 59266 1 10
2 59267 1 10
2 59268 1 10
2 59269 1 10
2 59270 1 10
2 59271 1 10
2 59272 1 10
2 59273 1 10
2 59274 1 10
2 59275 1 10
2 59276 1 10
2 59277 1 10
2 59278 1 10
2 59279 1 10
2 59280 1 10
2 59281 1 10
2 59282 1 10
2 59283 1 10
2 59284 1 10
2 59285 1 10
2 59286 1 10
2 59287 1 10
2 59288 1 10
2 59289 1 10
2 59290 1 10
2 59291 1 10
2 59292 1 10
2 59293 1 10
2 59294 1 10
2 59295 1 10
2 59296 1 10
2 59297 1 10
2 59298 1 10
2 59299 1 10
2 59300 1 10
2 59301 1 10
2 59302 1 10
2 59303 1 10
2 59304 1 10
2 59305 1 10
2 59306 1 10
2 59307 1 10
2 59308 1 10
2 59309 1 10
2 59310 1 10
2 59311 1 10
2 59312 1 10
2 59313 1 10
2 59314 1 10
2 59315 1 10
2 59316 1 10
2 59317 1 10
2 59318 1 10
2 59319 1 10
2 59320 1 10
2 59321 1 10
2 59322 1 10
2 59323 1 10
2 59324 1 10
2 59325 1 10
2 59326 1 10
2 59327 1 10
2 59328 1 10
2 59329 1 10
2 59330 1 10
2 59331 1 10
2 59332 1 10
2 59333 1 10
2 59334 1 10
2 59335 1 10
2 59336 1 10
2 59337 1 10
2 59338 1 10
2 59339 1 10
2 59340 1 10
2 59341 1 10
2 59342 1 10
2 59343 1 10
2 59344 1 10
2 59345 1 10
2 59346 1 10
2 59347 1 10
2 59348 1 10
2 59349 1 10
2 59350 1 10
2 59351 1 10
2 59352 1 10
2 59353 1 10
2 59354 1 10
2 59355 1 10
2 59356 1 10
2 59357 1 10
2 59358 1 10
2 59359 1 10
2 59360 1 10
2 59361 1 10
2 59362 1 10
2 59363 1 10
2 59364 1 10
2 59365 1 10
2 59366 1 10
2 59367 1 10
2 59368 1 10
2 59369 1 10
2 59370 1 10
2 59371 1 10
2 59372 1 10
2 59373 1 10
2 59374 1 10
2 59375 1 10
2 59376 1 10
2 59377 1 10
2 59378 1 10
2 59379 1 10
2 59380 1 10
2 59381 1 10
2 59382 1 10
2 59383 1 10
2 59384 1 10
2 59385 1 10
2 59386 1 10
2 59387 1 10
2 59388 1 10
2 59389 1 10
2 59390 1 10
2 59391 1 10
2 59392 1 10
2 59393 1 10
2 59394 1 10
2 59395 1 10
1 11 0 313 0
2 59396 1 11
2 59397 1 11
2 59398 1 11
2 59399 1 11
2 59400 1 11
2 59401 1 11
2 59402 1 11
2 59403 1 11
2 59404 1 11
2 59405 1 11
2 59406 1 11
2 59407 1 11
2 59408 1 11
2 59409 1 11
2 59410 1 11
2 59411 1 11
2 59412 1 11
2 59413 1 11
2 59414 1 11
2 59415 1 11
2 59416 1 11
2 59417 1 11
2 59418 1 11
2 59419 1 11
2 59420 1 11
2 59421 1 11
2 59422 1 11
2 59423 1 11
2 59424 1 11
2 59425 1 11
2 59426 1 11
2 59427 1 11
2 59428 1 11
2 59429 1 11
2 59430 1 11
2 59431 1 11
2 59432 1 11
2 59433 1 11
2 59434 1 11
2 59435 1 11
2 59436 1 11
2 59437 1 11
2 59438 1 11
2 59439 1 11
2 59440 1 11
2 59441 1 11
2 59442 1 11
2 59443 1 11
2 59444 1 11
2 59445 1 11
2 59446 1 11
2 59447 1 11
2 59448 1 11
2 59449 1 11
2 59450 1 11
2 59451 1 11
2 59452 1 11
2 59453 1 11
2 59454 1 11
2 59455 1 11
2 59456 1 11
2 59457 1 11
2 59458 1 11
2 59459 1 11
2 59460 1 11
2 59461 1 11
2 59462 1 11
2 59463 1 11
2 59464 1 11
2 59465 1 11
2 59466 1 11
2 59467 1 11
2 59468 1 11
2 59469 1 11
2 59470 1 11
2 59471 1 11
2 59472 1 11
2 59473 1 11
2 59474 1 11
2 59475 1 11
2 59476 1 11
2 59477 1 11
2 59478 1 11
2 59479 1 11
2 59480 1 11
2 59481 1 11
2 59482 1 11
2 59483 1 11
2 59484 1 11
2 59485 1 11
2 59486 1 11
2 59487 1 11
2 59488 1 11
2 59489 1 11
2 59490 1 11
2 59491 1 11
2 59492 1 11
2 59493 1 11
2 59494 1 11
2 59495 1 11
2 59496 1 11
2 59497 1 11
2 59498 1 11
2 59499 1 11
2 59500 1 11
2 59501 1 11
2 59502 1 11
2 59503 1 11
2 59504 1 11
2 59505 1 11
2 59506 1 11
2 59507 1 11
2 59508 1 11
2 59509 1 11
2 59510 1 11
2 59511 1 11
2 59512 1 11
2 59513 1 11
2 59514 1 11
2 59515 1 11
2 59516 1 11
2 59517 1 11
2 59518 1 11
2 59519 1 11
2 59520 1 11
2 59521 1 11
2 59522 1 11
2 59523 1 11
2 59524 1 11
2 59525 1 11
2 59526 1 11
2 59527 1 11
2 59528 1 11
2 59529 1 11
2 59530 1 11
2 59531 1 11
2 59532 1 11
2 59533 1 11
2 59534 1 11
2 59535 1 11
2 59536 1 11
2 59537 1 11
2 59538 1 11
2 59539 1 11
2 59540 1 11
2 59541 1 11
2 59542 1 11
2 59543 1 11
2 59544 1 11
2 59545 1 11
2 59546 1 11
2 59547 1 11
2 59548 1 11
2 59549 1 11
2 59550 1 11
2 59551 1 11
2 59552 1 11
2 59553 1 11
2 59554 1 11
2 59555 1 11
2 59556 1 11
2 59557 1 11
2 59558 1 11
2 59559 1 11
2 59560 1 11
2 59561 1 11
2 59562 1 11
2 59563 1 11
2 59564 1 11
2 59565 1 11
2 59566 1 11
2 59567 1 11
2 59568 1 11
2 59569 1 11
2 59570 1 11
2 59571 1 11
2 59572 1 11
2 59573 1 11
2 59574 1 11
2 59575 1 11
2 59576 1 11
2 59577 1 11
2 59578 1 11
2 59579 1 11
2 59580 1 11
2 59581 1 11
2 59582 1 11
2 59583 1 11
2 59584 1 11
2 59585 1 11
2 59586 1 11
2 59587 1 11
2 59588 1 11
2 59589 1 11
2 59590 1 11
2 59591 1 11
2 59592 1 11
2 59593 1 11
2 59594 1 11
2 59595 1 11
2 59596 1 11
2 59597 1 11
2 59598 1 11
2 59599 1 11
2 59600 1 11
2 59601 1 11
2 59602 1 11
2 59603 1 11
2 59604 1 11
2 59605 1 11
2 59606 1 11
2 59607 1 11
2 59608 1 11
2 59609 1 11
2 59610 1 11
2 59611 1 11
2 59612 1 11
2 59613 1 11
2 59614 1 11
2 59615 1 11
2 59616 1 11
2 59617 1 11
2 59618 1 11
2 59619 1 11
2 59620 1 11
2 59621 1 11
2 59622 1 11
2 59623 1 11
2 59624 1 11
2 59625 1 11
2 59626 1 11
2 59627 1 11
2 59628 1 11
2 59629 1 11
2 59630 1 11
2 59631 1 11
2 59632 1 11
2 59633 1 11
2 59634 1 11
2 59635 1 11
2 59636 1 11
2 59637 1 11
2 59638 1 11
2 59639 1 11
2 59640 1 11
2 59641 1 11
2 59642 1 11
2 59643 1 11
2 59644 1 11
2 59645 1 11
2 59646 1 11
2 59647 1 11
2 59648 1 11
2 59649 1 11
2 59650 1 11
2 59651 1 11
2 59652 1 11
2 59653 1 11
2 59654 1 11
2 59655 1 11
2 59656 1 11
2 59657 1 11
2 59658 1 11
2 59659 1 11
2 59660 1 11
2 59661 1 11
2 59662 1 11
2 59663 1 11
2 59664 1 11
2 59665 1 11
2 59666 1 11
2 59667 1 11
2 59668 1 11
2 59669 1 11
2 59670 1 11
2 59671 1 11
2 59672 1 11
2 59673 1 11
2 59674 1 11
2 59675 1 11
2 59676 1 11
2 59677 1 11
2 59678 1 11
2 59679 1 11
2 59680 1 11
2 59681 1 11
2 59682 1 11
2 59683 1 11
2 59684 1 11
2 59685 1 11
2 59686 1 11
2 59687 1 11
2 59688 1 11
2 59689 1 11
2 59690 1 11
2 59691 1 11
2 59692 1 11
2 59693 1 11
2 59694 1 11
2 59695 1 11
2 59696 1 11
2 59697 1 11
2 59698 1 11
2 59699 1 11
2 59700 1 11
2 59701 1 11
2 59702 1 11
2 59703 1 11
2 59704 1 11
2 59705 1 11
2 59706 1 11
2 59707 1 11
2 59708 1 11
1 12 0 246 0
2 59709 1 12
2 59710 1 12
2 59711 1 12
2 59712 1 12
2 59713 1 12
2 59714 1 12
2 59715 1 12
2 59716 1 12
2 59717 1 12
2 59718 1 12
2 59719 1 12
2 59720 1 12
2 59721 1 12
2 59722 1 12
2 59723 1 12
2 59724 1 12
2 59725 1 12
2 59726 1 12
2 59727 1 12
2 59728 1 12
2 59729 1 12
2 59730 1 12
2 59731 1 12
2 59732 1 12
2 59733 1 12
2 59734 1 12
2 59735 1 12
2 59736 1 12
2 59737 1 12
2 59738 1 12
2 59739 1 12
2 59740 1 12
2 59741 1 12
2 59742 1 12
2 59743 1 12
2 59744 1 12
2 59745 1 12
2 59746 1 12
2 59747 1 12
2 59748 1 12
2 59749 1 12
2 59750 1 12
2 59751 1 12
2 59752 1 12
2 59753 1 12
2 59754 1 12
2 59755 1 12
2 59756 1 12
2 59757 1 12
2 59758 1 12
2 59759 1 12
2 59760 1 12
2 59761 1 12
2 59762 1 12
2 59763 1 12
2 59764 1 12
2 59765 1 12
2 59766 1 12
2 59767 1 12
2 59768 1 12
2 59769 1 12
2 59770 1 12
2 59771 1 12
2 59772 1 12
2 59773 1 12
2 59774 1 12
2 59775 1 12
2 59776 1 12
2 59777 1 12
2 59778 1 12
2 59779 1 12
2 59780 1 12
2 59781 1 12
2 59782 1 12
2 59783 1 12
2 59784 1 12
2 59785 1 12
2 59786 1 12
2 59787 1 12
2 59788 1 12
2 59789 1 12
2 59790 1 12
2 59791 1 12
2 59792 1 12
2 59793 1 12
2 59794 1 12
2 59795 1 12
2 59796 1 12
2 59797 1 12
2 59798 1 12
2 59799 1 12
2 59800 1 12
2 59801 1 12
2 59802 1 12
2 59803 1 12
2 59804 1 12
2 59805 1 12
2 59806 1 12
2 59807 1 12
2 59808 1 12
2 59809 1 12
2 59810 1 12
2 59811 1 12
2 59812 1 12
2 59813 1 12
2 59814 1 12
2 59815 1 12
2 59816 1 12
2 59817 1 12
2 59818 1 12
2 59819 1 12
2 59820 1 12
2 59821 1 12
2 59822 1 12
2 59823 1 12
2 59824 1 12
2 59825 1 12
2 59826 1 12
2 59827 1 12
2 59828 1 12
2 59829 1 12
2 59830 1 12
2 59831 1 12
2 59832 1 12
2 59833 1 12
2 59834 1 12
2 59835 1 12
2 59836 1 12
2 59837 1 12
2 59838 1 12
2 59839 1 12
2 59840 1 12
2 59841 1 12
2 59842 1 12
2 59843 1 12
2 59844 1 12
2 59845 1 12
2 59846 1 12
2 59847 1 12
2 59848 1 12
2 59849 1 12
2 59850 1 12
2 59851 1 12
2 59852 1 12
2 59853 1 12
2 59854 1 12
2 59855 1 12
2 59856 1 12
2 59857 1 12
2 59858 1 12
2 59859 1 12
2 59860 1 12
2 59861 1 12
2 59862 1 12
2 59863 1 12
2 59864 1 12
2 59865 1 12
2 59866 1 12
2 59867 1 12
2 59868 1 12
2 59869 1 12
2 59870 1 12
2 59871 1 12
2 59872 1 12
2 59873 1 12
2 59874 1 12
2 59875 1 12
2 59876 1 12
2 59877 1 12
2 59878 1 12
2 59879 1 12
2 59880 1 12
2 59881 1 12
2 59882 1 12
2 59883 1 12
2 59884 1 12
2 59885 1 12
2 59886 1 12
2 59887 1 12
2 59888 1 12
2 59889 1 12
2 59890 1 12
2 59891 1 12
2 59892 1 12
2 59893 1 12
2 59894 1 12
2 59895 1 12
2 59896 1 12
2 59897 1 12
2 59898 1 12
2 59899 1 12
2 59900 1 12
2 59901 1 12
2 59902 1 12
2 59903 1 12
2 59904 1 12
2 59905 1 12
2 59906 1 12
2 59907 1 12
2 59908 1 12
2 59909 1 12
2 59910 1 12
2 59911 1 12
2 59912 1 12
2 59913 1 12
2 59914 1 12
2 59915 1 12
2 59916 1 12
2 59917 1 12
2 59918 1 12
2 59919 1 12
2 59920 1 12
2 59921 1 12
2 59922 1 12
2 59923 1 12
2 59924 1 12
2 59925 1 12
2 59926 1 12
2 59927 1 12
2 59928 1 12
2 59929 1 12
2 59930 1 12
2 59931 1 12
2 59932 1 12
2 59933 1 12
2 59934 1 12
2 59935 1 12
2 59936 1 12
2 59937 1 12
2 59938 1 12
2 59939 1 12
2 59940 1 12
2 59941 1 12
2 59942 1 12
2 59943 1 12
2 59944 1 12
2 59945 1 12
2 59946 1 12
2 59947 1 12
2 59948 1 12
2 59949 1 12
2 59950 1 12
2 59951 1 12
2 59952 1 12
2 59953 1 12
2 59954 1 12
1 13 0 128 0
2 59955 1 13
2 59956 1 13
2 59957 1 13
2 59958 1 13
2 59959 1 13
2 59960 1 13
2 59961 1 13
2 59962 1 13
2 59963 1 13
2 59964 1 13
2 59965 1 13
2 59966 1 13
2 59967 1 13
2 59968 1 13
2 59969 1 13
2 59970 1 13
2 59971 1 13
2 59972 1 13
2 59973 1 13
2 59974 1 13
2 59975 1 13
2 59976 1 13
2 59977 1 13
2 59978 1 13
2 59979 1 13
2 59980 1 13
2 59981 1 13
2 59982 1 13
2 59983 1 13
2 59984 1 13
2 59985 1 13
2 59986 1 13
2 59987 1 13
2 59988 1 13
2 59989 1 13
2 59990 1 13
2 59991 1 13
2 59992 1 13
2 59993 1 13
2 59994 1 13
2 59995 1 13
2 59996 1 13
2 59997 1 13
2 59998 1 13
2 59999 1 13
2 60000 1 13
2 60001 1 13
2 60002 1 13
2 60003 1 13
2 60004 1 13
2 60005 1 13
2 60006 1 13
2 60007 1 13
2 60008 1 13
2 60009 1 13
2 60010 1 13
2 60011 1 13
2 60012 1 13
2 60013 1 13
2 60014 1 13
2 60015 1 13
2 60016 1 13
2 60017 1 13
2 60018 1 13
2 60019 1 13
2 60020 1 13
2 60021 1 13
2 60022 1 13
2 60023 1 13
2 60024 1 13
2 60025 1 13
2 60026 1 13
2 60027 1 13
2 60028 1 13
2 60029 1 13
2 60030 1 13
2 60031 1 13
2 60032 1 13
2 60033 1 13
2 60034 1 13
2 60035 1 13
2 60036 1 13
2 60037 1 13
2 60038 1 13
2 60039 1 13
2 60040 1 13
2 60041 1 13
2 60042 1 13
2 60043 1 13
2 60044 1 13
2 60045 1 13
2 60046 1 13
2 60047 1 13
2 60048 1 13
2 60049 1 13
2 60050 1 13
2 60051 1 13
2 60052 1 13
2 60053 1 13
2 60054 1 13
2 60055 1 13
2 60056 1 13
2 60057 1 13
2 60058 1 13
2 60059 1 13
2 60060 1 13
2 60061 1 13
2 60062 1 13
2 60063 1 13
2 60064 1 13
2 60065 1 13
2 60066 1 13
2 60067 1 13
2 60068 1 13
2 60069 1 13
2 60070 1 13
2 60071 1 13
2 60072 1 13
2 60073 1 13
2 60074 1 13
2 60075 1 13
2 60076 1 13
2 60077 1 13
2 60078 1 13
2 60079 1 13
2 60080 1 13
2 60081 1 13
2 60082 1 13
1 14 0 87 0
2 60083 1 14
2 60084 1 14
2 60085 1 14
2 60086 1 14
2 60087 1 14
2 60088 1 14
2 60089 1 14
2 60090 1 14
2 60091 1 14
2 60092 1 14
2 60093 1 14
2 60094 1 14
2 60095 1 14
2 60096 1 14
2 60097 1 14
2 60098 1 14
2 60099 1 14
2 60100 1 14
2 60101 1 14
2 60102 1 14
2 60103 1 14
2 60104 1 14
2 60105 1 14
2 60106 1 14
2 60107 1 14
2 60108 1 14
2 60109 1 14
2 60110 1 14
2 60111 1 14
2 60112 1 14
2 60113 1 14
2 60114 1 14
2 60115 1 14
2 60116 1 14
2 60117 1 14
2 60118 1 14
2 60119 1 14
2 60120 1 14
2 60121 1 14
2 60122 1 14
2 60123 1 14
2 60124 1 14
2 60125 1 14
2 60126 1 14
2 60127 1 14
2 60128 1 14
2 60129 1 14
2 60130 1 14
2 60131 1 14
2 60132 1 14
2 60133 1 14
2 60134 1 14
2 60135 1 14
2 60136 1 14
2 60137 1 14
2 60138 1 14
2 60139 1 14
2 60140 1 14
2 60141 1 14
2 60142 1 14
2 60143 1 14
2 60144 1 14
2 60145 1 14
2 60146 1 14
2 60147 1 14
2 60148 1 14
2 60149 1 14
2 60150 1 14
2 60151 1 14
2 60152 1 14
2 60153 1 14
2 60154 1 14
2 60155 1 14
2 60156 1 14
2 60157 1 14
2 60158 1 14
2 60159 1 14
2 60160 1 14
2 60161 1 14
2 60162 1 14
2 60163 1 14
2 60164 1 14
2 60165 1 14
2 60166 1 14
2 60167 1 14
2 60168 1 14
2 60169 1 14
1 15 0 32 0
2 60170 1 15
2 60171 1 15
2 60172 1 15
2 60173 1 15
2 60174 1 15
2 60175 1 15
2 60176 1 15
2 60177 1 15
2 60178 1 15
2 60179 1 15
2 60180 1 15
2 60181 1 15
2 60182 1 15
2 60183 1 15
2 60184 1 15
2 60185 1 15
2 60186 1 15
2 60187 1 15
2 60188 1 15
2 60189 1 15
2 60190 1 15
2 60191 1 15
2 60192 1 15
2 60193 1 15
2 60194 1 15
2 60195 1 15
2 60196 1 15
2 60197 1 15
2 60198 1 15
2 60199 1 15
2 60200 1 15
2 60201 1 15
1 16 0 228 0
2 60202 1 16
2 60203 1 16
2 60204 1 16
2 60205 1 16
2 60206 1 16
2 60207 1 16
2 60208 1 16
2 60209 1 16
2 60210 1 16
2 60211 1 16
2 60212 1 16
2 60213 1 16
2 60214 1 16
2 60215 1 16
2 60216 1 16
2 60217 1 16
2 60218 1 16
2 60219 1 16
2 60220 1 16
2 60221 1 16
2 60222 1 16
2 60223 1 16
2 60224 1 16
2 60225 1 16
2 60226 1 16
2 60227 1 16
2 60228 1 16
2 60229 1 16
2 60230 1 16
2 60231 1 16
2 60232 1 16
2 60233 1 16
2 60234 1 16
2 60235 1 16
2 60236 1 16
2 60237 1 16
2 60238 1 16
2 60239 1 16
2 60240 1 16
2 60241 1 16
2 60242 1 16
2 60243 1 16
2 60244 1 16
2 60245 1 16
2 60246 1 16
2 60247 1 16
2 60248 1 16
2 60249 1 16
2 60250 1 16
2 60251 1 16
2 60252 1 16
2 60253 1 16
2 60254 1 16
2 60255 1 16
2 60256 1 16
2 60257 1 16
2 60258 1 16
2 60259 1 16
2 60260 1 16
2 60261 1 16
2 60262 1 16
2 60263 1 16
2 60264 1 16
2 60265 1 16
2 60266 1 16
2 60267 1 16
2 60268 1 16
2 60269 1 16
2 60270 1 16
2 60271 1 16
2 60272 1 16
2 60273 1 16
2 60274 1 16
2 60275 1 16
2 60276 1 16
2 60277 1 16
2 60278 1 16
2 60279 1 16
2 60280 1 16
2 60281 1 16
2 60282 1 16
2 60283 1 16
2 60284 1 16
2 60285 1 16
2 60286 1 16
2 60287 1 16
2 60288 1 16
2 60289 1 16
2 60290 1 16
2 60291 1 16
2 60292 1 16
2 60293 1 16
2 60294 1 16
2 60295 1 16
2 60296 1 16
2 60297 1 16
2 60298 1 16
2 60299 1 16
2 60300 1 16
2 60301 1 16
2 60302 1 16
2 60303 1 16
2 60304 1 16
2 60305 1 16
2 60306 1 16
2 60307 1 16
2 60308 1 16
2 60309 1 16
2 60310 1 16
2 60311 1 16
2 60312 1 16
2 60313 1 16
2 60314 1 16
2 60315 1 16
2 60316 1 16
2 60317 1 16
2 60318 1 16
2 60319 1 16
2 60320 1 16
2 60321 1 16
2 60322 1 16
2 60323 1 16
2 60324 1 16
2 60325 1 16
2 60326 1 16
2 60327 1 16
2 60328 1 16
2 60329 1 16
2 60330 1 16
2 60331 1 16
2 60332 1 16
2 60333 1 16
2 60334 1 16
2 60335 1 16
2 60336 1 16
2 60337 1 16
2 60338 1 16
2 60339 1 16
2 60340 1 16
2 60341 1 16
2 60342 1 16
2 60343 1 16
2 60344 1 16
2 60345 1 16
2 60346 1 16
2 60347 1 16
2 60348 1 16
2 60349 1 16
2 60350 1 16
2 60351 1 16
2 60352 1 16
2 60353 1 16
2 60354 1 16
2 60355 1 16
2 60356 1 16
2 60357 1 16
2 60358 1 16
2 60359 1 16
2 60360 1 16
2 60361 1 16
2 60362 1 16
2 60363 1 16
2 60364 1 16
2 60365 1 16
2 60366 1 16
2 60367 1 16
2 60368 1 16
2 60369 1 16
2 60370 1 16
2 60371 1 16
2 60372 1 16
2 60373 1 16
2 60374 1 16
2 60375 1 16
2 60376 1 16
2 60377 1 16
2 60378 1 16
2 60379 1 16
2 60380 1 16
2 60381 1 16
2 60382 1 16
2 60383 1 16
2 60384 1 16
2 60385 1 16
2 60386 1 16
2 60387 1 16
2 60388 1 16
2 60389 1 16
2 60390 1 16
2 60391 1 16
2 60392 1 16
2 60393 1 16
2 60394 1 16
2 60395 1 16
2 60396 1 16
2 60397 1 16
2 60398 1 16
2 60399 1 16
2 60400 1 16
2 60401 1 16
2 60402 1 16
2 60403 1 16
2 60404 1 16
2 60405 1 16
2 60406 1 16
2 60407 1 16
2 60408 1 16
2 60409 1 16
2 60410 1 16
2 60411 1 16
2 60412 1 16
2 60413 1 16
2 60414 1 16
2 60415 1 16
2 60416 1 16
2 60417 1 16
2 60418 1 16
2 60419 1 16
2 60420 1 16
2 60421 1 16
2 60422 1 16
2 60423 1 16
2 60424 1 16
2 60425 1 16
2 60426 1 16
2 60427 1 16
2 60428 1 16
2 60429 1 16
1 17 0 275 0
2 60430 1 17
2 60431 1 17
2 60432 1 17
2 60433 1 17
2 60434 1 17
2 60435 1 17
2 60436 1 17
2 60437 1 17
2 60438 1 17
2 60439 1 17
2 60440 1 17
2 60441 1 17
2 60442 1 17
2 60443 1 17
2 60444 1 17
2 60445 1 17
2 60446 1 17
2 60447 1 17
2 60448 1 17
2 60449 1 17
2 60450 1 17
2 60451 1 17
2 60452 1 17
2 60453 1 17
2 60454 1 17
2 60455 1 17
2 60456 1 17
2 60457 1 17
2 60458 1 17
2 60459 1 17
2 60460 1 17
2 60461 1 17
2 60462 1 17
2 60463 1 17
2 60464 1 17
2 60465 1 17
2 60466 1 17
2 60467 1 17
2 60468 1 17
2 60469 1 17
2 60470 1 17
2 60471 1 17
2 60472 1 17
2 60473 1 17
2 60474 1 17
2 60475 1 17
2 60476 1 17
2 60477 1 17
2 60478 1 17
2 60479 1 17
2 60480 1 17
2 60481 1 17
2 60482 1 17
2 60483 1 17
2 60484 1 17
2 60485 1 17
2 60486 1 17
2 60487 1 17
2 60488 1 17
2 60489 1 17
2 60490 1 17
2 60491 1 17
2 60492 1 17
2 60493 1 17
2 60494 1 17
2 60495 1 17
2 60496 1 17
2 60497 1 17
2 60498 1 17
2 60499 1 17
2 60500 1 17
2 60501 1 17
2 60502 1 17
2 60503 1 17
2 60504 1 17
2 60505 1 17
2 60506 1 17
2 60507 1 17
2 60508 1 17
2 60509 1 17
2 60510 1 17
2 60511 1 17
2 60512 1 17
2 60513 1 17
2 60514 1 17
2 60515 1 17
2 60516 1 17
2 60517 1 17
2 60518 1 17
2 60519 1 17
2 60520 1 17
2 60521 1 17
2 60522 1 17
2 60523 1 17
2 60524 1 17
2 60525 1 17
2 60526 1 17
2 60527 1 17
2 60528 1 17
2 60529 1 17
2 60530 1 17
2 60531 1 17
2 60532 1 17
2 60533 1 17
2 60534 1 17
2 60535 1 17
2 60536 1 17
2 60537 1 17
2 60538 1 17
2 60539 1 17
2 60540 1 17
2 60541 1 17
2 60542 1 17
2 60543 1 17
2 60544 1 17
2 60545 1 17
2 60546 1 17
2 60547 1 17
2 60548 1 17
2 60549 1 17
2 60550 1 17
2 60551 1 17
2 60552 1 17
2 60553 1 17
2 60554 1 17
2 60555 1 17
2 60556 1 17
2 60557 1 17
2 60558 1 17
2 60559 1 17
2 60560 1 17
2 60561 1 17
2 60562 1 17
2 60563 1 17
2 60564 1 17
2 60565 1 17
2 60566 1 17
2 60567 1 17
2 60568 1 17
2 60569 1 17
2 60570 1 17
2 60571 1 17
2 60572 1 17
2 60573 1 17
2 60574 1 17
2 60575 1 17
2 60576 1 17
2 60577 1 17
2 60578 1 17
2 60579 1 17
2 60580 1 17
2 60581 1 17
2 60582 1 17
2 60583 1 17
2 60584 1 17
2 60585 1 17
2 60586 1 17
2 60587 1 17
2 60588 1 17
2 60589 1 17
2 60590 1 17
2 60591 1 17
2 60592 1 17
2 60593 1 17
2 60594 1 17
2 60595 1 17
2 60596 1 17
2 60597 1 17
2 60598 1 17
2 60599 1 17
2 60600 1 17
2 60601 1 17
2 60602 1 17
2 60603 1 17
2 60604 1 17
2 60605 1 17
2 60606 1 17
2 60607 1 17
2 60608 1 17
2 60609 1 17
2 60610 1 17
2 60611 1 17
2 60612 1 17
2 60613 1 17
2 60614 1 17
2 60615 1 17
2 60616 1 17
2 60617 1 17
2 60618 1 17
2 60619 1 17
2 60620 1 17
2 60621 1 17
2 60622 1 17
2 60623 1 17
2 60624 1 17
2 60625 1 17
2 60626 1 17
2 60627 1 17
2 60628 1 17
2 60629 1 17
2 60630 1 17
2 60631 1 17
2 60632 1 17
2 60633 1 17
2 60634 1 17
2 60635 1 17
2 60636 1 17
2 60637 1 17
2 60638 1 17
2 60639 1 17
2 60640 1 17
2 60641 1 17
2 60642 1 17
2 60643 1 17
2 60644 1 17
2 60645 1 17
2 60646 1 17
2 60647 1 17
2 60648 1 17
2 60649 1 17
2 60650 1 17
2 60651 1 17
2 60652 1 17
2 60653 1 17
2 60654 1 17
2 60655 1 17
2 60656 1 17
2 60657 1 17
2 60658 1 17
2 60659 1 17
2 60660 1 17
2 60661 1 17
2 60662 1 17
2 60663 1 17
2 60664 1 17
2 60665 1 17
2 60666 1 17
2 60667 1 17
2 60668 1 17
2 60669 1 17
2 60670 1 17
2 60671 1 17
2 60672 1 17
2 60673 1 17
2 60674 1 17
2 60675 1 17
2 60676 1 17
2 60677 1 17
2 60678 1 17
2 60679 1 17
2 60680 1 17
2 60681 1 17
2 60682 1 17
2 60683 1 17
2 60684 1 17
2 60685 1 17
2 60686 1 17
2 60687 1 17
2 60688 1 17
2 60689 1 17
2 60690 1 17
2 60691 1 17
2 60692 1 17
2 60693 1 17
2 60694 1 17
2 60695 1 17
2 60696 1 17
2 60697 1 17
2 60698 1 17
2 60699 1 17
2 60700 1 17
2 60701 1 17
2 60702 1 17
2 60703 1 17
2 60704 1 17
1 18 0 431 0
2 60705 1 18
2 60706 1 18
2 60707 1 18
2 60708 1 18
2 60709 1 18
2 60710 1 18
2 60711 1 18
2 60712 1 18
2 60713 1 18
2 60714 1 18
2 60715 1 18
2 60716 1 18
2 60717 1 18
2 60718 1 18
2 60719 1 18
2 60720 1 18
2 60721 1 18
2 60722 1 18
2 60723 1 18
2 60724 1 18
2 60725 1 18
2 60726 1 18
2 60727 1 18
2 60728 1 18
2 60729 1 18
2 60730 1 18
2 60731 1 18
2 60732 1 18
2 60733 1 18
2 60734 1 18
2 60735 1 18
2 60736 1 18
2 60737 1 18
2 60738 1 18
2 60739 1 18
2 60740 1 18
2 60741 1 18
2 60742 1 18
2 60743 1 18
2 60744 1 18
2 60745 1 18
2 60746 1 18
2 60747 1 18
2 60748 1 18
2 60749 1 18
2 60750 1 18
2 60751 1 18
2 60752 1 18
2 60753 1 18
2 60754 1 18
2 60755 1 18
2 60756 1 18
2 60757 1 18
2 60758 1 18
2 60759 1 18
2 60760 1 18
2 60761 1 18
2 60762 1 18
2 60763 1 18
2 60764 1 18
2 60765 1 18
2 60766 1 18
2 60767 1 18
2 60768 1 18
2 60769 1 18
2 60770 1 18
2 60771 1 18
2 60772 1 18
2 60773 1 18
2 60774 1 18
2 60775 1 18
2 60776 1 18
2 60777 1 18
2 60778 1 18
2 60779 1 18
2 60780 1 18
2 60781 1 18
2 60782 1 18
2 60783 1 18
2 60784 1 18
2 60785 1 18
2 60786 1 18
2 60787 1 18
2 60788 1 18
2 60789 1 18
2 60790 1 18
2 60791 1 18
2 60792 1 18
2 60793 1 18
2 60794 1 18
2 60795 1 18
2 60796 1 18
2 60797 1 18
2 60798 1 18
2 60799 1 18
2 60800 1 18
2 60801 1 18
2 60802 1 18
2 60803 1 18
2 60804 1 18
2 60805 1 18
2 60806 1 18
2 60807 1 18
2 60808 1 18
2 60809 1 18
2 60810 1 18
2 60811 1 18
2 60812 1 18
2 60813 1 18
2 60814 1 18
2 60815 1 18
2 60816 1 18
2 60817 1 18
2 60818 1 18
2 60819 1 18
2 60820 1 18
2 60821 1 18
2 60822 1 18
2 60823 1 18
2 60824 1 18
2 60825 1 18
2 60826 1 18
2 60827 1 18
2 60828 1 18
2 60829 1 18
2 60830 1 18
2 60831 1 18
2 60832 1 18
2 60833 1 18
2 60834 1 18
2 60835 1 18
2 60836 1 18
2 60837 1 18
2 60838 1 18
2 60839 1 18
2 60840 1 18
2 60841 1 18
2 60842 1 18
2 60843 1 18
2 60844 1 18
2 60845 1 18
2 60846 1 18
2 60847 1 18
2 60848 1 18
2 60849 1 18
2 60850 1 18
2 60851 1 18
2 60852 1 18
2 60853 1 18
2 60854 1 18
2 60855 1 18
2 60856 1 18
2 60857 1 18
2 60858 1 18
2 60859 1 18
2 60860 1 18
2 60861 1 18
2 60862 1 18
2 60863 1 18
2 60864 1 18
2 60865 1 18
2 60866 1 18
2 60867 1 18
2 60868 1 18
2 60869 1 18
2 60870 1 18
2 60871 1 18
2 60872 1 18
2 60873 1 18
2 60874 1 18
2 60875 1 18
2 60876 1 18
2 60877 1 18
2 60878 1 18
2 60879 1 18
2 60880 1 18
2 60881 1 18
2 60882 1 18
2 60883 1 18
2 60884 1 18
2 60885 1 18
2 60886 1 18
2 60887 1 18
2 60888 1 18
2 60889 1 18
2 60890 1 18
2 60891 1 18
2 60892 1 18
2 60893 1 18
2 60894 1 18
2 60895 1 18
2 60896 1 18
2 60897 1 18
2 60898 1 18
2 60899 1 18
2 60900 1 18
2 60901 1 18
2 60902 1 18
2 60903 1 18
2 60904 1 18
2 60905 1 18
2 60906 1 18
2 60907 1 18
2 60908 1 18
2 60909 1 18
2 60910 1 18
2 60911 1 18
2 60912 1 18
2 60913 1 18
2 60914 1 18
2 60915 1 18
2 60916 1 18
2 60917 1 18
2 60918 1 18
2 60919 1 18
2 60920 1 18
2 60921 1 18
2 60922 1 18
2 60923 1 18
2 60924 1 18
2 60925 1 18
2 60926 1 18
2 60927 1 18
2 60928 1 18
2 60929 1 18
2 60930 1 18
2 60931 1 18
2 60932 1 18
2 60933 1 18
2 60934 1 18
2 60935 1 18
2 60936 1 18
2 60937 1 18
2 60938 1 18
2 60939 1 18
2 60940 1 18
2 60941 1 18
2 60942 1 18
2 60943 1 18
2 60944 1 18
2 60945 1 18
2 60946 1 18
2 60947 1 18
2 60948 1 18
2 60949 1 18
2 60950 1 18
2 60951 1 18
2 60952 1 18
2 60953 1 18
2 60954 1 18
2 60955 1 18
2 60956 1 18
2 60957 1 18
2 60958 1 18
2 60959 1 18
2 60960 1 18
2 60961 1 18
2 60962 1 18
2 60963 1 18
2 60964 1 18
2 60965 1 18
2 60966 1 18
2 60967 1 18
2 60968 1 18
2 60969 1 18
2 60970 1 18
2 60971 1 18
2 60972 1 18
2 60973 1 18
2 60974 1 18
2 60975 1 18
2 60976 1 18
2 60977 1 18
2 60978 1 18
2 60979 1 18
2 60980 1 18
2 60981 1 18
2 60982 1 18
2 60983 1 18
2 60984 1 18
2 60985 1 18
2 60986 1 18
2 60987 1 18
2 60988 1 18
2 60989 1 18
2 60990 1 18
2 60991 1 18
2 60992 1 18
2 60993 1 18
2 60994 1 18
2 60995 1 18
2 60996 1 18
2 60997 1 18
2 60998 1 18
2 60999 1 18
2 61000 1 18
2 61001 1 18
2 61002 1 18
2 61003 1 18
2 61004 1 18
2 61005 1 18
2 61006 1 18
2 61007 1 18
2 61008 1 18
2 61009 1 18
2 61010 1 18
2 61011 1 18
2 61012 1 18
2 61013 1 18
2 61014 1 18
2 61015 1 18
2 61016 1 18
2 61017 1 18
2 61018 1 18
2 61019 1 18
2 61020 1 18
2 61021 1 18
2 61022 1 18
2 61023 1 18
2 61024 1 18
2 61025 1 18
2 61026 1 18
2 61027 1 18
2 61028 1 18
2 61029 1 18
2 61030 1 18
2 61031 1 18
2 61032 1 18
2 61033 1 18
2 61034 1 18
2 61035 1 18
2 61036 1 18
2 61037 1 18
2 61038 1 18
2 61039 1 18
2 61040 1 18
2 61041 1 18
2 61042 1 18
2 61043 1 18
2 61044 1 18
2 61045 1 18
2 61046 1 18
2 61047 1 18
2 61048 1 18
2 61049 1 18
2 61050 1 18
2 61051 1 18
2 61052 1 18
2 61053 1 18
2 61054 1 18
2 61055 1 18
2 61056 1 18
2 61057 1 18
2 61058 1 18
2 61059 1 18
2 61060 1 18
2 61061 1 18
2 61062 1 18
2 61063 1 18
2 61064 1 18
2 61065 1 18
2 61066 1 18
2 61067 1 18
2 61068 1 18
2 61069 1 18
2 61070 1 18
2 61071 1 18
2 61072 1 18
2 61073 1 18
2 61074 1 18
2 61075 1 18
2 61076 1 18
2 61077 1 18
2 61078 1 18
2 61079 1 18
2 61080 1 18
2 61081 1 18
2 61082 1 18
2 61083 1 18
2 61084 1 18
2 61085 1 18
2 61086 1 18
2 61087 1 18
2 61088 1 18
2 61089 1 18
2 61090 1 18
2 61091 1 18
2 61092 1 18
2 61093 1 18
2 61094 1 18
2 61095 1 18
2 61096 1 18
2 61097 1 18
2 61098 1 18
2 61099 1 18
2 61100 1 18
2 61101 1 18
2 61102 1 18
2 61103 1 18
2 61104 1 18
2 61105 1 18
2 61106 1 18
2 61107 1 18
2 61108 1 18
2 61109 1 18
2 61110 1 18
2 61111 1 18
2 61112 1 18
2 61113 1 18
2 61114 1 18
2 61115 1 18
2 61116 1 18
2 61117 1 18
2 61118 1 18
2 61119 1 18
2 61120 1 18
2 61121 1 18
2 61122 1 18
2 61123 1 18
2 61124 1 18
2 61125 1 18
2 61126 1 18
2 61127 1 18
2 61128 1 18
2 61129 1 18
2 61130 1 18
2 61131 1 18
2 61132 1 18
2 61133 1 18
2 61134 1 18
2 61135 1 18
1 19 0 367 0
2 61136 1 19
2 61137 1 19
2 61138 1 19
2 61139 1 19
2 61140 1 19
2 61141 1 19
2 61142 1 19
2 61143 1 19
2 61144 1 19
2 61145 1 19
2 61146 1 19
2 61147 1 19
2 61148 1 19
2 61149 1 19
2 61150 1 19
2 61151 1 19
2 61152 1 19
2 61153 1 19
2 61154 1 19
2 61155 1 19
2 61156 1 19
2 61157 1 19
2 61158 1 19
2 61159 1 19
2 61160 1 19
2 61161 1 19
2 61162 1 19
2 61163 1 19
2 61164 1 19
2 61165 1 19
2 61166 1 19
2 61167 1 19
2 61168 1 19
2 61169 1 19
2 61170 1 19
2 61171 1 19
2 61172 1 19
2 61173 1 19
2 61174 1 19
2 61175 1 19
2 61176 1 19
2 61177 1 19
2 61178 1 19
2 61179 1 19
2 61180 1 19
2 61181 1 19
2 61182 1 19
2 61183 1 19
2 61184 1 19
2 61185 1 19
2 61186 1 19
2 61187 1 19
2 61188 1 19
2 61189 1 19
2 61190 1 19
2 61191 1 19
2 61192 1 19
2 61193 1 19
2 61194 1 19
2 61195 1 19
2 61196 1 19
2 61197 1 19
2 61198 1 19
2 61199 1 19
2 61200 1 19
2 61201 1 19
2 61202 1 19
2 61203 1 19
2 61204 1 19
2 61205 1 19
2 61206 1 19
2 61207 1 19
2 61208 1 19
2 61209 1 19
2 61210 1 19
2 61211 1 19
2 61212 1 19
2 61213 1 19
2 61214 1 19
2 61215 1 19
2 61216 1 19
2 61217 1 19
2 61218 1 19
2 61219 1 19
2 61220 1 19
2 61221 1 19
2 61222 1 19
2 61223 1 19
2 61224 1 19
2 61225 1 19
2 61226 1 19
2 61227 1 19
2 61228 1 19
2 61229 1 19
2 61230 1 19
2 61231 1 19
2 61232 1 19
2 61233 1 19
2 61234 1 19
2 61235 1 19
2 61236 1 19
2 61237 1 19
2 61238 1 19
2 61239 1 19
2 61240 1 19
2 61241 1 19
2 61242 1 19
2 61243 1 19
2 61244 1 19
2 61245 1 19
2 61246 1 19
2 61247 1 19
2 61248 1 19
2 61249 1 19
2 61250 1 19
2 61251 1 19
2 61252 1 19
2 61253 1 19
2 61254 1 19
2 61255 1 19
2 61256 1 19
2 61257 1 19
2 61258 1 19
2 61259 1 19
2 61260 1 19
2 61261 1 19
2 61262 1 19
2 61263 1 19
2 61264 1 19
2 61265 1 19
2 61266 1 19
2 61267 1 19
2 61268 1 19
2 61269 1 19
2 61270 1 19
2 61271 1 19
2 61272 1 19
2 61273 1 19
2 61274 1 19
2 61275 1 19
2 61276 1 19
2 61277 1 19
2 61278 1 19
2 61279 1 19
2 61280 1 19
2 61281 1 19
2 61282 1 19
2 61283 1 19
2 61284 1 19
2 61285 1 19
2 61286 1 19
2 61287 1 19
2 61288 1 19
2 61289 1 19
2 61290 1 19
2 61291 1 19
2 61292 1 19
2 61293 1 19
2 61294 1 19
2 61295 1 19
2 61296 1 19
2 61297 1 19
2 61298 1 19
2 61299 1 19
2 61300 1 19
2 61301 1 19
2 61302 1 19
2 61303 1 19
2 61304 1 19
2 61305 1 19
2 61306 1 19
2 61307 1 19
2 61308 1 19
2 61309 1 19
2 61310 1 19
2 61311 1 19
2 61312 1 19
2 61313 1 19
2 61314 1 19
2 61315 1 19
2 61316 1 19
2 61317 1 19
2 61318 1 19
2 61319 1 19
2 61320 1 19
2 61321 1 19
2 61322 1 19
2 61323 1 19
2 61324 1 19
2 61325 1 19
2 61326 1 19
2 61327 1 19
2 61328 1 19
2 61329 1 19
2 61330 1 19
2 61331 1 19
2 61332 1 19
2 61333 1 19
2 61334 1 19
2 61335 1 19
2 61336 1 19
2 61337 1 19
2 61338 1 19
2 61339 1 19
2 61340 1 19
2 61341 1 19
2 61342 1 19
2 61343 1 19
2 61344 1 19
2 61345 1 19
2 61346 1 19
2 61347 1 19
2 61348 1 19
2 61349 1 19
2 61350 1 19
2 61351 1 19
2 61352 1 19
2 61353 1 19
2 61354 1 19
2 61355 1 19
2 61356 1 19
2 61357 1 19
2 61358 1 19
2 61359 1 19
2 61360 1 19
2 61361 1 19
2 61362 1 19
2 61363 1 19
2 61364 1 19
2 61365 1 19
2 61366 1 19
2 61367 1 19
2 61368 1 19
2 61369 1 19
2 61370 1 19
2 61371 1 19
2 61372 1 19
2 61373 1 19
2 61374 1 19
2 61375 1 19
2 61376 1 19
2 61377 1 19
2 61378 1 19
2 61379 1 19
2 61380 1 19
2 61381 1 19
2 61382 1 19
2 61383 1 19
2 61384 1 19
2 61385 1 19
2 61386 1 19
2 61387 1 19
2 61388 1 19
2 61389 1 19
2 61390 1 19
2 61391 1 19
2 61392 1 19
2 61393 1 19
2 61394 1 19
2 61395 1 19
2 61396 1 19
2 61397 1 19
2 61398 1 19
2 61399 1 19
2 61400 1 19
2 61401 1 19
2 61402 1 19
2 61403 1 19
2 61404 1 19
2 61405 1 19
2 61406 1 19
2 61407 1 19
2 61408 1 19
2 61409 1 19
2 61410 1 19
2 61411 1 19
2 61412 1 19
2 61413 1 19
2 61414 1 19
2 61415 1 19
2 61416 1 19
2 61417 1 19
2 61418 1 19
2 61419 1 19
2 61420 1 19
2 61421 1 19
2 61422 1 19
2 61423 1 19
2 61424 1 19
2 61425 1 19
2 61426 1 19
2 61427 1 19
2 61428 1 19
2 61429 1 19
2 61430 1 19
2 61431 1 19
2 61432 1 19
2 61433 1 19
2 61434 1 19
2 61435 1 19
2 61436 1 19
2 61437 1 19
2 61438 1 19
2 61439 1 19
2 61440 1 19
2 61441 1 19
2 61442 1 19
2 61443 1 19
2 61444 1 19
2 61445 1 19
2 61446 1 19
2 61447 1 19
2 61448 1 19
2 61449 1 19
2 61450 1 19
2 61451 1 19
2 61452 1 19
2 61453 1 19
2 61454 1 19
2 61455 1 19
2 61456 1 19
2 61457 1 19
2 61458 1 19
2 61459 1 19
2 61460 1 19
2 61461 1 19
2 61462 1 19
2 61463 1 19
2 61464 1 19
2 61465 1 19
2 61466 1 19
2 61467 1 19
2 61468 1 19
2 61469 1 19
2 61470 1 19
2 61471 1 19
2 61472 1 19
2 61473 1 19
2 61474 1 19
2 61475 1 19
2 61476 1 19
2 61477 1 19
2 61478 1 19
2 61479 1 19
2 61480 1 19
2 61481 1 19
2 61482 1 19
2 61483 1 19
2 61484 1 19
2 61485 1 19
2 61486 1 19
2 61487 1 19
2 61488 1 19
2 61489 1 19
2 61490 1 19
2 61491 1 19
2 61492 1 19
2 61493 1 19
2 61494 1 19
2 61495 1 19
2 61496 1 19
2 61497 1 19
2 61498 1 19
2 61499 1 19
2 61500 1 19
2 61501 1 19
2 61502 1 19
1 20 0 257 0
2 61503 1 20
2 61504 1 20
2 61505 1 20
2 61506 1 20
2 61507 1 20
2 61508 1 20
2 61509 1 20
2 61510 1 20
2 61511 1 20
2 61512 1 20
2 61513 1 20
2 61514 1 20
2 61515 1 20
2 61516 1 20
2 61517 1 20
2 61518 1 20
2 61519 1 20
2 61520 1 20
2 61521 1 20
2 61522 1 20
2 61523 1 20
2 61524 1 20
2 61525 1 20
2 61526 1 20
2 61527 1 20
2 61528 1 20
2 61529 1 20
2 61530 1 20
2 61531 1 20
2 61532 1 20
2 61533 1 20
2 61534 1 20
2 61535 1 20
2 61536 1 20
2 61537 1 20
2 61538 1 20
2 61539 1 20
2 61540 1 20
2 61541 1 20
2 61542 1 20
2 61543 1 20
2 61544 1 20
2 61545 1 20
2 61546 1 20
2 61547 1 20
2 61548 1 20
2 61549 1 20
2 61550 1 20
2 61551 1 20
2 61552 1 20
2 61553 1 20
2 61554 1 20
2 61555 1 20
2 61556 1 20
2 61557 1 20
2 61558 1 20
2 61559 1 20
2 61560 1 20
2 61561 1 20
2 61562 1 20
2 61563 1 20
2 61564 1 20
2 61565 1 20
2 61566 1 20
2 61567 1 20
2 61568 1 20
2 61569 1 20
2 61570 1 20
2 61571 1 20
2 61572 1 20
2 61573 1 20
2 61574 1 20
2 61575 1 20
2 61576 1 20
2 61577 1 20
2 61578 1 20
2 61579 1 20
2 61580 1 20
2 61581 1 20
2 61582 1 20
2 61583 1 20
2 61584 1 20
2 61585 1 20
2 61586 1 20
2 61587 1 20
2 61588 1 20
2 61589 1 20
2 61590 1 20
2 61591 1 20
2 61592 1 20
2 61593 1 20
2 61594 1 20
2 61595 1 20
2 61596 1 20
2 61597 1 20
2 61598 1 20
2 61599 1 20
2 61600 1 20
2 61601 1 20
2 61602 1 20
2 61603 1 20
2 61604 1 20
2 61605 1 20
2 61606 1 20
2 61607 1 20
2 61608 1 20
2 61609 1 20
2 61610 1 20
2 61611 1 20
2 61612 1 20
2 61613 1 20
2 61614 1 20
2 61615 1 20
2 61616 1 20
2 61617 1 20
2 61618 1 20
2 61619 1 20
2 61620 1 20
2 61621 1 20
2 61622 1 20
2 61623 1 20
2 61624 1 20
2 61625 1 20
2 61626 1 20
2 61627 1 20
2 61628 1 20
2 61629 1 20
2 61630 1 20
2 61631 1 20
2 61632 1 20
2 61633 1 20
2 61634 1 20
2 61635 1 20
2 61636 1 20
2 61637 1 20
2 61638 1 20
2 61639 1 20
2 61640 1 20
2 61641 1 20
2 61642 1 20
2 61643 1 20
2 61644 1 20
2 61645 1 20
2 61646 1 20
2 61647 1 20
2 61648 1 20
2 61649 1 20
2 61650 1 20
2 61651 1 20
2 61652 1 20
2 61653 1 20
2 61654 1 20
2 61655 1 20
2 61656 1 20
2 61657 1 20
2 61658 1 20
2 61659 1 20
2 61660 1 20
2 61661 1 20
2 61662 1 20
2 61663 1 20
2 61664 1 20
2 61665 1 20
2 61666 1 20
2 61667 1 20
2 61668 1 20
2 61669 1 20
2 61670 1 20
2 61671 1 20
2 61672 1 20
2 61673 1 20
2 61674 1 20
2 61675 1 20
2 61676 1 20
2 61677 1 20
2 61678 1 20
2 61679 1 20
2 61680 1 20
2 61681 1 20
2 61682 1 20
2 61683 1 20
2 61684 1 20
2 61685 1 20
2 61686 1 20
2 61687 1 20
2 61688 1 20
2 61689 1 20
2 61690 1 20
2 61691 1 20
2 61692 1 20
2 61693 1 20
2 61694 1 20
2 61695 1 20
2 61696 1 20
2 61697 1 20
2 61698 1 20
2 61699 1 20
2 61700 1 20
2 61701 1 20
2 61702 1 20
2 61703 1 20
2 61704 1 20
2 61705 1 20
2 61706 1 20
2 61707 1 20
2 61708 1 20
2 61709 1 20
2 61710 1 20
2 61711 1 20
2 61712 1 20
2 61713 1 20
2 61714 1 20
2 61715 1 20
2 61716 1 20
2 61717 1 20
2 61718 1 20
2 61719 1 20
2 61720 1 20
2 61721 1 20
2 61722 1 20
2 61723 1 20
2 61724 1 20
2 61725 1 20
2 61726 1 20
2 61727 1 20
2 61728 1 20
2 61729 1 20
2 61730 1 20
2 61731 1 20
2 61732 1 20
2 61733 1 20
2 61734 1 20
2 61735 1 20
2 61736 1 20
2 61737 1 20
2 61738 1 20
2 61739 1 20
2 61740 1 20
2 61741 1 20
2 61742 1 20
2 61743 1 20
2 61744 1 20
2 61745 1 20
2 61746 1 20
2 61747 1 20
2 61748 1 20
2 61749 1 20
2 61750 1 20
2 61751 1 20
2 61752 1 20
2 61753 1 20
2 61754 1 20
2 61755 1 20
2 61756 1 20
2 61757 1 20
2 61758 1 20
2 61759 1 20
1 21 0 114 0
2 61760 1 21
2 61761 1 21
2 61762 1 21
2 61763 1 21
2 61764 1 21
2 61765 1 21
2 61766 1 21
2 61767 1 21
2 61768 1 21
2 61769 1 21
2 61770 1 21
2 61771 1 21
2 61772 1 21
2 61773 1 21
2 61774 1 21
2 61775 1 21
2 61776 1 21
2 61777 1 21
2 61778 1 21
2 61779 1 21
2 61780 1 21
2 61781 1 21
2 61782 1 21
2 61783 1 21
2 61784 1 21
2 61785 1 21
2 61786 1 21
2 61787 1 21
2 61788 1 21
2 61789 1 21
2 61790 1 21
2 61791 1 21
2 61792 1 21
2 61793 1 21
2 61794 1 21
2 61795 1 21
2 61796 1 21
2 61797 1 21
2 61798 1 21
2 61799 1 21
2 61800 1 21
2 61801 1 21
2 61802 1 21
2 61803 1 21
2 61804 1 21
2 61805 1 21
2 61806 1 21
2 61807 1 21
2 61808 1 21
2 61809 1 21
2 61810 1 21
2 61811 1 21
2 61812 1 21
2 61813 1 21
2 61814 1 21
2 61815 1 21
2 61816 1 21
2 61817 1 21
2 61818 1 21
2 61819 1 21
2 61820 1 21
2 61821 1 21
2 61822 1 21
2 61823 1 21
2 61824 1 21
2 61825 1 21
2 61826 1 21
2 61827 1 21
2 61828 1 21
2 61829 1 21
2 61830 1 21
2 61831 1 21
2 61832 1 21
2 61833 1 21
2 61834 1 21
2 61835 1 21
2 61836 1 21
2 61837 1 21
2 61838 1 21
2 61839 1 21
2 61840 1 21
2 61841 1 21
2 61842 1 21
2 61843 1 21
2 61844 1 21
2 61845 1 21
2 61846 1 21
2 61847 1 21
2 61848 1 21
2 61849 1 21
2 61850 1 21
2 61851 1 21
2 61852 1 21
2 61853 1 21
2 61854 1 21
2 61855 1 21
2 61856 1 21
2 61857 1 21
2 61858 1 21
2 61859 1 21
2 61860 1 21
2 61861 1 21
2 61862 1 21
2 61863 1 21
2 61864 1 21
2 61865 1 21
2 61866 1 21
2 61867 1 21
2 61868 1 21
2 61869 1 21
2 61870 1 21
2 61871 1 21
2 61872 1 21
2 61873 1 21
1 22 0 133 0
2 61874 1 22
2 61875 1 22
2 61876 1 22
2 61877 1 22
2 61878 1 22
2 61879 1 22
2 61880 1 22
2 61881 1 22
2 61882 1 22
2 61883 1 22
2 61884 1 22
2 61885 1 22
2 61886 1 22
2 61887 1 22
2 61888 1 22
2 61889 1 22
2 61890 1 22
2 61891 1 22
2 61892 1 22
2 61893 1 22
2 61894 1 22
2 61895 1 22
2 61896 1 22
2 61897 1 22
2 61898 1 22
2 61899 1 22
2 61900 1 22
2 61901 1 22
2 61902 1 22
2 61903 1 22
2 61904 1 22
2 61905 1 22
2 61906 1 22
2 61907 1 22
2 61908 1 22
2 61909 1 22
2 61910 1 22
2 61911 1 22
2 61912 1 22
2 61913 1 22
2 61914 1 22
2 61915 1 22
2 61916 1 22
2 61917 1 22
2 61918 1 22
2 61919 1 22
2 61920 1 22
2 61921 1 22
2 61922 1 22
2 61923 1 22
2 61924 1 22
2 61925 1 22
2 61926 1 22
2 61927 1 22
2 61928 1 22
2 61929 1 22
2 61930 1 22
2 61931 1 22
2 61932 1 22
2 61933 1 22
2 61934 1 22
2 61935 1 22
2 61936 1 22
2 61937 1 22
2 61938 1 22
2 61939 1 22
2 61940 1 22
2 61941 1 22
2 61942 1 22
2 61943 1 22
2 61944 1 22
2 61945 1 22
2 61946 1 22
2 61947 1 22
2 61948 1 22
2 61949 1 22
2 61950 1 22
2 61951 1 22
2 61952 1 22
2 61953 1 22
2 61954 1 22
2 61955 1 22
2 61956 1 22
2 61957 1 22
2 61958 1 22
2 61959 1 22
2 61960 1 22
2 61961 1 22
2 61962 1 22
2 61963 1 22
2 61964 1 22
2 61965 1 22
2 61966 1 22
2 61967 1 22
2 61968 1 22
2 61969 1 22
2 61970 1 22
2 61971 1 22
2 61972 1 22
2 61973 1 22
2 61974 1 22
2 61975 1 22
2 61976 1 22
2 61977 1 22
2 61978 1 22
2 61979 1 22
2 61980 1 22
2 61981 1 22
2 61982 1 22
2 61983 1 22
2 61984 1 22
2 61985 1 22
2 61986 1 22
2 61987 1 22
2 61988 1 22
2 61989 1 22
2 61990 1 22
2 61991 1 22
2 61992 1 22
2 61993 1 22
2 61994 1 22
2 61995 1 22
2 61996 1 22
2 61997 1 22
2 61998 1 22
2 61999 1 22
2 62000 1 22
2 62001 1 22
2 62002 1 22
2 62003 1 22
2 62004 1 22
2 62005 1 22
2 62006 1 22
1 23 0 135 0
2 62007 1 23
2 62008 1 23
2 62009 1 23
2 62010 1 23
2 62011 1 23
2 62012 1 23
2 62013 1 23
2 62014 1 23
2 62015 1 23
2 62016 1 23
2 62017 1 23
2 62018 1 23
2 62019 1 23
2 62020 1 23
2 62021 1 23
2 62022 1 23
2 62023 1 23
2 62024 1 23
2 62025 1 23
2 62026 1 23
2 62027 1 23
2 62028 1 23
2 62029 1 23
2 62030 1 23
2 62031 1 23
2 62032 1 23
2 62033 1 23
2 62034 1 23
2 62035 1 23
2 62036 1 23
2 62037 1 23
2 62038 1 23
2 62039 1 23
2 62040 1 23
2 62041 1 23
2 62042 1 23
2 62043 1 23
2 62044 1 23
2 62045 1 23
2 62046 1 23
2 62047 1 23
2 62048 1 23
2 62049 1 23
2 62050 1 23
2 62051 1 23
2 62052 1 23
2 62053 1 23
2 62054 1 23
2 62055 1 23
2 62056 1 23
2 62057 1 23
2 62058 1 23
2 62059 1 23
2 62060 1 23
2 62061 1 23
2 62062 1 23
2 62063 1 23
2 62064 1 23
2 62065 1 23
2 62066 1 23
2 62067 1 23
2 62068 1 23
2 62069 1 23
2 62070 1 23
2 62071 1 23
2 62072 1 23
2 62073 1 23
2 62074 1 23
2 62075 1 23
2 62076 1 23
2 62077 1 23
2 62078 1 23
2 62079 1 23
2 62080 1 23
2 62081 1 23
2 62082 1 23
2 62083 1 23
2 62084 1 23
2 62085 1 23
2 62086 1 23
2 62087 1 23
2 62088 1 23
2 62089 1 23
2 62090 1 23
2 62091 1 23
2 62092 1 23
2 62093 1 23
2 62094 1 23
2 62095 1 23
2 62096 1 23
2 62097 1 23
2 62098 1 23
2 62099 1 23
2 62100 1 23
2 62101 1 23
2 62102 1 23
2 62103 1 23
2 62104 1 23
2 62105 1 23
2 62106 1 23
2 62107 1 23
2 62108 1 23
2 62109 1 23
2 62110 1 23
2 62111 1 23
2 62112 1 23
2 62113 1 23
2 62114 1 23
2 62115 1 23
2 62116 1 23
2 62117 1 23
2 62118 1 23
2 62119 1 23
2 62120 1 23
2 62121 1 23
2 62122 1 23
2 62123 1 23
2 62124 1 23
2 62125 1 23
2 62126 1 23
2 62127 1 23
2 62128 1 23
2 62129 1 23
2 62130 1 23
2 62131 1 23
2 62132 1 23
2 62133 1 23
2 62134 1 23
2 62135 1 23
2 62136 1 23
2 62137 1 23
2 62138 1 23
2 62139 1 23
2 62140 1 23
2 62141 1 23
1 24 0 2 0
2 62142 1 24
2 62143 1 24
2 62144 1 27
2 62145 1 27
2 62146 1 27
2 62147 1 27
2 62148 1 27
2 62149 1 27
2 62150 1 27
2 62151 1 27
2 62152 1 27
2 62153 1 27
2 62154 1 27
2 62155 1 27
2 62156 1 27
2 62157 1 27
2 62158 1 27
2 62159 1 27
2 62160 1 27
2 62161 1 27
2 62162 1 27
2 62163 1 27
2 62164 1 27
2 62165 1 27
2 62166 1 27
2 62167 1 27
2 62168 1 27
2 62169 1 27
2 62170 1 27
2 62171 1 27
2 62172 1 27
2 62173 1 27
2 62174 1 27
2 62175 1 27
2 62176 1 27
2 62177 1 27
2 62178 1 27
2 62179 1 27
2 62180 1 27
2 62181 1 27
2 62182 1 27
2 62183 1 27
2 62184 1 27
2 62185 1 27
2 62186 1 27
2 62187 1 27
2 62188 1 27
2 62189 1 27
2 62190 1 27
2 62191 1 27
2 62192 1 27
2 62193 1 27
2 62194 1 27
2 62195 1 27
2 62196 1 27
2 62197 1 27
2 62198 1 27
2 62199 1 27
2 62200 1 27
2 62201 1 27
2 62202 1 27
2 62203 1 27
2 62204 1 27
2 62205 1 27
2 62206 1 27
2 62207 1 27
2 62208 1 27
2 62209 1 27
2 62210 1 27
2 62211 1 27
2 62212 1 27
2 62213 1 27
2 62214 1 27
2 62215 1 27
2 62216 1 27
2 62217 1 27
2 62218 1 27
2 62219 1 27
2 62220 1 27
2 62221 1 27
2 62222 1 27
2 62223 1 27
2 62224 1 27
2 62225 1 27
2 62226 1 27
2 62227 1 27
2 62228 1 27
2 62229 1 27
2 62230 1 27
2 62231 1 27
2 62232 1 27
2 62233 1 27
2 62234 1 27
2 62235 1 27
2 62236 1 27
2 62237 1 27
2 62238 1 27
2 62239 1 27
2 62240 1 27
2 62241 1 27
2 62242 1 27
2 62243 1 27
2 62244 1 27
2 62245 1 27
2 62246 1 27
2 62247 1 27
2 62248 1 27
2 62249 1 27
2 62250 1 27
2 62251 1 27
2 62252 1 27
2 62253 1 27
2 62254 1 27
2 62255 1 27
2 62256 1 27
2 62257 1 27
2 62258 1 27
2 62259 1 27
2 62260 1 27
2 62261 1 27
2 62262 1 27
2 62263 1 27
2 62264 1 27
2 62265 1 27
2 62266 1 27
2 62267 1 27
2 62268 1 27
2 62269 1 27
2 62270 1 27
2 62271 1 27
2 62272 1 27
2 62273 1 27
2 62274 1 27
2 62275 1 27
2 62276 1 27
2 62277 1 27
2 62278 1 27
2 62279 1 27
2 62280 1 27
2 62281 1 27
2 62282 1 27
2 62283 1 27
2 62284 1 28
2 62285 1 28
2 62286 1 28
2 62287 1 28
2 62288 1 28
2 62289 1 28
2 62290 1 28
2 62291 1 28
2 62292 1 28
2 62293 1 28
2 62294 1 28
2 62295 1 28
2 62296 1 28
2 62297 1 28
2 62298 1 28
2 62299 1 28
2 62300 1 28
2 62301 1 28
2 62302 1 28
2 62303 1 28
2 62304 1 28
2 62305 1 28
2 62306 1 28
2 62307 1 28
2 62308 1 28
2 62309 1 28
2 62310 1 28
2 62311 1 28
2 62312 1 28
2 62313 1 28
2 62314 1 28
2 62315 1 28
2 62316 1 28
2 62317 1 28
2 62318 1 28
2 62319 1 28
2 62320 1 28
2 62321 1 28
2 62322 1 28
2 62323 1 28
2 62324 1 28
2 62325 1 28
2 62326 1 28
2 62327 1 28
2 62328 1 28
2 62329 1 28
2 62330 1 28
2 62331 1 28
2 62332 1 28
2 62333 1 28
2 62334 1 28
2 62335 1 28
2 62336 1 28
2 62337 1 28
2 62338 1 28
2 62339 1 28
2 62340 1 28
2 62341 1 28
2 62342 1 28
2 62343 1 28
2 62344 1 28
2 62345 1 28
2 62346 1 28
2 62347 1 28
2 62348 1 28
2 62349 1 28
2 62350 1 28
2 62351 1 28
2 62352 1 28
2 62353 1 28
2 62354 1 28
2 62355 1 28
2 62356 1 28
2 62357 1 28
2 62358 1 28
2 62359 1 28
2 62360 1 28
2 62361 1 28
2 62362 1 28
2 62363 1 28
2 62364 1 28
2 62365 1 28
2 62366 1 28
2 62367 1 28
2 62368 1 28
2 62369 1 28
2 62370 1 28
2 62371 1 28
2 62372 1 28
2 62373 1 28
2 62374 1 28
2 62375 1 28
2 62376 1 28
2 62377 1 28
2 62378 1 28
2 62379 1 28
2 62380 1 28
2 62381 1 28
2 62382 1 28
2 62383 1 28
2 62384 1 28
2 62385 1 28
2 62386 1 28
2 62387 1 28
2 62388 1 28
2 62389 1 28
2 62390 1 28
2 62391 1 28
2 62392 1 28
2 62393 1 28
2 62394 1 28
2 62395 1 28
2 62396 1 28
2 62397 1 28
2 62398 1 28
2 62399 1 28
2 62400 1 28
2 62401 1 28
2 62402 1 28
2 62403 1 28
2 62404 1 28
2 62405 1 28
2 62406 1 28
2 62407 1 28
2 62408 1 28
2 62409 1 28
2 62410 1 28
2 62411 1 28
2 62412 1 28
2 62413 1 28
2 62414 1 28
2 62415 1 28
2 62416 1 28
2 62417 1 28
2 62418 1 28
2 62419 1 28
2 62420 1 28
2 62421 1 28
2 62422 1 28
2 62423 1 28
2 62424 1 28
2 62425 1 28
2 62426 1 28
2 62427 1 28
2 62428 1 28
2 62429 1 28
2 62430 1 28
2 62431 1 28
2 62432 1 28
2 62433 1 28
2 62434 1 28
2 62435 1 28
2 62436 1 28
2 62437 1 28
2 62438 1 28
2 62439 1 28
2 62440 1 28
2 62441 1 28
2 62442 1 28
2 62443 1 28
2 62444 1 28
2 62445 1 28
2 62446 1 28
2 62447 1 28
2 62448 1 28
2 62449 1 28
2 62450 1 28
2 62451 1 28
2 62452 1 28
2 62453 1 28
2 62454 1 28
2 62455 1 28
2 62456 1 28
2 62457 1 28
2 62458 1 28
2 62459 1 28
2 62460 1 28
2 62461 1 28
2 62462 1 28
2 62463 1 28
2 62464 1 28
2 62465 1 28
2 62466 1 28
2 62467 1 28
2 62468 1 28
2 62469 1 28
2 62470 1 28
2 62471 1 28
2 62472 1 28
2 62473 1 28
2 62474 1 28
2 62475 1 28
2 62476 1 28
2 62477 1 28
2 62478 1 28
2 62479 1 28
2 62480 1 28
2 62481 1 28
2 62482 1 28
2 62483 1 28
2 62484 1 28
2 62485 1 28
2 62486 1 28
2 62487 1 28
2 62488 1 28
2 62489 1 28
2 62490 1 28
2 62491 1 28
2 62492 1 28
2 62493 1 28
2 62494 1 28
2 62495 1 28
2 62496 1 28
2 62497 1 28
2 62498 1 28
2 62499 1 28
2 62500 1 28
2 62501 1 28
2 62502 1 28
2 62503 1 28
2 62504 1 28
2 62505 1 28
2 62506 1 28
2 62507 1 28
2 62508 1 28
2 62509 1 28
2 62510 1 28
2 62511 1 28
2 62512 1 28
2 62513 1 28
2 62514 1 28
2 62515 1 28
2 62516 1 28
2 62517 1 28
2 62518 1 28
2 62519 1 28
2 62520 1 28
2 62521 1 28
2 62522 1 28
2 62523 1 28
2 62524 1 28
2 62525 1 28
2 62526 1 28
2 62527 1 28
2 62528 1 28
2 62529 1 28
2 62530 1 28
2 62531 1 28
2 62532 1 28
2 62533 1 28
2 62534 1 28
2 62535 1 28
2 62536 1 28
2 62537 1 28
2 62538 1 28
2 62539 1 28
2 62540 1 28
2 62541 1 28
2 62542 1 28
2 62543 1 29
2 62544 1 29
2 62545 1 29
2 62546 1 29
2 62547 1 29
2 62548 1 29
2 62549 1 29
2 62550 1 29
2 62551 1 29
2 62552 1 29
2 62553 1 29
2 62554 1 29
2 62555 1 29
2 62556 1 29
2 62557 1 29
2 62558 1 29
2 62559 1 29
2 62560 1 29
2 62561 1 29
2 62562 1 29
2 62563 1 29
2 62564 1 29
2 62565 1 29
2 62566 1 29
2 62567 1 29
2 62568 1 29
2 62569 1 29
2 62570 1 29
2 62571 1 29
2 62572 1 29
2 62573 1 29
2 62574 1 29
2 62575 1 29
2 62576 1 29
2 62577 1 29
2 62578 1 29
2 62579 1 29
2 62580 1 29
2 62581 1 29
2 62582 1 29
2 62583 1 29
2 62584 1 29
2 62585 1 29
2 62586 1 29
2 62587 1 29
2 62588 1 29
2 62589 1 29
2 62590 1 29
2 62591 1 29
2 62592 1 29
2 62593 1 29
2 62594 1 29
2 62595 1 29
2 62596 1 29
2 62597 1 29
2 62598 1 29
2 62599 1 29
2 62600 1 29
2 62601 1 29
2 62602 1 29
2 62603 1 29
2 62604 1 29
2 62605 1 29
2 62606 1 29
2 62607 1 29
2 62608 1 29
2 62609 1 29
2 62610 1 29
2 62611 1 29
2 62612 1 29
2 62613 1 29
2 62614 1 29
2 62615 1 29
2 62616 1 29
2 62617 1 29
2 62618 1 29
2 62619 1 29
2 62620 1 29
2 62621 1 29
2 62622 1 29
2 62623 1 29
2 62624 1 29
2 62625 1 29
2 62626 1 29
2 62627 1 29
2 62628 1 29
2 62629 1 29
2 62630 1 29
2 62631 1 29
2 62632 1 29
2 62633 1 29
2 62634 1 29
2 62635 1 29
2 62636 1 29
2 62637 1 29
2 62638 1 29
2 62639 1 29
2 62640 1 29
2 62641 1 29
2 62642 1 29
2 62643 1 29
2 62644 1 29
2 62645 1 29
2 62646 1 29
2 62647 1 29
2 62648 1 29
2 62649 1 29
2 62650 1 29
2 62651 1 29
2 62652 1 29
2 62653 1 29
2 62654 1 29
2 62655 1 29
2 62656 1 29
2 62657 1 29
2 62658 1 29
2 62659 1 29
2 62660 1 29
2 62661 1 29
2 62662 1 29
2 62663 1 29
2 62664 1 29
2 62665 1 29
2 62666 1 29
2 62667 1 29
2 62668 1 29
2 62669 1 29
2 62670 1 29
2 62671 1 29
2 62672 1 29
2 62673 1 29
2 62674 1 29
2 62675 1 29
2 62676 1 29
2 62677 1 29
2 62678 1 29
2 62679 1 29
2 62680 1 29
2 62681 1 29
2 62682 1 29
2 62683 1 29
2 62684 1 29
2 62685 1 29
2 62686 1 29
2 62687 1 29
2 62688 1 29
2 62689 1 29
2 62690 1 29
2 62691 1 29
2 62692 1 29
2 62693 1 29
2 62694 1 29
2 62695 1 29
2 62696 1 29
2 62697 1 29
2 62698 1 29
2 62699 1 29
2 62700 1 29
2 62701 1 29
2 62702 1 29
2 62703 1 29
2 62704 1 29
2 62705 1 29
2 62706 1 29
2 62707 1 29
2 62708 1 29
2 62709 1 29
2 62710 1 29
2 62711 1 29
2 62712 1 29
2 62713 1 29
2 62714 1 29
2 62715 1 29
2 62716 1 29
2 62717 1 29
2 62718 1 29
2 62719 1 29
2 62720 1 29
2 62721 1 29
2 62722 1 29
2 62723 1 29
2 62724 1 29
2 62725 1 29
2 62726 1 29
2 62727 1 29
2 62728 1 29
2 62729 1 29
2 62730 1 29
2 62731 1 29
2 62732 1 29
2 62733 1 29
2 62734 1 29
2 62735 1 29
2 62736 1 29
2 62737 1 29
2 62738 1 29
2 62739 1 29
2 62740 1 29
2 62741 1 29
2 62742 1 29
2 62743 1 29
2 62744 1 29
2 62745 1 29
2 62746 1 29
2 62747 1 29
2 62748 1 29
2 62749 1 29
2 62750 1 29
2 62751 1 29
2 62752 1 29
2 62753 1 29
2 62754 1 29
2 62755 1 29
2 62756 1 29
2 62757 1 29
2 62758 1 29
2 62759 1 29
2 62760 1 29
2 62761 1 29
2 62762 1 29
2 62763 1 29
2 62764 1 29
2 62765 1 29
2 62766 1 29
2 62767 1 29
2 62768 1 29
2 62769 1 29
2 62770 1 29
2 62771 1 29
2 62772 1 29
2 62773 1 29
2 62774 1 29
2 62775 1 29
2 62776 1 29
2 62777 1 29
2 62778 1 29
2 62779 1 29
2 62780 1 29
2 62781 1 29
2 62782 1 29
2 62783 1 29
2 62784 1 29
2 62785 1 29
2 62786 1 29
2 62787 1 29
2 62788 1 29
2 62789 1 29
2 62790 1 29
2 62791 1 29
2 62792 1 29
2 62793 1 29
2 62794 1 29
2 62795 1 29
2 62796 1 29
2 62797 1 29
2 62798 1 29
2 62799 1 29
2 62800 1 29
2 62801 1 29
2 62802 1 29
2 62803 1 29
2 62804 1 29
2 62805 1 29
2 62806 1 29
2 62807 1 29
2 62808 1 29
2 62809 1 29
2 62810 1 29
2 62811 1 29
2 62812 1 29
2 62813 1 29
2 62814 1 29
2 62815 1 29
2 62816 1 29
2 62817 1 29
2 62818 1 29
2 62819 1 29
2 62820 1 29
2 62821 1 29
2 62822 1 29
2 62823 1 29
2 62824 1 30
2 62825 1 30
2 62826 1 30
2 62827 1 30
2 62828 1 30
2 62829 1 30
2 62830 1 30
2 62831 1 30
2 62832 1 30
2 62833 1 30
2 62834 1 30
2 62835 1 30
2 62836 1 30
2 62837 1 30
2 62838 1 30
2 62839 1 30
2 62840 1 30
2 62841 1 30
2 62842 1 30
2 62843 1 30
2 62844 1 30
2 62845 1 30
2 62846 1 30
2 62847 1 30
2 62848 1 30
2 62849 1 30
2 62850 1 30
2 62851 1 30
2 62852 1 30
2 62853 1 30
2 62854 1 30
2 62855 1 30
2 62856 1 30
2 62857 1 30
2 62858 1 30
2 62859 1 30
2 62860 1 30
2 62861 1 30
2 62862 1 30
2 62863 1 30
2 62864 1 30
2 62865 1 30
2 62866 1 30
2 62867 1 30
2 62868 1 30
2 62869 1 30
2 62870 1 30
2 62871 1 30
2 62872 1 30
2 62873 1 30
2 62874 1 30
2 62875 1 30
2 62876 1 30
2 62877 1 30
2 62878 1 30
2 62879 1 30
2 62880 1 30
2 62881 1 30
2 62882 1 30
2 62883 1 30
2 62884 1 30
2 62885 1 30
2 62886 1 30
2 62887 1 30
2 62888 1 30
2 62889 1 30
2 62890 1 30
2 62891 1 30
2 62892 1 30
2 62893 1 30
2 62894 1 30
2 62895 1 30
2 62896 1 30
2 62897 1 30
2 62898 1 30
2 62899 1 30
2 62900 1 30
2 62901 1 30
2 62902 1 30
2 62903 1 30
2 62904 1 30
2 62905 1 30
2 62906 1 30
2 62907 1 30
2 62908 1 30
2 62909 1 30
2 62910 1 30
2 62911 1 30
2 62912 1 30
2 62913 1 30
2 62914 1 30
2 62915 1 30
2 62916 1 30
2 62917 1 30
2 62918 1 30
2 62919 1 30
2 62920 1 30
2 62921 1 30
2 62922 1 30
2 62923 1 30
2 62924 1 30
2 62925 1 30
2 62926 1 30
2 62927 1 30
2 62928 1 30
2 62929 1 30
2 62930 1 30
2 62931 1 30
2 62932 1 30
2 62933 1 30
2 62934 1 30
2 62935 1 30
2 62936 1 30
2 62937 1 30
2 62938 1 30
2 62939 1 30
2 62940 1 30
2 62941 1 30
2 62942 1 30
2 62943 1 30
2 62944 1 30
2 62945 1 30
2 62946 1 30
2 62947 1 30
2 62948 1 30
2 62949 1 30
2 62950 1 30
2 62951 1 30
2 62952 1 30
2 62953 1 30
2 62954 1 30
2 62955 1 30
2 62956 1 30
2 62957 1 30
2 62958 1 30
2 62959 1 30
2 62960 1 30
2 62961 1 30
2 62962 1 30
2 62963 1 30
2 62964 1 30
2 62965 1 30
2 62966 1 30
2 62967 1 30
2 62968 1 30
2 62969 1 30
2 62970 1 30
2 62971 1 30
2 62972 1 30
2 62973 1 30
2 62974 1 30
2 62975 1 30
2 62976 1 30
2 62977 1 30
2 62978 1 30
2 62979 1 30
2 62980 1 30
2 62981 1 30
2 62982 1 30
2 62983 1 30
2 62984 1 30
2 62985 1 30
2 62986 1 30
2 62987 1 30
2 62988 1 30
2 62989 1 30
2 62990 1 30
2 62991 1 30
2 62992 1 30
2 62993 1 30
2 62994 1 30
2 62995 1 30
2 62996 1 30
2 62997 1 30
2 62998 1 30
2 62999 1 30
2 63000 1 30
2 63001 1 30
2 63002 1 30
2 63003 1 30
2 63004 1 30
2 63005 1 30
2 63006 1 30
2 63007 1 30
2 63008 1 30
2 63009 1 30
2 63010 1 30
2 63011 1 30
2 63012 1 30
2 63013 1 30
2 63014 1 30
2 63015 1 30
2 63016 1 30
2 63017 1 30
2 63018 1 30
2 63019 1 30
2 63020 1 30
2 63021 1 30
2 63022 1 30
2 63023 1 30
2 63024 1 30
2 63025 1 30
2 63026 1 30
2 63027 1 30
2 63028 1 30
2 63029 1 30
2 63030 1 30
2 63031 1 30
2 63032 1 30
2 63033 1 30
2 63034 1 30
2 63035 1 30
2 63036 1 30
2 63037 1 30
2 63038 1 30
2 63039 1 30
2 63040 1 30
2 63041 1 30
2 63042 1 30
2 63043 1 30
2 63044 1 30
2 63045 1 30
2 63046 1 30
2 63047 1 30
2 63048 1 30
2 63049 1 30
2 63050 1 30
2 63051 1 30
2 63052 1 30
2 63053 1 30
2 63054 1 30
2 63055 1 30
2 63056 1 30
2 63057 1 30
2 63058 1 30
2 63059 1 30
2 63060 1 30
2 63061 1 30
2 63062 1 30
2 63063 1 30
2 63064 1 30
2 63065 1 30
2 63066 1 30
2 63067 1 30
2 63068 1 30
2 63069 1 30
2 63070 1 30
2 63071 1 30
2 63072 1 30
2 63073 1 30
2 63074 1 30
2 63075 1 30
2 63076 1 30
2 63077 1 30
2 63078 1 30
2 63079 1 30
2 63080 1 30
2 63081 1 30
2 63082 1 30
2 63083 1 30
2 63084 1 30
2 63085 1 30
2 63086 1 30
2 63087 1 30
2 63088 1 30
2 63089 1 30
2 63090 1 30
2 63091 1 30
2 63092 1 30
2 63093 1 30
2 63094 1 30
2 63095 1 30
2 63096 1 30
2 63097 1 30
2 63098 1 30
2 63099 1 30
2 63100 1 30
2 63101 1 30
2 63102 1 30
2 63103 1 30
2 63104 1 30
2 63105 1 30
2 63106 1 30
2 63107 1 30
2 63108 1 30
2 63109 1 30
2 63110 1 30
2 63111 1 30
2 63112 1 30
2 63113 1 30
2 63114 1 30
2 63115 1 30
2 63116 1 30
2 63117 1 30
2 63118 1 30
2 63119 1 30
2 63120 1 30
2 63121 1 30
2 63122 1 30
2 63123 1 30
2 63124 1 30
2 63125 1 31
2 63126 1 31
2 63127 1 31
2 63128 1 31
2 63129 1 31
2 63130 1 31
2 63131 1 31
2 63132 1 31
2 63133 1 31
2 63134 1 31
2 63135 1 31
2 63136 1 31
2 63137 1 31
2 63138 1 31
2 63139 1 31
2 63140 1 31
2 63141 1 31
2 63142 1 31
2 63143 1 31
2 63144 1 31
2 63145 1 31
2 63146 1 31
2 63147 1 31
2 63148 1 31
2 63149 1 31
2 63150 1 31
2 63151 1 31
2 63152 1 31
2 63153 1 31
2 63154 1 31
2 63155 1 31
2 63156 1 31
2 63157 1 31
2 63158 1 31
2 63159 1 31
2 63160 1 31
2 63161 1 31
2 63162 1 31
2 63163 1 31
2 63164 1 31
2 63165 1 31
2 63166 1 31
2 63167 1 31
2 63168 1 31
2 63169 1 31
2 63170 1 31
2 63171 1 31
2 63172 1 31
2 63173 1 31
2 63174 1 31
2 63175 1 31
2 63176 1 31
2 63177 1 31
2 63178 1 31
2 63179 1 31
2 63180 1 31
2 63181 1 31
2 63182 1 31
2 63183 1 31
2 63184 1 31
2 63185 1 31
2 63186 1 31
2 63187 1 31
2 63188 1 31
2 63189 1 31
2 63190 1 31
2 63191 1 31
2 63192 1 31
2 63193 1 31
2 63194 1 31
2 63195 1 31
2 63196 1 31
2 63197 1 31
2 63198 1 31
2 63199 1 31
2 63200 1 31
2 63201 1 31
2 63202 1 31
2 63203 1 31
2 63204 1 31
2 63205 1 31
2 63206 1 31
2 63207 1 31
2 63208 1 31
2 63209 1 31
2 63210 1 31
2 63211 1 31
2 63212 1 31
2 63213 1 31
2 63214 1 31
2 63215 1 31
2 63216 1 31
2 63217 1 31
2 63218 1 31
2 63219 1 31
2 63220 1 31
2 63221 1 31
2 63222 1 31
2 63223 1 31
2 63224 1 31
2 63225 1 31
2 63226 1 31
2 63227 1 31
2 63228 1 31
2 63229 1 31
2 63230 1 31
2 63231 1 31
2 63232 1 31
2 63233 1 31
2 63234 1 31
2 63235 1 31
2 63236 1 31
2 63237 1 31
2 63238 1 31
2 63239 1 31
2 63240 1 31
2 63241 1 31
2 63242 1 31
2 63243 1 31
2 63244 1 31
2 63245 1 31
2 63246 1 31
2 63247 1 31
2 63248 1 31
2 63249 1 31
2 63250 1 31
2 63251 1 31
2 63252 1 31
2 63253 1 31
2 63254 1 31
2 63255 1 31
2 63256 1 31
2 63257 1 31
2 63258 1 31
2 63259 1 31
2 63260 1 31
2 63261 1 31
2 63262 1 31
2 63263 1 31
2 63264 1 31
2 63265 1 31
2 63266 1 31
2 63267 1 31
2 63268 1 31
2 63269 1 31
2 63270 1 31
2 63271 1 31
2 63272 1 31
2 63273 1 31
2 63274 1 31
2 63275 1 31
2 63276 1 31
2 63277 1 31
2 63278 1 31
2 63279 1 31
2 63280 1 31
2 63281 1 31
2 63282 1 31
2 63283 1 31
2 63284 1 31
2 63285 1 31
2 63286 1 31
2 63287 1 31
2 63288 1 31
2 63289 1 31
2 63290 1 31
2 63291 1 31
2 63292 1 31
2 63293 1 31
2 63294 1 31
2 63295 1 31
2 63296 1 31
2 63297 1 31
2 63298 1 31
2 63299 1 31
2 63300 1 31
2 63301 1 31
2 63302 1 31
2 63303 1 31
2 63304 1 31
2 63305 1 31
2 63306 1 31
2 63307 1 31
2 63308 1 31
2 63309 1 31
2 63310 1 31
2 63311 1 31
2 63312 1 31
2 63313 1 31
2 63314 1 31
2 63315 1 31
2 63316 1 31
2 63317 1 31
2 63318 1 31
2 63319 1 31
2 63320 1 31
2 63321 1 31
2 63322 1 31
2 63323 1 31
2 63324 1 31
2 63325 1 31
2 63326 1 31
2 63327 1 31
2 63328 1 31
2 63329 1 31
2 63330 1 31
2 63331 1 31
2 63332 1 31
2 63333 1 31
2 63334 1 31
2 63335 1 31
2 63336 1 31
2 63337 1 31
2 63338 1 31
2 63339 1 31
2 63340 1 31
2 63341 1 31
2 63342 1 31
2 63343 1 31
2 63344 1 31
2 63345 1 31
2 63346 1 31
2 63347 1 31
2 63348 1 31
2 63349 1 31
2 63350 1 31
2 63351 1 31
2 63352 1 31
2 63353 1 31
2 63354 1 31
2 63355 1 31
2 63356 1 31
2 63357 1 31
2 63358 1 31
2 63359 1 31
2 63360 1 31
2 63361 1 31
2 63362 1 31
2 63363 1 31
2 63364 1 31
2 63365 1 31
2 63366 1 31
2 63367 1 31
2 63368 1 31
2 63369 1 31
2 63370 1 31
2 63371 1 31
2 63372 1 31
2 63373 1 31
2 63374 1 31
2 63375 1 31
2 63376 1 31
2 63377 1 31
2 63378 1 31
2 63379 1 31
2 63380 1 31
2 63381 1 31
2 63382 1 31
2 63383 1 31
2 63384 1 31
2 63385 1 31
2 63386 1 31
2 63387 1 31
2 63388 1 31
2 63389 1 31
2 63390 1 31
2 63391 1 31
2 63392 1 31
2 63393 1 31
2 63394 1 31
2 63395 1 31
2 63396 1 31
2 63397 1 31
2 63398 1 31
2 63399 1 31
2 63400 1 31
2 63401 1 31
2 63402 1 31
2 63403 1 31
2 63404 1 31
2 63405 1 31
2 63406 1 31
2 63407 1 31
2 63408 1 31
2 63409 1 31
2 63410 1 31
2 63411 1 31
2 63412 1 31
2 63413 1 31
2 63414 1 31
2 63415 1 31
2 63416 1 31
2 63417 1 31
2 63418 1 31
2 63419 1 31
2 63420 1 31
2 63421 1 31
2 63422 1 31
2 63423 1 31
2 63424 1 31
2 63425 1 31
2 63426 1 31
2 63427 1 31
2 63428 1 31
2 63429 1 31
2 63430 1 31
2 63431 1 31
2 63432 1 31
2 63433 1 31
2 63434 1 31
2 63435 1 31
2 63436 1 31
2 63437 1 32
2 63438 1 32
2 63439 1 32
2 63440 1 32
2 63441 1 32
2 63442 1 32
2 63443 1 32
2 63444 1 32
2 63445 1 32
2 63446 1 32
2 63447 1 32
2 63448 1 32
2 63449 1 32
2 63450 1 32
2 63451 1 32
2 63452 1 32
2 63453 1 32
2 63454 1 32
2 63455 1 32
2 63456 1 32
2 63457 1 32
2 63458 1 32
2 63459 1 32
2 63460 1 32
2 63461 1 32
2 63462 1 32
2 63463 1 32
2 63464 1 32
2 63465 1 32
2 63466 1 32
2 63467 1 32
2 63468 1 32
2 63469 1 32
2 63470 1 32
2 63471 1 32
2 63472 1 32
2 63473 1 32
2 63474 1 32
2 63475 1 32
2 63476 1 32
2 63477 1 32
2 63478 1 32
2 63479 1 32
2 63480 1 32
2 63481 1 32
2 63482 1 32
2 63483 1 32
2 63484 1 32
2 63485 1 32
2 63486 1 32
2 63487 1 32
2 63488 1 32
2 63489 1 32
2 63490 1 32
2 63491 1 32
2 63492 1 32
2 63493 1 32
2 63494 1 32
2 63495 1 32
2 63496 1 32
2 63497 1 32
2 63498 1 32
2 63499 1 32
2 63500 1 32
2 63501 1 32
2 63502 1 32
2 63503 1 32
2 63504 1 32
2 63505 1 32
2 63506 1 32
2 63507 1 32
2 63508 1 32
2 63509 1 32
2 63510 1 32
2 63511 1 32
2 63512 1 32
2 63513 1 32
2 63514 1 32
2 63515 1 32
2 63516 1 32
2 63517 1 32
2 63518 1 32
2 63519 1 32
2 63520 1 32
2 63521 1 32
2 63522 1 32
2 63523 1 32
2 63524 1 32
2 63525 1 32
2 63526 1 32
2 63527 1 32
2 63528 1 32
2 63529 1 32
2 63530 1 32
2 63531 1 32
2 63532 1 32
2 63533 1 32
2 63534 1 32
2 63535 1 32
2 63536 1 32
2 63537 1 32
2 63538 1 32
2 63539 1 32
2 63540 1 32
2 63541 1 32
2 63542 1 32
2 63543 1 32
2 63544 1 32
2 63545 1 32
2 63546 1 32
2 63547 1 32
2 63548 1 32
2 63549 1 32
2 63550 1 32
2 63551 1 32
2 63552 1 32
2 63553 1 32
2 63554 1 32
2 63555 1 32
2 63556 1 32
2 63557 1 32
2 63558 1 32
2 63559 1 32
2 63560 1 32
2 63561 1 32
2 63562 1 33
2 63563 1 33
2 63564 1 33
2 63565 1 33
2 63566 1 33
2 63567 1 33
2 63568 1 33
2 63569 1 33
2 63570 1 33
2 63571 1 33
2 63572 1 33
2 63573 1 33
2 63574 1 33
2 63575 1 33
2 63576 1 33
2 63577 1 33
2 63578 1 33
2 63579 1 33
2 63580 1 33
2 63581 1 33
2 63582 1 33
2 63583 1 33
2 63584 1 33
2 63585 1 33
2 63586 1 33
2 63587 1 33
2 63588 1 33
2 63589 1 33
2 63590 1 33
2 63591 1 33
2 63592 1 33
2 63593 1 33
2 63594 1 33
2 63595 1 33
2 63596 1 33
2 63597 1 33
2 63598 1 33
2 63599 1 33
2 63600 1 33
2 63601 1 33
2 63602 1 33
2 63603 1 33
2 63604 1 33
2 63605 1 33
2 63606 1 33
2 63607 1 33
2 63608 1 33
2 63609 1 33
2 63610 1 33
2 63611 1 33
2 63612 1 33
2 63613 1 33
2 63614 1 33
2 63615 1 33
2 63616 1 33
2 63617 1 33
2 63618 1 33
2 63619 1 33
2 63620 1 33
2 63621 1 33
2 63622 1 33
2 63623 1 33
2 63624 1 33
2 63625 1 33
2 63626 1 33
2 63627 1 33
2 63628 1 33
2 63629 1 33
2 63630 1 33
2 63631 1 33
2 63632 1 33
2 63633 1 33
2 63634 1 33
2 63635 1 33
2 63636 1 33
2 63637 1 33
2 63638 1 33
2 63639 1 33
2 63640 1 33
2 63641 1 33
2 63642 1 33
2 63643 1 33
2 63644 1 33
2 63645 1 33
2 63646 1 33
2 63647 1 33
2 63648 1 33
2 63649 1 33
2 63650 1 33
2 63651 1 33
2 63652 1 33
2 63653 1 33
2 63654 1 33
2 63655 1 33
2 63656 1 33
2 63657 1 34
2 63658 1 34
2 63659 1 34
2 63660 1 34
2 63661 1 34
2 63662 1 34
2 63663 1 34
2 63664 1 34
2 63665 1 34
2 63666 1 34
2 63667 1 34
2 63668 1 34
2 63669 1 34
2 63670 1 34
2 63671 1 34
2 63672 1 34
2 63673 1 34
2 63674 1 34
2 63675 1 34
2 63676 1 34
2 63677 1 34
2 63678 1 34
2 63679 1 34
2 63680 1 34
2 63681 1 34
2 63682 1 34
2 63683 1 34
2 63684 1 34
2 63685 1 34
2 63686 1 34
2 63687 1 34
2 63688 1 34
2 63689 1 34
2 63690 1 34
2 63691 1 34
2 63692 1 34
2 63693 1 34
2 63694 1 34
2 63695 1 34
2 63696 1 34
2 63697 1 34
2 63698 1 34
2 63699 1 34
2 63700 1 34
2 63701 1 34
2 63702 1 34
2 63703 1 34
2 63704 1 34
2 63705 1 34
2 63706 1 34
2 63707 1 34
2 63708 1 34
2 63709 1 34
2 63710 1 34
2 63711 1 34
2 63712 1 34
2 63713 1 34
2 63714 1 34
2 63715 1 34
2 63716 1 34
2 63717 1 34
2 63718 1 34
2 63719 1 34
2 63720 1 34
2 63721 1 34
2 63722 1 34
2 63723 1 34
2 63724 1 34
2 63725 1 34
2 63726 1 34
2 63727 1 34
2 63728 1 34
2 63729 1 34
2 63730 1 34
2 63731 1 34
2 63732 1 34
2 63733 1 34
2 63734 1 35
2 63735 1 35
2 63736 1 35
2 63737 1 35
2 63738 1 35
2 63739 1 35
2 63740 1 35
2 63741 1 35
2 63742 1 35
2 63743 1 35
2 63744 1 35
2 63745 1 35
2 63746 1 35
2 63747 1 35
2 63748 1 35
2 63749 1 35
2 63750 1 35
2 63751 1 35
2 63752 1 35
2 63753 1 35
2 63754 1 35
2 63755 1 35
2 63756 1 35
2 63757 1 35
2 63758 1 35
2 63759 1 35
2 63760 1 35
2 63761 1 35
2 63762 1 35
2 63763 1 35
2 63764 1 35
2 63765 1 35
2 63766 1 35
2 63767 1 35
2 63768 1 35
2 63769 1 35
2 63770 1 35
2 63771 1 35
2 63772 1 35
2 63773 1 35
2 63774 1 35
2 63775 1 35
2 63776 1 35
2 63777 1 35
2 63778 1 35
2 63779 1 35
2 63780 1 35
2 63781 1 35
2 63782 1 35
2 63783 1 35
2 63784 1 35
2 63785 1 35
2 63786 1 35
2 63787 1 35
2 63788 1 35
2 63789 1 35
2 63790 1 35
2 63791 1 36
2 63792 1 36
2 63793 1 36
2 63794 1 36
2 63795 1 36
2 63796 1 36
2 63797 1 36
2 63798 1 36
2 63799 1 36
2 63800 1 36
2 63801 1 36
2 63802 1 36
2 63803 1 36
2 63804 1 36
2 63805 1 36
2 63806 1 36
2 63807 1 36
2 63808 1 36
2 63809 1 36
2 63810 1 36
2 63811 1 36
2 63812 1 36
2 63813 1 36
2 63814 1 36
2 63815 1 36
2 63816 1 36
2 63817 1 36
2 63818 1 36
2 63819 1 36
2 63820 1 36
2 63821 1 36
2 63822 1 36
2 63823 1 36
2 63824 1 36
2 63825 1 36
2 63826 1 36
2 63827 1 36
2 63828 1 36
2 63829 1 36
2 63830 1 36
2 63831 1 36
2 63832 1 36
2 63833 1 36
2 63834 1 36
2 63835 1 36
2 63836 1 36
2 63837 1 36
2 63838 1 36
2 63839 1 36
2 63840 1 36
2 63841 1 36
2 63842 1 36
2 63843 1 36
2 63844 1 36
2 63845 1 36
2 63846 1 36
2 63847 1 36
2 63848 1 36
2 63849 1 36
2 63850 1 36
2 63851 1 36
2 63852 1 36
2 63853 1 36
2 63854 1 36
2 63855 1 36
2 63856 1 36
2 63857 1 36
2 63858 1 36
2 63859 1 36
2 63860 1 36
2 63861 1 36
2 63862 1 36
2 63863 1 36
2 63864 1 36
2 63865 1 36
2 63866 1 36
2 63867 1 36
2 63868 1 36
2 63869 1 36
2 63870 1 36
2 63871 1 36
2 63872 1 36
2 63873 1 36
2 63874 1 36
2 63875 1 36
2 63876 1 36
2 63877 1 36
2 63878 1 36
2 63879 1 36
2 63880 1 36
2 63881 1 36
2 63882 1 36
2 63883 1 36
2 63884 1 36
2 63885 1 36
2 63886 1 36
2 63887 1 36
2 63888 1 36
2 63889 1 36
2 63890 1 36
2 63891 1 36
2 63892 1 36
2 63893 1 36
2 63894 1 36
2 63895 1 36
2 63896 1 36
2 63897 1 36
2 63898 1 36
2 63899 1 36
2 63900 1 36
2 63901 1 36
2 63902 1 36
2 63903 1 36
2 63904 1 36
2 63905 1 36
2 63906 1 36
2 63907 1 36
2 63908 1 36
2 63909 1 36
2 63910 1 36
2 63911 1 36
2 63912 1 36
2 63913 1 36
2 63914 1 36
2 63915 1 36
2 63916 1 36
2 63917 1 36
2 63918 1 36
2 63919 1 36
2 63920 1 36
2 63921 1 36
2 63922 1 36
2 63923 1 36
2 63924 1 36
2 63925 1 37
2 63926 1 37
2 63927 1 37
2 63928 1 37
2 63929 1 37
2 63930 1 37
2 63931 1 37
2 63932 1 37
2 63933 1 37
2 63934 1 37
2 63935 1 37
2 63936 1 37
2 63937 1 37
2 63938 1 37
2 63939 1 37
2 63940 1 37
2 63941 1 37
2 63942 1 37
2 63943 1 37
2 63944 1 37
2 63945 1 37
2 63946 1 37
2 63947 1 37
2 63948 1 37
2 63949 1 37
2 63950 1 37
2 63951 1 37
2 63952 1 37
2 63953 1 37
2 63954 1 37
2 63955 1 37
2 63956 1 37
2 63957 1 37
2 63958 1 37
2 63959 1 37
2 63960 1 37
2 63961 1 37
2 63962 1 37
2 63963 1 37
2 63964 1 37
2 63965 1 37
2 63966 1 37
2 63967 1 37
2 63968 1 37
2 63969 1 37
2 63970 1 37
2 63971 1 37
2 63972 1 37
2 63973 1 37
2 63974 1 37
2 63975 1 37
2 63976 1 37
2 63977 1 37
2 63978 1 37
2 63979 1 37
2 63980 1 37
2 63981 1 37
2 63982 1 37
2 63983 1 37
2 63984 1 37
2 63985 1 37
2 63986 1 37
2 63987 1 37
2 63988 1 37
2 63989 1 37
2 63990 1 37
2 63991 1 37
2 63992 1 37
2 63993 1 37
2 63994 1 37
2 63995 1 37
2 63996 1 37
2 63997 1 37
2 63998 1 37
2 63999 1 37
2 64000 1 37
2 64001 1 37
2 64002 1 37
2 64003 1 37
2 64004 1 37
2 64005 1 37
2 64006 1 37
2 64007 1 37
2 64008 1 37
2 64009 1 37
2 64010 1 37
2 64011 1 37
2 64012 1 37
2 64013 1 37
2 64014 1 37
2 64015 1 37
2 64016 1 37
2 64017 1 37
2 64018 1 37
2 64019 1 37
2 64020 1 37
2 64021 1 37
2 64022 1 37
2 64023 1 37
2 64024 1 37
2 64025 1 37
2 64026 1 37
2 64027 1 37
2 64028 1 37
2 64029 1 37
2 64030 1 37
2 64031 1 37
2 64032 1 37
2 64033 1 37
2 64034 1 37
2 64035 1 37
2 64036 1 37
2 64037 1 37
2 64038 1 37
2 64039 1 37
2 64040 1 37
2 64041 1 37
2 64042 1 37
2 64043 1 37
2 64044 1 37
2 64045 1 37
2 64046 1 37
2 64047 1 37
2 64048 1 37
2 64049 1 37
2 64050 1 37
2 64051 1 37
2 64052 1 37
2 64053 1 37
2 64054 1 37
2 64055 1 37
2 64056 1 37
2 64057 1 37
2 64058 1 37
2 64059 1 37
2 64060 1 37
2 64061 1 37
2 64062 1 37
2 64063 1 37
2 64064 1 37
2 64065 1 37
2 64066 1 37
2 64067 1 37
2 64068 1 37
2 64069 1 37
2 64070 1 37
2 64071 1 37
2 64072 1 37
2 64073 1 37
2 64074 1 37
2 64075 1 37
2 64076 1 37
2 64077 1 37
2 64078 1 37
2 64079 1 37
2 64080 1 37
2 64081 1 37
2 64082 1 37
2 64083 1 37
2 64084 1 37
2 64085 1 37
2 64086 1 37
2 64087 1 37
2 64088 1 37
2 64089 1 37
2 64090 1 37
2 64091 1 37
2 64092 1 37
2 64093 1 37
2 64094 1 37
2 64095 1 37
2 64096 1 37
2 64097 1 37
2 64098 1 37
2 64099 1 37
2 64100 1 37
2 64101 1 37
2 64102 1 37
2 64103 1 37
2 64104 1 37
2 64105 1 37
2 64106 1 37
2 64107 1 37
2 64108 1 37
2 64109 1 37
2 64110 1 37
2 64111 1 37
2 64112 1 37
2 64113 1 37
2 64114 1 37
2 64115 1 37
2 64116 1 37
2 64117 1 37
2 64118 1 37
2 64119 1 38
2 64120 1 38
2 64121 1 38
2 64122 1 38
2 64123 1 38
2 64124 1 38
2 64125 1 38
2 64126 1 38
2 64127 1 38
2 64128 1 38
2 64129 1 38
2 64130 1 38
2 64131 1 38
2 64132 1 38
2 64133 1 38
2 64134 1 38
2 64135 1 38
2 64136 1 38
2 64137 1 38
2 64138 1 38
2 64139 1 38
2 64140 1 38
2 64141 1 38
2 64142 1 38
2 64143 1 38
2 64144 1 38
2 64145 1 38
2 64146 1 38
2 64147 1 38
2 64148 1 38
2 64149 1 38
2 64150 1 38
2 64151 1 38
2 64152 1 38
2 64153 1 38
2 64154 1 38
2 64155 1 38
2 64156 1 38
2 64157 1 38
2 64158 1 38
2 64159 1 38
2 64160 1 38
2 64161 1 38
2 64162 1 38
2 64163 1 38
2 64164 1 38
2 64165 1 38
2 64166 1 38
2 64167 1 38
2 64168 1 38
2 64169 1 38
2 64170 1 38
2 64171 1 38
2 64172 1 38
2 64173 1 38
2 64174 1 38
2 64175 1 38
2 64176 1 38
2 64177 1 38
2 64178 1 38
2 64179 1 38
2 64180 1 38
2 64181 1 38
2 64182 1 38
2 64183 1 38
2 64184 1 38
2 64185 1 38
2 64186 1 38
2 64187 1 38
2 64188 1 38
2 64189 1 38
2 64190 1 38
2 64191 1 38
2 64192 1 38
2 64193 1 38
2 64194 1 38
2 64195 1 38
2 64196 1 38
2 64197 1 38
2 64198 1 38
2 64199 1 38
2 64200 1 38
2 64201 1 38
2 64202 1 38
2 64203 1 38
2 64204 1 38
2 64205 1 38
2 64206 1 38
2 64207 1 38
2 64208 1 38
2 64209 1 38
2 64210 1 38
2 64211 1 38
2 64212 1 38
2 64213 1 38
2 64214 1 38
2 64215 1 38
2 64216 1 38
2 64217 1 38
2 64218 1 38
2 64219 1 38
2 64220 1 38
2 64221 1 38
2 64222 1 38
2 64223 1 38
2 64224 1 38
2 64225 1 38
2 64226 1 38
2 64227 1 38
2 64228 1 38
2 64229 1 38
2 64230 1 38
2 64231 1 38
2 64232 1 38
2 64233 1 38
2 64234 1 38
2 64235 1 38
2 64236 1 38
2 64237 1 38
2 64238 1 38
2 64239 1 38
2 64240 1 38
2 64241 1 38
2 64242 1 38
2 64243 1 38
2 64244 1 38
2 64245 1 38
2 64246 1 38
2 64247 1 38
2 64248 1 38
2 64249 1 38
2 64250 1 38
2 64251 1 38
2 64252 1 38
2 64253 1 38
2 64254 1 38
2 64255 1 38
2 64256 1 38
2 64257 1 38
2 64258 1 38
2 64259 1 38
2 64260 1 38
2 64261 1 38
2 64262 1 38
2 64263 1 38
2 64264 1 38
2 64265 1 38
2 64266 1 38
2 64267 1 38
2 64268 1 38
2 64269 1 38
2 64270 1 38
2 64271 1 38
2 64272 1 38
2 64273 1 38
2 64274 1 38
2 64275 1 38
2 64276 1 38
2 64277 1 38
2 64278 1 38
2 64279 1 38
2 64280 1 38
2 64281 1 38
2 64282 1 38
2 64283 1 38
2 64284 1 38
2 64285 1 38
2 64286 1 38
2 64287 1 38
2 64288 1 38
2 64289 1 38
2 64290 1 38
2 64291 1 38
2 64292 1 38
2 64293 1 38
2 64294 1 38
2 64295 1 38
2 64296 1 38
2 64297 1 38
2 64298 1 38
2 64299 1 38
2 64300 1 38
2 64301 1 38
2 64302 1 38
2 64303 1 38
2 64304 1 38
2 64305 1 38
2 64306 1 38
2 64307 1 38
2 64308 1 38
2 64309 1 38
2 64310 1 38
2 64311 1 38
2 64312 1 38
2 64313 1 38
2 64314 1 38
2 64315 1 38
2 64316 1 38
2 64317 1 38
2 64318 1 38
2 64319 1 38
2 64320 1 38
2 64321 1 38
2 64322 1 38
2 64323 1 38
2 64324 1 38
2 64325 1 38
2 64326 1 38
2 64327 1 38
2 64328 1 38
2 64329 1 38
2 64330 1 38
2 64331 1 38
2 64332 1 38
2 64333 1 38
2 64334 1 38
2 64335 1 38
2 64336 1 38
2 64337 1 38
2 64338 1 38
2 64339 1 38
2 64340 1 38
2 64341 1 38
2 64342 1 38
2 64343 1 38
2 64344 1 38
2 64345 1 38
2 64346 1 38
2 64347 1 38
2 64348 1 38
2 64349 1 38
2 64350 1 38
2 64351 1 38
2 64352 1 38
2 64353 1 38
2 64354 1 38
2 64355 1 38
2 64356 1 38
2 64357 1 38
2 64358 1 38
2 64359 1 38
2 64360 1 38
2 64361 1 38
2 64362 1 38
2 64363 1 38
2 64364 1 38
2 64365 1 38
2 64366 1 38
2 64367 1 38
2 64368 1 38
2 64369 1 38
2 64370 1 38
2 64371 1 38
2 64372 1 38
2 64373 1 38
2 64374 1 38
2 64375 1 38
2 64376 1 38
2 64377 1 38
2 64378 1 38
2 64379 1 38
2 64380 1 38
2 64381 1 38
2 64382 1 38
2 64383 1 38
2 64384 1 38
2 64385 1 38
2 64386 1 38
2 64387 1 38
2 64388 1 38
2 64389 1 38
2 64390 1 38
2 64391 1 38
2 64392 1 38
2 64393 1 38
2 64394 1 38
2 64395 1 38
2 64396 1 38
2 64397 1 38
2 64398 1 38
2 64399 1 38
2 64400 1 38
2 64401 1 38
2 64402 1 38
2 64403 1 38
2 64404 1 38
2 64405 1 38
2 64406 1 38
2 64407 1 38
2 64408 1 38
2 64409 1 38
2 64410 1 38
2 64411 1 38
2 64412 1 38
2 64413 1 38
2 64414 1 38
2 64415 1 38
2 64416 1 38
2 64417 1 38
2 64418 1 38
2 64419 1 38
2 64420 1 38
2 64421 1 38
2 64422 1 38
2 64423 1 38
2 64424 1 38
2 64425 1 38
2 64426 1 38
2 64427 1 38
2 64428 1 38
2 64429 1 38
2 64430 1 38
2 64431 1 38
2 64432 1 38
2 64433 1 39
2 64434 1 39
2 64435 1 39
2 64436 1 39
2 64437 1 39
2 64438 1 39
2 64439 1 39
2 64440 1 39
2 64441 1 39
2 64442 1 39
2 64443 1 39
2 64444 1 39
2 64445 1 39
2 64446 1 39
2 64447 1 39
2 64448 1 39
2 64449 1 39
2 64450 1 39
2 64451 1 39
2 64452 1 39
2 64453 1 39
2 64454 1 39
2 64455 1 39
2 64456 1 39
2 64457 1 39
2 64458 1 39
2 64459 1 39
2 64460 1 39
2 64461 1 39
2 64462 1 39
2 64463 1 39
2 64464 1 39
2 64465 1 39
2 64466 1 39
2 64467 1 39
2 64468 1 39
2 64469 1 39
2 64470 1 39
2 64471 1 39
2 64472 1 39
2 64473 1 39
2 64474 1 39
2 64475 1 39
2 64476 1 39
2 64477 1 39
2 64478 1 39
2 64479 1 39
2 64480 1 39
2 64481 1 39
2 64482 1 39
2 64483 1 39
2 64484 1 39
2 64485 1 39
2 64486 1 39
2 64487 1 39
2 64488 1 39
2 64489 1 39
2 64490 1 39
2 64491 1 39
2 64492 1 39
2 64493 1 39
2 64494 1 39
2 64495 1 39
2 64496 1 39
2 64497 1 39
2 64498 1 39
2 64499 1 39
2 64500 1 39
2 64501 1 39
2 64502 1 39
2 64503 1 39
2 64504 1 39
2 64505 1 39
2 64506 1 39
2 64507 1 39
2 64508 1 39
2 64509 1 39
2 64510 1 39
2 64511 1 39
2 64512 1 39
2 64513 1 39
2 64514 1 39
2 64515 1 39
2 64516 1 39
2 64517 1 39
2 64518 1 39
2 64519 1 39
2 64520 1 39
2 64521 1 39
2 64522 1 39
2 64523 1 39
2 64524 1 39
2 64525 1 39
2 64526 1 39
2 64527 1 39
2 64528 1 39
2 64529 1 39
2 64530 1 39
2 64531 1 39
2 64532 1 39
2 64533 1 39
2 64534 1 39
2 64535 1 39
2 64536 1 39
2 64537 1 39
2 64538 1 39
2 64539 1 39
2 64540 1 39
2 64541 1 39
2 64542 1 39
2 64543 1 39
2 64544 1 39
2 64545 1 39
2 64546 1 39
2 64547 1 39
2 64548 1 39
2 64549 1 39
2 64550 1 39
2 64551 1 39
2 64552 1 39
2 64553 1 39
2 64554 1 39
2 64555 1 39
2 64556 1 39
2 64557 1 39
2 64558 1 39
2 64559 1 39
2 64560 1 39
2 64561 1 39
2 64562 1 39
2 64563 1 39
2 64564 1 39
2 64565 1 39
2 64566 1 39
2 64567 1 39
2 64568 1 39
2 64569 1 39
2 64570 1 39
2 64571 1 39
2 64572 1 39
2 64573 1 39
2 64574 1 39
2 64575 1 39
2 64576 1 39
2 64577 1 39
2 64578 1 39
2 64579 1 39
2 64580 1 39
2 64581 1 39
2 64582 1 39
2 64583 1 39
2 64584 1 39
2 64585 1 39
2 64586 1 39
2 64587 1 39
2 64588 1 39
2 64589 1 39
2 64590 1 39
2 64591 1 39
2 64592 1 39
2 64593 1 39
2 64594 1 39
2 64595 1 39
2 64596 1 39
2 64597 1 39
2 64598 1 39
2 64599 1 39
2 64600 1 39
2 64601 1 39
2 64602 1 39
2 64603 1 39
2 64604 1 39
2 64605 1 39
2 64606 1 39
2 64607 1 39
2 64608 1 39
2 64609 1 39
2 64610 1 39
2 64611 1 39
2 64612 1 39
2 64613 1 39
2 64614 1 39
2 64615 1 39
2 64616 1 39
2 64617 1 39
2 64618 1 39
2 64619 1 39
2 64620 1 39
2 64621 1 39
2 64622 1 39
2 64623 1 39
2 64624 1 39
2 64625 1 39
2 64626 1 39
2 64627 1 39
2 64628 1 39
2 64629 1 39
2 64630 1 39
2 64631 1 39
2 64632 1 39
2 64633 1 39
2 64634 1 39
2 64635 1 39
2 64636 1 39
2 64637 1 39
2 64638 1 39
2 64639 1 39
2 64640 1 39
2 64641 1 39
2 64642 1 39
2 64643 1 39
2 64644 1 39
2 64645 1 39
2 64646 1 39
2 64647 1 39
2 64648 1 39
2 64649 1 39
2 64650 1 39
2 64651 1 39
2 64652 1 39
2 64653 1 40
2 64654 1 40
2 64655 1 40
2 64656 1 40
2 64657 1 40
2 64658 1 40
2 64659 1 40
2 64660 1 40
2 64661 1 40
2 64662 1 40
2 64663 1 40
2 64664 1 40
2 64665 1 40
2 64666 1 40
2 64667 1 40
2 64668 1 40
2 64669 1 40
2 64670 1 40
2 64671 1 40
2 64672 1 40
2 64673 1 40
2 64674 1 40
2 64675 1 40
2 64676 1 40
2 64677 1 40
2 64678 1 40
2 64679 1 40
2 64680 1 40
2 64681 1 40
2 64682 1 40
2 64683 1 40
2 64684 1 40
2 64685 1 40
2 64686 1 40
2 64687 1 40
2 64688 1 40
2 64689 1 40
2 64690 1 40
2 64691 1 40
2 64692 1 40
2 64693 1 40
2 64694 1 40
2 64695 1 40
2 64696 1 40
2 64697 1 40
2 64698 1 40
2 64699 1 40
2 64700 1 40
2 64701 1 40
2 64702 1 40
2 64703 1 40
2 64704 1 40
2 64705 1 40
2 64706 1 40
2 64707 1 40
2 64708 1 40
2 64709 1 40
2 64710 1 40
2 64711 1 40
2 64712 1 40
2 64713 1 40
2 64714 1 40
2 64715 1 40
2 64716 1 40
2 64717 1 40
2 64718 1 40
2 64719 1 40
2 64720 1 40
2 64721 1 40
2 64722 1 40
2 64723 1 40
2 64724 1 40
2 64725 1 40
2 64726 1 40
2 64727 1 40
2 64728 1 40
2 64729 1 40
2 64730 1 40
2 64731 1 40
2 64732 1 40
2 64733 1 40
2 64734 1 40
2 64735 1 40
2 64736 1 40
2 64737 1 40
2 64738 1 40
2 64739 1 40
2 64740 1 40
2 64741 1 40
2 64742 1 40
2 64743 1 40
2 64744 1 40
2 64745 1 40
2 64746 1 40
2 64747 1 40
2 64748 1 40
2 64749 1 40
2 64750 1 40
2 64751 1 40
2 64752 1 40
2 64753 1 40
2 64754 1 40
2 64755 1 40
2 64756 1 40
2 64757 1 40
2 64758 1 40
2 64759 1 40
2 64760 1 41
2 64761 1 41
2 64762 1 41
2 64763 1 41
2 64764 1 41
2 64765 1 41
2 64766 1 41
2 64767 1 41
2 64768 1 41
2 64769 1 41
2 64770 1 41
2 64771 1 41
2 64772 1 41
2 64773 1 41
2 64774 1 41
2 64775 1 41
2 64776 1 41
2 64777 1 41
2 64778 1 41
2 64779 1 41
2 64780 1 41
2 64781 1 41
2 64782 1 41
2 64783 1 41
2 64784 1 41
2 64785 1 41
2 64786 1 41
2 64787 1 41
2 64788 1 41
2 64789 1 41
2 64790 1 41
2 64791 1 41
2 64792 1 41
2 64793 1 41
2 64794 1 41
2 64795 1 41
2 64796 1 41
2 64797 1 41
2 64798 1 41
2 64799 1 41
2 64800 1 41
2 64801 1 41
2 64802 1 41
2 64803 1 41
2 64804 1 41
2 64805 1 41
2 64806 1 41
2 64807 1 41
2 64808 1 41
2 64809 1 41
2 64810 1 41
2 64811 1 41
2 64812 1 41
2 64813 1 41
2 64814 1 41
2 64815 1 41
2 64816 1 41
2 64817 1 41
2 64818 1 41
2 64819 1 41
2 64820 1 41
2 64821 1 41
2 64822 1 41
2 64823 1 41
2 64824 1 41
2 64825 1 41
2 64826 1 41
2 64827 1 41
2 64828 1 41
2 64829 1 41
2 64830 1 41
2 64831 1 41
2 64832 1 41
2 64833 1 41
2 64834 1 41
2 64835 1 41
2 64836 1 41
2 64837 1 41
2 64838 1 41
2 64839 1 41
2 64840 1 41
2 64841 1 41
2 64842 1 41
2 64843 1 41
2 64844 1 41
2 64845 1 41
2 64846 1 42
2 64847 1 42
2 64848 1 42
2 64849 1 42
2 64850 1 42
2 64851 1 42
2 64852 1 42
2 64853 1 42
2 64854 1 42
2 64855 1 42
2 64856 1 42
2 64857 1 42
2 64858 1 42
2 64859 1 42
2 64860 1 42
2 64861 1 42
2 64862 1 42
2 64863 1 42
2 64864 1 42
2 64865 1 42
2 64866 1 42
2 64867 1 42
2 64868 1 42
2 64869 1 42
2 64870 1 42
2 64871 1 42
2 64872 1 42
2 64873 1 42
2 64874 1 42
2 64875 1 42
2 64876 1 42
2 64877 1 42
2 64878 1 42
2 64879 1 42
2 64880 1 42
2 64881 1 42
2 64882 1 42
2 64883 1 42
2 64884 1 42
2 64885 1 42
2 64886 1 42
2 64887 1 42
2 64888 1 42
2 64889 1 42
2 64890 1 42
2 64891 1 42
2 64892 1 42
2 64893 1 42
2 64894 1 42
2 64895 1 42
2 64896 1 42
2 64897 1 42
2 64898 1 42
2 64899 1 42
2 64900 1 42
2 64901 1 42
2 64902 1 42
2 64903 1 42
2 64904 1 42
2 64905 1 42
2 64906 1 43
2 64907 1 43
2 64908 1 43
2 64909 1 43
2 64910 1 43
2 64911 1 43
2 64912 1 43
2 64913 1 43
2 64914 1 43
2 64915 1 43
2 64916 1 43
2 64917 1 43
2 64918 1 43
2 64919 1 43
2 64920 1 43
2 64921 1 43
2 64922 1 43
2 64923 1 43
2 64924 1 43
2 64925 1 43
2 64926 1 43
2 64927 1 43
2 64928 1 43
2 64929 1 43
2 64930 1 43
2 64931 1 43
2 64932 1 43
2 64933 1 43
2 64934 1 43
2 64935 1 43
2 64936 1 43
2 64937 1 43
2 64938 1 43
2 64939 1 43
2 64940 1 43
2 64941 1 43
2 64942 1 43
2 64943 1 43
2 64944 1 43
2 64945 1 43
2 64946 1 43
2 64947 1 43
2 64948 1 43
2 64949 1 43
2 64950 1 43
2 64951 1 43
2 64952 1 43
2 64953 1 43
2 64954 1 43
2 64955 1 43
2 64956 1 43
2 64957 1 43
2 64958 1 43
2 64959 1 43
2 64960 1 43
2 64961 1 43
2 64962 1 43
2 64963 1 43
2 64964 1 43
2 64965 1 43
2 64966 1 43
2 64967 1 43
2 64968 1 43
2 64969 1 43
2 64970 1 43
2 64971 1 43
2 64972 1 43
2 64973 1 43
2 64974 1 43
2 64975 1 43
2 64976 1 43
2 64977 1 43
2 64978 1 43
2 64979 1 43
2 64980 1 43
2 64981 1 43
2 64982 1 43
2 64983 1 43
2 64984 1 43
2 64985 1 43
2 64986 1 43
2 64987 1 43
2 64988 1 43
2 64989 1 43
2 64990 1 43
2 64991 1 43
2 64992 1 43
2 64993 1 43
2 64994 1 43
2 64995 1 43
2 64996 1 43
2 64997 1 43
2 64998 1 43
2 64999 1 43
2 65000 1 43
2 65001 1 43
2 65002 1 43
2 65003 1 43
2 65004 1 43
2 65005 1 43
2 65006 1 43
2 65007 1 43
2 65008 1 43
2 65009 1 43
2 65010 1 43
2 65011 1 43
2 65012 1 43
2 65013 1 43
2 65014 1 43
2 65015 1 43
2 65016 1 43
2 65017 1 43
2 65018 1 43
2 65019 1 43
2 65020 1 43
2 65021 1 43
2 65022 1 43
2 65023 1 43
2 65024 1 43
2 65025 1 43
2 65026 1 43
2 65027 1 43
2 65028 1 43
2 65029 1 43
2 65030 1 43
2 65031 1 43
2 65032 1 43
2 65033 1 43
2 65034 1 43
2 65035 1 43
2 65036 1 43
2 65037 1 43
2 65038 1 43
2 65039 1 43
2 65040 1 43
2 65041 1 43
2 65042 1 43
2 65043 1 43
2 65044 1 43
2 65045 1 43
2 65046 1 43
2 65047 1 43
2 65048 1 43
2 65049 1 43
2 65050 1 43
2 65051 1 43
2 65052 1 43
2 65053 1 43
2 65054 1 43
2 65055 1 43
2 65056 1 43
2 65057 1 43
2 65058 1 43
2 65059 1 43
2 65060 1 43
2 65061 1 43
2 65062 1 43
2 65063 1 43
2 65064 1 43
2 65065 1 43
2 65066 1 43
2 65067 1 43
2 65068 1 43
2 65069 1 43
2 65070 1 43
2 65071 1 43
2 65072 1 43
2 65073 1 43
2 65074 1 43
2 65075 1 43
2 65076 1 43
2 65077 1 43
2 65078 1 43
2 65079 1 43
2 65080 1 43
2 65081 1 43
2 65082 1 43
2 65083 1 43
2 65084 1 43
2 65085 1 43
2 65086 1 43
2 65087 1 43
2 65088 1 43
2 65089 1 43
2 65090 1 43
2 65091 1 43
2 65092 1 43
2 65093 1 43
2 65094 1 43
2 65095 1 43
2 65096 1 43
2 65097 1 43
2 65098 1 43
2 65099 1 43
2 65100 1 43
2 65101 1 43
2 65102 1 43
2 65103 1 43
2 65104 1 43
2 65105 1 43
2 65106 1 44
2 65107 1 44
2 65108 1 44
2 65109 1 44
2 65110 1 44
2 65111 1 44
2 65112 1 44
2 65113 1 44
2 65114 1 44
2 65115 1 44
2 65116 1 44
2 65117 1 44
2 65118 1 44
2 65119 1 44
2 65120 1 44
2 65121 1 44
2 65122 1 44
2 65123 1 44
2 65124 1 44
2 65125 1 44
2 65126 1 44
2 65127 1 44
2 65128 1 44
2 65129 1 44
2 65130 1 44
2 65131 1 44
2 65132 1 44
2 65133 1 44
2 65134 1 44
2 65135 1 44
2 65136 1 44
2 65137 1 44
2 65138 1 44
2 65139 1 44
2 65140 1 44
2 65141 1 44
2 65142 1 44
2 65143 1 44
2 65144 1 44
2 65145 1 44
2 65146 1 44
2 65147 1 44
2 65148 1 44
2 65149 1 44
2 65150 1 44
2 65151 1 44
2 65152 1 44
2 65153 1 44
2 65154 1 44
2 65155 1 44
2 65156 1 44
2 65157 1 44
2 65158 1 44
2 65159 1 44
2 65160 1 44
2 65161 1 44
2 65162 1 44
2 65163 1 44
2 65164 1 44
2 65165 1 44
2 65166 1 44
2 65167 1 44
2 65168 1 44
2 65169 1 44
2 65170 1 44
2 65171 1 44
2 65172 1 44
2 65173 1 44
2 65174 1 44
2 65175 1 44
2 65176 1 44
2 65177 1 44
2 65178 1 44
2 65179 1 44
2 65180 1 44
2 65181 1 44
2 65182 1 44
2 65183 1 44
2 65184 1 44
2 65185 1 44
2 65186 1 44
2 65187 1 44
2 65188 1 44
2 65189 1 44
2 65190 1 44
2 65191 1 44
2 65192 1 44
2 65193 1 44
2 65194 1 44
2 65195 1 44
2 65196 1 44
2 65197 1 44
2 65198 1 44
2 65199 1 44
2 65200 1 44
2 65201 1 44
2 65202 1 44
2 65203 1 44
2 65204 1 44
2 65205 1 44
2 65206 1 44
2 65207 1 44
2 65208 1 44
2 65209 1 44
2 65210 1 44
2 65211 1 44
2 65212 1 44
2 65213 1 44
2 65214 1 44
2 65215 1 44
2 65216 1 44
2 65217 1 44
2 65218 1 44
2 65219 1 44
2 65220 1 44
2 65221 1 44
2 65222 1 44
2 65223 1 44
2 65224 1 44
2 65225 1 44
2 65226 1 44
2 65227 1 44
2 65228 1 44
2 65229 1 44
2 65230 1 44
2 65231 1 44
2 65232 1 44
2 65233 1 44
2 65234 1 44
2 65235 1 44
2 65236 1 44
2 65237 1 44
2 65238 1 44
2 65239 1 44
2 65240 1 44
2 65241 1 44
2 65242 1 44
2 65243 1 44
2 65244 1 44
2 65245 1 44
2 65246 1 44
2 65247 1 44
2 65248 1 44
2 65249 1 44
2 65250 1 44
2 65251 1 44
2 65252 1 44
2 65253 1 44
2 65254 1 44
2 65255 1 44
2 65256 1 44
2 65257 1 44
2 65258 1 44
2 65259 1 44
2 65260 1 44
2 65261 1 44
2 65262 1 44
2 65263 1 44
2 65264 1 44
2 65265 1 44
2 65266 1 44
2 65267 1 44
2 65268 1 44
2 65269 1 44
2 65270 1 44
2 65271 1 44
2 65272 1 44
2 65273 1 44
2 65274 1 44
2 65275 1 44
2 65276 1 44
2 65277 1 44
2 65278 1 44
2 65279 1 44
2 65280 1 44
2 65281 1 44
2 65282 1 44
2 65283 1 44
2 65284 1 44
2 65285 1 44
2 65286 1 44
2 65287 1 44
2 65288 1 44
2 65289 1 44
2 65290 1 44
2 65291 1 44
2 65292 1 44
2 65293 1 44
2 65294 1 44
2 65295 1 44
2 65296 1 44
2 65297 1 44
2 65298 1 44
2 65299 1 44
2 65300 1 44
2 65301 1 44
2 65302 1 44
2 65303 1 44
2 65304 1 44
2 65305 1 44
2 65306 1 44
2 65307 1 44
2 65308 1 44
2 65309 1 44
2 65310 1 44
2 65311 1 44
2 65312 1 44
2 65313 1 44
2 65314 1 44
2 65315 1 44
2 65316 1 44
2 65317 1 44
2 65318 1 44
2 65319 1 44
2 65320 1 44
2 65321 1 44
2 65322 1 44
2 65323 1 44
2 65324 1 44
2 65325 1 44
2 65326 1 44
2 65327 1 44
2 65328 1 44
2 65329 1 44
2 65330 1 44
2 65331 1 44
2 65332 1 44
2 65333 1 44
2 65334 1 44
2 65335 1 44
2 65336 1 44
2 65337 1 44
2 65338 1 44
2 65339 1 44
2 65340 1 44
2 65341 1 44
2 65342 1 44
2 65343 1 44
2 65344 1 44
2 65345 1 44
2 65346 1 44
2 65347 1 44
2 65348 1 44
2 65349 1 44
2 65350 1 44
2 65351 1 44
2 65352 1 44
2 65353 1 44
2 65354 1 44
2 65355 1 44
2 65356 1 44
2 65357 1 44
2 65358 1 44
2 65359 1 44
2 65360 1 44
2 65361 1 44
2 65362 1 44
2 65363 1 45
2 65364 1 45
2 65365 1 45
2 65366 1 45
2 65367 1 45
2 65368 1 45
2 65369 1 45
2 65370 1 45
2 65371 1 45
2 65372 1 45
2 65373 1 45
2 65374 1 45
2 65375 1 45
2 65376 1 45
2 65377 1 45
2 65378 1 45
2 65379 1 45
2 65380 1 45
2 65381 1 45
2 65382 1 45
2 65383 1 45
2 65384 1 45
2 65385 1 45
2 65386 1 45
2 65387 1 45
2 65388 1 45
2 65389 1 45
2 65390 1 45
2 65391 1 45
2 65392 1 45
2 65393 1 45
2 65394 1 45
2 65395 1 45
2 65396 1 45
2 65397 1 45
2 65398 1 45
2 65399 1 45
2 65400 1 45
2 65401 1 45
2 65402 1 45
2 65403 1 45
2 65404 1 45
2 65405 1 45
2 65406 1 45
2 65407 1 45
2 65408 1 45
2 65409 1 45
2 65410 1 45
2 65411 1 45
2 65412 1 45
2 65413 1 45
2 65414 1 45
2 65415 1 45
2 65416 1 45
2 65417 1 45
2 65418 1 45
2 65419 1 45
2 65420 1 45
2 65421 1 45
2 65422 1 45
2 65423 1 45
2 65424 1 45
2 65425 1 45
2 65426 1 45
2 65427 1 45
2 65428 1 45
2 65429 1 45
2 65430 1 45
2 65431 1 45
2 65432 1 45
2 65433 1 45
2 65434 1 45
2 65435 1 45
2 65436 1 45
2 65437 1 45
2 65438 1 45
2 65439 1 45
2 65440 1 45
2 65441 1 45
2 65442 1 45
2 65443 1 45
2 65444 1 45
2 65445 1 45
2 65446 1 45
2 65447 1 45
2 65448 1 45
2 65449 1 45
2 65450 1 45
2 65451 1 45
2 65452 1 45
2 65453 1 45
2 65454 1 45
2 65455 1 45
2 65456 1 45
2 65457 1 45
2 65458 1 45
2 65459 1 45
2 65460 1 45
2 65461 1 45
2 65462 1 45
2 65463 1 45
2 65464 1 45
2 65465 1 45
2 65466 1 45
2 65467 1 45
2 65468 1 45
2 65469 1 45
2 65470 1 45
2 65471 1 45
2 65472 1 45
2 65473 1 45
2 65474 1 45
2 65475 1 45
2 65476 1 45
2 65477 1 45
2 65478 1 45
2 65479 1 45
2 65480 1 45
2 65481 1 45
2 65482 1 45
2 65483 1 45
2 65484 1 45
2 65485 1 45
2 65486 1 45
2 65487 1 45
2 65488 1 45
2 65489 1 45
2 65490 1 45
2 65491 1 45
2 65492 1 45
2 65493 1 45
2 65494 1 45
2 65495 1 45
2 65496 1 45
2 65497 1 45
2 65498 1 45
2 65499 1 45
2 65500 1 45
2 65501 1 45
2 65502 1 45
2 65503 1 45
2 65504 1 45
2 65505 1 45
2 65506 1 45
2 65507 1 45
2 65508 1 45
2 65509 1 45
2 65510 1 45
2 65511 1 45
2 65512 1 45
2 65513 1 45
2 65514 1 45
2 65515 1 45
2 65516 1 45
2 65517 1 45
2 65518 1 45
2 65519 1 45
2 65520 1 45
2 65521 1 45
2 65522 1 45
2 65523 1 45
2 65524 1 45
2 65525 1 45
2 65526 1 45
2 65527 1 45
2 65528 1 45
2 65529 1 45
2 65530 1 45
2 65531 1 45
2 65532 1 45
2 65533 1 45
2 65534 1 45
2 65535 1 45
2 65536 1 45
2 65537 1 45
2 65538 1 45
2 65539 1 45
2 65540 1 45
2 65541 1 45
2 65542 1 45
2 65543 1 45
2 65544 1 45
2 65545 1 45
2 65546 1 45
2 65547 1 45
2 65548 1 45
2 65549 1 45
2 65550 1 45
2 65551 1 45
2 65552 1 45
2 65553 1 45
2 65554 1 45
2 65555 1 45
2 65556 1 45
2 65557 1 45
2 65558 1 45
2 65559 1 45
2 65560 1 45
2 65561 1 45
2 65562 1 45
2 65563 1 45
2 65564 1 45
2 65565 1 45
2 65566 1 45
2 65567 1 45
2 65568 1 45
2 65569 1 45
2 65570 1 45
2 65571 1 45
2 65572 1 45
2 65573 1 45
2 65574 1 45
2 65575 1 45
2 65576 1 45
2 65577 1 45
2 65578 1 45
2 65579 1 45
2 65580 1 45
2 65581 1 45
2 65582 1 45
2 65583 1 45
2 65584 1 45
2 65585 1 45
2 65586 1 45
2 65587 1 45
2 65588 1 45
2 65589 1 45
2 65590 1 45
2 65591 1 45
2 65592 1 45
2 65593 1 45
2 65594 1 45
2 65595 1 45
2 65596 1 45
2 65597 1 45
2 65598 1 45
2 65599 1 45
2 65600 1 45
2 65601 1 45
2 65602 1 45
2 65603 1 45
2 65604 1 45
2 65605 1 45
2 65606 1 45
2 65607 1 45
2 65608 1 45
2 65609 1 45
2 65610 1 45
2 65611 1 45
2 65612 1 45
2 65613 1 45
2 65614 1 45
2 65615 1 45
2 65616 1 45
2 65617 1 45
2 65618 1 45
2 65619 1 45
2 65620 1 45
2 65621 1 45
2 65622 1 45
2 65623 1 45
2 65624 1 45
2 65625 1 45
2 65626 1 45
2 65627 1 45
2 65628 1 45
2 65629 1 45
2 65630 1 45
2 65631 1 45
2 65632 1 45
2 65633 1 45
2 65634 1 45
2 65635 1 45
2 65636 1 45
2 65637 1 45
2 65638 1 45
2 65639 1 45
2 65640 1 45
2 65641 1 45
2 65642 1 45
2 65643 1 45
2 65644 1 45
2 65645 1 45
2 65646 1 45
2 65647 1 45
2 65648 1 45
2 65649 1 45
2 65650 1 45
2 65651 1 45
2 65652 1 45
2 65653 1 45
2 65654 1 45
2 65655 1 45
2 65656 1 45
2 65657 1 45
2 65658 1 45
2 65659 1 45
2 65660 1 45
2 65661 1 45
2 65662 1 45
2 65663 1 45
2 65664 1 45
2 65665 1 45
2 65666 1 45
2 65667 1 45
2 65668 1 45
2 65669 1 45
2 65670 1 45
2 65671 1 45
2 65672 1 45
2 65673 1 45
2 65674 1 45
2 65675 1 45
2 65676 1 45
2 65677 1 45
2 65678 1 45
2 65679 1 45
2 65680 1 45
2 65681 1 45
2 65682 1 45
2 65683 1 45
2 65684 1 45
2 65685 1 45
2 65686 1 45
2 65687 1 45
2 65688 1 45
2 65689 1 45
2 65690 1 45
2 65691 1 45
2 65692 1 45
2 65693 1 45
2 65694 1 45
2 65695 1 45
2 65696 1 45
2 65697 1 45
2 65698 1 45
2 65699 1 45
2 65700 1 45
2 65701 1 45
2 65702 1 45
2 65703 1 45
2 65704 1 45
2 65705 1 45
2 65706 1 45
2 65707 1 45
2 65708 1 45
2 65709 1 45
2 65710 1 45
2 65711 1 45
2 65712 1 45
2 65713 1 45
2 65714 1 45
2 65715 1 45
2 65716 1 45
2 65717 1 45
2 65718 1 45
2 65719 1 45
2 65720 1 45
2 65721 1 45
2 65722 1 45
2 65723 1 45
2 65724 1 45
2 65725 1 45
2 65726 1 45
2 65727 1 45
2 65728 1 45
2 65729 1 45
2 65730 1 45
2 65731 1 45
2 65732 1 45
2 65733 1 45
2 65734 1 45
2 65735 1 45
2 65736 1 45
2 65737 1 45
2 65738 1 45
2 65739 1 45
2 65740 1 45
2 65741 1 45
2 65742 1 45
2 65743 1 45
2 65744 1 45
2 65745 1 45
2 65746 1 45
2 65747 1 45
2 65748 1 45
2 65749 1 45
2 65750 1 45
2 65751 1 45
2 65752 1 45
2 65753 1 45
2 65754 1 45
2 65755 1 45
2 65756 1 45
2 65757 1 45
2 65758 1 45
2 65759 1 45
2 65760 1 46
2 65761 1 46
2 65762 1 46
2 65763 1 46
2 65764 1 46
2 65765 1 46
2 65766 1 46
2 65767 1 46
2 65768 1 46
2 65769 1 46
2 65770 1 46
2 65771 1 46
2 65772 1 46
2 65773 1 46
2 65774 1 46
2 65775 1 46
2 65776 1 46
2 65777 1 46
2 65778 1 46
2 65779 1 46
2 65780 1 46
2 65781 1 46
2 65782 1 46
2 65783 1 46
2 65784 1 46
2 65785 1 46
2 65786 1 46
2 65787 1 46
2 65788 1 46
2 65789 1 46
2 65790 1 46
2 65791 1 46
2 65792 1 46
2 65793 1 46
2 65794 1 46
2 65795 1 46
2 65796 1 46
2 65797 1 46
2 65798 1 46
2 65799 1 46
2 65800 1 46
2 65801 1 46
2 65802 1 46
2 65803 1 46
2 65804 1 46
2 65805 1 46
2 65806 1 46
2 65807 1 46
2 65808 1 46
2 65809 1 46
2 65810 1 46
2 65811 1 46
2 65812 1 46
2 65813 1 46
2 65814 1 46
2 65815 1 46
2 65816 1 46
2 65817 1 46
2 65818 1 46
2 65819 1 46
2 65820 1 46
2 65821 1 46
2 65822 1 46
2 65823 1 46
2 65824 1 46
2 65825 1 46
2 65826 1 46
2 65827 1 46
2 65828 1 46
2 65829 1 46
2 65830 1 46
2 65831 1 46
2 65832 1 46
2 65833 1 46
2 65834 1 46
2 65835 1 46
2 65836 1 46
2 65837 1 46
2 65838 1 46
2 65839 1 46
2 65840 1 46
2 65841 1 46
2 65842 1 46
2 65843 1 46
2 65844 1 46
2 65845 1 46
2 65846 1 46
2 65847 1 46
2 65848 1 46
2 65849 1 46
2 65850 1 46
2 65851 1 46
2 65852 1 46
2 65853 1 46
2 65854 1 46
2 65855 1 46
2 65856 1 46
2 65857 1 46
2 65858 1 46
2 65859 1 46
2 65860 1 46
2 65861 1 46
2 65862 1 46
2 65863 1 46
2 65864 1 46
2 65865 1 46
2 65866 1 46
2 65867 1 46
2 65868 1 46
2 65869 1 46
2 65870 1 46
2 65871 1 46
2 65872 1 46
2 65873 1 46
2 65874 1 46
2 65875 1 46
2 65876 1 46
2 65877 1 46
2 65878 1 46
2 65879 1 46
2 65880 1 46
2 65881 1 46
2 65882 1 46
2 65883 1 46
2 65884 1 46
2 65885 1 46
2 65886 1 46
2 65887 1 46
2 65888 1 46
2 65889 1 46
2 65890 1 46
2 65891 1 46
2 65892 1 46
2 65893 1 46
2 65894 1 46
2 65895 1 46
2 65896 1 46
2 65897 1 46
2 65898 1 46
2 65899 1 46
2 65900 1 46
2 65901 1 46
2 65902 1 46
2 65903 1 46
2 65904 1 46
2 65905 1 46
2 65906 1 46
2 65907 1 46
2 65908 1 46
2 65909 1 46
2 65910 1 46
2 65911 1 46
2 65912 1 46
2 65913 1 46
2 65914 1 46
2 65915 1 46
2 65916 1 46
2 65917 1 46
2 65918 1 46
2 65919 1 46
2 65920 1 46
2 65921 1 46
2 65922 1 46
2 65923 1 46
2 65924 1 46
2 65925 1 46
2 65926 1 46
2 65927 1 46
2 65928 1 46
2 65929 1 46
2 65930 1 46
2 65931 1 46
2 65932 1 46
2 65933 1 46
2 65934 1 46
2 65935 1 46
2 65936 1 46
2 65937 1 46
2 65938 1 46
2 65939 1 46
2 65940 1 46
2 65941 1 46
2 65942 1 46
2 65943 1 46
2 65944 1 46
2 65945 1 46
2 65946 1 46
2 65947 1 46
2 65948 1 46
2 65949 1 46
2 65950 1 46
2 65951 1 46
2 65952 1 46
2 65953 1 46
2 65954 1 46
2 65955 1 46
2 65956 1 46
2 65957 1 46
2 65958 1 46
2 65959 1 46
2 65960 1 46
2 65961 1 46
2 65962 1 46
2 65963 1 46
2 65964 1 46
2 65965 1 46
2 65966 1 46
2 65967 1 46
2 65968 1 46
2 65969 1 46
2 65970 1 46
2 65971 1 46
2 65972 1 46
2 65973 1 46
2 65974 1 46
2 65975 1 46
2 65976 1 46
2 65977 1 46
2 65978 1 46
2 65979 1 46
2 65980 1 46
2 65981 1 46
2 65982 1 46
2 65983 1 46
2 65984 1 46
2 65985 1 46
2 65986 1 46
2 65987 1 46
2 65988 1 46
2 65989 1 46
2 65990 1 46
2 65991 1 46
2 65992 1 46
2 65993 1 46
2 65994 1 46
2 65995 1 46
2 65996 1 46
2 65997 1 46
2 65998 1 46
2 65999 1 46
2 66000 1 46
2 66001 1 46
2 66002 1 46
2 66003 1 46
2 66004 1 46
2 66005 1 46
2 66006 1 46
2 66007 1 46
2 66008 1 46
2 66009 1 46
2 66010 1 46
2 66011 1 46
2 66012 1 46
2 66013 1 46
2 66014 1 46
2 66015 1 46
2 66016 1 46
2 66017 1 46
2 66018 1 46
2 66019 1 46
2 66020 1 46
2 66021 1 46
2 66022 1 46
2 66023 1 46
2 66024 1 46
2 66025 1 46
2 66026 1 46
2 66027 1 46
2 66028 1 46
2 66029 1 46
2 66030 1 46
2 66031 1 46
2 66032 1 46
2 66033 1 46
2 66034 1 46
2 66035 1 46
2 66036 1 46
2 66037 1 46
2 66038 1 46
2 66039 1 46
2 66040 1 46
2 66041 1 46
2 66042 1 46
2 66043 1 46
2 66044 1 46
2 66045 1 46
2 66046 1 46
2 66047 1 46
2 66048 1 46
2 66049 1 46
2 66050 1 46
2 66051 1 46
2 66052 1 46
2 66053 1 46
2 66054 1 46
2 66055 1 46
2 66056 1 46
2 66057 1 46
2 66058 1 46
2 66059 1 46
2 66060 1 46
2 66061 1 46
2 66062 1 46
2 66063 1 46
2 66064 1 46
2 66065 1 46
2 66066 1 46
2 66067 1 46
2 66068 1 46
2 66069 1 46
2 66070 1 46
2 66071 1 46
2 66072 1 46
2 66073 1 46
2 66074 1 46
2 66075 1 46
2 66076 1 46
2 66077 1 46
2 66078 1 46
2 66079 1 46
2 66080 1 46
2 66081 1 46
2 66082 1 46
2 66083 1 46
2 66084 1 46
2 66085 1 46
2 66086 1 46
2 66087 1 46
2 66088 1 46
2 66089 1 46
2 66090 1 46
2 66091 1 46
2 66092 1 46
2 66093 1 46
2 66094 1 46
2 66095 1 46
2 66096 1 46
2 66097 1 46
2 66098 1 46
2 66099 1 46
2 66100 1 46
2 66101 1 46
2 66102 1 46
2 66103 1 46
2 66104 1 46
2 66105 1 46
2 66106 1 46
2 66107 1 46
2 66108 1 46
2 66109 1 46
2 66110 1 47
2 66111 1 47
2 66112 1 47
2 66113 1 47
2 66114 1 47
2 66115 1 47
2 66116 1 47
2 66117 1 47
2 66118 1 47
2 66119 1 47
2 66120 1 47
2 66121 1 47
2 66122 1 47
2 66123 1 47
2 66124 1 47
2 66125 1 47
2 66126 1 47
2 66127 1 47
2 66128 1 47
2 66129 1 47
2 66130 1 47
2 66131 1 47
2 66132 1 47
2 66133 1 47
2 66134 1 47
2 66135 1 47
2 66136 1 47
2 66137 1 47
2 66138 1 47
2 66139 1 47
2 66140 1 47
2 66141 1 47
2 66142 1 47
2 66143 1 47
2 66144 1 47
2 66145 1 47
2 66146 1 47
2 66147 1 47
2 66148 1 47
2 66149 1 47
2 66150 1 47
2 66151 1 47
2 66152 1 47
2 66153 1 47
2 66154 1 47
2 66155 1 47
2 66156 1 47
2 66157 1 47
2 66158 1 47
2 66159 1 47
2 66160 1 47
2 66161 1 47
2 66162 1 47
2 66163 1 47
2 66164 1 47
2 66165 1 47
2 66166 1 47
2 66167 1 47
2 66168 1 47
2 66169 1 47
2 66170 1 47
2 66171 1 47
2 66172 1 47
2 66173 1 47
2 66174 1 47
2 66175 1 47
2 66176 1 47
2 66177 1 47
2 66178 1 47
2 66179 1 47
2 66180 1 47
2 66181 1 47
2 66182 1 47
2 66183 1 47
2 66184 1 47
2 66185 1 47
2 66186 1 47
2 66187 1 47
2 66188 1 47
2 66189 1 47
2 66190 1 47
2 66191 1 47
2 66192 1 47
2 66193 1 47
2 66194 1 47
2 66195 1 47
2 66196 1 47
2 66197 1 47
2 66198 1 47
2 66199 1 47
2 66200 1 47
2 66201 1 47
2 66202 1 47
2 66203 1 47
2 66204 1 47
2 66205 1 47
2 66206 1 47
2 66207 1 47
2 66208 1 47
2 66209 1 47
2 66210 1 47
2 66211 1 47
2 66212 1 47
2 66213 1 47
2 66214 1 47
2 66215 1 47
2 66216 1 47
2 66217 1 47
2 66218 1 47
2 66219 1 47
2 66220 1 47
2 66221 1 47
2 66222 1 47
2 66223 1 47
2 66224 1 47
2 66225 1 47
2 66226 1 47
2 66227 1 47
2 66228 1 47
2 66229 1 47
2 66230 1 47
2 66231 1 47
2 66232 1 47
2 66233 1 47
2 66234 1 47
2 66235 1 47
2 66236 1 47
2 66237 1 47
2 66238 1 47
2 66239 1 47
2 66240 1 47
2 66241 1 47
2 66242 1 47
2 66243 1 47
2 66244 1 47
2 66245 1 47
2 66246 1 47
2 66247 1 47
2 66248 1 47
2 66249 1 47
2 66250 1 47
2 66251 1 47
2 66252 1 47
2 66253 1 47
2 66254 1 47
2 66255 1 47
2 66256 1 47
2 66257 1 47
2 66258 1 47
2 66259 1 47
2 66260 1 47
2 66261 1 47
2 66262 1 47
2 66263 1 47
2 66264 1 47
2 66265 1 47
2 66266 1 47
2 66267 1 47
2 66268 1 47
2 66269 1 47
2 66270 1 47
2 66271 1 47
2 66272 1 47
2 66273 1 47
2 66274 1 47
2 66275 1 47
2 66276 1 47
2 66277 1 47
2 66278 1 47
2 66279 1 47
2 66280 1 47
2 66281 1 47
2 66282 1 47
2 66283 1 47
2 66284 1 47
2 66285 1 47
2 66286 1 47
2 66287 1 47
2 66288 1 47
2 66289 1 47
2 66290 1 47
2 66291 1 47
2 66292 1 47
2 66293 1 47
2 66294 1 47
2 66295 1 47
2 66296 1 47
2 66297 1 47
2 66298 1 47
2 66299 1 47
2 66300 1 47
2 66301 1 47
2 66302 1 47
2 66303 1 47
2 66304 1 47
2 66305 1 47
2 66306 1 47
2 66307 1 47
2 66308 1 47
2 66309 1 47
2 66310 1 47
2 66311 1 47
2 66312 1 47
2 66313 1 47
2 66314 1 47
2 66315 1 47
2 66316 1 47
2 66317 1 47
2 66318 1 47
2 66319 1 47
2 66320 1 47
2 66321 1 47
2 66322 1 47
2 66323 1 47
2 66324 1 47
2 66325 1 47
2 66326 1 47
2 66327 1 47
2 66328 1 47
2 66329 1 47
2 66330 1 47
2 66331 1 47
2 66332 1 47
2 66333 1 47
2 66334 1 47
2 66335 1 47
2 66336 1 47
2 66337 1 47
2 66338 1 47
2 66339 1 47
2 66340 1 47
2 66341 1 47
2 66342 1 47
2 66343 1 47
2 66344 1 47
2 66345 1 47
2 66346 1 47
2 66347 1 47
2 66348 1 47
2 66349 1 47
2 66350 1 47
2 66351 1 47
2 66352 1 47
2 66353 1 47
2 66354 1 47
2 66355 1 47
2 66356 1 47
2 66357 1 47
2 66358 1 47
2 66359 1 47
2 66360 1 47
2 66361 1 47
2 66362 1 47
2 66363 1 47
2 66364 1 47
2 66365 1 47
2 66366 1 47
2 66367 1 47
2 66368 1 47
2 66369 1 47
2 66370 1 47
2 66371 1 47
2 66372 1 47
2 66373 1 47
2 66374 1 47
2 66375 1 47
2 66376 1 47
2 66377 1 47
2 66378 1 47
2 66379 1 47
2 66380 1 47
2 66381 1 47
2 66382 1 47
2 66383 1 47
2 66384 1 47
2 66385 1 47
2 66386 1 47
2 66387 1 47
2 66388 1 47
2 66389 1 47
2 66390 1 47
2 66391 1 47
2 66392 1 47
2 66393 1 47
2 66394 1 47
2 66395 1 47
2 66396 1 47
2 66397 1 47
2 66398 1 47
2 66399 1 47
2 66400 1 47
2 66401 1 47
2 66402 1 47
2 66403 1 48
2 66404 1 48
2 66405 1 48
2 66406 1 48
2 66407 1 48
2 66408 1 48
2 66409 1 48
2 66410 1 48
2 66411 1 48
2 66412 1 48
2 66413 1 48
2 66414 1 48
2 66415 1 48
2 66416 1 48
2 66417 1 48
2 66418 1 48
2 66419 1 48
2 66420 1 48
2 66421 1 48
2 66422 1 48
2 66423 1 48
2 66424 1 48
2 66425 1 48
2 66426 1 48
2 66427 1 48
2 66428 1 48
2 66429 1 48
2 66430 1 48
2 66431 1 48
2 66432 1 48
2 66433 1 48
2 66434 1 48
2 66435 1 48
2 66436 1 48
2 66437 1 48
2 66438 1 48
2 66439 1 48
2 66440 1 48
2 66441 1 48
2 66442 1 48
2 66443 1 48
2 66444 1 48
2 66445 1 48
2 66446 1 48
2 66447 1 48
2 66448 1 48
2 66449 1 48
2 66450 1 48
2 66451 1 48
2 66452 1 48
2 66453 1 48
2 66454 1 48
2 66455 1 48
2 66456 1 48
2 66457 1 48
2 66458 1 48
2 66459 1 48
2 66460 1 48
2 66461 1 48
2 66462 1 48
2 66463 1 48
2 66464 1 48
2 66465 1 48
2 66466 1 48
2 66467 1 48
2 66468 1 48
2 66469 1 48
2 66470 1 48
2 66471 1 48
2 66472 1 48
2 66473 1 48
2 66474 1 48
2 66475 1 48
2 66476 1 48
2 66477 1 48
2 66478 1 48
2 66479 1 48
2 66480 1 48
2 66481 1 48
2 66482 1 48
2 66483 1 48
2 66484 1 48
2 66485 1 48
2 66486 1 48
2 66487 1 48
2 66488 1 48
2 66489 1 48
2 66490 1 48
2 66491 1 48
2 66492 1 48
2 66493 1 48
2 66494 1 48
2 66495 1 48
2 66496 1 48
2 66497 1 48
2 66498 1 48
2 66499 1 48
2 66500 1 48
2 66501 1 48
2 66502 1 48
2 66503 1 48
2 66504 1 48
2 66505 1 48
2 66506 1 48
2 66507 1 48
2 66508 1 48
2 66509 1 48
2 66510 1 48
2 66511 1 48
2 66512 1 48
2 66513 1 48
2 66514 1 48
2 66515 1 48
2 66516 1 48
2 66517 1 48
2 66518 1 48
2 66519 1 48
2 66520 1 48
2 66521 1 48
2 66522 1 48
2 66523 1 48
2 66524 1 48
2 66525 1 48
2 66526 1 48
2 66527 1 48
2 66528 1 48
2 66529 1 48
2 66530 1 48
2 66531 1 48
2 66532 1 48
2 66533 1 48
2 66534 1 48
2 66535 1 49
2 66536 1 49
2 66537 1 49
2 66538 1 49
2 66539 1 49
2 66540 1 49
2 66541 1 49
2 66542 1 49
2 66543 1 49
2 66544 1 49
2 66545 1 49
2 66546 1 49
2 66547 1 49
2 66548 1 49
2 66549 1 49
2 66550 1 49
2 66551 1 49
2 66552 1 49
2 66553 1 49
2 66554 1 49
2 66555 1 49
2 66556 1 49
2 66557 1 49
2 66558 1 49
2 66559 1 49
2 66560 1 49
2 66561 1 49
2 66562 1 49
2 66563 1 49
2 66564 1 49
2 66565 1 49
2 66566 1 49
2 66567 1 49
2 66568 1 49
2 66569 1 49
2 66570 1 49
2 66571 1 49
2 66572 1 49
2 66573 1 49
2 66574 1 49
2 66575 1 49
2 66576 1 49
2 66577 1 49
2 66578 1 49
2 66579 1 49
2 66580 1 49
2 66581 1 49
2 66582 1 49
2 66583 1 49
2 66584 1 49
2 66585 1 49
2 66586 1 49
2 66587 1 49
2 66588 1 49
2 66589 1 49
2 66590 1 49
2 66591 1 49
2 66592 1 49
2 66593 1 49
2 66594 1 49
2 66595 1 49
2 66596 1 49
2 66597 1 49
2 66598 1 49
2 66599 1 49
2 66600 1 49
2 66601 1 49
2 66602 1 49
2 66603 1 49
2 66604 1 49
2 66605 1 49
2 66606 1 49
2 66607 1 49
2 66608 1 49
2 66609 1 49
2 66610 1 49
2 66611 1 49
2 66612 1 49
2 66613 1 49
2 66614 1 49
2 66615 1 49
2 66616 1 49
2 66617 1 49
2 66618 1 49
2 66619 1 49
2 66620 1 49
2 66621 1 49
2 66622 1 49
2 66623 1 49
2 66624 1 49
2 66625 1 49
2 66626 1 49
2 66627 1 49
2 66628 1 49
2 66629 1 49
2 66630 1 49
2 66631 1 49
2 66632 1 49
2 66633 1 49
2 66634 1 49
2 66635 1 49
2 66636 1 49
2 66637 1 49
2 66638 1 49
2 66639 1 49
2 66640 1 49
2 66641 1 49
2 66642 1 49
2 66643 1 49
2 66644 1 49
2 66645 1 49
2 66646 1 49
2 66647 1 49
2 66648 1 49
2 66649 1 49
2 66650 1 49
2 66651 1 49
2 66652 1 49
2 66653 1 49
2 66654 1 50
2 66655 1 50
2 66656 1 50
2 66657 1 50
2 66658 1 50
2 66659 1 50
2 66660 1 50
2 66661 1 50
2 66662 1 50
2 66663 1 50
2 66664 1 50
2 66665 1 50
2 66666 1 50
2 66667 1 50
2 66668 1 50
2 66669 1 50
2 66670 1 50
2 66671 1 50
2 66672 1 50
2 66673 1 50
2 66674 1 50
2 66675 1 50
2 66676 1 50
2 66677 1 50
2 66678 1 50
2 66679 1 50
2 66680 1 50
2 66681 1 50
2 66682 1 50
2 66683 1 50
2 66684 1 50
2 66685 1 50
2 66686 1 50
2 66687 1 50
2 66688 1 50
2 66689 1 50
2 66690 1 50
2 66691 1 50
2 66692 1 50
2 66693 1 50
2 66694 1 50
2 66695 1 50
2 66696 1 50
2 66697 1 50
2 66698 1 50
2 66699 1 50
2 66700 1 50
2 66701 1 50
2 66702 1 50
2 66703 1 50
2 66704 1 50
2 66705 1 50
2 66706 1 50
2 66707 1 50
2 66708 1 50
2 66709 1 50
2 66710 1 50
2 66711 1 50
2 66712 1 50
2 66713 1 50
2 66714 1 50
2 66715 1 50
2 66716 1 50
2 66717 1 50
2 66718 1 50
2 66719 1 50
2 66720 1 50
2 66721 1 50
2 66722 1 50
2 66723 1 50
2 66724 1 50
2 66725 1 50
2 66726 1 50
2 66727 1 50
2 66728 1 50
2 66729 1 50
2 66730 1 50
2 66731 1 50
2 66732 1 50
2 66733 1 50
2 66734 1 50
2 66735 1 50
2 66736 1 50
2 66737 1 50
2 66738 1 52
2 66739 1 52
2 66740 1 52
2 66741 1 52
2 66742 1 52
2 66743 1 52
2 66744 1 52
2 66745 1 52
2 66746 1 52
2 66747 1 52
2 66748 1 52
2 66749 1 52
2 66750 1 52
2 66751 1 52
2 66752 1 52
2 66753 1 52
2 66754 1 52
2 66755 1 52
2 66756 1 52
2 66757 1 52
2 66758 1 52
2 66759 1 52
2 66760 1 52
2 66761 1 52
2 66762 1 52
2 66763 1 52
2 66764 1 52
2 66765 1 52
2 66766 1 52
2 66767 1 52
2 66768 1 52
2 66769 1 52
2 66770 1 52
2 66771 1 52
2 66772 1 52
2 66773 1 52
2 66774 1 52
2 66775 1 52
2 66776 1 52
2 66777 1 52
2 66778 1 52
2 66779 1 52
2 66780 1 52
2 66781 1 52
2 66782 1 52
2 66783 1 52
2 66784 1 52
2 66785 1 52
2 66786 1 52
2 66787 1 52
2 66788 1 52
2 66789 1 52
2 66790 1 52
2 66791 1 52
2 66792 1 52
2 66793 1 52
2 66794 1 52
2 66795 1 52
2 66796 1 52
2 66797 1 52
2 66798 1 53
2 66799 1 53
2 66800 1 53
2 66801 1 53
2 66802 1 53
2 66803 1 53
2 66804 1 53
2 66805 1 53
2 66806 1 54
2 66807 1 54
2 66808 1 54
2 66809 1 54
2 66810 1 54
2 66811 1 54
2 66812 1 54
2 66813 1 54
2 66814 1 54
2 66815 1 54
2 66816 1 54
2 66817 1 54
2 66818 1 54
2 66819 1 54
2 66820 1 54
2 66821 1 54
2 66822 1 54
2 66823 1 54
2 66824 1 54
2 66825 1 54
2 66826 1 54
2 66827 1 54
2 66828 1 54
2 66829 1 54
2 66830 1 54
2 66831 1 54
2 66832 1 54
2 66833 1 54
2 66834 1 54
2 66835 1 54
2 66836 1 54
2 66837 1 54
2 66838 1 54
2 66839 1 54
2 66840 1 54
2 66841 1 54
2 66842 1 54
2 66843 1 54
2 66844 1 54
2 66845 1 54
2 66846 1 54
2 66847 1 54
2 66848 1 54
2 66849 1 54
2 66850 1 54
2 66851 1 54
2 66852 1 54
2 66853 1 54
2 66854 1 54
2 66855 1 54
2 66856 1 54
2 66857 1 54
2 66858 1 54
2 66859 1 54
2 66860 1 54
2 66861 1 54
2 66862 1 54
2 66863 1 54
2 66864 1 54
2 66865 1 54
2 66866 1 54
2 66867 1 54
2 66868 1 54
2 66869 1 54
2 66870 1 54
2 66871 1 54
2 66872 1 54
2 66873 1 54
2 66874 1 54
2 66875 1 54
2 66876 1 54
2 66877 1 54
2 66878 1 54
2 66879 1 55
2 66880 1 55
2 66881 1 55
2 66882 1 56
2 66883 1 56
2 66884 1 56
2 66885 1 56
2 66886 1 56
2 66887 1 56
2 66888 1 56
2 66889 1 56
2 66890 1 56
2 66891 1 56
2 66892 1 56
2 66893 1 56
2 66894 1 56
2 66895 1 56
2 66896 1 56
2 66897 1 56
2 66898 1 56
2 66899 1 56
2 66900 1 56
2 66901 1 56
2 66902 1 56
2 66903 1 56
2 66904 1 56
2 66905 1 56
2 66906 1 56
2 66907 1 56
2 66908 1 56
2 66909 1 56
2 66910 1 56
2 66911 1 56
2 66912 1 56
2 66913 1 56
2 66914 1 56
2 66915 1 56
2 66916 1 56
2 66917 1 56
2 66918 1 56
2 66919 1 56
2 66920 1 56
2 66921 1 56
2 66922 1 56
2 66923 1 56
2 66924 1 56
2 66925 1 56
2 66926 1 56
2 66927 1 56
2 66928 1 56
2 66929 1 56
2 66930 1 56
2 66931 1 56
2 66932 1 56
2 66933 1 56
2 66934 1 56
2 66935 1 56
2 66936 1 56
2 66937 1 56
2 66938 1 56
2 66939 1 56
2 66940 1 56
2 66941 1 56
2 66942 1 56
2 66943 1 56
2 66944 1 56
2 66945 1 56
2 66946 1 56
2 66947 1 56
2 66948 1 56
2 66949 1 56
2 66950 1 56
2 66951 1 56
2 66952 1 57
2 66953 1 57
2 66954 1 58
2 66955 1 58
2 66956 1 58
2 66957 1 58
2 66958 1 58
2 66959 1 58
2 66960 1 58
2 66961 1 58
2 66962 1 58
2 66963 1 58
2 66964 1 58
2 66965 1 58
2 66966 1 58
2 66967 1 58
2 66968 1 58
2 66969 1 58
2 66970 1 58
2 66971 1 58
2 66972 1 58
2 66973 1 58
2 66974 1 58
2 66975 1 58
2 66976 1 58
2 66977 1 58
2 66978 1 58
2 66979 1 58
2 66980 1 58
2 66981 1 58
2 66982 1 58
2 66983 1 58
2 66984 1 58
2 66985 1 58
2 66986 1 58
2 66987 1 58
2 66988 1 58
2 66989 1 58
2 66990 1 58
2 66991 1 58
2 66992 1 58
2 66993 1 58
2 66994 1 58
2 66995 1 58
2 66996 1 58
2 66997 1 58
2 66998 1 58
2 66999 1 58
2 67000 1 58
2 67001 1 60
2 67002 1 60
2 67003 1 60
2 67004 1 60
2 67005 1 60
2 67006 1 60
2 67007 1 60
2 67008 1 60
2 67009 1 60
2 67010 1 60
2 67011 1 60
2 67012 1 60
2 67013 1 60
2 67014 1 60
2 67015 1 60
2 67016 1 61
2 67017 1 61
2 67018 1 61
2 67019 1 61
2 67020 1 61
2 67021 1 61
2 67022 1 61
2 67023 1 61
2 67024 1 61
2 67025 1 61
2 67026 1 61
2 67027 1 63
2 67028 1 63
2 67029 1 63
2 67030 1 66
2 67031 1 66
2 67032 1 66
2 67033 1 66
2 67034 1 66
2 67035 1 66
2 67036 1 66
2 67037 1 66
2 67038 1 66
2 67039 1 66
2 67040 1 66
2 67041 1 66
2 67042 1 66
2 67043 1 66
2 67044 1 66
2 67045 1 66
2 67046 1 66
2 67047 1 66
2 67048 1 66
2 67049 1 66
2 67050 1 66
2 67051 1 66
2 67052 1 66
2 67053 1 66
2 67054 1 66
2 67055 1 66
2 67056 1 66
2 67057 1 66
2 67058 1 66
2 67059 1 66
2 67060 1 66
2 67061 1 66
2 67062 1 66
2 67063 1 66
2 67064 1 66
2 67065 1 66
2 67066 1 66
2 67067 1 66
2 67068 1 66
2 67069 1 66
2 67070 1 66
2 67071 1 66
2 67072 1 66
2 67073 1 66
2 67074 1 66
2 67075 1 66
2 67076 1 66
2 67077 1 66
2 67078 1 66
2 67079 1 66
2 67080 1 66
2 67081 1 67
2 67082 1 67
2 67083 1 67
2 67084 1 67
2 67085 1 67
2 67086 1 67
2 67087 1 67
2 67088 1 67
2 67089 1 69
2 67090 1 69
2 67091 1 69
2 67092 1 74
2 67093 1 74
2 67094 1 74
2 67095 1 74
2 67096 1 74
2 67097 1 74
2 67098 1 74
2 67099 1 74
2 67100 1 74
2 67101 1 75
2 67102 1 75
2 67103 1 75
2 67104 1 75
2 67105 1 76
2 67106 1 76
2 67107 1 76
2 67108 1 76
2 67109 1 76
2 67110 1 76
2 67111 1 77
2 67112 1 77
2 67113 1 77
2 67114 1 77
2 67115 1 77
2 67116 1 80
2 67117 1 80
2 67118 1 80
2 67119 1 80
2 67120 1 80
2 67121 1 80
2 67122 1 80
2 67123 1 81
2 67124 1 81
2 67125 1 81
2 67126 1 90
2 67127 1 90
2 67128 1 90
2 67129 1 90
2 67130 1 90
2 67131 1 90
2 67132 1 90
2 67133 1 90
2 67134 1 90
2 67135 1 90
2 67136 1 90
2 67137 1 90
2 67138 1 90
2 67139 1 90
2 67140 1 90
2 67141 1 90
2 67142 1 90
2 67143 1 90
2 67144 1 90
2 67145 1 90
2 67146 1 90
2 67147 1 90
2 67148 1 90
2 67149 1 90
2 67150 1 90
2 67151 1 90
2 67152 1 90
2 67153 1 90
2 67154 1 90
2 67155 1 90
2 67156 1 90
2 67157 1 90
2 67158 1 90
2 67159 1 90
2 67160 1 90
2 67161 1 90
2 67162 1 90
2 67163 1 90
2 67164 1 90
2 67165 1 90
2 67166 1 90
2 67167 1 90
2 67168 1 90
2 67169 1 90
2 67170 1 90
2 67171 1 90
2 67172 1 90
2 67173 1 90
2 67174 1 90
2 67175 1 90
2 67176 1 90
2 67177 1 90
2 67178 1 90
2 67179 1 90
2 67180 1 90
2 67181 1 90
2 67182 1 90
2 67183 1 90
2 67184 1 90
2 67185 1 90
2 67186 1 90
2 67187 1 90
2 67188 1 90
2 67189 1 90
2 67190 1 90
2 67191 1 90
2 67192 1 90
2 67193 1 90
2 67194 1 90
2 67195 1 90
2 67196 1 90
2 67197 1 90
2 67198 1 90
2 67199 1 90
2 67200 1 90
2 67201 1 90
2 67202 1 90
2 67203 1 90
2 67204 1 90
2 67205 1 90
2 67206 1 90
2 67207 1 90
2 67208 1 90
2 67209 1 90
2 67210 1 90
2 67211 1 90
2 67212 1 90
2 67213 1 90
2 67214 1 90
2 67215 1 90
2 67216 1 90
2 67217 1 90
2 67218 1 90
2 67219 1 90
2 67220 1 90
2 67221 1 90
2 67222 1 90
2 67223 1 90
2 67224 1 90
2 67225 1 90
2 67226 1 90
2 67227 1 90
2 67228 1 90
2 67229 1 90
2 67230 1 90
2 67231 1 90
2 67232 1 90
2 67233 1 90
2 67234 1 90
2 67235 1 90
2 67236 1 91
2 67237 1 91
2 67238 1 91
2 67239 1 91
2 67240 1 91
2 67241 1 91
2 67242 1 91
2 67243 1 91
2 67244 1 91
2 67245 1 91
2 67246 1 91
2 67247 1 91
2 67248 1 91
2 67249 1 91
2 67250 1 91
2 67251 1 91
2 67252 1 91
2 67253 1 91
2 67254 1 91
2 67255 1 91
2 67256 1 91
2 67257 1 91
2 67258 1 91
2 67259 1 91
2 67260 1 91
2 67261 1 91
2 67262 1 91
2 67263 1 91
2 67264 1 91
2 67265 1 91
2 67266 1 91
2 67267 1 91
2 67268 1 91
2 67269 1 91
2 67270 1 91
2 67271 1 91
2 67272 1 91
2 67273 1 91
2 67274 1 91
2 67275 1 91
2 67276 1 91
2 67277 1 91
2 67278 1 91
2 67279 1 91
2 67280 1 91
2 67281 1 91
2 67282 1 91
2 67283 1 91
2 67284 1 91
2 67285 1 91
2 67286 1 91
2 67287 1 91
2 67288 1 91
2 67289 1 91
2 67290 1 91
2 67291 1 91
2 67292 1 91
2 67293 1 91
2 67294 1 91
2 67295 1 91
2 67296 1 91
2 67297 1 91
2 67298 1 91
2 67299 1 91
2 67300 1 91
2 67301 1 91
2 67302 1 91
2 67303 1 91
2 67304 1 91
2 67305 1 91
2 67306 1 91
2 67307 1 91
2 67308 1 91
2 67309 1 91
2 67310 1 91
2 67311 1 91
2 67312 1 91
2 67313 1 91
2 67314 1 91
2 67315 1 91
2 67316 1 91
2 67317 1 91
2 67318 1 91
2 67319 1 91
2 67320 1 91
2 67321 1 91
2 67322 1 91
2 67323 1 91
2 67324 1 91
2 67325 1 91
2 67326 1 91
2 67327 1 91
2 67328 1 91
2 67329 1 91
2 67330 1 91
2 67331 1 91
2 67332 1 91
2 67333 1 91
2 67334 1 91
2 67335 1 91
2 67336 1 91
2 67337 1 91
2 67338 1 91
2 67339 1 91
2 67340 1 91
2 67341 1 91
2 67342 1 91
2 67343 1 91
2 67344 1 91
2 67345 1 91
2 67346 1 91
2 67347 1 91
2 67348 1 91
2 67349 1 91
2 67350 1 91
2 67351 1 91
2 67352 1 91
2 67353 1 91
2 67354 1 91
2 67355 1 91
2 67356 1 91
2 67357 1 91
2 67358 1 91
2 67359 1 91
2 67360 1 91
2 67361 1 91
2 67362 1 91
2 67363 1 91
2 67364 1 91
2 67365 1 91
2 67366 1 91
2 67367 1 91
2 67368 1 91
2 67369 1 91
2 67370 1 91
2 67371 1 91
2 67372 1 91
2 67373 1 91
2 67374 1 91
2 67375 1 91
2 67376 1 91
2 67377 1 91
2 67378 1 91
2 67379 1 91
2 67380 1 91
2 67381 1 91
2 67382 1 91
2 67383 1 91
2 67384 1 91
2 67385 1 91
2 67386 1 91
2 67387 1 91
2 67388 1 91
2 67389 1 91
2 67390 1 91
2 67391 1 91
2 67392 1 91
2 67393 1 91
2 67394 1 91
2 67395 1 91
2 67396 1 91
2 67397 1 91
2 67398 1 91
2 67399 1 91
2 67400 1 91
2 67401 1 91
2 67402 1 91
2 67403 1 91
2 67404 1 91
2 67405 1 91
2 67406 1 91
2 67407 1 91
2 67408 1 91
2 67409 1 91
2 67410 1 91
2 67411 1 91
2 67412 1 91
2 67413 1 91
2 67414 1 91
2 67415 1 91
2 67416 1 91
2 67417 1 92
2 67418 1 92
2 67419 1 92
2 67420 1 92
2 67421 1 92
2 67422 1 92
2 67423 1 93
2 67424 1 93
2 67425 1 93
2 67426 1 94
2 67427 1 94
2 67428 1 94
2 67429 1 94
2 67430 1 95
2 67431 1 95
2 67432 1 95
2 67433 1 95
2 67434 1 95
2 67435 1 95
2 67436 1 95
2 67437 1 95
2 67438 1 103
2 67439 1 103
2 67440 1 103
2 67441 1 103
2 67442 1 103
2 67443 1 103
2 67444 1 103
2 67445 1 103
2 67446 1 103
2 67447 1 104
2 67448 1 104
2 67449 1 105
2 67450 1 105
2 67451 1 105
2 67452 1 105
2 67453 1 105
2 67454 1 105
2 67455 1 105
2 67456 1 105
2 67457 1 105
2 67458 1 105
2 67459 1 105
2 67460 1 105
2 67461 1 105
2 67462 1 105
2 67463 1 105
2 67464 1 105
2 67465 1 105
2 67466 1 105
2 67467 1 105
2 67468 1 105
2 67469 1 105
2 67470 1 105
2 67471 1 105
2 67472 1 105
2 67473 1 105
2 67474 1 105
2 67475 1 105
2 67476 1 105
2 67477 1 105
2 67478 1 105
2 67479 1 105
2 67480 1 105
2 67481 1 105
2 67482 1 105
2 67483 1 105
2 67484 1 105
2 67485 1 105
2 67486 1 105
2 67487 1 105
2 67488 1 105
2 67489 1 105
2 67490 1 105
2 67491 1 105
2 67492 1 106
2 67493 1 106
2 67494 1 106
2 67495 1 107
2 67496 1 107
2 67497 1 107
2 67498 1 107
2 67499 1 108
2 67500 1 108
2 67501 1 108
2 67502 1 108
2 67503 1 108
2 67504 1 108
2 67505 1 108
2 67506 1 108
2 67507 1 108
2 67508 1 108
2 67509 1 108
2 67510 1 108
2 67511 1 108
2 67512 1 108
2 67513 1 108
2 67514 1 108
2 67515 1 108
2 67516 1 108
2 67517 1 108
2 67518 1 108
2 67519 1 108
2 67520 1 108
2 67521 1 108
2 67522 1 108
2 67523 1 108
2 67524 1 108
2 67525 1 108
2 67526 1 108
2 67527 1 108
2 67528 1 108
2 67529 1 108
2 67530 1 108
2 67531 1 108
2 67532 1 108
2 67533 1 108
2 67534 1 108
2 67535 1 108
2 67536 1 108
2 67537 1 108
2 67538 1 108
2 67539 1 108
2 67540 1 108
2 67541 1 108
2 67542 1 109
2 67543 1 109
2 67544 1 109
2 67545 1 109
2 67546 1 109
2 67547 1 109
2 67548 1 109
2 67549 1 109
2 67550 1 109
2 67551 1 109
2 67552 1 109
2 67553 1 109
2 67554 1 109
2 67555 1 110
2 67556 1 110
2 67557 1 110
2 67558 1 110
2 67559 1 110
2 67560 1 110
2 67561 1 110
2 67562 1 110
2 67563 1 110
2 67564 1 110
2 67565 1 110
2 67566 1 110
2 67567 1 110
2 67568 1 110
2 67569 1 110
2 67570 1 110
2 67571 1 111
2 67572 1 111
2 67573 1 111
2 67574 1 111
2 67575 1 111
2 67576 1 111
2 67577 1 111
2 67578 1 111
2 67579 1 111
2 67580 1 111
2 67581 1 111
2 67582 1 111
2 67583 1 111
2 67584 1 111
2 67585 1 123
2 67586 1 123
2 67587 1 124
2 67588 1 124
2 67589 1 124
2 67590 1 124
2 67591 1 124
2 67592 1 124
2 67593 1 124
2 67594 1 124
2 67595 1 124
2 67596 1 124
2 67597 1 124
2 67598 1 124
2 67599 1 124
2 67600 1 124
2 67601 1 124
2 67602 1 124
2 67603 1 125
2 67604 1 125
2 67605 1 125
2 67606 1 125
2 67607 1 125
2 67608 1 125
2 67609 1 125
2 67610 1 126
2 67611 1 126
2 67612 1 126
2 67613 1 126
2 67614 1 126
2 67615 1 126
2 67616 1 126
2 67617 1 126
2 67618 1 126
2 67619 1 126
2 67620 1 126
2 67621 1 126
2 67622 1 135
2 67623 1 135
2 67624 1 135
2 67625 1 135
2 67626 1 135
2 67627 1 135
2 67628 1 135
2 67629 1 135
2 67630 1 135
2 67631 1 135
2 67632 1 135
2 67633 1 135
2 67634 1 135
2 67635 1 135
2 67636 1 135
2 67637 1 135
2 67638 1 135
2 67639 1 135
2 67640 1 135
2 67641 1 135
2 67642 1 135
2 67643 1 135
2 67644 1 135
2 67645 1 135
2 67646 1 135
2 67647 1 135
2 67648 1 135
2 67649 1 135
2 67650 1 135
2 67651 1 135
2 67652 1 135
2 67653 1 135
2 67654 1 135
2 67655 1 135
2 67656 1 135
2 67657 1 135
2 67658 1 135
2 67659 1 135
2 67660 1 135
2 67661 1 135
2 67662 1 135
2 67663 1 135
2 67664 1 135
2 67665 1 135
2 67666 1 135
2 67667 1 135
2 67668 1 135
2 67669 1 135
2 67670 1 135
2 67671 1 135
2 67672 1 135
2 67673 1 135
2 67674 1 135
2 67675 1 135
2 67676 1 135
2 67677 1 135
2 67678 1 135
2 67679 1 135
2 67680 1 135
2 67681 1 135
2 67682 1 135
2 67683 1 135
2 67684 1 135
2 67685 1 135
2 67686 1 135
2 67687 1 135
2 67688 1 135
2 67689 1 135
2 67690 1 135
2 67691 1 135
2 67692 1 135
2 67693 1 135
2 67694 1 135
2 67695 1 135
2 67696 1 135
2 67697 1 135
2 67698 1 135
2 67699 1 135
2 67700 1 135
2 67701 1 135
2 67702 1 135
2 67703 1 135
2 67704 1 135
2 67705 1 135
2 67706 1 136
2 67707 1 136
2 67708 1 136
2 67709 1 136
2 67710 1 136
2 67711 1 136
2 67712 1 136
2 67713 1 136
2 67714 1 136
2 67715 1 136
2 67716 1 136
2 67717 1 136
2 67718 1 136
2 67719 1 136
2 67720 1 136
2 67721 1 136
2 67722 1 136
2 67723 1 136
2 67724 1 136
2 67725 1 136
2 67726 1 136
2 67727 1 136
2 67728 1 136
2 67729 1 136
2 67730 1 136
2 67731 1 136
2 67732 1 136
2 67733 1 136
2 67734 1 136
2 67735 1 136
2 67736 1 136
2 67737 1 136
2 67738 1 136
2 67739 1 136
2 67740 1 136
2 67741 1 136
2 67742 1 136
2 67743 1 136
2 67744 1 136
2 67745 1 136
2 67746 1 136
2 67747 1 136
2 67748 1 136
2 67749 1 136
2 67750 1 136
2 67751 1 136
2 67752 1 136
2 67753 1 136
2 67754 1 136
2 67755 1 136
2 67756 1 136
2 67757 1 136
2 67758 1 136
2 67759 1 136
2 67760 1 136
2 67761 1 136
2 67762 1 136
2 67763 1 136
2 67764 1 136
2 67765 1 136
2 67766 1 136
2 67767 1 136
2 67768 1 136
2 67769 1 136
2 67770 1 136
2 67771 1 136
2 67772 1 136
2 67773 1 136
2 67774 1 136
2 67775 1 136
2 67776 1 136
2 67777 1 136
2 67778 1 136
2 67779 1 136
2 67780 1 136
2 67781 1 136
2 67782 1 136
2 67783 1 136
2 67784 1 136
2 67785 1 136
2 67786 1 136
2 67787 1 136
2 67788 1 136
2 67789 1 136
2 67790 1 136
2 67791 1 136
2 67792 1 136
2 67793 1 136
2 67794 1 136
2 67795 1 136
2 67796 1 136
2 67797 1 136
2 67798 1 136
2 67799 1 136
2 67800 1 136
2 67801 1 136
2 67802 1 136
2 67803 1 136
2 67804 1 136
2 67805 1 136
2 67806 1 136
2 67807 1 136
2 67808 1 136
2 67809 1 137
2 67810 1 137
2 67811 1 137
2 67812 1 137
2 67813 1 137
2 67814 1 137
2 67815 1 137
2 67816 1 137
2 67817 1 137
2 67818 1 137
2 67819 1 137
2 67820 1 137
2 67821 1 138
2 67822 1 138
2 67823 1 138
2 67824 1 138
2 67825 1 138
2 67826 1 138
2 67827 1 138
2 67828 1 138
2 67829 1 138
2 67830 1 138
2 67831 1 138
2 67832 1 138
2 67833 1 138
2 67834 1 138
2 67835 1 138
2 67836 1 138
2 67837 1 138
2 67838 1 138
2 67839 1 138
2 67840 1 138
2 67841 1 138
2 67842 1 138
2 67843 1 138
2 67844 1 138
2 67845 1 138
2 67846 1 138
2 67847 1 138
2 67848 1 138
2 67849 1 138
2 67850 1 138
2 67851 1 138
2 67852 1 138
2 67853 1 138
2 67854 1 138
2 67855 1 138
2 67856 1 138
2 67857 1 138
2 67858 1 138
2 67859 1 138
2 67860 1 138
2 67861 1 138
2 67862 1 138
2 67863 1 138
2 67864 1 139
2 67865 1 139
2 67866 1 140
2 67867 1 140
2 67868 1 140
2 67869 1 140
2 67870 1 140
2 67871 1 140
2 67872 1 140
2 67873 1 141
2 67874 1 141
2 67875 1 141
2 67876 1 141
2 67877 1 141
2 67878 1 141
2 67879 1 142
2 67880 1 142
2 67881 1 143
2 67882 1 143
2 67883 1 143
2 67884 1 143
2 67885 1 143
2 67886 1 143
2 67887 1 143
2 67888 1 143
2 67889 1 143
2 67890 1 143
2 67891 1 143
2 67892 1 143
2 67893 1 143
2 67894 1 143
2 67895 1 143
2 67896 1 143
2 67897 1 143
2 67898 1 143
2 67899 1 143
2 67900 1 144
2 67901 1 144
2 67902 1 145
2 67903 1 145
2 67904 1 145
2 67905 1 145
2 67906 1 145
2 67907 1 145
2 67908 1 145
2 67909 1 145
2 67910 1 145
2 67911 1 145
2 67912 1 145
2 67913 1 145
2 67914 1 145
2 67915 1 145
2 67916 1 145
2 67917 1 145
2 67918 1 145
2 67919 1 145
2 67920 1 145
2 67921 1 145
2 67922 1 145
2 67923 1 145
2 67924 1 145
2 67925 1 145
2 67926 1 145
2 67927 1 145
2 67928 1 145
2 67929 1 145
2 67930 1 145
2 67931 1 145
2 67932 1 145
2 67933 1 145
2 67934 1 145
2 67935 1 145
2 67936 1 145
2 67937 1 145
2 67938 1 145
2 67939 1 145
2 67940 1 145
2 67941 1 145
2 67942 1 145
2 67943 1 145
2 67944 1 145
2 67945 1 145
2 67946 1 146
2 67947 1 146
2 67948 1 147
2 67949 1 147
2 67950 1 147
2 67951 1 147
2 67952 1 147
2 67953 1 147
2 67954 1 147
2 67955 1 147
2 67956 1 147
2 67957 1 147
2 67958 1 147
2 67959 1 147
2 67960 1 147
2 67961 1 147
2 67962 1 148
2 67963 1 148
2 67964 1 148
2 67965 1 148
2 67966 1 148
2 67967 1 155
2 67968 1 155
2 67969 1 155
2 67970 1 155
2 67971 1 156
2 67972 1 156
2 67973 1 156
2 67974 1 156
2 67975 1 156
2 67976 1 156
2 67977 1 156
2 67978 1 156
2 67979 1 156
2 67980 1 156
2 67981 1 156
2 67982 1 156
2 67983 1 156
2 67984 1 156
2 67985 1 156
2 67986 1 156
2 67987 1 156
2 67988 1 156
2 67989 1 156
2 67990 1 156
2 67991 1 156
2 67992 1 156
2 67993 1 156
2 67994 1 156
2 67995 1 156
2 67996 1 156
2 67997 1 156
2 67998 1 156
2 67999 1 156
2 68000 1 156
2 68001 1 156
2 68002 1 156
2 68003 1 156
2 68004 1 156
2 68005 1 156
2 68006 1 156
2 68007 1 156
2 68008 1 156
2 68009 1 156
2 68010 1 156
2 68011 1 156
2 68012 1 156
2 68013 1 156
2 68014 1 156
2 68015 1 156
2 68016 1 156
2 68017 1 156
2 68018 1 156
2 68019 1 156
2 68020 1 156
2 68021 1 156
2 68022 1 156
2 68023 1 156
2 68024 1 156
2 68025 1 156
2 68026 1 156
2 68027 1 156
2 68028 1 156
2 68029 1 156
2 68030 1 156
2 68031 1 156
2 68032 1 156
2 68033 1 156
2 68034 1 156
2 68035 1 156
2 68036 1 156
2 68037 1 156
2 68038 1 156
2 68039 1 156
2 68040 1 156
2 68041 1 156
2 68042 1 156
2 68043 1 156
2 68044 1 156
2 68045 1 156
2 68046 1 156
2 68047 1 156
2 68048 1 156
2 68049 1 156
2 68050 1 156
2 68051 1 156
2 68052 1 156
2 68053 1 156
2 68054 1 156
2 68055 1 156
2 68056 1 156
2 68057 1 156
2 68058 1 156
2 68059 1 156
2 68060 1 156
2 68061 1 156
2 68062 1 156
2 68063 1 156
2 68064 1 156
2 68065 1 157
2 68066 1 157
2 68067 1 157
2 68068 1 157
2 68069 1 157
2 68070 1 157
2 68071 1 157
2 68072 1 157
2 68073 1 157
2 68074 1 157
2 68075 1 157
2 68076 1 157
2 68077 1 157
2 68078 1 157
2 68079 1 157
2 68080 1 157
2 68081 1 157
2 68082 1 157
2 68083 1 157
2 68084 1 157
2 68085 1 157
2 68086 1 157
2 68087 1 157
2 68088 1 157
2 68089 1 157
2 68090 1 157
2 68091 1 157
2 68092 1 157
2 68093 1 157
2 68094 1 157
2 68095 1 157
2 68096 1 157
2 68097 1 157
2 68098 1 157
2 68099 1 157
2 68100 1 157
2 68101 1 157
2 68102 1 157
2 68103 1 157
2 68104 1 157
2 68105 1 157
2 68106 1 157
2 68107 1 157
2 68108 1 157
2 68109 1 157
2 68110 1 157
2 68111 1 157
2 68112 1 157
2 68113 1 157
2 68114 1 157
2 68115 1 157
2 68116 1 157
2 68117 1 157
2 68118 1 157
2 68119 1 157
2 68120 1 157
2 68121 1 157
2 68122 1 157
2 68123 1 157
2 68124 1 157
2 68125 1 157
2 68126 1 157
2 68127 1 157
2 68128 1 157
2 68129 1 157
2 68130 1 157
2 68131 1 157
2 68132 1 157
2 68133 1 157
2 68134 1 157
2 68135 1 157
2 68136 1 157
2 68137 1 157
2 68138 1 157
2 68139 1 157
2 68140 1 157
2 68141 1 157
2 68142 1 157
2 68143 1 157
2 68144 1 157
2 68145 1 157
2 68146 1 157
2 68147 1 157
2 68148 1 157
2 68149 1 157
2 68150 1 157
2 68151 1 157
2 68152 1 157
2 68153 1 157
2 68154 1 157
2 68155 1 157
2 68156 1 157
2 68157 1 157
2 68158 1 157
2 68159 1 157
2 68160 1 157
2 68161 1 157
2 68162 1 157
2 68163 1 157
2 68164 1 157
2 68165 1 157
2 68166 1 157
2 68167 1 157
2 68168 1 157
2 68169 1 157
2 68170 1 157
2 68171 1 157
2 68172 1 157
2 68173 1 157
2 68174 1 157
2 68175 1 157
2 68176 1 157
2 68177 1 157
2 68178 1 157
2 68179 1 157
2 68180 1 157
2 68181 1 157
2 68182 1 157
2 68183 1 157
2 68184 1 157
2 68185 1 157
2 68186 1 157
2 68187 1 157
2 68188 1 157
2 68189 1 157
2 68190 1 157
2 68191 1 157
2 68192 1 157
2 68193 1 158
2 68194 1 158
2 68195 1 160
2 68196 1 160
2 68197 1 160
2 68198 1 160
2 68199 1 160
2 68200 1 160
2 68201 1 160
2 68202 1 161
2 68203 1 161
2 68204 1 161
2 68205 1 161
2 68206 1 161
2 68207 1 161
2 68208 1 182
2 68209 1 182
2 68210 1 185
2 68211 1 185
2 68212 1 185
2 68213 1 185
2 68214 1 185
2 68215 1 185
2 68216 1 185
2 68217 1 185
2 68218 1 185
2 68219 1 185
2 68220 1 185
2 68221 1 185
2 68222 1 185
2 68223 1 185
2 68224 1 185
2 68225 1 185
2 68226 1 185
2 68227 1 185
2 68228 1 185
2 68229 1 185
2 68230 1 185
2 68231 1 185
2 68232 1 185
2 68233 1 185
2 68234 1 185
2 68235 1 185
2 68236 1 185
2 68237 1 185
2 68238 1 185
2 68239 1 185
2 68240 1 185
2 68241 1 185
2 68242 1 185
2 68243 1 185
2 68244 1 185
2 68245 1 185
2 68246 1 185
2 68247 1 185
2 68248 1 185
2 68249 1 185
2 68250 1 185
2 68251 1 185
2 68252 1 185
2 68253 1 185
2 68254 1 185
2 68255 1 185
2 68256 1 185
2 68257 1 185
2 68258 1 185
2 68259 1 185
2 68260 1 185
2 68261 1 185
2 68262 1 185
2 68263 1 185
2 68264 1 185
2 68265 1 185
2 68266 1 185
2 68267 1 185
2 68268 1 185
2 68269 1 185
2 68270 1 185
2 68271 1 185
2 68272 1 185
2 68273 1 185
2 68274 1 185
2 68275 1 185
2 68276 1 185
2 68277 1 185
2 68278 1 185
2 68279 1 185
2 68280 1 185
2 68281 1 185
2 68282 1 185
2 68283 1 185
2 68284 1 185
2 68285 1 185
2 68286 1 185
2 68287 1 185
2 68288 1 185
2 68289 1 185
2 68290 1 185
2 68291 1 186
2 68292 1 186
2 68293 1 186
2 68294 1 186
2 68295 1 186
2 68296 1 186
2 68297 1 186
2 68298 1 186
2 68299 1 186
2 68300 1 186
2 68301 1 186
2 68302 1 186
2 68303 1 186
2 68304 1 186
2 68305 1 186
2 68306 1 186
2 68307 1 186
2 68308 1 186
2 68309 1 186
2 68310 1 186
2 68311 1 186
2 68312 1 186
2 68313 1 186
2 68314 1 186
2 68315 1 186
2 68316 1 186
2 68317 1 186
2 68318 1 186
2 68319 1 186
2 68320 1 186
2 68321 1 186
2 68322 1 186
2 68323 1 186
2 68324 1 186
2 68325 1 186
2 68326 1 186
2 68327 1 186
2 68328 1 186
2 68329 1 186
2 68330 1 186
2 68331 1 186
2 68332 1 186
2 68333 1 186
2 68334 1 186
2 68335 1 186
2 68336 1 186
2 68337 1 186
2 68338 1 186
2 68339 1 186
2 68340 1 186
2 68341 1 186
2 68342 1 186
2 68343 1 186
2 68344 1 186
2 68345 1 186
2 68346 1 186
2 68347 1 186
2 68348 1 186
2 68349 1 186
2 68350 1 186
2 68351 1 186
2 68352 1 186
2 68353 1 186
2 68354 1 186
2 68355 1 186
2 68356 1 186
2 68357 1 186
2 68358 1 186
2 68359 1 186
2 68360 1 186
2 68361 1 186
2 68362 1 186
2 68363 1 186
2 68364 1 186
2 68365 1 186
2 68366 1 186
2 68367 1 186
2 68368 1 186
2 68369 1 186
2 68370 1 186
2 68371 1 186
2 68372 1 186
2 68373 1 186
2 68374 1 186
2 68375 1 186
2 68376 1 186
2 68377 1 186
2 68378 1 186
2 68379 1 186
2 68380 1 186
2 68381 1 186
2 68382 1 186
2 68383 1 186
2 68384 1 186
2 68385 1 186
2 68386 1 186
2 68387 1 186
2 68388 1 186
2 68389 1 186
2 68390 1 186
2 68391 1 186
2 68392 1 186
2 68393 1 186
2 68394 1 186
2 68395 1 186
2 68396 1 186
2 68397 1 186
2 68398 1 186
2 68399 1 186
2 68400 1 186
2 68401 1 186
2 68402 1 186
2 68403 1 186
2 68404 1 186
2 68405 1 186
2 68406 1 186
2 68407 1 186
2 68408 1 186
2 68409 1 186
2 68410 1 186
2 68411 1 186
2 68412 1 186
2 68413 1 186
2 68414 1 186
2 68415 1 186
2 68416 1 186
2 68417 1 186
2 68418 1 186
2 68419 1 186
2 68420 1 186
2 68421 1 186
2 68422 1 186
2 68423 1 186
2 68424 1 186
2 68425 1 187
2 68426 1 187
2 68427 1 187
2 68428 1 188
2 68429 1 188
2 68430 1 188
2 68431 1 188
2 68432 1 188
2 68433 1 188
2 68434 1 188
2 68435 1 188
2 68436 1 188
2 68437 1 188
2 68438 1 188
2 68439 1 188
2 68440 1 188
2 68441 1 188
2 68442 1 188
2 68443 1 188
2 68444 1 189
2 68445 1 189
2 68446 1 189
2 68447 1 189
2 68448 1 189
2 68449 1 189
2 68450 1 189
2 68451 1 189
2 68452 1 189
2 68453 1 189
2 68454 1 189
2 68455 1 189
2 68456 1 189
2 68457 1 189
2 68458 1 189
2 68459 1 189
2 68460 1 189
2 68461 1 189
2 68462 1 189
2 68463 1 189
2 68464 1 189
2 68465 1 189
2 68466 1 189
2 68467 1 189
2 68468 1 189
2 68469 1 189
2 68470 1 189
2 68471 1 189
2 68472 1 189
2 68473 1 189
2 68474 1 189
2 68475 1 189
2 68476 1 189
2 68477 1 189
2 68478 1 189
2 68479 1 189
2 68480 1 189
2 68481 1 189
2 68482 1 189
2 68483 1 189
2 68484 1 189
2 68485 1 189
2 68486 1 189
2 68487 1 189
2 68488 1 189
2 68489 1 189
2 68490 1 189
2 68491 1 189
2 68492 1 189
2 68493 1 189
2 68494 1 189
2 68495 1 189
2 68496 1 189
2 68497 1 189
2 68498 1 189
2 68499 1 189
2 68500 1 189
2 68501 1 189
2 68502 1 189
2 68503 1 189
2 68504 1 189
2 68505 1 189
2 68506 1 189
2 68507 1 189
2 68508 1 189
2 68509 1 189
2 68510 1 189
2 68511 1 189
2 68512 1 189
2 68513 1 189
2 68514 1 189
2 68515 1 189
2 68516 1 189
2 68517 1 189
2 68518 1 189
2 68519 1 189
2 68520 1 189
2 68521 1 189
2 68522 1 189
2 68523 1 189
2 68524 1 189
2 68525 1 189
2 68526 1 189
2 68527 1 189
2 68528 1 189
2 68529 1 189
2 68530 1 189
2 68531 1 189
2 68532 1 189
2 68533 1 189
2 68534 1 189
2 68535 1 189
2 68536 1 189
2 68537 1 189
2 68538 1 189
2 68539 1 189
2 68540 1 189
2 68541 1 189
2 68542 1 189
2 68543 1 189
2 68544 1 189
2 68545 1 189
2 68546 1 189
2 68547 1 190
2 68548 1 190
2 68549 1 190
2 68550 1 190
2 68551 1 190
2 68552 1 190
2 68553 1 190
2 68554 1 190
2 68555 1 190
2 68556 1 190
2 68557 1 190
2 68558 1 190
2 68559 1 190
2 68560 1 190
2 68561 1 190
2 68562 1 190
2 68563 1 190
2 68564 1 190
2 68565 1 190
2 68566 1 190
2 68567 1 190
2 68568 1 190
2 68569 1 190
2 68570 1 190
2 68571 1 190
2 68572 1 190
2 68573 1 190
2 68574 1 190
2 68575 1 190
2 68576 1 190
2 68577 1 190
2 68578 1 190
2 68579 1 190
2 68580 1 190
2 68581 1 190
2 68582 1 190
2 68583 1 190
2 68584 1 190
2 68585 1 190
2 68586 1 190
2 68587 1 190
2 68588 1 190
2 68589 1 190
2 68590 1 190
2 68591 1 190
2 68592 1 190
2 68593 1 190
2 68594 1 190
2 68595 1 190
2 68596 1 190
2 68597 1 190
2 68598 1 190
2 68599 1 190
2 68600 1 190
2 68601 1 190
2 68602 1 190
2 68603 1 190
2 68604 1 190
2 68605 1 190
2 68606 1 190
2 68607 1 190
2 68608 1 190
2 68609 1 190
2 68610 1 190
2 68611 1 190
2 68612 1 190
2 68613 1 190
2 68614 1 190
2 68615 1 190
2 68616 1 190
2 68617 1 190
2 68618 1 190
2 68619 1 190
2 68620 1 190
2 68621 1 190
2 68622 1 190
2 68623 1 190
2 68624 1 190
2 68625 1 190
2 68626 1 190
2 68627 1 190
2 68628 1 190
2 68629 1 190
2 68630 1 190
2 68631 1 190
2 68632 1 190
2 68633 1 190
2 68634 1 190
2 68635 1 190
2 68636 1 190
2 68637 1 190
2 68638 1 190
2 68639 1 190
2 68640 1 190
2 68641 1 190
2 68642 1 190
2 68643 1 190
2 68644 1 190
2 68645 1 190
2 68646 1 190
2 68647 1 190
2 68648 1 190
2 68649 1 190
2 68650 1 194
2 68651 1 194
2 68652 1 194
2 68653 1 194
2 68654 1 194
2 68655 1 194
2 68656 1 194
2 68657 1 195
2 68658 1 195
2 68659 1 195
2 68660 1 195
2 68661 1 195
2 68662 1 195
2 68663 1 195
2 68664 1 195
2 68665 1 195
2 68666 1 195
2 68667 1 195
2 68668 1 196
2 68669 1 196
2 68670 1 196
2 68671 1 196
2 68672 1 196
2 68673 1 196
2 68674 1 196
2 68675 1 196
2 68676 1 196
2 68677 1 196
2 68678 1 196
2 68679 1 196
2 68680 1 196
2 68681 1 196
2 68682 1 196
2 68683 1 196
2 68684 1 196
2 68685 1 196
2 68686 1 196
2 68687 1 196
2 68688 1 196
2 68689 1 196
2 68690 1 196
2 68691 1 197
2 68692 1 197
2 68693 1 197
2 68694 1 197
2 68695 1 197
2 68696 1 197
2 68697 1 197
2 68698 1 197
2 68699 1 197
2 68700 1 197
2 68701 1 197
2 68702 1 198
2 68703 1 198
2 68704 1 198
2 68705 1 198
2 68706 1 198
2 68707 1 198
2 68708 1 198
2 68709 1 198
2 68710 1 198
2 68711 1 199
2 68712 1 199
2 68713 1 202
2 68714 1 202
2 68715 1 207
2 68716 1 207
2 68717 1 207
2 68718 1 207
2 68719 1 207
2 68720 1 207
2 68721 1 207
2 68722 1 207
2 68723 1 207
2 68724 1 207
2 68725 1 207
2 68726 1 207
2 68727 1 207
2 68728 1 207
2 68729 1 207
2 68730 1 207
2 68731 1 207
2 68732 1 207
2 68733 1 207
2 68734 1 207
2 68735 1 207
2 68736 1 207
2 68737 1 207
2 68738 1 207
2 68739 1 207
2 68740 1 207
2 68741 1 207
2 68742 1 207
2 68743 1 207
2 68744 1 207
2 68745 1 207
2 68746 1 207
2 68747 1 207
2 68748 1 207
2 68749 1 207
2 68750 1 207
2 68751 1 207
2 68752 1 207
2 68753 1 207
2 68754 1 207
2 68755 1 207
2 68756 1 207
2 68757 1 207
2 68758 1 207
2 68759 1 207
2 68760 1 207
2 68761 1 207
2 68762 1 207
2 68763 1 207
2 68764 1 207
2 68765 1 207
2 68766 1 207
2 68767 1 207
2 68768 1 207
2 68769 1 207
2 68770 1 207
2 68771 1 207
2 68772 1 207
2 68773 1 207
2 68774 1 207
2 68775 1 207
2 68776 1 207
2 68777 1 207
2 68778 1 207
2 68779 1 207
2 68780 1 207
2 68781 1 207
2 68782 1 207
2 68783 1 207
2 68784 1 207
2 68785 1 207
2 68786 1 207
2 68787 1 207
2 68788 1 207
2 68789 1 207
2 68790 1 207
2 68791 1 207
2 68792 1 207
2 68793 1 207
2 68794 1 207
2 68795 1 207
2 68796 1 207
2 68797 1 207
2 68798 1 207
2 68799 1 207
2 68800 1 207
2 68801 1 207
2 68802 1 207
2 68803 1 207
2 68804 1 207
2 68805 1 207
2 68806 1 207
2 68807 1 207
2 68808 1 207
2 68809 1 207
2 68810 1 207
2 68811 1 207
2 68812 1 207
2 68813 1 207
2 68814 1 208
2 68815 1 208
2 68816 1 208
2 68817 1 208
2 68818 1 208
2 68819 1 208
2 68820 1 208
2 68821 1 208
2 68822 1 208
2 68823 1 208
2 68824 1 208
2 68825 1 208
2 68826 1 208
2 68827 1 208
2 68828 1 208
2 68829 1 208
2 68830 1 208
2 68831 1 208
2 68832 1 208
2 68833 1 208
2 68834 1 208
2 68835 1 208
2 68836 1 208
2 68837 1 208
2 68838 1 208
2 68839 1 208
2 68840 1 208
2 68841 1 208
2 68842 1 208
2 68843 1 208
2 68844 1 208
2 68845 1 208
2 68846 1 208
2 68847 1 208
2 68848 1 208
2 68849 1 208
2 68850 1 208
2 68851 1 208
2 68852 1 208
2 68853 1 208
2 68854 1 208
2 68855 1 208
2 68856 1 208
2 68857 1 208
2 68858 1 208
2 68859 1 208
2 68860 1 208
2 68861 1 208
2 68862 1 208
2 68863 1 208
2 68864 1 208
2 68865 1 208
2 68866 1 208
2 68867 1 208
2 68868 1 208
2 68869 1 208
2 68870 1 208
2 68871 1 208
2 68872 1 208
2 68873 1 208
2 68874 1 208
2 68875 1 208
2 68876 1 208
2 68877 1 208
2 68878 1 208
2 68879 1 208
2 68880 1 208
2 68881 1 208
2 68882 1 208
2 68883 1 208
2 68884 1 208
2 68885 1 208
2 68886 1 208
2 68887 1 208
2 68888 1 208
2 68889 1 208
2 68890 1 208
2 68891 1 208
2 68892 1 208
2 68893 1 208
2 68894 1 208
2 68895 1 208
2 68896 1 208
2 68897 1 209
2 68898 1 209
2 68899 1 209
2 68900 1 209
2 68901 1 209
2 68902 1 209
2 68903 1 209
2 68904 1 209
2 68905 1 210
2 68906 1 210
2 68907 1 211
2 68908 1 211
2 68909 1 211
2 68910 1 211
2 68911 1 211
2 68912 1 212
2 68913 1 212
2 68914 1 212
2 68915 1 212
2 68916 1 212
2 68917 1 212
2 68918 1 212
2 68919 1 212
2 68920 1 212
2 68921 1 212
2 68922 1 212
2 68923 1 212
2 68924 1 213
2 68925 1 213
2 68926 1 214
2 68927 1 214
2 68928 1 214
2 68929 1 214
2 68930 1 214
2 68931 1 214
2 68932 1 214
2 68933 1 214
2 68934 1 214
2 68935 1 215
2 68936 1 215
2 68937 1 215
2 68938 1 215
2 68939 1 215
2 68940 1 215
2 68941 1 215
2 68942 1 216
2 68943 1 216
2 68944 1 216
2 68945 1 218
2 68946 1 218
2 68947 1 219
2 68948 1 219
2 68949 1 220
2 68950 1 220
2 68951 1 220
2 68952 1 220
2 68953 1 220
2 68954 1 220
2 68955 1 220
2 68956 1 220
2 68957 1 220
2 68958 1 220
2 68959 1 220
2 68960 1 220
2 68961 1 220
2 68962 1 220
2 68963 1 220
2 68964 1 220
2 68965 1 220
2 68966 1 221
2 68967 1 221
2 68968 1 222
2 68969 1 222
2 68970 1 222
2 68971 1 222
2 68972 1 222
2 68973 1 222
2 68974 1 222
2 68975 1 222
2 68976 1 222
2 68977 1 222
2 68978 1 222
2 68979 1 222
2 68980 1 222
2 68981 1 222
2 68982 1 222
2 68983 1 222
2 68984 1 222
2 68985 1 222
2 68986 1 222
2 68987 1 222
2 68988 1 222
2 68989 1 222
2 68990 1 222
2 68991 1 222
2 68992 1 222
2 68993 1 222
2 68994 1 222
2 68995 1 222
2 68996 1 222
2 68997 1 222
2 68998 1 222
2 68999 1 222
2 69000 1 222
2 69001 1 222
2 69002 1 222
2 69003 1 222
2 69004 1 222
2 69005 1 222
2 69006 1 222
2 69007 1 222
2 69008 1 222
2 69009 1 222
2 69010 1 222
2 69011 1 222
2 69012 1 222
2 69013 1 222
2 69014 1 222
2 69015 1 223
2 69016 1 223
2 69017 1 223
2 69018 1 223
2 69019 1 223
2 69020 1 223
2 69021 1 223
2 69022 1 223
2 69023 1 223
2 69024 1 223
2 69025 1 223
2 69026 1 223
2 69027 1 223
2 69028 1 223
2 69029 1 223
2 69030 1 223
2 69031 1 223
2 69032 1 223
2 69033 1 223
2 69034 1 223
2 69035 1 223
2 69036 1 223
2 69037 1 223
2 69038 1 223
2 69039 1 223
2 69040 1 223
2 69041 1 223
2 69042 1 223
2 69043 1 223
2 69044 1 223
2 69045 1 223
2 69046 1 223
2 69047 1 223
2 69048 1 223
2 69049 1 223
2 69050 1 223
2 69051 1 223
2 69052 1 223
2 69053 1 223
2 69054 1 223
2 69055 1 223
2 69056 1 223
2 69057 1 223
2 69058 1 223
2 69059 1 223
2 69060 1 223
2 69061 1 223
2 69062 1 223
2 69063 1 223
2 69064 1 223
2 69065 1 223
2 69066 1 223
2 69067 1 223
2 69068 1 223
2 69069 1 223
2 69070 1 223
2 69071 1 223
2 69072 1 223
2 69073 1 223
2 69074 1 223
2 69075 1 223
2 69076 1 223
2 69077 1 223
2 69078 1 223
2 69079 1 223
2 69080 1 223
2 69081 1 223
2 69082 1 223
2 69083 1 223
2 69084 1 224
2 69085 1 224
2 69086 1 224
2 69087 1 225
2 69088 1 225
2 69089 1 225
2 69090 1 225
2 69091 1 227
2 69092 1 227
2 69093 1 227
2 69094 1 227
2 69095 1 227
2 69096 1 229
2 69097 1 229
2 69098 1 229
2 69099 1 231
2 69100 1 231
2 69101 1 233
2 69102 1 233
2 69103 1 234
2 69104 1 234
2 69105 1 234
2 69106 1 234
2 69107 1 234
2 69108 1 234
2 69109 1 234
2 69110 1 234
2 69111 1 234
2 69112 1 234
2 69113 1 234
2 69114 1 234
2 69115 1 234
2 69116 1 234
2 69117 1 234
2 69118 1 234
2 69119 1 234
2 69120 1 234
2 69121 1 234
2 69122 1 235
2 69123 1 235
2 69124 1 236
2 69125 1 236
2 69126 1 236
2 69127 1 236
2 69128 1 236
2 69129 1 236
2 69130 1 236
2 69131 1 236
2 69132 1 237
2 69133 1 237
2 69134 1 237
2 69135 1 238
2 69136 1 238
2 69137 1 238
2 69138 1 238
2 69139 1 238
2 69140 1 238
2 69141 1 238
2 69142 1 246
2 69143 1 246
2 69144 1 246
2 69145 1 246
2 69146 1 246
2 69147 1 246
2 69148 1 248
2 69149 1 248
2 69150 1 263
2 69151 1 263
2 69152 1 270
2 69153 1 270
2 69154 1 270
2 69155 1 270
2 69156 1 270
2 69157 1 270
2 69158 1 271
2 69159 1 271
2 69160 1 271
2 69161 1 271
2 69162 1 271
2 69163 1 271
2 69164 1 271
2 69165 1 271
2 69166 1 271
2 69167 1 271
2 69168 1 272
2 69169 1 272
2 69170 1 272
2 69171 1 272
2 69172 1 272
2 69173 1 273
2 69174 1 273
2 69175 1 273
2 69176 1 273
2 69177 1 273
2 69178 1 273
2 69179 1 273
2 69180 1 273
2 69181 1 273
2 69182 1 273
2 69183 1 273
2 69184 1 273
2 69185 1 273
2 69186 1 273
2 69187 1 273
2 69188 1 273
2 69189 1 273
2 69190 1 273
2 69191 1 273
2 69192 1 273
2 69193 1 273
2 69194 1 273
2 69195 1 273
2 69196 1 273
2 69197 1 273
2 69198 1 273
2 69199 1 274
2 69200 1 274
2 69201 1 274
2 69202 1 275
2 69203 1 275
2 69204 1 275
2 69205 1 276
2 69206 1 276
2 69207 1 277
2 69208 1 277
2 69209 1 278
2 69210 1 278
2 69211 1 278
2 69212 1 278
2 69213 1 286
2 69214 1 286
2 69215 1 286
2 69216 1 286
2 69217 1 286
2 69218 1 286
2 69219 1 286
2 69220 1 286
2 69221 1 287
2 69222 1 287
2 69223 1 287
2 69224 1 288
2 69225 1 288
2 69226 1 288
2 69227 1 288
2 69228 1 289
2 69229 1 289
2 69230 1 289
2 69231 1 289
2 69232 1 289
2 69233 1 289
2 69234 1 289
2 69235 1 289
2 69236 1 289
2 69237 1 289
2 69238 1 289
2 69239 1 289
2 69240 1 289
2 69241 1 289
2 69242 1 289
2 69243 1 289
2 69244 1 289
2 69245 1 289
2 69246 1 289
2 69247 1 289
2 69248 1 289
2 69249 1 289
2 69250 1 289
2 69251 1 290
2 69252 1 290
2 69253 1 290
2 69254 1 290
2 69255 1 290
2 69256 1 290
2 69257 1 290
2 69258 1 290
2 69259 1 290
2 69260 1 290
2 69261 1 290
2 69262 1 290
2 69263 1 290
2 69264 1 290
2 69265 1 290
2 69266 1 290
2 69267 1 290
2 69268 1 290
2 69269 1 290
2 69270 1 290
2 69271 1 290
2 69272 1 290
2 69273 1 290
2 69274 1 290
2 69275 1 290
2 69276 1 290
2 69277 1 290
2 69278 1 290
2 69279 1 290
2 69280 1 290
2 69281 1 290
2 69282 1 290
2 69283 1 290
2 69284 1 290
2 69285 1 290
2 69286 1 290
2 69287 1 290
2 69288 1 290
2 69289 1 290
2 69290 1 290
2 69291 1 290
2 69292 1 290
2 69293 1 290
2 69294 1 290
2 69295 1 290
2 69296 1 290
2 69297 1 290
2 69298 1 290
2 69299 1 290
2 69300 1 290
2 69301 1 290
2 69302 1 290
2 69303 1 291
2 69304 1 291
2 69305 1 291
2 69306 1 291
2 69307 1 291
2 69308 1 291
2 69309 1 291
2 69310 1 291
2 69311 1 291
2 69312 1 291
2 69313 1 291
2 69314 1 291
2 69315 1 291
2 69316 1 299
2 69317 1 299
2 69318 1 299
2 69319 1 299
2 69320 1 299
2 69321 1 299
2 69322 1 299
2 69323 1 299
2 69324 1 299
2 69325 1 307
2 69326 1 307
2 69327 1 307
2 69328 1 307
2 69329 1 307
2 69330 1 307
2 69331 1 307
2 69332 1 307
2 69333 1 307
2 69334 1 307
2 69335 1 307
2 69336 1 307
2 69337 1 307
2 69338 1 307
2 69339 1 307
2 69340 1 307
2 69341 1 308
2 69342 1 308
2 69343 1 308
2 69344 1 308
2 69345 1 308
2 69346 1 308
2 69347 1 308
2 69348 1 308
2 69349 1 308
2 69350 1 308
2 69351 1 308
2 69352 1 308
2 69353 1 308
2 69354 1 308
2 69355 1 309
2 69356 1 309
2 69357 1 309
2 69358 1 310
2 69359 1 310
2 69360 1 310
2 69361 1 310
2 69362 1 310
2 69363 1 310
2 69364 1 311
2 69365 1 311
2 69366 1 313
2 69367 1 313
2 69368 1 318
2 69369 1 318
2 69370 1 318
2 69371 1 318
2 69372 1 318
2 69373 1 318
2 69374 1 318
2 69375 1 318
2 69376 1 318
2 69377 1 318
2 69378 1 318
2 69379 1 318
2 69380 1 318
2 69381 1 318
2 69382 1 318
2 69383 1 318
2 69384 1 318
2 69385 1 318
2 69386 1 318
2 69387 1 318
2 69388 1 318
2 69389 1 318
2 69390 1 318
2 69391 1 318
2 69392 1 318
2 69393 1 318
2 69394 1 318
2 69395 1 318
2 69396 1 318
2 69397 1 318
2 69398 1 318
2 69399 1 318
2 69400 1 318
2 69401 1 318
2 69402 1 318
2 69403 1 318
2 69404 1 319
2 69405 1 319
2 69406 1 319
2 69407 1 319
2 69408 1 319
2 69409 1 319
2 69410 1 319
2 69411 1 319
2 69412 1 319
2 69413 1 319
2 69414 1 319
2 69415 1 319
2 69416 1 319
2 69417 1 319
2 69418 1 319
2 69419 1 319
2 69420 1 319
2 69421 1 319
2 69422 1 319
2 69423 1 319
2 69424 1 319
2 69425 1 319
2 69426 1 319
2 69427 1 319
2 69428 1 319
2 69429 1 319
2 69430 1 319
2 69431 1 319
2 69432 1 319
2 69433 1 319
2 69434 1 319
2 69435 1 319
2 69436 1 319
2 69437 1 321
2 69438 1 321
2 69439 1 322
2 69440 1 322
2 69441 1 322
2 69442 1 322
2 69443 1 322
2 69444 1 322
2 69445 1 323
2 69446 1 323
2 69447 1 323
2 69448 1 323
2 69449 1 323
2 69450 1 323
2 69451 1 323
2 69452 1 323
2 69453 1 323
2 69454 1 323
2 69455 1 323
2 69456 1 323
2 69457 1 323
2 69458 1 323
2 69459 1 323
2 69460 1 323
2 69461 1 323
2 69462 1 323
2 69463 1 323
2 69464 1 323
2 69465 1 323
2 69466 1 323
2 69467 1 323
2 69468 1 323
2 69469 1 323
2 69470 1 323
2 69471 1 323
2 69472 1 323
2 69473 1 323
2 69474 1 323
2 69475 1 324
2 69476 1 324
2 69477 1 324
2 69478 1 324
2 69479 1 325
2 69480 1 325
2 69481 1 325
2 69482 1 325
2 69483 1 325
2 69484 1 325
2 69485 1 325
2 69486 1 328
2 69487 1 328
2 69488 1 328
2 69489 1 328
2 69490 1 335
2 69491 1 335
2 69492 1 335
2 69493 1 335
2 69494 1 335
2 69495 1 335
2 69496 1 335
2 69497 1 335
2 69498 1 336
2 69499 1 336
2 69500 1 336
2 69501 1 339
2 69502 1 339
2 69503 1 339
2 69504 1 339
2 69505 1 339
2 69506 1 339
2 69507 1 339
2 69508 1 339
2 69509 1 340
2 69510 1 340
2 69511 1 341
2 69512 1 341
2 69513 1 341
2 69514 1 341
2 69515 1 341
2 69516 1 341
2 69517 1 341
2 69518 1 341
2 69519 1 341
2 69520 1 341
2 69521 1 341
2 69522 1 341
2 69523 1 341
2 69524 1 341
2 69525 1 341
2 69526 1 341
2 69527 1 341
2 69528 1 341
2 69529 1 341
2 69530 1 341
2 69531 1 341
2 69532 1 341
2 69533 1 341
2 69534 1 341
2 69535 1 341
2 69536 1 341
2 69537 1 341
2 69538 1 341
2 69539 1 341
2 69540 1 341
2 69541 1 341
2 69542 1 341
2 69543 1 341
2 69544 1 341
2 69545 1 341
2 69546 1 341
2 69547 1 341
2 69548 1 341
2 69549 1 341
2 69550 1 341
2 69551 1 341
2 69552 1 341
2 69553 1 341
2 69554 1 341
2 69555 1 341
2 69556 1 341
2 69557 1 341
2 69558 1 341
2 69559 1 341
2 69560 1 341
2 69561 1 341
2 69562 1 341
2 69563 1 341
2 69564 1 342
2 69565 1 342
2 69566 1 342
2 69567 1 343
2 69568 1 343
2 69569 1 343
2 69570 1 343
2 69571 1 343
2 69572 1 343
2 69573 1 343
2 69574 1 343
2 69575 1 343
2 69576 1 343
2 69577 1 343
2 69578 1 343
2 69579 1 343
2 69580 1 343
2 69581 1 343
2 69582 1 343
2 69583 1 343
2 69584 1 343
2 69585 1 343
2 69586 1 343
2 69587 1 345
2 69588 1 345
2 69589 1 358
2 69590 1 358
2 69591 1 358
2 69592 1 358
2 69593 1 358
2 69594 1 358
2 69595 1 358
2 69596 1 358
2 69597 1 358
2 69598 1 358
2 69599 1 358
2 69600 1 358
2 69601 1 358
2 69602 1 358
2 69603 1 358
2 69604 1 358
2 69605 1 358
2 69606 1 358
2 69607 1 358
2 69608 1 358
2 69609 1 358
2 69610 1 358
2 69611 1 358
2 69612 1 358
2 69613 1 358
2 69614 1 358
2 69615 1 358
2 69616 1 358
2 69617 1 358
2 69618 1 358
2 69619 1 358
2 69620 1 358
2 69621 1 358
2 69622 1 358
2 69623 1 358
2 69624 1 358
2 69625 1 358
2 69626 1 358
2 69627 1 358
2 69628 1 358
2 69629 1 358
2 69630 1 358
2 69631 1 358
2 69632 1 358
2 69633 1 358
2 69634 1 358
2 69635 1 358
2 69636 1 358
2 69637 1 358
2 69638 1 358
2 69639 1 358
2 69640 1 358
2 69641 1 358
2 69642 1 358
2 69643 1 358
2 69644 1 358
2 69645 1 358
2 69646 1 358
2 69647 1 358
2 69648 1 358
2 69649 1 358
2 69650 1 358
2 69651 1 358
2 69652 1 358
2 69653 1 358
2 69654 1 358
2 69655 1 358
2 69656 1 358
2 69657 1 358
2 69658 1 358
2 69659 1 358
2 69660 1 358
2 69661 1 358
2 69662 1 358
2 69663 1 358
2 69664 1 358
2 69665 1 358
2 69666 1 358
2 69667 1 358
2 69668 1 358
2 69669 1 358
2 69670 1 358
2 69671 1 358
2 69672 1 358
2 69673 1 358
2 69674 1 358
2 69675 1 358
2 69676 1 358
2 69677 1 358
2 69678 1 358
2 69679 1 358
2 69680 1 358
2 69681 1 358
2 69682 1 358
2 69683 1 358
2 69684 1 358
2 69685 1 358
2 69686 1 358
2 69687 1 358
2 69688 1 358
2 69689 1 358
2 69690 1 358
2 69691 1 358
2 69692 1 358
2 69693 1 358
2 69694 1 358
2 69695 1 358
2 69696 1 358
2 69697 1 358
2 69698 1 358
2 69699 1 358
2 69700 1 359
2 69701 1 359
2 69702 1 359
2 69703 1 359
2 69704 1 359
2 69705 1 359
2 69706 1 359
2 69707 1 360
2 69708 1 360
2 69709 1 360
2 69710 1 360
2 69711 1 360
2 69712 1 360
2 69713 1 360
2 69714 1 360
2 69715 1 360
2 69716 1 360
2 69717 1 360
2 69718 1 361
2 69719 1 361
2 69720 1 361
2 69721 1 361
2 69722 1 361
2 69723 1 361
2 69724 1 361
2 69725 1 362
2 69726 1 362
2 69727 1 362
2 69728 1 362
2 69729 1 362
2 69730 1 362
2 69731 1 362
2 69732 1 362
2 69733 1 362
2 69734 1 362
2 69735 1 362
2 69736 1 362
2 69737 1 362
2 69738 1 362
2 69739 1 362
2 69740 1 362
2 69741 1 362
2 69742 1 362
2 69743 1 362
2 69744 1 362
2 69745 1 362
2 69746 1 362
2 69747 1 362
2 69748 1 362
2 69749 1 363
2 69750 1 363
2 69751 1 363
2 69752 1 363
2 69753 1 363
2 69754 1 363
2 69755 1 363
2 69756 1 363
2 69757 1 363
2 69758 1 363
2 69759 1 363
2 69760 1 364
2 69761 1 364
2 69762 1 365
2 69763 1 365
2 69764 1 365
2 69765 1 371
2 69766 1 371
2 69767 1 371
2 69768 1 371
2 69769 1 372
2 69770 1 372
2 69771 1 372
2 69772 1 372
2 69773 1 372
2 69774 1 372
2 69775 1 372
2 69776 1 372
2 69777 1 372
2 69778 1 373
2 69779 1 373
2 69780 1 380
2 69781 1 380
2 69782 1 380
2 69783 1 380
2 69784 1 380
2 69785 1 380
2 69786 1 380
2 69787 1 380
2 69788 1 380
2 69789 1 380
2 69790 1 380
2 69791 1 380
2 69792 1 381
2 69793 1 381
2 69794 1 381
2 69795 1 381
2 69796 1 381
2 69797 1 382
2 69798 1 382
2 69799 1 382
2 69800 1 383
2 69801 1 383
2 69802 1 383
2 69803 1 383
2 69804 1 383
2 69805 1 384
2 69806 1 384
2 69807 1 385
2 69808 1 385
2 69809 1 385
2 69810 1 386
2 69811 1 386
2 69812 1 386
2 69813 1 386
2 69814 1 386
2 69815 1 386
2 69816 1 386
2 69817 1 386
2 69818 1 386
2 69819 1 386
2 69820 1 386
2 69821 1 386
2 69822 1 386
2 69823 1 386
2 69824 1 386
2 69825 1 386
2 69826 1 387
2 69827 1 387
2 69828 1 387
2 69829 1 387
2 69830 1 387
2 69831 1 388
2 69832 1 388
2 69833 1 388
2 69834 1 388
2 69835 1 388
2 69836 1 388
2 69837 1 388
2 69838 1 388
2 69839 1 388
2 69840 1 388
2 69841 1 388
2 69842 1 388
2 69843 1 388
2 69844 1 388
2 69845 1 388
2 69846 1 388
2 69847 1 388
2 69848 1 388
2 69849 1 388
2 69850 1 388
2 69851 1 388
2 69852 1 388
2 69853 1 388
2 69854 1 389
2 69855 1 389
2 69856 1 389
2 69857 1 389
2 69858 1 393
2 69859 1 393
2 69860 1 393
2 69861 1 394
2 69862 1 394
2 69863 1 399
2 69864 1 399
2 69865 1 399
2 69866 1 399
2 69867 1 399
2 69868 1 399
2 69869 1 399
2 69870 1 399
2 69871 1 399
2 69872 1 399
2 69873 1 399
2 69874 1 399
2 69875 1 399
2 69876 1 399
2 69877 1 399
2 69878 1 399
2 69879 1 399
2 69880 1 399
2 69881 1 399
2 69882 1 399
2 69883 1 400
2 69884 1 400
2 69885 1 400
2 69886 1 400
2 69887 1 400
2 69888 1 400
2 69889 1 400
2 69890 1 400
2 69891 1 400
2 69892 1 400
2 69893 1 400
2 69894 1 400
2 69895 1 401
2 69896 1 401
2 69897 1 401
2 69898 1 401
2 69899 1 401
2 69900 1 402
2 69901 1 402
2 69902 1 403
2 69903 1 403
2 69904 1 405
2 69905 1 405
2 69906 1 405
2 69907 1 405
2 69908 1 405
2 69909 1 405
2 69910 1 407
2 69911 1 407
2 69912 1 408
2 69913 1 408
2 69914 1 408
2 69915 1 408
2 69916 1 408
2 69917 1 408
2 69918 1 408
2 69919 1 408
2 69920 1 408
2 69921 1 408
2 69922 1 408
2 69923 1 408
2 69924 1 408
2 69925 1 408
2 69926 1 408
2 69927 1 408
2 69928 1 409
2 69929 1 409
2 69930 1 409
2 69931 1 409
2 69932 1 409
2 69933 1 411
2 69934 1 411
2 69935 1 421
2 69936 1 421
2 69937 1 421
2 69938 1 421
2 69939 1 421
2 69940 1 421
2 69941 1 422
2 69942 1 422
2 69943 1 422
2 69944 1 422
2 69945 1 422
2 69946 1 422
2 69947 1 424
2 69948 1 424
2 69949 1 424
2 69950 1 424
2 69951 1 424
2 69952 1 424
2 69953 1 424
2 69954 1 424
2 69955 1 424
2 69956 1 424
2 69957 1 424
2 69958 1 424
2 69959 1 424
2 69960 1 424
2 69961 1 424
2 69962 1 424
2 69963 1 424
2 69964 1 424
2 69965 1 424
2 69966 1 424
2 69967 1 424
2 69968 1 424
2 69969 1 424
2 69970 1 424
2 69971 1 424
2 69972 1 424
2 69973 1 424
2 69974 1 424
2 69975 1 425
2 69976 1 425
2 69977 1 425
2 69978 1 425
2 69979 1 425
2 69980 1 425
2 69981 1 426
2 69982 1 426
2 69983 1 426
2 69984 1 426
2 69985 1 426
2 69986 1 426
2 69987 1 426
2 69988 1 426
2 69989 1 427
2 69990 1 427
2 69991 1 429
2 69992 1 429
2 69993 1 429
2 69994 1 429
2 69995 1 429
2 69996 1 429
2 69997 1 429
2 69998 1 429
2 69999 1 429
2 70000 1 430
2 70001 1 430
2 70002 1 430
2 70003 1 430
2 70004 1 431
2 70005 1 431
2 70006 1 431
2 70007 1 431
2 70008 1 432
2 70009 1 432
2 70010 1 441
2 70011 1 441
2 70012 1 441
2 70013 1 441
2 70014 1 441
2 70015 1 442
2 70016 1 442
2 70017 1 443
2 70018 1 443
2 70019 1 443
2 70020 1 443
2 70021 1 443
2 70022 1 443
2 70023 1 443
2 70024 1 443
2 70025 1 444
2 70026 1 444
2 70027 1 444
2 70028 1 444
2 70029 1 446
2 70030 1 446
2 70031 1 449
2 70032 1 449
2 70033 1 449
2 70034 1 449
2 70035 1 450
2 70036 1 450
2 70037 1 450
2 70038 1 450
2 70039 1 450
2 70040 1 451
2 70041 1 451
2 70042 1 451
2 70043 1 457
2 70044 1 457
2 70045 1 457
2 70046 1 458
2 70047 1 458
2 70048 1 458
2 70049 1 458
2 70050 1 458
2 70051 1 467
2 70052 1 467
2 70053 1 467
2 70054 1 467
2 70055 1 467
2 70056 1 467
2 70057 1 467
2 70058 1 467
2 70059 1 467
2 70060 1 467
2 70061 1 467
2 70062 1 467
2 70063 1 468
2 70064 1 468
2 70065 1 468
2 70066 1 468
2 70067 1 468
2 70068 1 468
2 70069 1 468
2 70070 1 469
2 70071 1 469
2 70072 1 472
2 70073 1 472
2 70074 1 483
2 70075 1 483
2 70076 1 483
2 70077 1 483
2 70078 1 483
2 70079 1 483
2 70080 1 483
2 70081 1 483
2 70082 1 483
2 70083 1 483
2 70084 1 483
2 70085 1 483
2 70086 1 483
2 70087 1 484
2 70088 1 484
2 70089 1 484
2 70090 1 484
2 70091 1 484
2 70092 1 484
2 70093 1 484
2 70094 1 484
2 70095 1 484
2 70096 1 489
2 70097 1 489
2 70098 1 489
2 70099 1 489
2 70100 1 489
2 70101 1 489
2 70102 1 489
2 70103 1 489
2 70104 1 490
2 70105 1 490
2 70106 1 490
2 70107 1 490
2 70108 1 490
2 70109 1 490
2 70110 1 490
2 70111 1 490
2 70112 1 490
2 70113 1 490
2 70114 1 490
2 70115 1 490
2 70116 1 490
2 70117 1 490
2 70118 1 491
2 70119 1 491
2 70120 1 491
2 70121 1 491
2 70122 1 491
2 70123 1 492
2 70124 1 492
2 70125 1 492
2 70126 1 492
2 70127 1 494
2 70128 1 494
2 70129 1 494
2 70130 1 506
2 70131 1 506
2 70132 1 506
2 70133 1 506
2 70134 1 506
2 70135 1 506
2 70136 1 506
2 70137 1 506
2 70138 1 506
2 70139 1 506
2 70140 1 506
2 70141 1 506
2 70142 1 506
2 70143 1 506
2 70144 1 506
2 70145 1 506
2 70146 1 506
2 70147 1 506
2 70148 1 506
2 70149 1 506
2 70150 1 506
2 70151 1 506
2 70152 1 506
2 70153 1 506
2 70154 1 506
2 70155 1 506
2 70156 1 506
2 70157 1 506
2 70158 1 506
2 70159 1 506
2 70160 1 506
2 70161 1 506
2 70162 1 506
2 70163 1 506
2 70164 1 506
2 70165 1 506
2 70166 1 506
2 70167 1 506
2 70168 1 506
2 70169 1 506
2 70170 1 506
2 70171 1 506
2 70172 1 506
2 70173 1 506
2 70174 1 506
2 70175 1 506
2 70176 1 506
2 70177 1 506
2 70178 1 507
2 70179 1 507
2 70180 1 507
2 70181 1 507
2 70182 1 507
2 70183 1 507
2 70184 1 507
2 70185 1 507
2 70186 1 507
2 70187 1 507
2 70188 1 507
2 70189 1 507
2 70190 1 507
2 70191 1 507
2 70192 1 507
2 70193 1 507
2 70194 1 507
2 70195 1 507
2 70196 1 507
2 70197 1 507
2 70198 1 507
2 70199 1 507
2 70200 1 507
2 70201 1 507
2 70202 1 507
2 70203 1 507
2 70204 1 507
2 70205 1 507
2 70206 1 507
2 70207 1 507
2 70208 1 507
2 70209 1 507
2 70210 1 507
2 70211 1 507
2 70212 1 507
2 70213 1 507
2 70214 1 507
2 70215 1 507
2 70216 1 507
2 70217 1 507
2 70218 1 507
2 70219 1 507
2 70220 1 507
2 70221 1 507
2 70222 1 507
2 70223 1 507
2 70224 1 507
2 70225 1 507
2 70226 1 507
2 70227 1 507
2 70228 1 507
2 70229 1 507
2 70230 1 507
2 70231 1 507
2 70232 1 507
2 70233 1 507
2 70234 1 507
2 70235 1 507
2 70236 1 508
2 70237 1 508
2 70238 1 509
2 70239 1 509
2 70240 1 509
2 70241 1 509
2 70242 1 509
2 70243 1 510
2 70244 1 510
2 70245 1 510
2 70246 1 510
2 70247 1 510
2 70248 1 511
2 70249 1 511
2 70250 1 511
2 70251 1 511
2 70252 1 511
2 70253 1 511
2 70254 1 511
2 70255 1 511
2 70256 1 511
2 70257 1 511
2 70258 1 511
2 70259 1 511
2 70260 1 511
2 70261 1 511
2 70262 1 511
2 70263 1 511
2 70264 1 511
2 70265 1 512
2 70266 1 512
2 70267 1 512
2 70268 1 520
2 70269 1 520
2 70270 1 520
2 70271 1 520
2 70272 1 520
2 70273 1 520
2 70274 1 520
2 70275 1 520
2 70276 1 520
2 70277 1 520
2 70278 1 520
2 70279 1 520
2 70280 1 520
2 70281 1 520
2 70282 1 520
2 70283 1 520
2 70284 1 520
2 70285 1 520
2 70286 1 520
2 70287 1 520
2 70288 1 520
2 70289 1 520
2 70290 1 520
2 70291 1 520
2 70292 1 520
2 70293 1 520
2 70294 1 520
2 70295 1 520
2 70296 1 520
2 70297 1 520
2 70298 1 520
2 70299 1 520
2 70300 1 520
2 70301 1 520
2 70302 1 520
2 70303 1 520
2 70304 1 520
2 70305 1 520
2 70306 1 520
2 70307 1 520
2 70308 1 520
2 70309 1 520
2 70310 1 520
2 70311 1 521
2 70312 1 521
2 70313 1 521
2 70314 1 521
2 70315 1 521
2 70316 1 521
2 70317 1 521
2 70318 1 521
2 70319 1 521
2 70320 1 521
2 70321 1 521
2 70322 1 521
2 70323 1 521
2 70324 1 521
2 70325 1 521
2 70326 1 521
2 70327 1 521
2 70328 1 521
2 70329 1 521
2 70330 1 521
2 70331 1 521
2 70332 1 521
2 70333 1 521
2 70334 1 521
2 70335 1 521
2 70336 1 521
2 70337 1 522
2 70338 1 522
2 70339 1 524
2 70340 1 524
2 70341 1 524
2 70342 1 524
2 70343 1 524
2 70344 1 524
2 70345 1 524
2 70346 1 524
2 70347 1 524
2 70348 1 524
2 70349 1 524
2 70350 1 524
2 70351 1 524
2 70352 1 524
2 70353 1 524
2 70354 1 524
2 70355 1 524
2 70356 1 525
2 70357 1 525
2 70358 1 525
2 70359 1 525
2 70360 1 526
2 70361 1 526
2 70362 1 526
2 70363 1 526
2 70364 1 526
2 70365 1 534
2 70366 1 534
2 70367 1 534
2 70368 1 534
2 70369 1 534
2 70370 1 534
2 70371 1 534
2 70372 1 534
2 70373 1 534
2 70374 1 534
2 70375 1 534
2 70376 1 534
2 70377 1 534
2 70378 1 534
2 70379 1 535
2 70380 1 535
2 70381 1 535
2 70382 1 535
2 70383 1 535
2 70384 1 535
2 70385 1 535
2 70386 1 535
2 70387 1 535
2 70388 1 535
2 70389 1 535
2 70390 1 535
2 70391 1 535
2 70392 1 535
2 70393 1 535
2 70394 1 535
2 70395 1 535
2 70396 1 535
2 70397 1 535
2 70398 1 535
2 70399 1 535
2 70400 1 535
2 70401 1 535
2 70402 1 535
2 70403 1 535
2 70404 1 535
2 70405 1 535
2 70406 1 535
2 70407 1 535
2 70408 1 535
2 70409 1 535
2 70410 1 535
2 70411 1 535
2 70412 1 535
2 70413 1 535
2 70414 1 535
2 70415 1 535
2 70416 1 535
2 70417 1 535
2 70418 1 535
2 70419 1 535
2 70420 1 535
2 70421 1 535
2 70422 1 535
2 70423 1 535
2 70424 1 535
2 70425 1 535
2 70426 1 535
2 70427 1 535
2 70428 1 535
2 70429 1 535
2 70430 1 535
2 70431 1 535
2 70432 1 535
2 70433 1 535
2 70434 1 535
2 70435 1 535
2 70436 1 535
2 70437 1 535
2 70438 1 535
2 70439 1 535
2 70440 1 535
2 70441 1 536
2 70442 1 536
2 70443 1 536
2 70444 1 537
2 70445 1 537
2 70446 1 538
2 70447 1 538
2 70448 1 547
2 70449 1 547
2 70450 1 547
2 70451 1 547
2 70452 1 547
2 70453 1 547
2 70454 1 547
2 70455 1 547
2 70456 1 547
2 70457 1 547
2 70458 1 547
2 70459 1 547
2 70460 1 549
2 70461 1 549
2 70462 1 549
2 70463 1 549
2 70464 1 551
2 70465 1 551
2 70466 1 552
2 70467 1 552
2 70468 1 552
2 70469 1 552
2 70470 1 552
2 70471 1 552
2 70472 1 552
2 70473 1 552
2 70474 1 552
2 70475 1 552
2 70476 1 552
2 70477 1 552
2 70478 1 552
2 70479 1 552
2 70480 1 552
2 70481 1 552
2 70482 1 552
2 70483 1 552
2 70484 1 552
2 70485 1 552
2 70486 1 552
2 70487 1 552
2 70488 1 552
2 70489 1 552
2 70490 1 552
2 70491 1 552
2 70492 1 552
2 70493 1 552
2 70494 1 552
2 70495 1 552
2 70496 1 552
2 70497 1 552
2 70498 1 552
2 70499 1 552
2 70500 1 552
2 70501 1 552
2 70502 1 552
2 70503 1 552
2 70504 1 552
2 70505 1 552
2 70506 1 552
2 70507 1 552
2 70508 1 552
2 70509 1 552
2 70510 1 552
2 70511 1 552
2 70512 1 552
2 70513 1 552
2 70514 1 552
2 70515 1 552
2 70516 1 552
2 70517 1 552
2 70518 1 552
2 70519 1 552
2 70520 1 552
2 70521 1 552
2 70522 1 552
2 70523 1 552
2 70524 1 552
2 70525 1 552
2 70526 1 552
2 70527 1 552
2 70528 1 552
2 70529 1 552
2 70530 1 552
2 70531 1 552
2 70532 1 552
2 70533 1 552
2 70534 1 552
2 70535 1 552
2 70536 1 552
2 70537 1 552
2 70538 1 552
2 70539 1 552
2 70540 1 552
2 70541 1 552
2 70542 1 552
2 70543 1 552
2 70544 1 552
2 70545 1 553
2 70546 1 553
2 70547 1 553
2 70548 1 553
2 70549 1 553
2 70550 1 554
2 70551 1 554
2 70552 1 554
2 70553 1 554
2 70554 1 554
2 70555 1 554
2 70556 1 554
2 70557 1 554
2 70558 1 554
2 70559 1 554
2 70560 1 554
2 70561 1 554
2 70562 1 557
2 70563 1 557
2 70564 1 557
2 70565 1 557
2 70566 1 557
2 70567 1 557
2 70568 1 557
2 70569 1 557
2 70570 1 557
2 70571 1 557
2 70572 1 557
2 70573 1 557
2 70574 1 557
2 70575 1 557
2 70576 1 557
2 70577 1 557
2 70578 1 557
2 70579 1 557
2 70580 1 557
2 70581 1 557
2 70582 1 557
2 70583 1 558
2 70584 1 558
2 70585 1 558
2 70586 1 558
2 70587 1 558
2 70588 1 558
2 70589 1 558
2 70590 1 558
2 70591 1 558
2 70592 1 559
2 70593 1 559
2 70594 1 559
2 70595 1 559
2 70596 1 559
2 70597 1 559
2 70598 1 559
2 70599 1 559
2 70600 1 559
2 70601 1 559
2 70602 1 559
2 70603 1 559
2 70604 1 559
2 70605 1 559
2 70606 1 559
2 70607 1 559
2 70608 1 559
2 70609 1 559
2 70610 1 559
2 70611 1 559
2 70612 1 559
2 70613 1 559
2 70614 1 559
2 70615 1 559
2 70616 1 559
2 70617 1 559
2 70618 1 559
2 70619 1 559
2 70620 1 559
2 70621 1 559
2 70622 1 559
2 70623 1 559
2 70624 1 559
2 70625 1 559
2 70626 1 559
2 70627 1 559
2 70628 1 559
2 70629 1 559
2 70630 1 559
2 70631 1 559
2 70632 1 559
2 70633 1 559
2 70634 1 559
2 70635 1 559
2 70636 1 559
2 70637 1 559
2 70638 1 559
2 70639 1 559
2 70640 1 559
2 70641 1 559
2 70642 1 559
2 70643 1 559
2 70644 1 559
2 70645 1 559
2 70646 1 559
2 70647 1 559
2 70648 1 559
2 70649 1 559
2 70650 1 559
2 70651 1 559
2 70652 1 560
2 70653 1 560
2 70654 1 560
2 70655 1 560
2 70656 1 560
2 70657 1 560
2 70658 1 560
2 70659 1 560
2 70660 1 561
2 70661 1 561
2 70662 1 561
2 70663 1 562
2 70664 1 562
2 70665 1 562
2 70666 1 562
2 70667 1 562
2 70668 1 562
2 70669 1 562
2 70670 1 562
2 70671 1 562
2 70672 1 562
2 70673 1 562
2 70674 1 562
2 70675 1 562
2 70676 1 562
2 70677 1 562
2 70678 1 563
2 70679 1 563
2 70680 1 563
2 70681 1 563
2 70682 1 564
2 70683 1 564
2 70684 1 564
2 70685 1 564
2 70686 1 564
2 70687 1 564
2 70688 1 564
2 70689 1 564
2 70690 1 566
2 70691 1 566
2 70692 1 566
2 70693 1 571
2 70694 1 571
2 70695 1 571
2 70696 1 571
2 70697 1 571
2 70698 1 571
2 70699 1 571
2 70700 1 571
2 70701 1 571
2 70702 1 571
2 70703 1 572
2 70704 1 572
2 70705 1 572
2 70706 1 572
2 70707 1 572
2 70708 1 572
2 70709 1 572
2 70710 1 573
2 70711 1 573
2 70712 1 573
2 70713 1 574
2 70714 1 574
2 70715 1 577
2 70716 1 577
2 70717 1 577
2 70718 1 577
2 70719 1 577
2 70720 1 577
2 70721 1 577
2 70722 1 577
2 70723 1 578
2 70724 1 578
2 70725 1 578
2 70726 1 579
2 70727 1 579
2 70728 1 588
2 70729 1 588
2 70730 1 588
2 70731 1 589
2 70732 1 589
2 70733 1 589
2 70734 1 589
2 70735 1 589
2 70736 1 589
2 70737 1 589
2 70738 1 589
2 70739 1 589
2 70740 1 589
2 70741 1 591
2 70742 1 591
2 70743 1 594
2 70744 1 594
2 70745 1 594
2 70746 1 594
2 70747 1 595
2 70748 1 595
2 70749 1 595
2 70750 1 595
2 70751 1 595
2 70752 1 595
2 70753 1 595
2 70754 1 595
2 70755 1 595
2 70756 1 595
2 70757 1 595
2 70758 1 595
2 70759 1 595
2 70760 1 595
2 70761 1 595
2 70762 1 595
2 70763 1 595
2 70764 1 595
2 70765 1 595
2 70766 1 595
2 70767 1 595
2 70768 1 595
2 70769 1 595
2 70770 1 595
2 70771 1 595
2 70772 1 595
2 70773 1 595
2 70774 1 595
2 70775 1 595
2 70776 1 595
2 70777 1 595
2 70778 1 595
2 70779 1 595
2 70780 1 595
2 70781 1 595
2 70782 1 595
2 70783 1 595
2 70784 1 595
2 70785 1 595
2 70786 1 595
2 70787 1 595
2 70788 1 595
2 70789 1 595
2 70790 1 595
2 70791 1 595
2 70792 1 595
2 70793 1 595
2 70794 1 595
2 70795 1 595
2 70796 1 595
2 70797 1 595
2 70798 1 595
2 70799 1 595
2 70800 1 595
2 70801 1 595
2 70802 1 596
2 70803 1 596
2 70804 1 596
2 70805 1 596
2 70806 1 596
2 70807 1 596
2 70808 1 596
2 70809 1 596
2 70810 1 596
2 70811 1 596
2 70812 1 596
2 70813 1 596
2 70814 1 596
2 70815 1 596
2 70816 1 596
2 70817 1 596
2 70818 1 596
2 70819 1 596
2 70820 1 596
2 70821 1 596
2 70822 1 596
2 70823 1 596
2 70824 1 596
2 70825 1 596
2 70826 1 596
2 70827 1 596
2 70828 1 596
2 70829 1 596
2 70830 1 596
2 70831 1 596
2 70832 1 596
2 70833 1 596
2 70834 1 596
2 70835 1 596
2 70836 1 596
2 70837 1 596
2 70838 1 596
2 70839 1 596
2 70840 1 596
2 70841 1 596
2 70842 1 596
2 70843 1 596
2 70844 1 596
2 70845 1 596
2 70846 1 596
2 70847 1 596
2 70848 1 596
2 70849 1 596
2 70850 1 596
2 70851 1 596
2 70852 1 596
2 70853 1 596
2 70854 1 596
2 70855 1 596
2 70856 1 596
2 70857 1 598
2 70858 1 598
2 70859 1 599
2 70860 1 599
2 70861 1 603
2 70862 1 603
2 70863 1 606
2 70864 1 606
2 70865 1 606
2 70866 1 606
2 70867 1 606
2 70868 1 606
2 70869 1 606
2 70870 1 606
2 70871 1 606
2 70872 1 606
2 70873 1 606
2 70874 1 606
2 70875 1 606
2 70876 1 606
2 70877 1 606
2 70878 1 606
2 70879 1 606
2 70880 1 606
2 70881 1 607
2 70882 1 607
2 70883 1 607
2 70884 1 607
2 70885 1 609
2 70886 1 609
2 70887 1 609
2 70888 1 610
2 70889 1 610
2 70890 1 610
2 70891 1 611
2 70892 1 611
2 70893 1 621
2 70894 1 621
2 70895 1 621
2 70896 1 622
2 70897 1 622
2 70898 1 625
2 70899 1 625
2 70900 1 625
2 70901 1 625
2 70902 1 625
2 70903 1 625
2 70904 1 625
2 70905 1 625
2 70906 1 625
2 70907 1 625
2 70908 1 625
2 70909 1 626
2 70910 1 626
2 70911 1 626
2 70912 1 626
2 70913 1 626
2 70914 1 627
2 70915 1 627
2 70916 1 627
2 70917 1 627
2 70918 1 627
2 70919 1 627
2 70920 1 627
2 70921 1 627
2 70922 1 627
2 70923 1 627
2 70924 1 627
2 70925 1 627
2 70926 1 627
2 70927 1 627
2 70928 1 627
2 70929 1 627
2 70930 1 627
2 70931 1 628
2 70932 1 628
2 70933 1 628
2 70934 1 628
2 70935 1 628
2 70936 1 628
2 70937 1 628
2 70938 1 628
2 70939 1 628
2 70940 1 628
2 70941 1 630
2 70942 1 630
2 70943 1 630
2 70944 1 646
2 70945 1 646
2 70946 1 646
2 70947 1 646
2 70948 1 646
2 70949 1 646
2 70950 1 646
2 70951 1 646
2 70952 1 646
2 70953 1 646
2 70954 1 647
2 70955 1 647
2 70956 1 647
2 70957 1 647
2 70958 1 647
2 70959 1 647
2 70960 1 647
2 70961 1 647
2 70962 1 647
2 70963 1 647
2 70964 1 647
2 70965 1 647
2 70966 1 647
2 70967 1 647
2 70968 1 647
2 70969 1 647
2 70970 1 647
2 70971 1 647
2 70972 1 647
2 70973 1 647
2 70974 1 647
2 70975 1 648
2 70976 1 648
2 70977 1 649
2 70978 1 649
2 70979 1 650
2 70980 1 650
2 70981 1 651
2 70982 1 651
2 70983 1 651
2 70984 1 651
2 70985 1 651
2 70986 1 653
2 70987 1 653
2 70988 1 655
2 70989 1 655
2 70990 1 657
2 70991 1 657
2 70992 1 658
2 70993 1 658
2 70994 1 658
2 70995 1 660
2 70996 1 660
2 70997 1 660
2 70998 1 660
2 70999 1 662
2 71000 1 662
2 71001 1 663
2 71002 1 663
2 71003 1 663
2 71004 1 663
2 71005 1 663
2 71006 1 663
2 71007 1 663
2 71008 1 663
2 71009 1 663
2 71010 1 664
2 71011 1 664
2 71012 1 667
2 71013 1 667
2 71014 1 672
2 71015 1 672
2 71016 1 673
2 71017 1 673
2 71018 1 674
2 71019 1 674
2 71020 1 675
2 71021 1 675
2 71022 1 675
2 71023 1 675
2 71024 1 675
2 71025 1 675
2 71026 1 675
2 71027 1 675
2 71028 1 675
2 71029 1 675
2 71030 1 675
2 71031 1 675
2 71032 1 675
2 71033 1 676
2 71034 1 676
2 71035 1 676
2 71036 1 676
2 71037 1 676
2 71038 1 676
2 71039 1 676
2 71040 1 676
2 71041 1 676
2 71042 1 676
2 71043 1 677
2 71044 1 677
2 71045 1 680
2 71046 1 680
2 71047 1 680
2 71048 1 686
2 71049 1 686
2 71050 1 693
2 71051 1 693
2 71052 1 693
2 71053 1 693
2 71054 1 693
2 71055 1 693
2 71056 1 693
2 71057 1 693
2 71058 1 693
2 71059 1 693
2 71060 1 693
2 71061 1 693
2 71062 1 693
2 71063 1 694
2 71064 1 694
2 71065 1 694
2 71066 1 694
2 71067 1 694
2 71068 1 695
2 71069 1 695
2 71070 1 695
2 71071 1 695
2 71072 1 695
2 71073 1 695
2 71074 1 695
2 71075 1 695
2 71076 1 695
2 71077 1 695
2 71078 1 695
2 71079 1 695
2 71080 1 695
2 71081 1 695
2 71082 1 695
2 71083 1 695
2 71084 1 695
2 71085 1 695
2 71086 1 695
2 71087 1 696
2 71088 1 696
2 71089 1 699
2 71090 1 699
2 71091 1 699
2 71092 1 700
2 71093 1 700
2 71094 1 700
2 71095 1 702
2 71096 1 702
2 71097 1 705
2 71098 1 705
2 71099 1 705
2 71100 1 706
2 71101 1 706
2 71102 1 706
2 71103 1 706
2 71104 1 706
2 71105 1 707
2 71106 1 707
2 71107 1 708
2 71108 1 708
2 71109 1 708
2 71110 1 708
2 71111 1 708
2 71112 1 708
2 71113 1 709
2 71114 1 709
2 71115 1 709
2 71116 1 709
2 71117 1 710
2 71118 1 710
2 71119 1 728
2 71120 1 728
2 71121 1 728
2 71122 1 728
2 71123 1 728
2 71124 1 728
2 71125 1 729
2 71126 1 729
2 71127 1 729
2 71128 1 730
2 71129 1 730
2 71130 1 731
2 71131 1 731
2 71132 1 731
2 71133 1 731
2 71134 1 731
2 71135 1 731
2 71136 1 733
2 71137 1 733
2 71138 1 741
2 71139 1 741
2 71140 1 741
2 71141 1 741
2 71142 1 741
2 71143 1 741
2 71144 1 741
2 71145 1 741
2 71146 1 741
2 71147 1 741
2 71148 1 741
2 71149 1 741
2 71150 1 741
2 71151 1 741
2 71152 1 741
2 71153 1 741
2 71154 1 741
2 71155 1 741
2 71156 1 741
2 71157 1 741
2 71158 1 741
2 71159 1 741
2 71160 1 741
2 71161 1 741
2 71162 1 741
2 71163 1 741
2 71164 1 741
2 71165 1 741
2 71166 1 741
2 71167 1 741
2 71168 1 741
2 71169 1 741
2 71170 1 741
2 71171 1 741
2 71172 1 741
2 71173 1 741
2 71174 1 741
2 71175 1 741
2 71176 1 741
2 71177 1 741
2 71178 1 741
2 71179 1 741
2 71180 1 741
2 71181 1 741
2 71182 1 741
2 71183 1 741
2 71184 1 741
2 71185 1 741
2 71186 1 741
2 71187 1 741
2 71188 1 741
2 71189 1 741
2 71190 1 741
2 71191 1 741
2 71192 1 741
2 71193 1 741
2 71194 1 741
2 71195 1 741
2 71196 1 741
2 71197 1 741
2 71198 1 741
2 71199 1 741
2 71200 1 741
2 71201 1 741
2 71202 1 741
2 71203 1 741
2 71204 1 741
2 71205 1 741
2 71206 1 741
2 71207 1 741
2 71208 1 741
2 71209 1 741
2 71210 1 741
2 71211 1 741
2 71212 1 741
2 71213 1 741
2 71214 1 741
2 71215 1 741
2 71216 1 741
2 71217 1 741
2 71218 1 741
2 71219 1 741
2 71220 1 741
2 71221 1 741
2 71222 1 741
2 71223 1 741
2 71224 1 741
2 71225 1 741
2 71226 1 741
2 71227 1 741
2 71228 1 741
2 71229 1 741
2 71230 1 741
2 71231 1 741
2 71232 1 741
2 71233 1 741
2 71234 1 741
2 71235 1 741
2 71236 1 741
2 71237 1 741
2 71238 1 742
2 71239 1 742
2 71240 1 742
2 71241 1 742
2 71242 1 742
2 71243 1 742
2 71244 1 742
2 71245 1 742
2 71246 1 742
2 71247 1 742
2 71248 1 742
2 71249 1 742
2 71250 1 742
2 71251 1 742
2 71252 1 742
2 71253 1 742
2 71254 1 742
2 71255 1 742
2 71256 1 742
2 71257 1 742
2 71258 1 742
2 71259 1 742
2 71260 1 742
2 71261 1 742
2 71262 1 742
2 71263 1 742
2 71264 1 742
2 71265 1 742
2 71266 1 742
2 71267 1 742
2 71268 1 742
2 71269 1 742
2 71270 1 742
2 71271 1 742
2 71272 1 742
2 71273 1 742
2 71274 1 742
2 71275 1 742
2 71276 1 742
2 71277 1 742
2 71278 1 742
2 71279 1 742
2 71280 1 742
2 71281 1 742
2 71282 1 742
2 71283 1 742
2 71284 1 742
2 71285 1 742
2 71286 1 742
2 71287 1 742
2 71288 1 742
2 71289 1 742
2 71290 1 742
2 71291 1 742
2 71292 1 742
2 71293 1 742
2 71294 1 742
2 71295 1 742
2 71296 1 742
2 71297 1 742
2 71298 1 742
2 71299 1 742
2 71300 1 742
2 71301 1 742
2 71302 1 742
2 71303 1 742
2 71304 1 742
2 71305 1 742
2 71306 1 742
2 71307 1 742
2 71308 1 742
2 71309 1 742
2 71310 1 742
2 71311 1 742
2 71312 1 742
2 71313 1 742
2 71314 1 742
2 71315 1 742
2 71316 1 742
2 71317 1 742
2 71318 1 742
2 71319 1 742
2 71320 1 742
2 71321 1 742
2 71322 1 742
2 71323 1 742
2 71324 1 742
2 71325 1 742
2 71326 1 742
2 71327 1 742
2 71328 1 742
2 71329 1 742
2 71330 1 742
2 71331 1 742
2 71332 1 742
2 71333 1 742
2 71334 1 742
2 71335 1 742
2 71336 1 742
2 71337 1 742
2 71338 1 742
2 71339 1 742
2 71340 1 742
2 71341 1 742
2 71342 1 749
2 71343 1 749
2 71344 1 749
2 71345 1 749
2 71346 1 751
2 71347 1 751
2 71348 1 751
2 71349 1 751
2 71350 1 751
2 71351 1 751
2 71352 1 751
2 71353 1 752
2 71354 1 752
2 71355 1 752
2 71356 1 752
2 71357 1 752
2 71358 1 752
2 71359 1 752
2 71360 1 752
2 71361 1 752
2 71362 1 752
2 71363 1 752
2 71364 1 752
2 71365 1 752
2 71366 1 760
2 71367 1 760
2 71368 1 760
2 71369 1 761
2 71370 1 761
2 71371 1 761
2 71372 1 761
2 71373 1 761
2 71374 1 761
2 71375 1 761
2 71376 1 761
2 71377 1 761
2 71378 1 762
2 71379 1 762
2 71380 1 777
2 71381 1 777
2 71382 1 777
2 71383 1 777
2 71384 1 777
2 71385 1 777
2 71386 1 777
2 71387 1 777
2 71388 1 777
2 71389 1 777
2 71390 1 777
2 71391 1 777
2 71392 1 777
2 71393 1 777
2 71394 1 777
2 71395 1 777
2 71396 1 777
2 71397 1 777
2 71398 1 777
2 71399 1 777
2 71400 1 777
2 71401 1 777
2 71402 1 777
2 71403 1 777
2 71404 1 777
2 71405 1 777
2 71406 1 777
2 71407 1 777
2 71408 1 777
2 71409 1 777
2 71410 1 777
2 71411 1 777
2 71412 1 777
2 71413 1 777
2 71414 1 777
2 71415 1 777
2 71416 1 777
2 71417 1 777
2 71418 1 777
2 71419 1 777
2 71420 1 777
2 71421 1 777
2 71422 1 777
2 71423 1 777
2 71424 1 777
2 71425 1 777
2 71426 1 777
2 71427 1 777
2 71428 1 777
2 71429 1 777
2 71430 1 777
2 71431 1 777
2 71432 1 777
2 71433 1 777
2 71434 1 777
2 71435 1 777
2 71436 1 777
2 71437 1 777
2 71438 1 777
2 71439 1 777
2 71440 1 777
2 71441 1 777
2 71442 1 777
2 71443 1 777
2 71444 1 777
2 71445 1 777
2 71446 1 777
2 71447 1 777
2 71448 1 777
2 71449 1 777
2 71450 1 777
2 71451 1 777
2 71452 1 777
2 71453 1 777
2 71454 1 777
2 71455 1 777
2 71456 1 777
2 71457 1 778
2 71458 1 778
2 71459 1 778
2 71460 1 778
2 71461 1 778
2 71462 1 778
2 71463 1 778
2 71464 1 778
2 71465 1 778
2 71466 1 778
2 71467 1 778
2 71468 1 778
2 71469 1 778
2 71470 1 778
2 71471 1 778
2 71472 1 778
2 71473 1 778
2 71474 1 778
2 71475 1 778
2 71476 1 778
2 71477 1 778
2 71478 1 778
2 71479 1 778
2 71480 1 778
2 71481 1 778
2 71482 1 778
2 71483 1 778
2 71484 1 778
2 71485 1 778
2 71486 1 778
2 71487 1 778
2 71488 1 778
2 71489 1 778
2 71490 1 778
2 71491 1 778
2 71492 1 778
2 71493 1 778
2 71494 1 778
2 71495 1 778
2 71496 1 778
2 71497 1 778
2 71498 1 778
2 71499 1 778
2 71500 1 778
2 71501 1 778
2 71502 1 778
2 71503 1 778
2 71504 1 778
2 71505 1 778
2 71506 1 778
2 71507 1 778
2 71508 1 778
2 71509 1 778
2 71510 1 778
2 71511 1 778
2 71512 1 778
2 71513 1 778
2 71514 1 778
2 71515 1 778
2 71516 1 778
2 71517 1 778
2 71518 1 778
2 71519 1 778
2 71520 1 778
2 71521 1 778
2 71522 1 778
2 71523 1 778
2 71524 1 778
2 71525 1 778
2 71526 1 778
2 71527 1 778
2 71528 1 778
2 71529 1 778
2 71530 1 778
2 71531 1 778
2 71532 1 778
2 71533 1 778
2 71534 1 778
2 71535 1 778
2 71536 1 778
2 71537 1 778
2 71538 1 778
2 71539 1 778
2 71540 1 778
2 71541 1 778
2 71542 1 778
2 71543 1 778
2 71544 1 778
2 71545 1 778
2 71546 1 778
2 71547 1 778
2 71548 1 778
2 71549 1 778
2 71550 1 778
2 71551 1 778
2 71552 1 778
2 71553 1 778
2 71554 1 778
2 71555 1 778
2 71556 1 778
2 71557 1 778
2 71558 1 778
2 71559 1 778
2 71560 1 778
2 71561 1 778
2 71562 1 778
2 71563 1 778
2 71564 1 778
2 71565 1 778
2 71566 1 778
2 71567 1 778
2 71568 1 778
2 71569 1 778
2 71570 1 778
2 71571 1 778
2 71572 1 779
2 71573 1 779
2 71574 1 779
2 71575 1 792
2 71576 1 792
2 71577 1 792
2 71578 1 792
2 71579 1 792
2 71580 1 792
2 71581 1 792
2 71582 1 792
2 71583 1 792
2 71584 1 792
2 71585 1 792
2 71586 1 792
2 71587 1 792
2 71588 1 792
2 71589 1 792
2 71590 1 792
2 71591 1 792
2 71592 1 793
2 71593 1 793
2 71594 1 793
2 71595 1 793
2 71596 1 793
2 71597 1 793
2 71598 1 793
2 71599 1 793
2 71600 1 793
2 71601 1 793
2 71602 1 796
2 71603 1 796
2 71604 1 796
2 71605 1 796
2 71606 1 796
2 71607 1 796
2 71608 1 798
2 71609 1 798
2 71610 1 798
2 71611 1 800
2 71612 1 800
2 71613 1 800
2 71614 1 800
2 71615 1 800
2 71616 1 800
2 71617 1 801
2 71618 1 801
2 71619 1 801
2 71620 1 801
2 71621 1 801
2 71622 1 801
2 71623 1 801
2 71624 1 801
2 71625 1 801
2 71626 1 801
2 71627 1 801
2 71628 1 801
2 71629 1 801
2 71630 1 802
2 71631 1 802
2 71632 1 802
2 71633 1 802
2 71634 1 804
2 71635 1 804
2 71636 1 805
2 71637 1 805
2 71638 1 805
2 71639 1 805
2 71640 1 806
2 71641 1 806
2 71642 1 806
2 71643 1 806
2 71644 1 807
2 71645 1 807
2 71646 1 807
2 71647 1 807
2 71648 1 807
2 71649 1 807
2 71650 1 808
2 71651 1 808
2 71652 1 809
2 71653 1 809
2 71654 1 809
2 71655 1 809
2 71656 1 809
2 71657 1 810
2 71658 1 810
2 71659 1 810
2 71660 1 811
2 71661 1 811
2 71662 1 811
2 71663 1 811
2 71664 1 811
2 71665 1 811
2 71666 1 811
2 71667 1 812
2 71668 1 812
2 71669 1 815
2 71670 1 815
2 71671 1 815
2 71672 1 815
2 71673 1 815
2 71674 1 815
2 71675 1 815
2 71676 1 815
2 71677 1 815
2 71678 1 815
2 71679 1 815
2 71680 1 815
2 71681 1 815
2 71682 1 815
2 71683 1 815
2 71684 1 815
2 71685 1 815
2 71686 1 815
2 71687 1 815
2 71688 1 815
2 71689 1 815
2 71690 1 815
2 71691 1 815
2 71692 1 815
2 71693 1 815
2 71694 1 815
2 71695 1 815
2 71696 1 815
2 71697 1 815
2 71698 1 815
2 71699 1 815
2 71700 1 815
2 71701 1 816
2 71702 1 816
2 71703 1 816
2 71704 1 816
2 71705 1 816
2 71706 1 816
2 71707 1 816
2 71708 1 816
2 71709 1 816
2 71710 1 816
2 71711 1 816
2 71712 1 816
2 71713 1 816
2 71714 1 816
2 71715 1 816
2 71716 1 816
2 71717 1 816
2 71718 1 816
2 71719 1 816
2 71720 1 816
2 71721 1 816
2 71722 1 816
2 71723 1 816
2 71724 1 816
2 71725 1 816
2 71726 1 816
2 71727 1 816
2 71728 1 816
2 71729 1 816
2 71730 1 816
2 71731 1 816
2 71732 1 816
2 71733 1 816
2 71734 1 816
2 71735 1 816
2 71736 1 816
2 71737 1 816
2 71738 1 816
2 71739 1 816
2 71740 1 816
2 71741 1 816
2 71742 1 816
2 71743 1 816
2 71744 1 816
2 71745 1 816
2 71746 1 816
2 71747 1 816
2 71748 1 816
2 71749 1 816
2 71750 1 816
2 71751 1 816
2 71752 1 816
2 71753 1 816
2 71754 1 816
2 71755 1 816
2 71756 1 816
2 71757 1 816
2 71758 1 816
2 71759 1 816
2 71760 1 816
2 71761 1 816
2 71762 1 816
2 71763 1 816
2 71764 1 816
2 71765 1 816
2 71766 1 816
2 71767 1 816
2 71768 1 817
2 71769 1 817
2 71770 1 817
2 71771 1 817
2 71772 1 817
2 71773 1 818
2 71774 1 818
2 71775 1 818
2 71776 1 818
2 71777 1 818
2 71778 1 819
2 71779 1 819
2 71780 1 819
2 71781 1 819
2 71782 1 819
2 71783 1 819
2 71784 1 819
2 71785 1 819
2 71786 1 830
2 71787 1 830
2 71788 1 830
2 71789 1 830
2 71790 1 830
2 71791 1 830
2 71792 1 830
2 71793 1 830
2 71794 1 830
2 71795 1 830
2 71796 1 830
2 71797 1 830
2 71798 1 830
2 71799 1 830
2 71800 1 830
2 71801 1 830
2 71802 1 830
2 71803 1 830
2 71804 1 830
2 71805 1 830
2 71806 1 830
2 71807 1 830
2 71808 1 830
2 71809 1 830
2 71810 1 830
2 71811 1 830
2 71812 1 830
2 71813 1 830
2 71814 1 830
2 71815 1 830
2 71816 1 830
2 71817 1 830
2 71818 1 830
2 71819 1 830
2 71820 1 830
2 71821 1 830
2 71822 1 830
2 71823 1 830
2 71824 1 830
2 71825 1 830
2 71826 1 830
2 71827 1 830
2 71828 1 830
2 71829 1 830
2 71830 1 830
2 71831 1 830
2 71832 1 830
2 71833 1 830
2 71834 1 830
2 71835 1 830
2 71836 1 830
2 71837 1 830
2 71838 1 830
2 71839 1 831
2 71840 1 831
2 71841 1 831
2 71842 1 831
2 71843 1 831
2 71844 1 831
2 71845 1 831
2 71846 1 831
2 71847 1 831
2 71848 1 831
2 71849 1 831
2 71850 1 831
2 71851 1 831
2 71852 1 831
2 71853 1 831
2 71854 1 831
2 71855 1 831
2 71856 1 831
2 71857 1 831
2 71858 1 831
2 71859 1 831
2 71860 1 831
2 71861 1 831
2 71862 1 831
2 71863 1 831
2 71864 1 831
2 71865 1 831
2 71866 1 831
2 71867 1 831
2 71868 1 831
2 71869 1 831
2 71870 1 831
2 71871 1 831
2 71872 1 831
2 71873 1 831
2 71874 1 831
2 71875 1 831
2 71876 1 831
2 71877 1 831
2 71878 1 831
2 71879 1 831
2 71880 1 831
2 71881 1 831
2 71882 1 831
2 71883 1 831
2 71884 1 831
2 71885 1 831
2 71886 1 831
2 71887 1 831
2 71888 1 831
2 71889 1 831
2 71890 1 831
2 71891 1 831
2 71892 1 831
2 71893 1 831
2 71894 1 831
2 71895 1 831
2 71896 1 831
2 71897 1 831
2 71898 1 831
2 71899 1 831
2 71900 1 831
2 71901 1 831
2 71902 1 831
2 71903 1 831
2 71904 1 831
2 71905 1 831
2 71906 1 831
2 71907 1 831
2 71908 1 831
2 71909 1 831
2 71910 1 831
2 71911 1 831
2 71912 1 831
2 71913 1 831
2 71914 1 831
2 71915 1 831
2 71916 1 831
2 71917 1 831
2 71918 1 831
2 71919 1 831
2 71920 1 831
2 71921 1 831
2 71922 1 831
2 71923 1 831
2 71924 1 831
2 71925 1 831
2 71926 1 831
2 71927 1 831
2 71928 1 831
2 71929 1 831
2 71930 1 831
2 71931 1 831
2 71932 1 831
2 71933 1 831
2 71934 1 831
2 71935 1 831
2 71936 1 831
2 71937 1 832
2 71938 1 832
2 71939 1 833
2 71940 1 833
2 71941 1 835
2 71942 1 835
2 71943 1 838
2 71944 1 838
2 71945 1 838
2 71946 1 838
2 71947 1 838
2 71948 1 838
2 71949 1 838
2 71950 1 838
2 71951 1 838
2 71952 1 838
2 71953 1 838
2 71954 1 838
2 71955 1 838
2 71956 1 845
2 71957 1 845
2 71958 1 845
2 71959 1 845
2 71960 1 845
2 71961 1 845
2 71962 1 849
2 71963 1 849
2 71964 1 849
2 71965 1 849
2 71966 1 849
2 71967 1 849
2 71968 1 857
2 71969 1 857
2 71970 1 857
2 71971 1 858
2 71972 1 858
2 71973 1 858
2 71974 1 858
2 71975 1 860
2 71976 1 860
2 71977 1 864
2 71978 1 864
2 71979 1 864
2 71980 1 864
2 71981 1 878
2 71982 1 878
2 71983 1 878
2 71984 1 878
2 71985 1 878
2 71986 1 878
2 71987 1 878
2 71988 1 878
2 71989 1 878
2 71990 1 878
2 71991 1 878
2 71992 1 878
2 71993 1 878
2 71994 1 878
2 71995 1 878
2 71996 1 878
2 71997 1 878
2 71998 1 878
2 71999 1 878
2 72000 1 878
2 72001 1 878
2 72002 1 878
2 72003 1 880
2 72004 1 880
2 72005 1 880
2 72006 1 880
2 72007 1 880
2 72008 1 881
2 72009 1 881
2 72010 1 884
2 72011 1 884
2 72012 1 884
2 72013 1 884
2 72014 1 884
2 72015 1 884
2 72016 1 884
2 72017 1 884
2 72018 1 884
2 72019 1 884
2 72020 1 884
2 72021 1 884
2 72022 1 884
2 72023 1 884
2 72024 1 884
2 72025 1 884
2 72026 1 884
2 72027 1 884
2 72028 1 884
2 72029 1 884
2 72030 1 884
2 72031 1 884
2 72032 1 884
2 72033 1 884
2 72034 1 884
2 72035 1 884
2 72036 1 884
2 72037 1 884
2 72038 1 885
2 72039 1 885
2 72040 1 885
2 72041 1 885
2 72042 1 885
2 72043 1 885
2 72044 1 885
2 72045 1 885
2 72046 1 885
2 72047 1 885
2 72048 1 885
2 72049 1 885
2 72050 1 885
2 72051 1 897
2 72052 1 897
2 72053 1 897
2 72054 1 897
2 72055 1 897
2 72056 1 897
2 72057 1 897
2 72058 1 897
2 72059 1 897
2 72060 1 897
2 72061 1 897
2 72062 1 897
2 72063 1 898
2 72064 1 898
2 72065 1 898
2 72066 1 898
2 72067 1 898
2 72068 1 898
2 72069 1 898
2 72070 1 898
2 72071 1 898
2 72072 1 898
2 72073 1 898
2 72074 1 898
2 72075 1 898
2 72076 1 898
2 72077 1 898
2 72078 1 898
2 72079 1 898
2 72080 1 898
2 72081 1 898
2 72082 1 898
2 72083 1 898
2 72084 1 898
2 72085 1 898
2 72086 1 898
2 72087 1 898
2 72088 1 898
2 72089 1 898
2 72090 1 898
2 72091 1 898
2 72092 1 898
2 72093 1 898
2 72094 1 898
2 72095 1 898
2 72096 1 898
2 72097 1 898
2 72098 1 898
2 72099 1 898
2 72100 1 898
2 72101 1 898
2 72102 1 899
2 72103 1 899
2 72104 1 899
2 72105 1 899
2 72106 1 899
2 72107 1 899
2 72108 1 899
2 72109 1 899
2 72110 1 900
2 72111 1 900
2 72112 1 900
2 72113 1 901
2 72114 1 901
2 72115 1 901
2 72116 1 905
2 72117 1 905
2 72118 1 905
2 72119 1 905
2 72120 1 905
2 72121 1 905
2 72122 1 906
2 72123 1 906
2 72124 1 906
2 72125 1 906
2 72126 1 906
2 72127 1 906
2 72128 1 907
2 72129 1 907
2 72130 1 907
2 72131 1 907
2 72132 1 907
2 72133 1 907
2 72134 1 907
2 72135 1 907
2 72136 1 907
2 72137 1 907
2 72138 1 907
2 72139 1 907
2 72140 1 907
2 72141 1 907
2 72142 1 907
2 72143 1 907
2 72144 1 907
2 72145 1 907
2 72146 1 907
2 72147 1 907
2 72148 1 907
2 72149 1 907
2 72150 1 907
2 72151 1 907
2 72152 1 907
2 72153 1 907
2 72154 1 907
2 72155 1 907
2 72156 1 907
2 72157 1 908
2 72158 1 908
2 72159 1 908
2 72160 1 908
2 72161 1 909
2 72162 1 909
2 72163 1 909
2 72164 1 909
2 72165 1 909
2 72166 1 909
2 72167 1 909
2 72168 1 909
2 72169 1 909
2 72170 1 909
2 72171 1 909
2 72172 1 922
2 72173 1 922
2 72174 1 922
2 72175 1 922
2 72176 1 922
2 72177 1 923
2 72178 1 923
2 72179 1 923
2 72180 1 924
2 72181 1 924
2 72182 1 924
2 72183 1 924
2 72184 1 924
2 72185 1 924
2 72186 1 925
2 72187 1 925
2 72188 1 925
2 72189 1 925
2 72190 1 925
2 72191 1 925
2 72192 1 925
2 72193 1 925
2 72194 1 925
2 72195 1 925
2 72196 1 926
2 72197 1 926
2 72198 1 926
2 72199 1 926
2 72200 1 926
2 72201 1 926
2 72202 1 926
2 72203 1 926
2 72204 1 926
2 72205 1 926
2 72206 1 934
2 72207 1 934
2 72208 1 936
2 72209 1 936
2 72210 1 936
2 72211 1 936
2 72212 1 936
2 72213 1 936
2 72214 1 937
2 72215 1 937
2 72216 1 938
2 72217 1 938
2 72218 1 938
2 72219 1 939
2 72220 1 939
2 72221 1 942
2 72222 1 942
2 72223 1 942
2 72224 1 942
2 72225 1 942
2 72226 1 943
2 72227 1 943
2 72228 1 943
2 72229 1 943
2 72230 1 943
2 72231 1 943
2 72232 1 943
2 72233 1 943
2 72234 1 943
2 72235 1 943
2 72236 1 943
2 72237 1 943
2 72238 1 943
2 72239 1 943
2 72240 1 943
2 72241 1 943
2 72242 1 943
2 72243 1 943
2 72244 1 943
2 72245 1 943
2 72246 1 943
2 72247 1 943
2 72248 1 943
2 72249 1 943
2 72250 1 943
2 72251 1 943
2 72252 1 943
2 72253 1 943
2 72254 1 943
2 72255 1 943
2 72256 1 944
2 72257 1 944
2 72258 1 944
2 72259 1 944
2 72260 1 944
2 72261 1 946
2 72262 1 946
2 72263 1 946
2 72264 1 946
2 72265 1 946
2 72266 1 956
2 72267 1 956
2 72268 1 956
2 72269 1 956
2 72270 1 957
2 72271 1 957
2 72272 1 957
2 72273 1 957
2 72274 1 957
2 72275 1 957
2 72276 1 957
2 72277 1 957
2 72278 1 958
2 72279 1 958
2 72280 1 958
2 72281 1 958
2 72282 1 958
2 72283 1 958
2 72284 1 958
2 72285 1 958
2 72286 1 958
2 72287 1 958
2 72288 1 958
2 72289 1 959
2 72290 1 959
2 72291 1 959
2 72292 1 959
2 72293 1 959
2 72294 1 959
2 72295 1 960
2 72296 1 960
2 72297 1 963
2 72298 1 963
2 72299 1 965
2 72300 1 965
2 72301 1 972
2 72302 1 972
2 72303 1 973
2 72304 1 973
2 72305 1 973
2 72306 1 973
2 72307 1 973
2 72308 1 973
2 72309 1 973
2 72310 1 973
2 72311 1 973
2 72312 1 973
2 72313 1 973
2 72314 1 973
2 72315 1 974
2 72316 1 974
2 72317 1 974
2 72318 1 974
2 72319 1 974
2 72320 1 981
2 72321 1 981
2 72322 1 982
2 72323 1 982
2 72324 1 983
2 72325 1 983
2 72326 1 983
2 72327 1 983
2 72328 1 983
2 72329 1 994
2 72330 1 994
2 72331 1 994
2 72332 1 994
2 72333 1 994
2 72334 1 994
2 72335 1 994
2 72336 1 994
2 72337 1 994
2 72338 1 994
2 72339 1 994
2 72340 1 994
2 72341 1 994
2 72342 1 994
2 72343 1 995
2 72344 1 995
2 72345 1 995
2 72346 1 995
2 72347 1 995
2 72348 1 995
2 72349 1 995
2 72350 1 995
2 72351 1 995
2 72352 1 995
2 72353 1 995
2 72354 1 995
2 72355 1 995
2 72356 1 995
2 72357 1 995
2 72358 1 995
2 72359 1 995
2 72360 1 995
2 72361 1 996
2 72362 1 996
2 72363 1 996
2 72364 1 997
2 72365 1 997
2 72366 1 999
2 72367 1 999
2 72368 1 1002
2 72369 1 1002
2 72370 1 1003
2 72371 1 1003
2 72372 1 1004
2 72373 1 1004
2 72374 1 1004
2 72375 1 1004
2 72376 1 1004
2 72377 1 1004
2 72378 1 1004
2 72379 1 1004
2 72380 1 1004
2 72381 1 1005
2 72382 1 1005
2 72383 1 1005
2 72384 1 1005
2 72385 1 1005
2 72386 1 1005
2 72387 1 1005
2 72388 1 1005
2 72389 1 1005
2 72390 1 1005
2 72391 1 1005
2 72392 1 1005
2 72393 1 1005
2 72394 1 1005
2 72395 1 1005
2 72396 1 1005
2 72397 1 1006
2 72398 1 1006
2 72399 1 1006
2 72400 1 1006
2 72401 1 1006
2 72402 1 1006
2 72403 1 1006
2 72404 1 1006
2 72405 1 1006
2 72406 1 1006
2 72407 1 1007
2 72408 1 1007
2 72409 1 1007
2 72410 1 1007
2 72411 1 1007
2 72412 1 1007
2 72413 1 1007
2 72414 1 1007
2 72415 1 1008
2 72416 1 1008
2 72417 1 1023
2 72418 1 1023
2 72419 1 1023
2 72420 1 1023
2 72421 1 1023
2 72422 1 1023
2 72423 1 1025
2 72424 1 1025
2 72425 1 1030
2 72426 1 1030
2 72427 1 1030
2 72428 1 1030
2 72429 1 1030
2 72430 1 1030
2 72431 1 1037
2 72432 1 1037
2 72433 1 1037
2 72434 1 1038
2 72435 1 1038
2 72436 1 1038
2 72437 1 1038
2 72438 1 1038
2 72439 1 1038
2 72440 1 1038
2 72441 1 1038
2 72442 1 1038
2 72443 1 1038
2 72444 1 1038
2 72445 1 1046
2 72446 1 1046
2 72447 1 1046
2 72448 1 1046
2 72449 1 1046
2 72450 1 1046
2 72451 1 1046
2 72452 1 1046
2 72453 1 1047
2 72454 1 1047
2 72455 1 1054
2 72456 1 1054
2 72457 1 1054
2 72458 1 1054
2 72459 1 1054
2 72460 1 1054
2 72461 1 1054
2 72462 1 1054
2 72463 1 1054
2 72464 1 1054
2 72465 1 1054
2 72466 1 1054
2 72467 1 1054
2 72468 1 1054
2 72469 1 1054
2 72470 1 1054
2 72471 1 1054
2 72472 1 1054
2 72473 1 1054
2 72474 1 1054
2 72475 1 1054
2 72476 1 1054
2 72477 1 1054
2 72478 1 1054
2 72479 1 1054
2 72480 1 1054
2 72481 1 1054
2 72482 1 1054
2 72483 1 1054
2 72484 1 1054
2 72485 1 1054
2 72486 1 1054
2 72487 1 1054
2 72488 1 1055
2 72489 1 1055
2 72490 1 1055
2 72491 1 1055
2 72492 1 1055
2 72493 1 1055
2 72494 1 1055
2 72495 1 1055
2 72496 1 1055
2 72497 1 1055
2 72498 1 1055
2 72499 1 1056
2 72500 1 1056
2 72501 1 1056
2 72502 1 1056
2 72503 1 1056
2 72504 1 1057
2 72505 1 1057
2 72506 1 1057
2 72507 1 1065
2 72508 1 1065
2 72509 1 1065
2 72510 1 1065
2 72511 1 1065
2 72512 1 1065
2 72513 1 1065
2 72514 1 1065
2 72515 1 1065
2 72516 1 1066
2 72517 1 1066
2 72518 1 1066
2 72519 1 1066
2 72520 1 1066
2 72521 1 1066
2 72522 1 1066
2 72523 1 1066
2 72524 1 1066
2 72525 1 1066
2 72526 1 1066
2 72527 1 1066
2 72528 1 1067
2 72529 1 1067
2 72530 1 1067
2 72531 1 1067
2 72532 1 1067
2 72533 1 1068
2 72534 1 1068
2 72535 1 1069
2 72536 1 1069
2 72537 1 1069
2 72538 1 1070
2 72539 1 1070
2 72540 1 1070
2 72541 1 1070
2 72542 1 1070
2 72543 1 1070
2 72544 1 1070
2 72545 1 1070
2 72546 1 1071
2 72547 1 1071
2 72548 1 1071
2 72549 1 1071
2 72550 1 1071
2 72551 1 1071
2 72552 1 1071
2 72553 1 1071
2 72554 1 1071
2 72555 1 1071
2 72556 1 1071
2 72557 1 1071
2 72558 1 1071
2 72559 1 1076
2 72560 1 1076
2 72561 1 1076
2 72562 1 1076
2 72563 1 1076
2 72564 1 1076
2 72565 1 1076
2 72566 1 1076
2 72567 1 1077
2 72568 1 1077
2 72569 1 1077
2 72570 1 1077
2 72571 1 1077
2 72572 1 1078
2 72573 1 1078
2 72574 1 1088
2 72575 1 1088
2 72576 1 1088
2 72577 1 1088
2 72578 1 1088
2 72579 1 1088
2 72580 1 1088
2 72581 1 1088
2 72582 1 1088
2 72583 1 1088
2 72584 1 1088
2 72585 1 1088
2 72586 1 1089
2 72587 1 1089
2 72588 1 1089
2 72589 1 1089
2 72590 1 1090
2 72591 1 1090
2 72592 1 1095
2 72593 1 1095
2 72594 1 1095
2 72595 1 1095
2 72596 1 1095
2 72597 1 1095
2 72598 1 1095
2 72599 1 1095
2 72600 1 1095
2 72601 1 1095
2 72602 1 1095
2 72603 1 1095
2 72604 1 1095
2 72605 1 1095
2 72606 1 1095
2 72607 1 1095
2 72608 1 1095
2 72609 1 1106
2 72610 1 1106
2 72611 1 1106
2 72612 1 1107
2 72613 1 1107
2 72614 1 1110
2 72615 1 1110
2 72616 1 1111
2 72617 1 1111
2 72618 1 1111
2 72619 1 1112
2 72620 1 1112
2 72621 1 1113
2 72622 1 1113
2 72623 1 1113
2 72624 1 1115
2 72625 1 1115
2 72626 1 1115
2 72627 1 1115
2 72628 1 1115
2 72629 1 1121
2 72630 1 1121
2 72631 1 1121
2 72632 1 1121
2 72633 1 1137
2 72634 1 1137
2 72635 1 1137
2 72636 1 1139
2 72637 1 1139
2 72638 1 1139
2 72639 1 1139
2 72640 1 1140
2 72641 1 1140
2 72642 1 1157
2 72643 1 1157
2 72644 1 1157
2 72645 1 1158
2 72646 1 1158
2 72647 1 1158
2 72648 1 1158
2 72649 1 1158
2 72650 1 1158
2 72651 1 1158
2 72652 1 1158
2 72653 1 1158
2 72654 1 1158
2 72655 1 1158
2 72656 1 1158
2 72657 1 1158
2 72658 1 1158
2 72659 1 1158
2 72660 1 1158
2 72661 1 1158
2 72662 1 1159
2 72663 1 1159
2 72664 1 1159
2 72665 1 1159
2 72666 1 1160
2 72667 1 1160
2 72668 1 1160
2 72669 1 1160
2 72670 1 1160
2 72671 1 1161
2 72672 1 1161
2 72673 1 1162
2 72674 1 1162
2 72675 1 1162
2 72676 1 1162
2 72677 1 1162
2 72678 1 1162
2 72679 1 1162
2 72680 1 1163
2 72681 1 1163
2 72682 1 1168
2 72683 1 1168
2 72684 1 1168
2 72685 1 1168
2 72686 1 1168
2 72687 1 1168
2 72688 1 1168
2 72689 1 1168
2 72690 1 1168
2 72691 1 1171
2 72692 1 1171
2 72693 1 1171
2 72694 1 1171
2 72695 1 1171
2 72696 1 1178
2 72697 1 1178
2 72698 1 1178
2 72699 1 1178
2 72700 1 1178
2 72701 1 1178
2 72702 1 1178
2 72703 1 1178
2 72704 1 1178
2 72705 1 1178
2 72706 1 1178
2 72707 1 1178
2 72708 1 1178
2 72709 1 1178
2 72710 1 1178
2 72711 1 1178
2 72712 1 1179
2 72713 1 1179
2 72714 1 1179
2 72715 1 1179
2 72716 1 1179
2 72717 1 1179
2 72718 1 1179
2 72719 1 1179
2 72720 1 1179
2 72721 1 1179
2 72722 1 1179
2 72723 1 1179
2 72724 1 1179
2 72725 1 1179
2 72726 1 1179
2 72727 1 1179
2 72728 1 1179
2 72729 1 1179
2 72730 1 1179
2 72731 1 1180
2 72732 1 1180
2 72733 1 1180
2 72734 1 1180
2 72735 1 1180
2 72736 1 1180
2 72737 1 1180
2 72738 1 1180
2 72739 1 1180
2 72740 1 1180
2 72741 1 1180
2 72742 1 1180
2 72743 1 1180
2 72744 1 1180
2 72745 1 1180
2 72746 1 1180
2 72747 1 1180
2 72748 1 1180
2 72749 1 1180
2 72750 1 1180
2 72751 1 1181
2 72752 1 1181
2 72753 1 1184
2 72754 1 1184
2 72755 1 1184
2 72756 1 1184
2 72757 1 1189
2 72758 1 1189
2 72759 1 1189
2 72760 1 1189
2 72761 1 1189
2 72762 1 1189
2 72763 1 1189
2 72764 1 1189
2 72765 1 1189
2 72766 1 1189
2 72767 1 1190
2 72768 1 1190
2 72769 1 1190
2 72770 1 1196
2 72771 1 1196
2 72772 1 1196
2 72773 1 1196
2 72774 1 1196
2 72775 1 1196
2 72776 1 1196
2 72777 1 1196
2 72778 1 1196
2 72779 1 1196
2 72780 1 1196
2 72781 1 1196
2 72782 1 1196
2 72783 1 1196
2 72784 1 1197
2 72785 1 1197
2 72786 1 1197
2 72787 1 1197
2 72788 1 1198
2 72789 1 1198
2 72790 1 1198
2 72791 1 1198
2 72792 1 1198
2 72793 1 1198
2 72794 1 1198
2 72795 1 1198
2 72796 1 1198
2 72797 1 1198
2 72798 1 1198
2 72799 1 1198
2 72800 1 1198
2 72801 1 1198
2 72802 1 1198
2 72803 1 1199
2 72804 1 1199
2 72805 1 1199
2 72806 1 1199
2 72807 1 1199
2 72808 1 1199
2 72809 1 1200
2 72810 1 1200
2 72811 1 1208
2 72812 1 1208
2 72813 1 1208
2 72814 1 1208
2 72815 1 1208
2 72816 1 1208
2 72817 1 1208
2 72818 1 1208
2 72819 1 1208
2 72820 1 1208
2 72821 1 1208
2 72822 1 1208
2 72823 1 1208
2 72824 1 1208
2 72825 1 1210
2 72826 1 1210
2 72827 1 1210
2 72828 1 1210
2 72829 1 1210
2 72830 1 1210
2 72831 1 1210
2 72832 1 1210
2 72833 1 1212
2 72834 1 1212
2 72835 1 1212
2 72836 1 1213
2 72837 1 1213
2 72838 1 1213
2 72839 1 1214
2 72840 1 1214
2 72841 1 1215
2 72842 1 1215
2 72843 1 1215
2 72844 1 1215
2 72845 1 1215
2 72846 1 1215
2 72847 1 1215
2 72848 1 1215
2 72849 1 1215
2 72850 1 1225
2 72851 1 1225
2 72852 1 1225
2 72853 1 1225
2 72854 1 1225
2 72855 1 1225
2 72856 1 1225
2 72857 1 1225
2 72858 1 1225
2 72859 1 1225
2 72860 1 1225
2 72861 1 1225
2 72862 1 1225
2 72863 1 1225
2 72864 1 1225
2 72865 1 1225
2 72866 1 1225
2 72867 1 1225
2 72868 1 1225
2 72869 1 1225
2 72870 1 1225
2 72871 1 1225
2 72872 1 1225
2 72873 1 1225
2 72874 1 1225
2 72875 1 1225
2 72876 1 1225
2 72877 1 1225
2 72878 1 1225
2 72879 1 1225
2 72880 1 1225
2 72881 1 1225
2 72882 1 1225
2 72883 1 1225
2 72884 1 1225
2 72885 1 1225
2 72886 1 1226
2 72887 1 1226
2 72888 1 1226
2 72889 1 1226
2 72890 1 1226
2 72891 1 1226
2 72892 1 1226
2 72893 1 1226
2 72894 1 1226
2 72895 1 1226
2 72896 1 1226
2 72897 1 1226
2 72898 1 1226
2 72899 1 1226
2 72900 1 1226
2 72901 1 1226
2 72902 1 1226
2 72903 1 1226
2 72904 1 1226
2 72905 1 1226
2 72906 1 1226
2 72907 1 1226
2 72908 1 1226
2 72909 1 1226
2 72910 1 1226
2 72911 1 1226
2 72912 1 1226
2 72913 1 1226
2 72914 1 1226
2 72915 1 1226
2 72916 1 1226
2 72917 1 1226
2 72918 1 1226
2 72919 1 1226
2 72920 1 1226
2 72921 1 1226
2 72922 1 1226
2 72923 1 1226
2 72924 1 1226
2 72925 1 1226
2 72926 1 1227
2 72927 1 1227
2 72928 1 1227
2 72929 1 1228
2 72930 1 1228
2 72931 1 1228
2 72932 1 1228
2 72933 1 1228
2 72934 1 1228
2 72935 1 1228
2 72936 1 1228
2 72937 1 1228
2 72938 1 1229
2 72939 1 1229
2 72940 1 1229
2 72941 1 1229
2 72942 1 1229
2 72943 1 1229
2 72944 1 1230
2 72945 1 1230
2 72946 1 1230
2 72947 1 1230
2 72948 1 1230
2 72949 1 1231
2 72950 1 1231
2 72951 1 1232
2 72952 1 1232
2 72953 1 1232
2 72954 1 1234
2 72955 1 1234
2 72956 1 1235
2 72957 1 1235
2 72958 1 1235
2 72959 1 1235
2 72960 1 1235
2 72961 1 1235
2 72962 1 1235
2 72963 1 1235
2 72964 1 1238
2 72965 1 1238
2 72966 1 1241
2 72967 1 1241
2 72968 1 1241
2 72969 1 1241
2 72970 1 1241
2 72971 1 1241
2 72972 1 1241
2 72973 1 1241
2 72974 1 1241
2 72975 1 1241
2 72976 1 1241
2 72977 1 1241
2 72978 1 1242
2 72979 1 1242
2 72980 1 1242
2 72981 1 1242
2 72982 1 1242
2 72983 1 1242
2 72984 1 1242
2 72985 1 1242
2 72986 1 1242
2 72987 1 1242
2 72988 1 1242
2 72989 1 1242
2 72990 1 1242
2 72991 1 1242
2 72992 1 1242
2 72993 1 1251
2 72994 1 1251
2 72995 1 1251
2 72996 1 1251
2 72997 1 1251
2 72998 1 1251
2 72999 1 1251
2 73000 1 1251
2 73001 1 1251
2 73002 1 1251
2 73003 1 1251
2 73004 1 1251
2 73005 1 1251
2 73006 1 1251
2 73007 1 1251
2 73008 1 1251
2 73009 1 1251
2 73010 1 1251
2 73011 1 1251
2 73012 1 1251
2 73013 1 1251
2 73014 1 1251
2 73015 1 1251
2 73016 1 1251
2 73017 1 1251
2 73018 1 1251
2 73019 1 1251
2 73020 1 1251
2 73021 1 1252
2 73022 1 1252
2 73023 1 1252
2 73024 1 1252
2 73025 1 1252
2 73026 1 1252
2 73027 1 1252
2 73028 1 1252
2 73029 1 1254
2 73030 1 1254
2 73031 1 1255
2 73032 1 1255
2 73033 1 1255
2 73034 1 1255
2 73035 1 1255
2 73036 1 1255
2 73037 1 1255
2 73038 1 1255
2 73039 1 1255
2 73040 1 1255
2 73041 1 1255
2 73042 1 1255
2 73043 1 1255
2 73044 1 1255
2 73045 1 1255
2 73046 1 1255
2 73047 1 1255
2 73048 1 1255
2 73049 1 1255
2 73050 1 1255
2 73051 1 1255
2 73052 1 1255
2 73053 1 1255
2 73054 1 1255
2 73055 1 1255
2 73056 1 1255
2 73057 1 1255
2 73058 1 1256
2 73059 1 1256
2 73060 1 1256
2 73061 1 1256
2 73062 1 1256
2 73063 1 1256
2 73064 1 1256
2 73065 1 1256
2 73066 1 1256
2 73067 1 1256
2 73068 1 1256
2 73069 1 1256
2 73070 1 1256
2 73071 1 1256
2 73072 1 1256
2 73073 1 1256
2 73074 1 1257
2 73075 1 1257
2 73076 1 1257
2 73077 1 1258
2 73078 1 1258
2 73079 1 1258
2 73080 1 1258
2 73081 1 1258
2 73082 1 1258
2 73083 1 1258
2 73084 1 1258
2 73085 1 1258
2 73086 1 1258
2 73087 1 1258
2 73088 1 1258
2 73089 1 1258
2 73090 1 1258
2 73091 1 1258
2 73092 1 1258
2 73093 1 1258
2 73094 1 1258
2 73095 1 1258
2 73096 1 1258
2 73097 1 1258
2 73098 1 1258
2 73099 1 1259
2 73100 1 1259
2 73101 1 1259
2 73102 1 1259
2 73103 1 1259
2 73104 1 1259
2 73105 1 1259
2 73106 1 1259
2 73107 1 1259
2 73108 1 1259
2 73109 1 1259
2 73110 1 1259
2 73111 1 1259
2 73112 1 1259
2 73113 1 1259
2 73114 1 1259
2 73115 1 1259
2 73116 1 1259
2 73117 1 1259
2 73118 1 1259
2 73119 1 1259
2 73120 1 1259
2 73121 1 1259
2 73122 1 1259
2 73123 1 1259
2 73124 1 1259
2 73125 1 1259
2 73126 1 1259
2 73127 1 1259
2 73128 1 1259
2 73129 1 1259
2 73130 1 1259
2 73131 1 1259
2 73132 1 1259
2 73133 1 1259
2 73134 1 1259
2 73135 1 1259
2 73136 1 1259
2 73137 1 1260
2 73138 1 1260
2 73139 1 1260
2 73140 1 1260
2 73141 1 1260
2 73142 1 1260
2 73143 1 1260
2 73144 1 1260
2 73145 1 1260
2 73146 1 1260
2 73147 1 1260
2 73148 1 1260
2 73149 1 1260
2 73150 1 1260
2 73151 1 1260
2 73152 1 1260
2 73153 1 1260
2 73154 1 1260
2 73155 1 1260
2 73156 1 1260
2 73157 1 1260
2 73158 1 1260
2 73159 1 1260
2 73160 1 1260
2 73161 1 1260
2 73162 1 1260
2 73163 1 1260
2 73164 1 1260
2 73165 1 1260
2 73166 1 1260
2 73167 1 1260
2 73168 1 1260
2 73169 1 1260
2 73170 1 1260
2 73171 1 1260
2 73172 1 1260
2 73173 1 1260
2 73174 1 1260
2 73175 1 1260
2 73176 1 1260
2 73177 1 1260
2 73178 1 1260
2 73179 1 1260
2 73180 1 1260
2 73181 1 1260
2 73182 1 1260
2 73183 1 1260
2 73184 1 1261
2 73185 1 1261
2 73186 1 1274
2 73187 1 1274
2 73188 1 1276
2 73189 1 1276
2 73190 1 1276
2 73191 1 1276
2 73192 1 1285
2 73193 1 1285
2 73194 1 1285
2 73195 1 1285
2 73196 1 1285
2 73197 1 1285
2 73198 1 1286
2 73199 1 1286
2 73200 1 1288
2 73201 1 1288
2 73202 1 1288
2 73203 1 1288
2 73204 1 1288
2 73205 1 1288
2 73206 1 1288
2 73207 1 1288
2 73208 1 1288
2 73209 1 1288
2 73210 1 1288
2 73211 1 1288
2 73212 1 1289
2 73213 1 1289
2 73214 1 1289
2 73215 1 1289
2 73216 1 1289
2 73217 1 1289
2 73218 1 1289
2 73219 1 1289
2 73220 1 1289
2 73221 1 1289
2 73222 1 1292
2 73223 1 1292
2 73224 1 1292
2 73225 1 1292
2 73226 1 1292
2 73227 1 1292
2 73228 1 1292
2 73229 1 1292
2 73230 1 1292
2 73231 1 1294
2 73232 1 1294
2 73233 1 1294
2 73234 1 1294
2 73235 1 1305
2 73236 1 1305
2 73237 1 1305
2 73238 1 1305
2 73239 1 1305
2 73240 1 1305
2 73241 1 1305
2 73242 1 1305
2 73243 1 1305
2 73244 1 1305
2 73245 1 1305
2 73246 1 1305
2 73247 1 1305
2 73248 1 1305
2 73249 1 1305
2 73250 1 1305
2 73251 1 1305
2 73252 1 1305
2 73253 1 1305
2 73254 1 1305
2 73255 1 1305
2 73256 1 1305
2 73257 1 1305
2 73258 1 1305
2 73259 1 1305
2 73260 1 1305
2 73261 1 1305
2 73262 1 1305
2 73263 1 1305
2 73264 1 1305
2 73265 1 1305
2 73266 1 1305
2 73267 1 1305
2 73268 1 1305
2 73269 1 1305
2 73270 1 1305
2 73271 1 1305
2 73272 1 1305
2 73273 1 1306
2 73274 1 1306
2 73275 1 1306
2 73276 1 1308
2 73277 1 1308
2 73278 1 1308
2 73279 1 1310
2 73280 1 1310
2 73281 1 1311
2 73282 1 1311
2 73283 1 1311
2 73284 1 1311
2 73285 1 1312
2 73286 1 1312
2 73287 1 1312
2 73288 1 1312
2 73289 1 1312
2 73290 1 1312
2 73291 1 1312
2 73292 1 1312
2 73293 1 1312
2 73294 1 1312
2 73295 1 1312
2 73296 1 1312
2 73297 1 1327
2 73298 1 1327
2 73299 1 1327
2 73300 1 1327
2 73301 1 1327
2 73302 1 1327
2 73303 1 1327
2 73304 1 1327
2 73305 1 1327
2 73306 1 1327
2 73307 1 1327
2 73308 1 1327
2 73309 1 1327
2 73310 1 1327
2 73311 1 1327
2 73312 1 1327
2 73313 1 1327
2 73314 1 1327
2 73315 1 1327
2 73316 1 1327
2 73317 1 1327
2 73318 1 1327
2 73319 1 1327
2 73320 1 1327
2 73321 1 1327
2 73322 1 1327
2 73323 1 1327
2 73324 1 1327
2 73325 1 1327
2 73326 1 1327
2 73327 1 1327
2 73328 1 1328
2 73329 1 1328
2 73330 1 1328
2 73331 1 1328
2 73332 1 1328
2 73333 1 1328
2 73334 1 1328
2 73335 1 1328
2 73336 1 1329
2 73337 1 1329
2 73338 1 1329
2 73339 1 1330
2 73340 1 1330
2 73341 1 1330
2 73342 1 1330
2 73343 1 1331
2 73344 1 1331
2 73345 1 1332
2 73346 1 1332
2 73347 1 1332
2 73348 1 1332
2 73349 1 1332
2 73350 1 1333
2 73351 1 1333
2 73352 1 1341
2 73353 1 1341
2 73354 1 1341
2 73355 1 1341
2 73356 1 1341
2 73357 1 1341
2 73358 1 1341
2 73359 1 1342
2 73360 1 1342
2 73361 1 1342
2 73362 1 1342
2 73363 1 1342
2 73364 1 1342
2 73365 1 1342
2 73366 1 1342
2 73367 1 1342
2 73368 1 1342
2 73369 1 1342
2 73370 1 1343
2 73371 1 1343
2 73372 1 1344
2 73373 1 1344
2 73374 1 1344
2 73375 1 1344
2 73376 1 1344
2 73377 1 1344
2 73378 1 1344
2 73379 1 1344
2 73380 1 1344
2 73381 1 1344
2 73382 1 1344
2 73383 1 1344
2 73384 1 1344
2 73385 1 1344
2 73386 1 1344
2 73387 1 1344
2 73388 1 1344
2 73389 1 1344
2 73390 1 1344
2 73391 1 1345
2 73392 1 1345
2 73393 1 1345
2 73394 1 1346
2 73395 1 1346
2 73396 1 1346
2 73397 1 1346
2 73398 1 1346
2 73399 1 1346
2 73400 1 1346
2 73401 1 1346
2 73402 1 1346
2 73403 1 1346
2 73404 1 1346
2 73405 1 1346
2 73406 1 1346
2 73407 1 1346
2 73408 1 1346
2 73409 1 1346
2 73410 1 1347
2 73411 1 1347
2 73412 1 1347
2 73413 1 1347
2 73414 1 1347
2 73415 1 1350
2 73416 1 1350
2 73417 1 1350
2 73418 1 1352
2 73419 1 1352
2 73420 1 1352
2 73421 1 1352
2 73422 1 1352
2 73423 1 1352
2 73424 1 1352
2 73425 1 1353
2 73426 1 1353
2 73427 1 1355
2 73428 1 1355
2 73429 1 1358
2 73430 1 1358
2 73431 1 1358
2 73432 1 1358
2 73433 1 1358
2 73434 1 1359
2 73435 1 1359
2 73436 1 1359
2 73437 1 1359
2 73438 1 1359
2 73439 1 1359
2 73440 1 1359
2 73441 1 1361
2 73442 1 1361
2 73443 1 1361
2 73444 1 1361
2 73445 1 1361
2 73446 1 1361
2 73447 1 1361
2 73448 1 1362
2 73449 1 1362
2 73450 1 1365
2 73451 1 1365
2 73452 1 1365
2 73453 1 1365
2 73454 1 1365
2 73455 1 1365
2 73456 1 1365
2 73457 1 1366
2 73458 1 1366
2 73459 1 1366
2 73460 1 1366
2 73461 1 1366
2 73462 1 1366
2 73463 1 1366
2 73464 1 1366
2 73465 1 1366
2 73466 1 1366
2 73467 1 1366
2 73468 1 1366
2 73469 1 1366
2 73470 1 1366
2 73471 1 1366
2 73472 1 1366
2 73473 1 1366
2 73474 1 1366
2 73475 1 1366
2 73476 1 1366
2 73477 1 1366
2 73478 1 1366
2 73479 1 1373
2 73480 1 1373
2 73481 1 1373
2 73482 1 1373
2 73483 1 1373
2 73484 1 1374
2 73485 1 1374
2 73486 1 1374
2 73487 1 1374
2 73488 1 1374
2 73489 1 1374
2 73490 1 1374
2 73491 1 1374
2 73492 1 1376
2 73493 1 1376
2 73494 1 1376
2 73495 1 1376
2 73496 1 1376
2 73497 1 1376
2 73498 1 1376
2 73499 1 1376
2 73500 1 1376
2 73501 1 1376
2 73502 1 1376
2 73503 1 1376
2 73504 1 1377
2 73505 1 1377
2 73506 1 1377
2 73507 1 1378
2 73508 1 1378
2 73509 1 1378
2 73510 1 1378
2 73511 1 1378
2 73512 1 1378
2 73513 1 1378
2 73514 1 1378
2 73515 1 1378
2 73516 1 1378
2 73517 1 1378
2 73518 1 1378
2 73519 1 1378
2 73520 1 1378
2 73521 1 1379
2 73522 1 1379
2 73523 1 1379
2 73524 1 1381
2 73525 1 1381
2 73526 1 1383
2 73527 1 1383
2 73528 1 1386
2 73529 1 1386
2 73530 1 1386
2 73531 1 1386
2 73532 1 1386
2 73533 1 1386
2 73534 1 1386
2 73535 1 1393
2 73536 1 1393
2 73537 1 1393
2 73538 1 1394
2 73539 1 1394
2 73540 1 1394
2 73541 1 1394
2 73542 1 1394
2 73543 1 1394
2 73544 1 1394
2 73545 1 1394
2 73546 1 1394
2 73547 1 1394
2 73548 1 1394
2 73549 1 1394
2 73550 1 1394
2 73551 1 1394
2 73552 1 1394
2 73553 1 1394
2 73554 1 1394
2 73555 1 1394
2 73556 1 1396
2 73557 1 1396
2 73558 1 1396
2 73559 1 1396
2 73560 1 1396
2 73561 1 1396
2 73562 1 1396
2 73563 1 1396
2 73564 1 1396
2 73565 1 1396
2 73566 1 1396
2 73567 1 1396
2 73568 1 1396
2 73569 1 1396
2 73570 1 1397
2 73571 1 1397
2 73572 1 1397
2 73573 1 1397
2 73574 1 1397
2 73575 1 1398
2 73576 1 1398
2 73577 1 1406
2 73578 1 1406
2 73579 1 1406
2 73580 1 1406
2 73581 1 1406
2 73582 1 1407
2 73583 1 1407
2 73584 1 1407
2 73585 1 1407
2 73586 1 1407
2 73587 1 1407
2 73588 1 1407
2 73589 1 1407
2 73590 1 1407
2 73591 1 1407
2 73592 1 1407
2 73593 1 1407
2 73594 1 1407
2 73595 1 1407
2 73596 1 1407
2 73597 1 1407
2 73598 1 1407
2 73599 1 1407
2 73600 1 1415
2 73601 1 1415
2 73602 1 1415
2 73603 1 1416
2 73604 1 1416
2 73605 1 1416
2 73606 1 1416
2 73607 1 1416
2 73608 1 1416
2 73609 1 1416
2 73610 1 1416
2 73611 1 1416
2 73612 1 1416
2 73613 1 1416
2 73614 1 1416
2 73615 1 1416
2 73616 1 1416
2 73617 1 1416
2 73618 1 1416
2 73619 1 1416
2 73620 1 1416
2 73621 1 1416
2 73622 1 1416
2 73623 1 1416
2 73624 1 1416
2 73625 1 1416
2 73626 1 1416
2 73627 1 1416
2 73628 1 1416
2 73629 1 1416
2 73630 1 1416
2 73631 1 1416
2 73632 1 1416
2 73633 1 1416
2 73634 1 1416
2 73635 1 1416
2 73636 1 1417
2 73637 1 1417
2 73638 1 1417
2 73639 1 1417
2 73640 1 1419
2 73641 1 1419
2 73642 1 1421
2 73643 1 1421
2 73644 1 1421
2 73645 1 1428
2 73646 1 1428
2 73647 1 1428
2 73648 1 1428
2 73649 1 1428
2 73650 1 1428
2 73651 1 1428
2 73652 1 1428
2 73653 1 1428
2 73654 1 1428
2 73655 1 1428
2 73656 1 1428
2 73657 1 1428
2 73658 1 1428
2 73659 1 1428
2 73660 1 1428
2 73661 1 1428
2 73662 1 1428
2 73663 1 1428
2 73664 1 1428
2 73665 1 1428
2 73666 1 1428
2 73667 1 1428
2 73668 1 1428
2 73669 1 1428
2 73670 1 1428
2 73671 1 1428
2 73672 1 1428
2 73673 1 1428
2 73674 1 1428
2 73675 1 1428
2 73676 1 1428
2 73677 1 1428
2 73678 1 1428
2 73679 1 1428
2 73680 1 1428
2 73681 1 1428
2 73682 1 1428
2 73683 1 1428
2 73684 1 1428
2 73685 1 1429
2 73686 1 1429
2 73687 1 1429
2 73688 1 1429
2 73689 1 1429
2 73690 1 1429
2 73691 1 1429
2 73692 1 1429
2 73693 1 1429
2 73694 1 1429
2 73695 1 1429
2 73696 1 1429
2 73697 1 1429
2 73698 1 1429
2 73699 1 1429
2 73700 1 1429
2 73701 1 1429
2 73702 1 1429
2 73703 1 1429
2 73704 1 1429
2 73705 1 1435
2 73706 1 1435
2 73707 1 1438
2 73708 1 1438
2 73709 1 1438
2 73710 1 1438
2 73711 1 1438
2 73712 1 1438
2 73713 1 1438
2 73714 1 1438
2 73715 1 1438
2 73716 1 1438
2 73717 1 1438
2 73718 1 1438
2 73719 1 1438
2 73720 1 1438
2 73721 1 1438
2 73722 1 1438
2 73723 1 1438
2 73724 1 1438
2 73725 1 1438
2 73726 1 1438
2 73727 1 1438
2 73728 1 1438
2 73729 1 1438
2 73730 1 1438
2 73731 1 1439
2 73732 1 1439
2 73733 1 1440
2 73734 1 1440
2 73735 1 1440
2 73736 1 1440
2 73737 1 1440
2 73738 1 1442
2 73739 1 1442
2 73740 1 1443
2 73741 1 1443
2 73742 1 1443
2 73743 1 1443
2 73744 1 1443
2 73745 1 1443
2 73746 1 1451
2 73747 1 1451
2 73748 1 1466
2 73749 1 1466
2 73750 1 1468
2 73751 1 1468
2 73752 1 1468
2 73753 1 1468
2 73754 1 1468
2 73755 1 1468
2 73756 1 1468
2 73757 1 1468
2 73758 1 1468
2 73759 1 1468
2 73760 1 1468
2 73761 1 1468
2 73762 1 1468
2 73763 1 1468
2 73764 1 1468
2 73765 1 1468
2 73766 1 1468
2 73767 1 1468
2 73768 1 1469
2 73769 1 1469
2 73770 1 1469
2 73771 1 1480
2 73772 1 1480
2 73773 1 1480
2 73774 1 1480
2 73775 1 1480
2 73776 1 1480
2 73777 1 1480
2 73778 1 1480
2 73779 1 1480
2 73780 1 1480
2 73781 1 1480
2 73782 1 1480
2 73783 1 1480
2 73784 1 1480
2 73785 1 1481
2 73786 1 1481
2 73787 1 1482
2 73788 1 1482
2 73789 1 1485
2 73790 1 1485
2 73791 1 1485
2 73792 1 1485
2 73793 1 1485
2 73794 1 1485
2 73795 1 1485
2 73796 1 1485
2 73797 1 1486
2 73798 1 1486
2 73799 1 1486
2 73800 1 1486
2 73801 1 1486
2 73802 1 1488
2 73803 1 1488
2 73804 1 1496
2 73805 1 1496
2 73806 1 1496
2 73807 1 1496
2 73808 1 1497
2 73809 1 1497
2 73810 1 1498
2 73811 1 1498
2 73812 1 1499
2 73813 1 1499
2 73814 1 1499
2 73815 1 1499
2 73816 1 1507
2 73817 1 1507
2 73818 1 1507
2 73819 1 1507
2 73820 1 1507
2 73821 1 1508
2 73822 1 1508
2 73823 1 1508
2 73824 1 1508
2 73825 1 1509
2 73826 1 1509
2 73827 1 1509
2 73828 1 1509
2 73829 1 1509
2 73830 1 1509
2 73831 1 1509
2 73832 1 1509
2 73833 1 1509
2 73834 1 1509
2 73835 1 1509
2 73836 1 1509
2 73837 1 1509
2 73838 1 1509
2 73839 1 1509
2 73840 1 1509
2 73841 1 1509
2 73842 1 1509
2 73843 1 1509
2 73844 1 1509
2 73845 1 1509
2 73846 1 1510
2 73847 1 1510
2 73848 1 1517
2 73849 1 1517
2 73850 1 1517
2 73851 1 1517
2 73852 1 1517
2 73853 1 1517
2 73854 1 1517
2 73855 1 1517
2 73856 1 1517
2 73857 1 1517
2 73858 1 1517
2 73859 1 1517
2 73860 1 1518
2 73861 1 1518
2 73862 1 1518
2 73863 1 1520
2 73864 1 1520
2 73865 1 1523
2 73866 1 1523
2 73867 1 1523
2 73868 1 1523
2 73869 1 1523
2 73870 1 1523
2 73871 1 1523
2 73872 1 1523
2 73873 1 1523
2 73874 1 1523
2 73875 1 1523
2 73876 1 1523
2 73877 1 1523
2 73878 1 1523
2 73879 1 1523
2 73880 1 1523
2 73881 1 1523
2 73882 1 1524
2 73883 1 1524
2 73884 1 1524
2 73885 1 1524
2 73886 1 1524
2 73887 1 1524
2 73888 1 1524
2 73889 1 1531
2 73890 1 1531
2 73891 1 1531
2 73892 1 1532
2 73893 1 1532
2 73894 1 1532
2 73895 1 1532
2 73896 1 1532
2 73897 1 1532
2 73898 1 1532
2 73899 1 1532
2 73900 1 1532
2 73901 1 1532
2 73902 1 1534
2 73903 1 1534
2 73904 1 1534
2 73905 1 1534
2 73906 1 1534
2 73907 1 1534
2 73908 1 1534
2 73909 1 1534
2 73910 1 1534
2 73911 1 1534
2 73912 1 1534
2 73913 1 1534
2 73914 1 1534
2 73915 1 1541
2 73916 1 1541
2 73917 1 1541
2 73918 1 1541
2 73919 1 1541
2 73920 1 1542
2 73921 1 1542
2 73922 1 1542
2 73923 1 1542
2 73924 1 1542
2 73925 1 1542
2 73926 1 1542
2 73927 1 1543
2 73928 1 1543
2 73929 1 1543
2 73930 1 1543
2 73931 1 1543
2 73932 1 1543
2 73933 1 1543
2 73934 1 1543
2 73935 1 1543
2 73936 1 1543
2 73937 1 1543
2 73938 1 1543
2 73939 1 1543
2 73940 1 1543
2 73941 1 1543
2 73942 1 1543
2 73943 1 1543
2 73944 1 1543
2 73945 1 1543
2 73946 1 1543
2 73947 1 1543
2 73948 1 1545
2 73949 1 1545
2 73950 1 1545
2 73951 1 1545
2 73952 1 1545
2 73953 1 1545
2 73954 1 1545
2 73955 1 1545
2 73956 1 1546
2 73957 1 1546
2 73958 1 1546
2 73959 1 1567
2 73960 1 1567
2 73961 1 1567
2 73962 1 1567
2 73963 1 1567
2 73964 1 1567
2 73965 1 1567
2 73966 1 1567
2 73967 1 1567
2 73968 1 1567
2 73969 1 1567
2 73970 1 1567
2 73971 1 1567
2 73972 1 1569
2 73973 1 1569
2 73974 1 1572
2 73975 1 1572
2 73976 1 1572
2 73977 1 1572
2 73978 1 1572
2 73979 1 1572
2 73980 1 1572
2 73981 1 1572
2 73982 1 1572
2 73983 1 1572
2 73984 1 1579
2 73985 1 1579
2 73986 1 1582
2 73987 1 1582
2 73988 1 1582
2 73989 1 1582
2 73990 1 1582
2 73991 1 1583
2 73992 1 1583
2 73993 1 1584
2 73994 1 1584
2 73995 1 1584
2 73996 1 1584
2 73997 1 1584
2 73998 1 1584
2 73999 1 1584
2 74000 1 1584
2 74001 1 1584
2 74002 1 1584
2 74003 1 1595
2 74004 1 1595
2 74005 1 1595
2 74006 1 1595
2 74007 1 1595
2 74008 1 1595
2 74009 1 1595
2 74010 1 1596
2 74011 1 1596
2 74012 1 1601
2 74013 1 1601
2 74014 1 1601
2 74015 1 1601
2 74016 1 1601
2 74017 1 1601
2 74018 1 1601
2 74019 1 1609
2 74020 1 1609
2 74021 1 1621
2 74022 1 1621
2 74023 1 1621
2 74024 1 1621
2 74025 1 1621
2 74026 1 1621
2 74027 1 1621
2 74028 1 1622
2 74029 1 1622
2 74030 1 1622
2 74031 1 1622
2 74032 1 1622
2 74033 1 1622
2 74034 1 1622
2 74035 1 1622
2 74036 1 1622
2 74037 1 1622
2 74038 1 1622
2 74039 1 1622
2 74040 1 1622
2 74041 1 1622
2 74042 1 1622
2 74043 1 1623
2 74044 1 1623
2 74045 1 1623
2 74046 1 1632
2 74047 1 1632
2 74048 1 1632
2 74049 1 1632
2 74050 1 1632
2 74051 1 1632
2 74052 1 1632
2 74053 1 1634
2 74054 1 1634
2 74055 1 1634
2 74056 1 1634
2 74057 1 1641
2 74058 1 1641
2 74059 1 1642
2 74060 1 1642
2 74061 1 1643
2 74062 1 1643
2 74063 1 1654
2 74064 1 1654
2 74065 1 1655
2 74066 1 1655
2 74067 1 1655
2 74068 1 1660
2 74069 1 1660
2 74070 1 1665
2 74071 1 1665
2 74072 1 1665
2 74073 1 1665
2 74074 1 1665
2 74075 1 1665
2 74076 1 1665
2 74077 1 1665
2 74078 1 1666
2 74079 1 1666
2 74080 1 1666
2 74081 1 1668
2 74082 1 1668
2 74083 1 1668
2 74084 1 1673
2 74085 1 1673
2 74086 1 1676
2 74087 1 1676
2 74088 1 1677
2 74089 1 1677
2 74090 1 1677
2 74091 1 1677
2 74092 1 1677
2 74093 1 1677
2 74094 1 1677
2 74095 1 1677
2 74096 1 1677
2 74097 1 1677
2 74098 1 1677
2 74099 1 1677
2 74100 1 1677
2 74101 1 1678
2 74102 1 1678
2 74103 1 1678
2 74104 1 1678
2 74105 1 1682
2 74106 1 1682
2 74107 1 1693
2 74108 1 1693
2 74109 1 1712
2 74110 1 1712
2 74111 1 1712
2 74112 1 1719
2 74113 1 1719
2 74114 1 1720
2 74115 1 1720
2 74116 1 1720
2 74117 1 1721
2 74118 1 1721
2 74119 1 1721
2 74120 1 1721
2 74121 1 1721
2 74122 1 1721
2 74123 1 1721
2 74124 1 1721
2 74125 1 1721
2 74126 1 1721
2 74127 1 1721
2 74128 1 1721
2 74129 1 1721
2 74130 1 1721
2 74131 1 1721
2 74132 1 1721
2 74133 1 1721
2 74134 1 1721
2 74135 1 1721
2 74136 1 1721
2 74137 1 1721
2 74138 1 1721
2 74139 1 1721
2 74140 1 1722
2 74141 1 1722
2 74142 1 1722
2 74143 1 1722
2 74144 1 1722
2 74145 1 1722
2 74146 1 1722
2 74147 1 1722
2 74148 1 1722
2 74149 1 1722
2 74150 1 1722
2 74151 1 1722
2 74152 1 1723
2 74153 1 1723
2 74154 1 1723
2 74155 1 1723
2 74156 1 1723
2 74157 1 1723
2 74158 1 1723
2 74159 1 1723
2 74160 1 1734
2 74161 1 1734
2 74162 1 1734
2 74163 1 1734
2 74164 1 1755
2 74165 1 1755
2 74166 1 1755
2 74167 1 1755
2 74168 1 1755
2 74169 1 1756
2 74170 1 1756
2 74171 1 1756
2 74172 1 1757
2 74173 1 1757
2 74174 1 1757
2 74175 1 1757
2 74176 1 1757
2 74177 1 1769
2 74178 1 1769
2 74179 1 1769
2 74180 1 1769
2 74181 1 1769
2 74182 1 1769
2 74183 1 1772
2 74184 1 1772
2 74185 1 1772
2 74186 1 1772
2 74187 1 1772
2 74188 1 1772
2 74189 1 1772
2 74190 1 1772
2 74191 1 1772
2 74192 1 1772
2 74193 1 1772
2 74194 1 1772
2 74195 1 1772
2 74196 1 1772
2 74197 1 1772
2 74198 1 1773
2 74199 1 1773
2 74200 1 1773
2 74201 1 1773
2 74202 1 1773
2 74203 1 1773
2 74204 1 1781
2 74205 1 1781
2 74206 1 1781
2 74207 1 1781
2 74208 1 1781
2 74209 1 1797
2 74210 1 1797
2 74211 1 1797
2 74212 1 1797
2 74213 1 1797
2 74214 1 1797
2 74215 1 1797
2 74216 1 1797
2 74217 1 1797
2 74218 1 1797
2 74219 1 1797
2 74220 1 1797
2 74221 1 1797
2 74222 1 1797
2 74223 1 1797
2 74224 1 1797
2 74225 1 1797
2 74226 1 1797
2 74227 1 1797
2 74228 1 1798
2 74229 1 1798
2 74230 1 1798
2 74231 1 1798
2 74232 1 1799
2 74233 1 1799
2 74234 1 1799
2 74235 1 1799
2 74236 1 1817
2 74237 1 1817
2 74238 1 1817
2 74239 1 1818
2 74240 1 1818
2 74241 1 1818
2 74242 1 1818
2 74243 1 1821
2 74244 1 1821
2 74245 1 1821
2 74246 1 1821
2 74247 1 1821
2 74248 1 1821
2 74249 1 1821
2 74250 1 1821
2 74251 1 1821
2 74252 1 1822
2 74253 1 1822
2 74254 1 1822
2 74255 1 1822
2 74256 1 1822
2 74257 1 1822
2 74258 1 1822
2 74259 1 1822
2 74260 1 1822
2 74261 1 1822
2 74262 1 1822
2 74263 1 1822
2 74264 1 1822
2 74265 1 1822
2 74266 1 1822
2 74267 1 1822
2 74268 1 1822
2 74269 1 1822
2 74270 1 1822
2 74271 1 1822
2 74272 1 1822
2 74273 1 1822
2 74274 1 1822
2 74275 1 1822
2 74276 1 1822
2 74277 1 1822
2 74278 1 1822
2 74279 1 1822
2 74280 1 1822
2 74281 1 1822
2 74282 1 1822
2 74283 1 1822
2 74284 1 1823
2 74285 1 1823
2 74286 1 1823
2 74287 1 1830
2 74288 1 1830
2 74289 1 1830
2 74290 1 1830
2 74291 1 1830
2 74292 1 1830
2 74293 1 1830
2 74294 1 1830
2 74295 1 1830
2 74296 1 1830
2 74297 1 1830
2 74298 1 1830
2 74299 1 1830
2 74300 1 1830
2 74301 1 1830
2 74302 1 1830
2 74303 1 1830
2 74304 1 1831
2 74305 1 1831
2 74306 1 1831
2 74307 1 1831
2 74308 1 1831
2 74309 1 1831
2 74310 1 1832
2 74311 1 1832
2 74312 1 1832
2 74313 1 1834
2 74314 1 1834
2 74315 1 1834
2 74316 1 1834
2 74317 1 1834
2 74318 1 1834
2 74319 1 1834
2 74320 1 1834
2 74321 1 1834
2 74322 1 1834
2 74323 1 1834
2 74324 1 1834
2 74325 1 1834
2 74326 1 1834
2 74327 1 1834
2 74328 1 1834
2 74329 1 1834
2 74330 1 1834
2 74331 1 1834
2 74332 1 1834
2 74333 1 1834
2 74334 1 1834
2 74335 1 1834
2 74336 1 1834
2 74337 1 1834
2 74338 1 1834
2 74339 1 1834
2 74340 1 1834
2 74341 1 1834
2 74342 1 1834
2 74343 1 1834
2 74344 1 1834
2 74345 1 1834
2 74346 1 1834
2 74347 1 1834
2 74348 1 1834
2 74349 1 1834
2 74350 1 1835
2 74351 1 1835
2 74352 1 1835
2 74353 1 1835
2 74354 1 1835
2 74355 1 1835
2 74356 1 1835
2 74357 1 1835
2 74358 1 1835
2 74359 1 1835
2 74360 1 1835
2 74361 1 1835
2 74362 1 1835
2 74363 1 1835
2 74364 1 1835
2 74365 1 1835
2 74366 1 1835
2 74367 1 1835
2 74368 1 1835
2 74369 1 1835
2 74370 1 1835
2 74371 1 1835
2 74372 1 1835
2 74373 1 1835
2 74374 1 1835
2 74375 1 1835
2 74376 1 1835
2 74377 1 1835
2 74378 1 1835
2 74379 1 1835
2 74380 1 1835
2 74381 1 1835
2 74382 1 1835
2 74383 1 1835
2 74384 1 1835
2 74385 1 1835
2 74386 1 1844
2 74387 1 1844
2 74388 1 1844
2 74389 1 1848
2 74390 1 1848
2 74391 1 1848
2 74392 1 1848
2 74393 1 1848
2 74394 1 1848
2 74395 1 1848
2 74396 1 1848
2 74397 1 1849
2 74398 1 1849
2 74399 1 1849
2 74400 1 1849
2 74401 1 1849
2 74402 1 1849
2 74403 1 1849
2 74404 1 1849
2 74405 1 1849
2 74406 1 1849
2 74407 1 1849
2 74408 1 1849
2 74409 1 1849
2 74410 1 1849
2 74411 1 1849
2 74412 1 1849
2 74413 1 1849
2 74414 1 1853
2 74415 1 1853
2 74416 1 1853
2 74417 1 1854
2 74418 1 1854
2 74419 1 1854
2 74420 1 1854
2 74421 1 1854
2 74422 1 1854
2 74423 1 1863
2 74424 1 1863
2 74425 1 1869
2 74426 1 1869
2 74427 1 1869
2 74428 1 1869
2 74429 1 1869
2 74430 1 1870
2 74431 1 1870
2 74432 1 1870
2 74433 1 1870
2 74434 1 1871
2 74435 1 1871
2 74436 1 1871
2 74437 1 1871
2 74438 1 1871
2 74439 1 1871
2 74440 1 1871
2 74441 1 1871
2 74442 1 1872
2 74443 1 1872
2 74444 1 1880
2 74445 1 1880
2 74446 1 1881
2 74447 1 1881
2 74448 1 1887
2 74449 1 1887
2 74450 1 1887
2 74451 1 1887
2 74452 1 1887
2 74453 1 1887
2 74454 1 1887
2 74455 1 1887
2 74456 1 1888
2 74457 1 1888
2 74458 1 1888
2 74459 1 1888
2 74460 1 1888
2 74461 1 1888
2 74462 1 1890
2 74463 1 1890
2 74464 1 1893
2 74465 1 1893
2 74466 1 1893
2 74467 1 1893
2 74468 1 1893
2 74469 1 1893
2 74470 1 1893
2 74471 1 1893
2 74472 1 1894
2 74473 1 1894
2 74474 1 1894
2 74475 1 1895
2 74476 1 1895
2 74477 1 1895
2 74478 1 1895
2 74479 1 1895
2 74480 1 1895
2 74481 1 1895
2 74482 1 1895
2 74483 1 1895
2 74484 1 1895
2 74485 1 1904
2 74486 1 1904
2 74487 1 1904
2 74488 1 1904
2 74489 1 1907
2 74490 1 1907
2 74491 1 1907
2 74492 1 1907
2 74493 1 1908
2 74494 1 1908
2 74495 1 1909
2 74496 1 1909
2 74497 1 1909
2 74498 1 1909
2 74499 1 1909
2 74500 1 1910
2 74501 1 1910
2 74502 1 1910
2 74503 1 1910
2 74504 1 1918
2 74505 1 1918
2 74506 1 1918
2 74507 1 1918
2 74508 1 1918
2 74509 1 1918
2 74510 1 1918
2 74511 1 1918
2 74512 1 1918
2 74513 1 1918
2 74514 1 1918
2 74515 1 1918
2 74516 1 1918
2 74517 1 1918
2 74518 1 1918
2 74519 1 1918
2 74520 1 1918
2 74521 1 1919
2 74522 1 1919
2 74523 1 1920
2 74524 1 1920
2 74525 1 1935
2 74526 1 1935
2 74527 1 1935
2 74528 1 1935
2 74529 1 1935
2 74530 1 1935
2 74531 1 1935
2 74532 1 1935
2 74533 1 1935
2 74534 1 1935
2 74535 1 1935
2 74536 1 1935
2 74537 1 1935
2 74538 1 1935
2 74539 1 1935
2 74540 1 1935
2 74541 1 1935
2 74542 1 1935
2 74543 1 1935
2 74544 1 1935
2 74545 1 1935
2 74546 1 1935
2 74547 1 1936
2 74548 1 1936
2 74549 1 1936
2 74550 1 1936
2 74551 1 1936
2 74552 1 1936
2 74553 1 1936
2 74554 1 1937
2 74555 1 1937
2 74556 1 1937
2 74557 1 1937
2 74558 1 1947
2 74559 1 1947
2 74560 1 1947
2 74561 1 1947
2 74562 1 1969
2 74563 1 1969
2 74564 1 1969
2 74565 1 1979
2 74566 1 1979
2 74567 1 1979
2 74568 1 1979
2 74569 1 1979
2 74570 1 1979
2 74571 1 1981
2 74572 1 1981
2 74573 1 1982
2 74574 1 1982
2 74575 1 1991
2 74576 1 1991
2 74577 1 1991
2 74578 1 1991
2 74579 1 1991
2 74580 1 1991
2 74581 1 1991
2 74582 1 1993
2 74583 1 1993
2 74584 1 1994
2 74585 1 1994
2 74586 1 1994
2 74587 1 1994
2 74588 1 1994
2 74589 1 1994
2 74590 1 1994
2 74591 1 1994
2 74592 1 1994
2 74593 1 1997
2 74594 1 1997
2 74595 1 2004
2 74596 1 2004
2 74597 1 2004
2 74598 1 2004
2 74599 1 2004
2 74600 1 2005
2 74601 1 2005
2 74602 1 2005
2 74603 1 2005
2 74604 1 2006
2 74605 1 2006
2 74606 1 2012
2 74607 1 2012
2 74608 1 2012
2 74609 1 2013
2 74610 1 2013
2 74611 1 2013
2 74612 1 2013
2 74613 1 2013
2 74614 1 2030
2 74615 1 2030
2 74616 1 2030
2 74617 1 2030
2 74618 1 2032
2 74619 1 2032
2 74620 1 2033
2 74621 1 2033
2 74622 1 2033
2 74623 1 2042
2 74624 1 2042
2 74625 1 2045
2 74626 1 2045
2 74627 1 2045
2 74628 1 2045
2 74629 1 2045
2 74630 1 2045
2 74631 1 2045
2 74632 1 2046
2 74633 1 2046
2 74634 1 2046
2 74635 1 2046
2 74636 1 2046
2 74637 1 2046
2 74638 1 2046
2 74639 1 2048
2 74640 1 2048
2 74641 1 2063
2 74642 1 2063
2 74643 1 2063
2 74644 1 2063
2 74645 1 2069
2 74646 1 2069
2 74647 1 2072
2 74648 1 2072
2 74649 1 2072
2 74650 1 2072
2 74651 1 2076
2 74652 1 2076
2 74653 1 2076
2 74654 1 2076
2 74655 1 2076
2 74656 1 2076
2 74657 1 2076
2 74658 1 2076
2 74659 1 2076
2 74660 1 2078
2 74661 1 2078
2 74662 1 2078
2 74663 1 2078
2 74664 1 2078
2 74665 1 2078
2 74666 1 2078
2 74667 1 2078
2 74668 1 2078
2 74669 1 2078
2 74670 1 2096
2 74671 1 2096
2 74672 1 2099
2 74673 1 2099
2 74674 1 2099
2 74675 1 2099
2 74676 1 2099
2 74677 1 2100
2 74678 1 2100
2 74679 1 2100
2 74680 1 2102
2 74681 1 2102
2 74682 1 2105
2 74683 1 2105
2 74684 1 2105
2 74685 1 2105
2 74686 1 2105
2 74687 1 2105
2 74688 1 2105
2 74689 1 2105
2 74690 1 2105
2 74691 1 2105
2 74692 1 2106
2 74693 1 2106
2 74694 1 2106
2 74695 1 2106
2 74696 1 2106
2 74697 1 2106
2 74698 1 2108
2 74699 1 2108
2 74700 1 2108
2 74701 1 2108
2 74702 1 2108
2 74703 1 2108
2 74704 1 2109
2 74705 1 2109
2 74706 1 2111
2 74707 1 2111
2 74708 1 2112
2 74709 1 2112
2 74710 1 2115
2 74711 1 2115
2 74712 1 2123
2 74713 1 2123
2 74714 1 2138
2 74715 1 2138
2 74716 1 2139
2 74717 1 2139
2 74718 1 2143
2 74719 1 2143
2 74720 1 2149
2 74721 1 2149
2 74722 1 2165
2 74723 1 2165
2 74724 1 2165
2 74725 1 2165
2 74726 1 2165
2 74727 1 2165
2 74728 1 2165
2 74729 1 2165
2 74730 1 2166
2 74731 1 2166
2 74732 1 2166
2 74733 1 2173
2 74734 1 2173
2 74735 1 2175
2 74736 1 2175
2 74737 1 2175
2 74738 1 2175
2 74739 1 2176
2 74740 1 2176
2 74741 1 2176
2 74742 1 2178
2 74743 1 2178
2 74744 1 2178
2 74745 1 2178
2 74746 1 2179
2 74747 1 2179
2 74748 1 2179
2 74749 1 2179
2 74750 1 2179
2 74751 1 2179
2 74752 1 2180
2 74753 1 2180
2 74754 1 2205
2 74755 1 2205
2 74756 1 2205
2 74757 1 2216
2 74758 1 2216
2 74759 1 2216
2 74760 1 2216
2 74761 1 2216
2 74762 1 2216
2 74763 1 2216
2 74764 1 2216
2 74765 1 2226
2 74766 1 2226
2 74767 1 2231
2 74768 1 2231
2 74769 1 2232
2 74770 1 2232
2 74771 1 2232
2 74772 1 2232
2 74773 1 2232
2 74774 1 2232
2 74775 1 2233
2 74776 1 2233
2 74777 1 2234
2 74778 1 2234
2 74779 1 2235
2 74780 1 2235
2 74781 1 2235
2 74782 1 2235
2 74783 1 2235
2 74784 1 2236
2 74785 1 2236
2 74786 1 2236
2 74787 1 2237
2 74788 1 2237
2 74789 1 2240
2 74790 1 2240
2 74791 1 2248
2 74792 1 2248
2 74793 1 2248
2 74794 1 2248
2 74795 1 2248
2 74796 1 2248
2 74797 1 2248
2 74798 1 2249
2 74799 1 2249
2 74800 1 2249
2 74801 1 2250
2 74802 1 2250
2 74803 1 2250
2 74804 1 2250
2 74805 1 2250
2 74806 1 2250
2 74807 1 2250
2 74808 1 2250
2 74809 1 2250
2 74810 1 2250
2 74811 1 2250
2 74812 1 2250
2 74813 1 2250
2 74814 1 2250
2 74815 1 2250
2 74816 1 2251
2 74817 1 2251
2 74818 1 2251
2 74819 1 2251
2 74820 1 2251
2 74821 1 2252
2 74822 1 2252
2 74823 1 2252
2 74824 1 2252
2 74825 1 2252
2 74826 1 2252
2 74827 1 2252
2 74828 1 2253
2 74829 1 2253
2 74830 1 2260
2 74831 1 2260
2 74832 1 2260
2 74833 1 2260
2 74834 1 2260
2 74835 1 2260
2 74836 1 2260
2 74837 1 2260
2 74838 1 2260
2 74839 1 2260
2 74840 1 2260
2 74841 1 2260
2 74842 1 2261
2 74843 1 2261
2 74844 1 2262
2 74845 1 2262
2 74846 1 2262
2 74847 1 2262
2 74848 1 2262
2 74849 1 2262
2 74850 1 2262
2 74851 1 2264
2 74852 1 2264
2 74853 1 2265
2 74854 1 2265
2 74855 1 2265
2 74856 1 2270
2 74857 1 2270
2 74858 1 2270
2 74859 1 2270
2 74860 1 2270
2 74861 1 2270
2 74862 1 2270
2 74863 1 2271
2 74864 1 2271
2 74865 1 2271
2 74866 1 2271
2 74867 1 2271
2 74868 1 2271
2 74869 1 2271
2 74870 1 2271
2 74871 1 2271
2 74872 1 2271
2 74873 1 2271
2 74874 1 2271
2 74875 1 2271
2 74876 1 2271
2 74877 1 2271
2 74878 1 2271
2 74879 1 2272
2 74880 1 2272
2 74881 1 2272
2 74882 1 2272
2 74883 1 2273
2 74884 1 2273
2 74885 1 2282
2 74886 1 2282
2 74887 1 2282
2 74888 1 2282
2 74889 1 2282
2 74890 1 2282
2 74891 1 2282
2 74892 1 2282
2 74893 1 2283
2 74894 1 2283
2 74895 1 2283
2 74896 1 2283
2 74897 1 2283
2 74898 1 2283
2 74899 1 2284
2 74900 1 2284
2 74901 1 2287
2 74902 1 2287
2 74903 1 2287
2 74904 1 2287
2 74905 1 2287
2 74906 1 2287
2 74907 1 2287
2 74908 1 2287
2 74909 1 2287
2 74910 1 2287
2 74911 1 2289
2 74912 1 2289
2 74913 1 2289
2 74914 1 2289
2 74915 1 2289
2 74916 1 2289
2 74917 1 2289
2 74918 1 2303
2 74919 1 2303
2 74920 1 2303
2 74921 1 2303
2 74922 1 2314
2 74923 1 2314
2 74924 1 2329
2 74925 1 2329
2 74926 1 2329
2 74927 1 2329
2 74928 1 2329
2 74929 1 2329
2 74930 1 2330
2 74931 1 2330
2 74932 1 2331
2 74933 1 2331
2 74934 1 2331
2 74935 1 2332
2 74936 1 2332
2 74937 1 2332
2 74938 1 2332
2 74939 1 2332
2 74940 1 2332
2 74941 1 2332
2 74942 1 2332
2 74943 1 2332
2 74944 1 2332
2 74945 1 2332
2 74946 1 2333
2 74947 1 2333
2 74948 1 2334
2 74949 1 2334
2 74950 1 2334
2 74951 1 2334
2 74952 1 2336
2 74953 1 2336
2 74954 1 2340
2 74955 1 2340
2 74956 1 2340
2 74957 1 2347
2 74958 1 2347
2 74959 1 2354
2 74960 1 2354
2 74961 1 2354
2 74962 1 2354
2 74963 1 2354
2 74964 1 2354
2 74965 1 2354
2 74966 1 2355
2 74967 1 2355
2 74968 1 2356
2 74969 1 2356
2 74970 1 2356
2 74971 1 2356
2 74972 1 2356
2 74973 1 2356
2 74974 1 2356
2 74975 1 2356
2 74976 1 2356
2 74977 1 2356
2 74978 1 2356
2 74979 1 2356
2 74980 1 2356
2 74981 1 2356
2 74982 1 2356
2 74983 1 2356
2 74984 1 2356
2 74985 1 2356
2 74986 1 2356
2 74987 1 2356
2 74988 1 2356
2 74989 1 2356
2 74990 1 2356
2 74991 1 2356
2 74992 1 2356
2 74993 1 2356
2 74994 1 2356
2 74995 1 2356
2 74996 1 2356
2 74997 1 2356
2 74998 1 2356
2 74999 1 2357
2 75000 1 2357
2 75001 1 2357
2 75002 1 2357
2 75003 1 2357
2 75004 1 2357
2 75005 1 2357
2 75006 1 2357
2 75007 1 2357
2 75008 1 2357
2 75009 1 2357
2 75010 1 2357
2 75011 1 2357
2 75012 1 2357
2 75013 1 2359
2 75014 1 2359
2 75015 1 2360
2 75016 1 2360
2 75017 1 2360
2 75018 1 2360
2 75019 1 2360
2 75020 1 2360
2 75021 1 2360
2 75022 1 2360
2 75023 1 2360
2 75024 1 2360
2 75025 1 2360
2 75026 1 2361
2 75027 1 2361
2 75028 1 2361
2 75029 1 2361
2 75030 1 2362
2 75031 1 2362
2 75032 1 2362
2 75033 1 2362
2 75034 1 2363
2 75035 1 2363
2 75036 1 2363
2 75037 1 2363
2 75038 1 2363
2 75039 1 2363
2 75040 1 2363
2 75041 1 2368
2 75042 1 2368
2 75043 1 2368
2 75044 1 2368
2 75045 1 2369
2 75046 1 2369
2 75047 1 2370
2 75048 1 2370
2 75049 1 2370
2 75050 1 2370
2 75051 1 2371
2 75052 1 2371
2 75053 1 2372
2 75054 1 2372
2 75055 1 2372
2 75056 1 2386
2 75057 1 2386
2 75058 1 2386
2 75059 1 2386
2 75060 1 2389
2 75061 1 2389
2 75062 1 2389
2 75063 1 2389
2 75064 1 2389
2 75065 1 2389
2 75066 1 2390
2 75067 1 2390
2 75068 1 2392
2 75069 1 2392
2 75070 1 2393
2 75071 1 2393
2 75072 1 2393
2 75073 1 2393
2 75074 1 2393
2 75075 1 2393
2 75076 1 2393
2 75077 1 2394
2 75078 1 2394
2 75079 1 2395
2 75080 1 2395
2 75081 1 2395
2 75082 1 2397
2 75083 1 2397
2 75084 1 2397
2 75085 1 2411
2 75086 1 2411
2 75087 1 2411
2 75088 1 2411
2 75089 1 2411
2 75090 1 2411
2 75091 1 2415
2 75092 1 2415
2 75093 1 2416
2 75094 1 2416
2 75095 1 2416
2 75096 1 2417
2 75097 1 2417
2 75098 1 2417
2 75099 1 2417
2 75100 1 2417
2 75101 1 2417
2 75102 1 2417
2 75103 1 2417
2 75104 1 2418
2 75105 1 2418
2 75106 1 2418
2 75107 1 2418
2 75108 1 2418
2 75109 1 2419
2 75110 1 2419
2 75111 1 2419
2 75112 1 2419
2 75113 1 2419
2 75114 1 2419
2 75115 1 2420
2 75116 1 2420
2 75117 1 2428
2 75118 1 2428
2 75119 1 2428
2 75120 1 2434
2 75121 1 2434
2 75122 1 2434
2 75123 1 2434
2 75124 1 2434
2 75125 1 2434
2 75126 1 2434
2 75127 1 2434
2 75128 1 2434
2 75129 1 2434
2 75130 1 2434
2 75131 1 2434
2 75132 1 2434
2 75133 1 2434
2 75134 1 2443
2 75135 1 2443
2 75136 1 2443
2 75137 1 2443
2 75138 1 2443
2 75139 1 2443
2 75140 1 2443
2 75141 1 2443
2 75142 1 2443
2 75143 1 2443
2 75144 1 2443
2 75145 1 2443
2 75146 1 2443
2 75147 1 2443
2 75148 1 2443
2 75149 1 2443
2 75150 1 2444
2 75151 1 2444
2 75152 1 2444
2 75153 1 2444
2 75154 1 2444
2 75155 1 2444
2 75156 1 2455
2 75157 1 2455
2 75158 1 2456
2 75159 1 2456
2 75160 1 2456
2 75161 1 2464
2 75162 1 2464
2 75163 1 2476
2 75164 1 2476
2 75165 1 2476
2 75166 1 2476
2 75167 1 2476
2 75168 1 2476
2 75169 1 2476
2 75170 1 2476
2 75171 1 2476
2 75172 1 2476
2 75173 1 2476
2 75174 1 2476
2 75175 1 2476
2 75176 1 2476
2 75177 1 2476
2 75178 1 2477
2 75179 1 2477
2 75180 1 2477
2 75181 1 2477
2 75182 1 2477
2 75183 1 2477
2 75184 1 2477
2 75185 1 2477
2 75186 1 2477
2 75187 1 2477
2 75188 1 2477
2 75189 1 2477
2 75190 1 2477
2 75191 1 2477
2 75192 1 2477
2 75193 1 2477
2 75194 1 2477
2 75195 1 2478
2 75196 1 2478
2 75197 1 2479
2 75198 1 2479
2 75199 1 2479
2 75200 1 2479
2 75201 1 2479
2 75202 1 2479
2 75203 1 2479
2 75204 1 2479
2 75205 1 2479
2 75206 1 2479
2 75207 1 2479
2 75208 1 2480
2 75209 1 2480
2 75210 1 2480
2 75211 1 2480
2 75212 1 2495
2 75213 1 2495
2 75214 1 2495
2 75215 1 2495
2 75216 1 2495
2 75217 1 2495
2 75218 1 2495
2 75219 1 2495
2 75220 1 2496
2 75221 1 2496
2 75222 1 2498
2 75223 1 2498
2 75224 1 2499
2 75225 1 2499
2 75226 1 2501
2 75227 1 2501
2 75228 1 2503
2 75229 1 2503
2 75230 1 2503
2 75231 1 2503
2 75232 1 2503
2 75233 1 2503
2 75234 1 2503
2 75235 1 2505
2 75236 1 2505
2 75237 1 2505
2 75238 1 2505
2 75239 1 2505
2 75240 1 2505
2 75241 1 2505
2 75242 1 2505
2 75243 1 2508
2 75244 1 2508
2 75245 1 2508
2 75246 1 2508
2 75247 1 2508
2 75248 1 2512
2 75249 1 2512
2 75250 1 2530
2 75251 1 2530
2 75252 1 2530
2 75253 1 2530
2 75254 1 2530
2 75255 1 2530
2 75256 1 2530
2 75257 1 2530
2 75258 1 2531
2 75259 1 2531
2 75260 1 2531
2 75261 1 2531
2 75262 1 2531
2 75263 1 2531
2 75264 1 2531
2 75265 1 2531
2 75266 1 2531
2 75267 1 2532
2 75268 1 2532
2 75269 1 2532
2 75270 1 2532
2 75271 1 2532
2 75272 1 2532
2 75273 1 2532
2 75274 1 2532
2 75275 1 2532
2 75276 1 2532
2 75277 1 2532
2 75278 1 2532
2 75279 1 2533
2 75280 1 2533
2 75281 1 2533
2 75282 1 2533
2 75283 1 2533
2 75284 1 2533
2 75285 1 2533
2 75286 1 2533
2 75287 1 2533
2 75288 1 2533
2 75289 1 2535
2 75290 1 2535
2 75291 1 2535
2 75292 1 2535
2 75293 1 2538
2 75294 1 2538
2 75295 1 2543
2 75296 1 2543
2 75297 1 2543
2 75298 1 2543
2 75299 1 2543
2 75300 1 2543
2 75301 1 2545
2 75302 1 2545
2 75303 1 2545
2 75304 1 2545
2 75305 1 2545
2 75306 1 2546
2 75307 1 2546
2 75308 1 2546
2 75309 1 2553
2 75310 1 2553
2 75311 1 2553
2 75312 1 2555
2 75313 1 2555
2 75314 1 2564
2 75315 1 2564
2 75316 1 2564
2 75317 1 2564
2 75318 1 2564
2 75319 1 2564
2 75320 1 2564
2 75321 1 2564
2 75322 1 2564
2 75323 1 2564
2 75324 1 2564
2 75325 1 2564
2 75326 1 2564
2 75327 1 2564
2 75328 1 2564
2 75329 1 2564
2 75330 1 2564
2 75331 1 2564
2 75332 1 2564
2 75333 1 2564
2 75334 1 2564
2 75335 1 2564
2 75336 1 2564
2 75337 1 2564
2 75338 1 2564
2 75339 1 2564
2 75340 1 2564
2 75341 1 2564
2 75342 1 2564
2 75343 1 2568
2 75344 1 2568
2 75345 1 2575
2 75346 1 2575
2 75347 1 2577
2 75348 1 2577
2 75349 1 2582
2 75350 1 2582
2 75351 1 2582
2 75352 1 2582
2 75353 1 2583
2 75354 1 2583
2 75355 1 2584
2 75356 1 2584
2 75357 1 2584
2 75358 1 2584
2 75359 1 2584
2 75360 1 2584
2 75361 1 2585
2 75362 1 2585
2 75363 1 2592
2 75364 1 2592
2 75365 1 2597
2 75366 1 2597
2 75367 1 2603
2 75368 1 2603
2 75369 1 2603
2 75370 1 2603
2 75371 1 2604
2 75372 1 2604
2 75373 1 2604
2 75374 1 2604
2 75375 1 2604
2 75376 1 2604
2 75377 1 2604
2 75378 1 2608
2 75379 1 2608
2 75380 1 2622
2 75381 1 2622
2 75382 1 2622
2 75383 1 2626
2 75384 1 2626
2 75385 1 2627
2 75386 1 2627
2 75387 1 2627
2 75388 1 2628
2 75389 1 2628
2 75390 1 2628
2 75391 1 2628
2 75392 1 2628
2 75393 1 2628
2 75394 1 2628
2 75395 1 2628
2 75396 1 2628
2 75397 1 2628
2 75398 1 2628
2 75399 1 2628
2 75400 1 2628
2 75401 1 2628
2 75402 1 2628
2 75403 1 2628
2 75404 1 2628
2 75405 1 2629
2 75406 1 2629
2 75407 1 2629
2 75408 1 2629
2 75409 1 2630
2 75410 1 2630
2 75411 1 2630
2 75412 1 2631
2 75413 1 2631
2 75414 1 2646
2 75415 1 2646
2 75416 1 2649
2 75417 1 2649
2 75418 1 2649
2 75419 1 2649
2 75420 1 2649
2 75421 1 2650
2 75422 1 2650
2 75423 1 2650
2 75424 1 2650
2 75425 1 2650
2 75426 1 2662
2 75427 1 2662
2 75428 1 2662
2 75429 1 2662
2 75430 1 2662
2 75431 1 2662
2 75432 1 2662
2 75433 1 2662
2 75434 1 2662
2 75435 1 2662
2 75436 1 2662
2 75437 1 2662
2 75438 1 2662
2 75439 1 2662
2 75440 1 2662
2 75441 1 2662
2 75442 1 2662
2 75443 1 2662
2 75444 1 2662
2 75445 1 2662
2 75446 1 2662
2 75447 1 2662
2 75448 1 2662
2 75449 1 2662
2 75450 1 2662
2 75451 1 2663
2 75452 1 2663
2 75453 1 2663
2 75454 1 2663
2 75455 1 2663
2 75456 1 2663
2 75457 1 2663
2 75458 1 2663
2 75459 1 2664
2 75460 1 2664
2 75461 1 2664
2 75462 1 2664
2 75463 1 2664
2 75464 1 2664
2 75465 1 2664
2 75466 1 2664
2 75467 1 2664
2 75468 1 2664
2 75469 1 2664
2 75470 1 2664
2 75471 1 2666
2 75472 1 2666
2 75473 1 2666
2 75474 1 2667
2 75475 1 2667
2 75476 1 2669
2 75477 1 2669
2 75478 1 2669
2 75479 1 2669
2 75480 1 2669
2 75481 1 2669
2 75482 1 2669
2 75483 1 2669
2 75484 1 2669
2 75485 1 2669
2 75486 1 2669
2 75487 1 2669
2 75488 1 2669
2 75489 1 2669
2 75490 1 2670
2 75491 1 2670
2 75492 1 2670
2 75493 1 2670
2 75494 1 2670
2 75495 1 2694
2 75496 1 2694
2 75497 1 2694
2 75498 1 2694
2 75499 1 2694
2 75500 1 2694
2 75501 1 2694
2 75502 1 2694
2 75503 1 2694
2 75504 1 2694
2 75505 1 2694
2 75506 1 2694
2 75507 1 2694
2 75508 1 2694
2 75509 1 2694
2 75510 1 2694
2 75511 1 2694
2 75512 1 2694
2 75513 1 2694
2 75514 1 2694
2 75515 1 2694
2 75516 1 2694
2 75517 1 2694
2 75518 1 2694
2 75519 1 2694
2 75520 1 2694
2 75521 1 2694
2 75522 1 2694
2 75523 1 2694
2 75524 1 2694
2 75525 1 2694
2 75526 1 2694
2 75527 1 2694
2 75528 1 2694
2 75529 1 2694
2 75530 1 2694
2 75531 1 2694
2 75532 1 2694
2 75533 1 2694
2 75534 1 2694
2 75535 1 2694
2 75536 1 2694
2 75537 1 2694
2 75538 1 2694
2 75539 1 2694
2 75540 1 2694
2 75541 1 2694
2 75542 1 2694
2 75543 1 2694
2 75544 1 2694
2 75545 1 2694
2 75546 1 2694
2 75547 1 2694
2 75548 1 2694
2 75549 1 2694
2 75550 1 2694
2 75551 1 2694
2 75552 1 2694
2 75553 1 2694
2 75554 1 2694
2 75555 1 2694
2 75556 1 2694
2 75557 1 2694
2 75558 1 2694
2 75559 1 2694
2 75560 1 2694
2 75561 1 2694
2 75562 1 2694
2 75563 1 2694
2 75564 1 2694
2 75565 1 2694
2 75566 1 2695
2 75567 1 2695
2 75568 1 2695
2 75569 1 2695
2 75570 1 2695
2 75571 1 2695
2 75572 1 2695
2 75573 1 2695
2 75574 1 2695
2 75575 1 2695
2 75576 1 2695
2 75577 1 2695
2 75578 1 2695
2 75579 1 2695
2 75580 1 2695
2 75581 1 2695
2 75582 1 2695
2 75583 1 2695
2 75584 1 2695
2 75585 1 2695
2 75586 1 2695
2 75587 1 2695
2 75588 1 2695
2 75589 1 2695
2 75590 1 2695
2 75591 1 2695
2 75592 1 2695
2 75593 1 2695
2 75594 1 2695
2 75595 1 2695
2 75596 1 2695
2 75597 1 2695
2 75598 1 2695
2 75599 1 2695
2 75600 1 2695
2 75601 1 2695
2 75602 1 2695
2 75603 1 2695
2 75604 1 2695
2 75605 1 2695
2 75606 1 2695
2 75607 1 2696
2 75608 1 2696
2 75609 1 2696
2 75610 1 2696
2 75611 1 2696
2 75612 1 2696
2 75613 1 2696
2 75614 1 2696
2 75615 1 2696
2 75616 1 2696
2 75617 1 2696
2 75618 1 2696
2 75619 1 2696
2 75620 1 2696
2 75621 1 2696
2 75622 1 2696
2 75623 1 2696
2 75624 1 2696
2 75625 1 2696
2 75626 1 2696
2 75627 1 2696
2 75628 1 2696
2 75629 1 2696
2 75630 1 2696
2 75631 1 2696
2 75632 1 2696
2 75633 1 2696
2 75634 1 2696
2 75635 1 2696
2 75636 1 2696
2 75637 1 2696
2 75638 1 2696
2 75639 1 2696
2 75640 1 2696
2 75641 1 2696
2 75642 1 2696
2 75643 1 2696
2 75644 1 2696
2 75645 1 2696
2 75646 1 2696
2 75647 1 2696
2 75648 1 2696
2 75649 1 2696
2 75650 1 2696
2 75651 1 2696
2 75652 1 2696
2 75653 1 2696
2 75654 1 2696
2 75655 1 2696
2 75656 1 2696
2 75657 1 2696
2 75658 1 2696
2 75659 1 2696
2 75660 1 2696
2 75661 1 2696
2 75662 1 2696
2 75663 1 2696
2 75664 1 2696
2 75665 1 2696
2 75666 1 2696
2 75667 1 2696
2 75668 1 2697
2 75669 1 2697
2 75670 1 2697
2 75671 1 2697
2 75672 1 2697
2 75673 1 2698
2 75674 1 2698
2 75675 1 2699
2 75676 1 2699
2 75677 1 2706
2 75678 1 2706
2 75679 1 2706
2 75680 1 2706
2 75681 1 2706
2 75682 1 2706
2 75683 1 2706
2 75684 1 2706
2 75685 1 2706
2 75686 1 2706
2 75687 1 2706
2 75688 1 2706
2 75689 1 2707
2 75690 1 2707
2 75691 1 2707
2 75692 1 2707
2 75693 1 2707
2 75694 1 2707
2 75695 1 2708
2 75696 1 2708
2 75697 1 2708
2 75698 1 2708
2 75699 1 2709
2 75700 1 2709
2 75701 1 2709
2 75702 1 2709
2 75703 1 2709
2 75704 1 2709
2 75705 1 2709
2 75706 1 2710
2 75707 1 2710
2 75708 1 2710
2 75709 1 2710
2 75710 1 2710
2 75711 1 2710
2 75712 1 2710
2 75713 1 2710
2 75714 1 2710
2 75715 1 2710
2 75716 1 2710
2 75717 1 2710
2 75718 1 2710
2 75719 1 2710
2 75720 1 2710
2 75721 1 2711
2 75722 1 2711
2 75723 1 2711
2 75724 1 2712
2 75725 1 2712
2 75726 1 2712
2 75727 1 2712
2 75728 1 2712
2 75729 1 2712
2 75730 1 2712
2 75731 1 2712
2 75732 1 2712
2 75733 1 2712
2 75734 1 2712
2 75735 1 2712
2 75736 1 2712
2 75737 1 2712
2 75738 1 2712
2 75739 1 2712
2 75740 1 2712
2 75741 1 2712
2 75742 1 2712
2 75743 1 2713
2 75744 1 2713
2 75745 1 2713
2 75746 1 2713
2 75747 1 2713
2 75748 1 2713
2 75749 1 2713
2 75750 1 2713
2 75751 1 2713
2 75752 1 2713
2 75753 1 2713
2 75754 1 2713
2 75755 1 2713
2 75756 1 2713
2 75757 1 2713
2 75758 1 2713
2 75759 1 2713
2 75760 1 2713
2 75761 1 2713
2 75762 1 2713
2 75763 1 2713
2 75764 1 2713
2 75765 1 2713
2 75766 1 2713
2 75767 1 2713
2 75768 1 2713
2 75769 1 2713
2 75770 1 2713
2 75771 1 2720
2 75772 1 2720
2 75773 1 2720
2 75774 1 2720
2 75775 1 2720
2 75776 1 2720
2 75777 1 2721
2 75778 1 2721
2 75779 1 2721
2 75780 1 2721
2 75781 1 2721
2 75782 1 2721
2 75783 1 2721
2 75784 1 2721
2 75785 1 2721
2 75786 1 2721
2 75787 1 2721
2 75788 1 2721
2 75789 1 2721
2 75790 1 2721
2 75791 1 2721
2 75792 1 2721
2 75793 1 2721
2 75794 1 2722
2 75795 1 2722
2 75796 1 2722
2 75797 1 2723
2 75798 1 2723
2 75799 1 2723
2 75800 1 2724
2 75801 1 2724
2 75802 1 2724
2 75803 1 2724
2 75804 1 2724
2 75805 1 2724
2 75806 1 2724
2 75807 1 2724
2 75808 1 2724
2 75809 1 2724
2 75810 1 2724
2 75811 1 2725
2 75812 1 2725
2 75813 1 2726
2 75814 1 2726
2 75815 1 2728
2 75816 1 2728
2 75817 1 2728
2 75818 1 2731
2 75819 1 2731
2 75820 1 2731
2 75821 1 2731
2 75822 1 2731
2 75823 1 2732
2 75824 1 2732
2 75825 1 2732
2 75826 1 2732
2 75827 1 2733
2 75828 1 2733
2 75829 1 2733
2 75830 1 2736
2 75831 1 2736
2 75832 1 2744
2 75833 1 2744
2 75834 1 2745
2 75835 1 2745
2 75836 1 2745
2 75837 1 2745
2 75838 1 2745
2 75839 1 2745
2 75840 1 2745
2 75841 1 2745
2 75842 1 2745
2 75843 1 2745
2 75844 1 2746
2 75845 1 2746
2 75846 1 2746
2 75847 1 2746
2 75848 1 2746
2 75849 1 2746
2 75850 1 2746
2 75851 1 2746
2 75852 1 2746
2 75853 1 2747
2 75854 1 2747
2 75855 1 2747
2 75856 1 2747
2 75857 1 2747
2 75858 1 2747
2 75859 1 2747
2 75860 1 2747
2 75861 1 2747
2 75862 1 2747
2 75863 1 2747
2 75864 1 2747
2 75865 1 2747
2 75866 1 2747
2 75867 1 2747
2 75868 1 2747
2 75869 1 2747
2 75870 1 2747
2 75871 1 2747
2 75872 1 2747
2 75873 1 2747
2 75874 1 2747
2 75875 1 2747
2 75876 1 2747
2 75877 1 2747
2 75878 1 2747
2 75879 1 2747
2 75880 1 2747
2 75881 1 2747
2 75882 1 2747
2 75883 1 2747
2 75884 1 2747
2 75885 1 2747
2 75886 1 2747
2 75887 1 2747
2 75888 1 2749
2 75889 1 2749
2 75890 1 2749
2 75891 1 2749
2 75892 1 2751
2 75893 1 2751
2 75894 1 2751
2 75895 1 2751
2 75896 1 2752
2 75897 1 2752
2 75898 1 2752
2 75899 1 2752
2 75900 1 2752
2 75901 1 2752
2 75902 1 2752
2 75903 1 2752
2 75904 1 2752
2 75905 1 2752
2 75906 1 2752
2 75907 1 2752
2 75908 1 2752
2 75909 1 2752
2 75910 1 2752
2 75911 1 2752
2 75912 1 2752
2 75913 1 2752
2 75914 1 2752
2 75915 1 2752
2 75916 1 2753
2 75917 1 2753
2 75918 1 2753
2 75919 1 2753
2 75920 1 2754
2 75921 1 2754
2 75922 1 2756
2 75923 1 2756
2 75924 1 2756
2 75925 1 2756
2 75926 1 2756
2 75927 1 2756
2 75928 1 2756
2 75929 1 2760
2 75930 1 2760
2 75931 1 2771
2 75932 1 2771
2 75933 1 2771
2 75934 1 2771
2 75935 1 2771
2 75936 1 2772
2 75937 1 2772
2 75938 1 2772
2 75939 1 2772
2 75940 1 2772
2 75941 1 2772
2 75942 1 2772
2 75943 1 2772
2 75944 1 2772
2 75945 1 2772
2 75946 1 2772
2 75947 1 2772
2 75948 1 2781
2 75949 1 2781
2 75950 1 2781
2 75951 1 2781
2 75952 1 2781
2 75953 1 2781
2 75954 1 2781
2 75955 1 2781
2 75956 1 2781
2 75957 1 2781
2 75958 1 2781
2 75959 1 2781
2 75960 1 2781
2 75961 1 2781
2 75962 1 2781
2 75963 1 2781
2 75964 1 2781
2 75965 1 2781
2 75966 1 2781
2 75967 1 2782
2 75968 1 2782
2 75969 1 2782
2 75970 1 2782
2 75971 1 2782
2 75972 1 2782
2 75973 1 2782
2 75974 1 2782
2 75975 1 2782
2 75976 1 2782
2 75977 1 2782
2 75978 1 2782
2 75979 1 2782
2 75980 1 2782
2 75981 1 2782
2 75982 1 2782
2 75983 1 2782
2 75984 1 2782
2 75985 1 2782
2 75986 1 2782
2 75987 1 2782
2 75988 1 2782
2 75989 1 2783
2 75990 1 2783
2 75991 1 2783
2 75992 1 2783
2 75993 1 2783
2 75994 1 2783
2 75995 1 2783
2 75996 1 2783
2 75997 1 2783
2 75998 1 2783
2 75999 1 2783
2 76000 1 2783
2 76001 1 2783
2 76002 1 2783
2 76003 1 2783
2 76004 1 2783
2 76005 1 2783
2 76006 1 2785
2 76007 1 2785
2 76008 1 2787
2 76009 1 2787
2 76010 1 2792
2 76011 1 2792
2 76012 1 2792
2 76013 1 2792
2 76014 1 2792
2 76015 1 2793
2 76016 1 2793
2 76017 1 2793
2 76018 1 2793
2 76019 1 2795
2 76020 1 2795
2 76021 1 2800
2 76022 1 2800
2 76023 1 2800
2 76024 1 2800
2 76025 1 2800
2 76026 1 2800
2 76027 1 2800
2 76028 1 2800
2 76029 1 2800
2 76030 1 2800
2 76031 1 2800
2 76032 1 2800
2 76033 1 2800
2 76034 1 2800
2 76035 1 2800
2 76036 1 2800
2 76037 1 2800
2 76038 1 2800
2 76039 1 2801
2 76040 1 2801
2 76041 1 2801
2 76042 1 2802
2 76043 1 2802
2 76044 1 2803
2 76045 1 2803
2 76046 1 2803
2 76047 1 2803
2 76048 1 2805
2 76049 1 2805
2 76050 1 2805
2 76051 1 2805
2 76052 1 2805
2 76053 1 2805
2 76054 1 2814
2 76055 1 2814
2 76056 1 2814
2 76057 1 2814
2 76058 1 2814
2 76059 1 2814
2 76060 1 2814
2 76061 1 2814
2 76062 1 2814
2 76063 1 2814
2 76064 1 2814
2 76065 1 2814
2 76066 1 2815
2 76067 1 2815
2 76068 1 2815
2 76069 1 2815
2 76070 1 2818
2 76071 1 2818
2 76072 1 2818
2 76073 1 2818
2 76074 1 2818
2 76075 1 2818
2 76076 1 2818
2 76077 1 2818
2 76078 1 2819
2 76079 1 2819
2 76080 1 2819
2 76081 1 2819
2 76082 1 2819
2 76083 1 2820
2 76084 1 2820
2 76085 1 2820
2 76086 1 2829
2 76087 1 2829
2 76088 1 2829
2 76089 1 2829
2 76090 1 2829
2 76091 1 2829
2 76092 1 2829
2 76093 1 2830
2 76094 1 2830
2 76095 1 2830
2 76096 1 2830
2 76097 1 2830
2 76098 1 2831
2 76099 1 2831
2 76100 1 2831
2 76101 1 2831
2 76102 1 2839
2 76103 1 2839
2 76104 1 2839
2 76105 1 2839
2 76106 1 2839
2 76107 1 2839
2 76108 1 2839
2 76109 1 2839
2 76110 1 2839
2 76111 1 2839
2 76112 1 2839
2 76113 1 2839
2 76114 1 2839
2 76115 1 2839
2 76116 1 2842
2 76117 1 2842
2 76118 1 2842
2 76119 1 2842
2 76120 1 2843
2 76121 1 2843
2 76122 1 2844
2 76123 1 2844
2 76124 1 2854
2 76125 1 2854
2 76126 1 2854
2 76127 1 2854
2 76128 1 2854
2 76129 1 2854
2 76130 1 2854
2 76131 1 2854
2 76132 1 2854
2 76133 1 2854
2 76134 1 2854
2 76135 1 2854
2 76136 1 2855
2 76137 1 2855
2 76138 1 2855
2 76139 1 2855
2 76140 1 2855
2 76141 1 2855
2 76142 1 2856
2 76143 1 2856
2 76144 1 2856
2 76145 1 2856
2 76146 1 2856
2 76147 1 2856
2 76148 1 2856
2 76149 1 2856
2 76150 1 2856
2 76151 1 2856
2 76152 1 2856
2 76153 1 2856
2 76154 1 2856
2 76155 1 2856
2 76156 1 2856
2 76157 1 2857
2 76158 1 2857
2 76159 1 2857
2 76160 1 2857
2 76161 1 2857
2 76162 1 2857
2 76163 1 2857
2 76164 1 2857
2 76165 1 2857
2 76166 1 2857
2 76167 1 2857
2 76168 1 2857
2 76169 1 2857
2 76170 1 2857
2 76171 1 2857
2 76172 1 2857
2 76173 1 2857
2 76174 1 2857
2 76175 1 2857
2 76176 1 2857
2 76177 1 2857
2 76178 1 2857
2 76179 1 2857
2 76180 1 2857
2 76181 1 2857
2 76182 1 2857
2 76183 1 2857
2 76184 1 2857
2 76185 1 2857
2 76186 1 2857
2 76187 1 2857
2 76188 1 2857
2 76189 1 2857
2 76190 1 2857
2 76191 1 2857
2 76192 1 2857
2 76193 1 2857
2 76194 1 2857
2 76195 1 2857
2 76196 1 2857
2 76197 1 2857
2 76198 1 2857
2 76199 1 2857
2 76200 1 2857
2 76201 1 2857
2 76202 1 2857
2 76203 1 2857
2 76204 1 2857
2 76205 1 2857
2 76206 1 2857
2 76207 1 2857
2 76208 1 2857
2 76209 1 2857
2 76210 1 2857
2 76211 1 2857
2 76212 1 2857
2 76213 1 2857
2 76214 1 2857
2 76215 1 2857
2 76216 1 2857
2 76217 1 2857
2 76218 1 2857
2 76219 1 2857
2 76220 1 2857
2 76221 1 2857
2 76222 1 2857
2 76223 1 2857
2 76224 1 2857
2 76225 1 2857
2 76226 1 2857
2 76227 1 2857
2 76228 1 2857
2 76229 1 2857
2 76230 1 2857
2 76231 1 2857
2 76232 1 2857
2 76233 1 2857
2 76234 1 2857
2 76235 1 2857
2 76236 1 2857
2 76237 1 2859
2 76238 1 2859
2 76239 1 2859
2 76240 1 2859
2 76241 1 2860
2 76242 1 2860
2 76243 1 2860
2 76244 1 2860
2 76245 1 2860
2 76246 1 2861
2 76247 1 2861
2 76248 1 2861
2 76249 1 2861
2 76250 1 2861
2 76251 1 2861
2 76252 1 2861
2 76253 1 2863
2 76254 1 2863
2 76255 1 2863
2 76256 1 2863
2 76257 1 2866
2 76258 1 2866
2 76259 1 2866
2 76260 1 2866
2 76261 1 2866
2 76262 1 2867
2 76263 1 2867
2 76264 1 2867
2 76265 1 2867
2 76266 1 2867
2 76267 1 2867
2 76268 1 2867
2 76269 1 2867
2 76270 1 2867
2 76271 1 2867
2 76272 1 2867
2 76273 1 2867
2 76274 1 2868
2 76275 1 2868
2 76276 1 2868
2 76277 1 2868
2 76278 1 2868
2 76279 1 2869
2 76280 1 2869
2 76281 1 2869
2 76282 1 2869
2 76283 1 2869
2 76284 1 2869
2 76285 1 2869
2 76286 1 2871
2 76287 1 2871
2 76288 1 2871
2 76289 1 2887
2 76290 1 2887
2 76291 1 2893
2 76292 1 2893
2 76293 1 2894
2 76294 1 2894
2 76295 1 2894
2 76296 1 2894
2 76297 1 2894
2 76298 1 2894
2 76299 1 2894
2 76300 1 2894
2 76301 1 2894
2 76302 1 2894
2 76303 1 2894
2 76304 1 2894
2 76305 1 2894
2 76306 1 2894
2 76307 1 2895
2 76308 1 2895
2 76309 1 2897
2 76310 1 2897
2 76311 1 2899
2 76312 1 2899
2 76313 1 2903
2 76314 1 2903
2 76315 1 2905
2 76316 1 2905
2 76317 1 2905
2 76318 1 2907
2 76319 1 2907
2 76320 1 2913
2 76321 1 2913
2 76322 1 2913
2 76323 1 2913
2 76324 1 2913
2 76325 1 2913
2 76326 1 2913
2 76327 1 2913
2 76328 1 2913
2 76329 1 2913
2 76330 1 2913
2 76331 1 2913
2 76332 1 2913
2 76333 1 2913
2 76334 1 2913
2 76335 1 2914
2 76336 1 2914
2 76337 1 2914
2 76338 1 2914
2 76339 1 2914
2 76340 1 2914
2 76341 1 2914
2 76342 1 2914
2 76343 1 2914
2 76344 1 2914
2 76345 1 2916
2 76346 1 2916
2 76347 1 2918
2 76348 1 2918
2 76349 1 2926
2 76350 1 2926
2 76351 1 2926
2 76352 1 2926
2 76353 1 2927
2 76354 1 2927
2 76355 1 2927
2 76356 1 2927
2 76357 1 2927
2 76358 1 2927
2 76359 1 2928
2 76360 1 2928
2 76361 1 2928
2 76362 1 2928
2 76363 1 2929
2 76364 1 2929
2 76365 1 2929
2 76366 1 2929
2 76367 1 2929
2 76368 1 2929
2 76369 1 2929
2 76370 1 2929
2 76371 1 2929
2 76372 1 2930
2 76373 1 2930
2 76374 1 2930
2 76375 1 2931
2 76376 1 2931
2 76377 1 2934
2 76378 1 2934
2 76379 1 2934
2 76380 1 2934
2 76381 1 2934
2 76382 1 2934
2 76383 1 2934
2 76384 1 2934
2 76385 1 2934
2 76386 1 2935
2 76387 1 2935
2 76388 1 2936
2 76389 1 2936
2 76390 1 2936
2 76391 1 2936
2 76392 1 2937
2 76393 1 2937
2 76394 1 2937
2 76395 1 2937
2 76396 1 2937
2 76397 1 2940
2 76398 1 2940
2 76399 1 2941
2 76400 1 2941
2 76401 1 2946
2 76402 1 2946
2 76403 1 2946
2 76404 1 2946
2 76405 1 2947
2 76406 1 2947
2 76407 1 2955
2 76408 1 2955
2 76409 1 2965
2 76410 1 2965
2 76411 1 2965
2 76412 1 2966
2 76413 1 2966
2 76414 1 2968
2 76415 1 2968
2 76416 1 2969
2 76417 1 2969
2 76418 1 2970
2 76419 1 2970
2 76420 1 2970
2 76421 1 2975
2 76422 1 2975
2 76423 1 2975
2 76424 1 2983
2 76425 1 2983
2 76426 1 2983
2 76427 1 2983
2 76428 1 2983
2 76429 1 2983
2 76430 1 2983
2 76431 1 2984
2 76432 1 2984
2 76433 1 2984
2 76434 1 2984
2 76435 1 2987
2 76436 1 2987
2 76437 1 2987
2 76438 1 2990
2 76439 1 2990
2 76440 1 2999
2 76441 1 2999
2 76442 1 2999
2 76443 1 2999
2 76444 1 3000
2 76445 1 3000
2 76446 1 3000
2 76447 1 3007
2 76448 1 3007
2 76449 1 3007
2 76450 1 3007
2 76451 1 3007
2 76452 1 3007
2 76453 1 3007
2 76454 1 3007
2 76455 1 3008
2 76456 1 3008
2 76457 1 3008
2 76458 1 3008
2 76459 1 3008
2 76460 1 3008
2 76461 1 3008
2 76462 1 3008
2 76463 1 3008
2 76464 1 3008
2 76465 1 3008
2 76466 1 3008
2 76467 1 3008
2 76468 1 3008
2 76469 1 3008
2 76470 1 3008
2 76471 1 3008
2 76472 1 3008
2 76473 1 3008
2 76474 1 3008
2 76475 1 3008
2 76476 1 3008
2 76477 1 3008
2 76478 1 3008
2 76479 1 3008
2 76480 1 3008
2 76481 1 3008
2 76482 1 3008
2 76483 1 3008
2 76484 1 3008
2 76485 1 3008
2 76486 1 3009
2 76487 1 3009
2 76488 1 3009
2 76489 1 3009
2 76490 1 3009
2 76491 1 3009
2 76492 1 3009
2 76493 1 3009
2 76494 1 3009
2 76495 1 3009
2 76496 1 3010
2 76497 1 3010
2 76498 1 3010
2 76499 1 3010
2 76500 1 3010
2 76501 1 3010
2 76502 1 3010
2 76503 1 3010
2 76504 1 3010
2 76505 1 3010
2 76506 1 3010
2 76507 1 3010
2 76508 1 3010
2 76509 1 3010
2 76510 1 3010
2 76511 1 3010
2 76512 1 3010
2 76513 1 3010
2 76514 1 3010
2 76515 1 3010
2 76516 1 3010
2 76517 1 3010
2 76518 1 3011
2 76519 1 3011
2 76520 1 3011
2 76521 1 3012
2 76522 1 3012
2 76523 1 3012
2 76524 1 3012
2 76525 1 3034
2 76526 1 3034
2 76527 1 3034
2 76528 1 3034
2 76529 1 3034
2 76530 1 3034
2 76531 1 3034
2 76532 1 3034
2 76533 1 3034
2 76534 1 3034
2 76535 1 3036
2 76536 1 3036
2 76537 1 3051
2 76538 1 3051
2 76539 1 3051
2 76540 1 3051
2 76541 1 3051
2 76542 1 3052
2 76543 1 3052
2 76544 1 3052
2 76545 1 3052
2 76546 1 3052
2 76547 1 3052
2 76548 1 3052
2 76549 1 3052
2 76550 1 3052
2 76551 1 3067
2 76552 1 3067
2 76553 1 3067
2 76554 1 3067
2 76555 1 3089
2 76556 1 3089
2 76557 1 3089
2 76558 1 3089
2 76559 1 3089
2 76560 1 3090
2 76561 1 3090
2 76562 1 3090
2 76563 1 3090
2 76564 1 3090
2 76565 1 3090
2 76566 1 3090
2 76567 1 3090
2 76568 1 3090
2 76569 1 3090
2 76570 1 3090
2 76571 1 3092
2 76572 1 3092
2 76573 1 3092
2 76574 1 3093
2 76575 1 3093
2 76576 1 3093
2 76577 1 3093
2 76578 1 3093
2 76579 1 3093
2 76580 1 3095
2 76581 1 3095
2 76582 1 3106
2 76583 1 3106
2 76584 1 3106
2 76585 1 3106
2 76586 1 3107
2 76587 1 3107
2 76588 1 3107
2 76589 1 3108
2 76590 1 3108
2 76591 1 3108
2 76592 1 3124
2 76593 1 3124
2 76594 1 3124
2 76595 1 3124
2 76596 1 3124
2 76597 1 3125
2 76598 1 3125
2 76599 1 3126
2 76600 1 3126
2 76601 1 3127
2 76602 1 3127
2 76603 1 3127
2 76604 1 3127
2 76605 1 3127
2 76606 1 3127
2 76607 1 3127
2 76608 1 3127
2 76609 1 3127
2 76610 1 3127
2 76611 1 3127
2 76612 1 3127
2 76613 1 3136
2 76614 1 3136
2 76615 1 3136
2 76616 1 3136
2 76617 1 3136
2 76618 1 3136
2 76619 1 3136
2 76620 1 3136
2 76621 1 3136
2 76622 1 3136
2 76623 1 3136
2 76624 1 3136
2 76625 1 3136
2 76626 1 3136
2 76627 1 3136
2 76628 1 3136
2 76629 1 3136
2 76630 1 3136
2 76631 1 3136
2 76632 1 3136
2 76633 1 3136
2 76634 1 3136
2 76635 1 3136
2 76636 1 3136
2 76637 1 3136
2 76638 1 3136
2 76639 1 3136
2 76640 1 3136
2 76641 1 3136
2 76642 1 3136
2 76643 1 3136
2 76644 1 3136
2 76645 1 3136
2 76646 1 3136
2 76647 1 3136
2 76648 1 3136
2 76649 1 3136
2 76650 1 3136
2 76651 1 3136
2 76652 1 3136
2 76653 1 3136
2 76654 1 3136
2 76655 1 3136
2 76656 1 3136
2 76657 1 3136
2 76658 1 3136
2 76659 1 3136
2 76660 1 3136
2 76661 1 3136
2 76662 1 3136
2 76663 1 3136
2 76664 1 3136
2 76665 1 3137
2 76666 1 3137
2 76667 1 3137
2 76668 1 3137
2 76669 1 3137
2 76670 1 3137
2 76671 1 3137
2 76672 1 3137
2 76673 1 3137
2 76674 1 3137
2 76675 1 3137
2 76676 1 3137
2 76677 1 3137
2 76678 1 3137
2 76679 1 3137
2 76680 1 3137
2 76681 1 3137
2 76682 1 3137
2 76683 1 3137
2 76684 1 3137
2 76685 1 3137
2 76686 1 3137
2 76687 1 3137
2 76688 1 3137
2 76689 1 3137
2 76690 1 3137
2 76691 1 3137
2 76692 1 3137
2 76693 1 3137
2 76694 1 3137
2 76695 1 3137
2 76696 1 3137
2 76697 1 3137
2 76698 1 3137
2 76699 1 3137
2 76700 1 3137
2 76701 1 3137
2 76702 1 3137
2 76703 1 3137
2 76704 1 3137
2 76705 1 3137
2 76706 1 3137
2 76707 1 3137
2 76708 1 3137
2 76709 1 3137
2 76710 1 3137
2 76711 1 3137
2 76712 1 3137
2 76713 1 3137
2 76714 1 3137
2 76715 1 3137
2 76716 1 3137
2 76717 1 3137
2 76718 1 3137
2 76719 1 3137
2 76720 1 3137
2 76721 1 3137
2 76722 1 3137
2 76723 1 3138
2 76724 1 3138
2 76725 1 3138
2 76726 1 3138
2 76727 1 3138
2 76728 1 3138
2 76729 1 3138
2 76730 1 3138
2 76731 1 3138
2 76732 1 3138
2 76733 1 3138
2 76734 1 3138
2 76735 1 3138
2 76736 1 3138
2 76737 1 3138
2 76738 1 3138
2 76739 1 3138
2 76740 1 3138
2 76741 1 3138
2 76742 1 3138
2 76743 1 3138
2 76744 1 3138
2 76745 1 3138
2 76746 1 3138
2 76747 1 3138
2 76748 1 3138
2 76749 1 3138
2 76750 1 3138
2 76751 1 3138
2 76752 1 3138
2 76753 1 3138
2 76754 1 3138
2 76755 1 3138
2 76756 1 3138
2 76757 1 3138
2 76758 1 3138
2 76759 1 3138
2 76760 1 3138
2 76761 1 3138
2 76762 1 3138
2 76763 1 3139
2 76764 1 3139
2 76765 1 3142
2 76766 1 3142
2 76767 1 3145
2 76768 1 3145
2 76769 1 3150
2 76770 1 3150
2 76771 1 3150
2 76772 1 3157
2 76773 1 3157
2 76774 1 3157
2 76775 1 3157
2 76776 1 3157
2 76777 1 3160
2 76778 1 3160
2 76779 1 3161
2 76780 1 3161
2 76781 1 3161
2 76782 1 3168
2 76783 1 3168
2 76784 1 3168
2 76785 1 3179
2 76786 1 3179
2 76787 1 3179
2 76788 1 3179
2 76789 1 3179
2 76790 1 3179
2 76791 1 3181
2 76792 1 3181
2 76793 1 3188
2 76794 1 3188
2 76795 1 3192
2 76796 1 3192
2 76797 1 3192
2 76798 1 3192
2 76799 1 3192
2 76800 1 3192
2 76801 1 3192
2 76802 1 3192
2 76803 1 3192
2 76804 1 3193
2 76805 1 3193
2 76806 1 3193
2 76807 1 3193
2 76808 1 3193
2 76809 1 3193
2 76810 1 3193
2 76811 1 3193
2 76812 1 3193
2 76813 1 3193
2 76814 1 3193
2 76815 1 3193
2 76816 1 3193
2 76817 1 3193
2 76818 1 3193
2 76819 1 3193
2 76820 1 3194
2 76821 1 3194
2 76822 1 3194
2 76823 1 3195
2 76824 1 3195
2 76825 1 3197
2 76826 1 3197
2 76827 1 3198
2 76828 1 3198
2 76829 1 3198
2 76830 1 3199
2 76831 1 3199
2 76832 1 3212
2 76833 1 3212
2 76834 1 3212
2 76835 1 3212
2 76836 1 3212
2 76837 1 3212
2 76838 1 3229
2 76839 1 3229
2 76840 1 3229
2 76841 1 3230
2 76842 1 3230
2 76843 1 3230
2 76844 1 3230
2 76845 1 3230
2 76846 1 3230
2 76847 1 3230
2 76848 1 3246
2 76849 1 3246
2 76850 1 3246
2 76851 1 3247
2 76852 1 3247
2 76853 1 3249
2 76854 1 3249
2 76855 1 3250
2 76856 1 3250
2 76857 1 3250
2 76858 1 3250
2 76859 1 3250
2 76860 1 3250
2 76861 1 3250
2 76862 1 3250
2 76863 1 3259
2 76864 1 3259
2 76865 1 3259
2 76866 1 3259
2 76867 1 3266
2 76868 1 3266
2 76869 1 3266
2 76870 1 3266
2 76871 1 3267
2 76872 1 3267
2 76873 1 3267
2 76874 1 3267
2 76875 1 3289
2 76876 1 3289
2 76877 1 3289
2 76878 1 3289
2 76879 1 3289
2 76880 1 3289
2 76881 1 3289
2 76882 1 3289
2 76883 1 3289
2 76884 1 3289
2 76885 1 3289
2 76886 1 3289
2 76887 1 3289
2 76888 1 3289
2 76889 1 3290
2 76890 1 3290
2 76891 1 3290
2 76892 1 3290
2 76893 1 3291
2 76894 1 3291
2 76895 1 3291
2 76896 1 3291
2 76897 1 3291
2 76898 1 3291
2 76899 1 3291
2 76900 1 3291
2 76901 1 3291
2 76902 1 3292
2 76903 1 3292
2 76904 1 3292
2 76905 1 3292
2 76906 1 3292
2 76907 1 3292
2 76908 1 3292
2 76909 1 3292
2 76910 1 3292
2 76911 1 3293
2 76912 1 3293
2 76913 1 3294
2 76914 1 3294
2 76915 1 3302
2 76916 1 3302
2 76917 1 3302
2 76918 1 3302
2 76919 1 3302
2 76920 1 3302
2 76921 1 3302
2 76922 1 3302
2 76923 1 3302
2 76924 1 3302
2 76925 1 3302
2 76926 1 3302
2 76927 1 3302
2 76928 1 3302
2 76929 1 3302
2 76930 1 3303
2 76931 1 3303
2 76932 1 3306
2 76933 1 3306
2 76934 1 3306
2 76935 1 3306
2 76936 1 3306
2 76937 1 3307
2 76938 1 3307
2 76939 1 3308
2 76940 1 3308
2 76941 1 3312
2 76942 1 3312
2 76943 1 3319
2 76944 1 3319
2 76945 1 3319
2 76946 1 3319
2 76947 1 3320
2 76948 1 3320
2 76949 1 3320
2 76950 1 3320
2 76951 1 3320
2 76952 1 3320
2 76953 1 3320
2 76954 1 3320
2 76955 1 3320
2 76956 1 3320
2 76957 1 3320
2 76958 1 3320
2 76959 1 3320
2 76960 1 3320
2 76961 1 3320
2 76962 1 3320
2 76963 1 3320
2 76964 1 3320
2 76965 1 3320
2 76966 1 3320
2 76967 1 3320
2 76968 1 3320
2 76969 1 3320
2 76970 1 3321
2 76971 1 3321
2 76972 1 3321
2 76973 1 3321
2 76974 1 3322
2 76975 1 3322
2 76976 1 3329
2 76977 1 3329
2 76978 1 3329
2 76979 1 3329
2 76980 1 3329
2 76981 1 3330
2 76982 1 3330
2 76983 1 3330
2 76984 1 3331
2 76985 1 3331
2 76986 1 3331
2 76987 1 3331
2 76988 1 3331
2 76989 1 3331
2 76990 1 3331
2 76991 1 3331
2 76992 1 3331
2 76993 1 3332
2 76994 1 3332
2 76995 1 3332
2 76996 1 3335
2 76997 1 3335
2 76998 1 3338
2 76999 1 3338
2 77000 1 3338
2 77001 1 3339
2 77002 1 3339
2 77003 1 3339
2 77004 1 3339
2 77005 1 3339
2 77006 1 3339
2 77007 1 3339
2 77008 1 3339
2 77009 1 3339
2 77010 1 3340
2 77011 1 3340
2 77012 1 3340
2 77013 1 3340
2 77014 1 3340
2 77015 1 3354
2 77016 1 3354
2 77017 1 3354
2 77018 1 3354
2 77019 1 3354
2 77020 1 3354
2 77021 1 3355
2 77022 1 3355
2 77023 1 3355
2 77024 1 3355
2 77025 1 3355
2 77026 1 3357
2 77027 1 3357
2 77028 1 3357
2 77029 1 3357
2 77030 1 3357
2 77031 1 3357
2 77032 1 3357
2 77033 1 3357
2 77034 1 3357
2 77035 1 3357
2 77036 1 3357
2 77037 1 3357
2 77038 1 3358
2 77039 1 3358
2 77040 1 3358
2 77041 1 3358
2 77042 1 3362
2 77043 1 3362
2 77044 1 3362
2 77045 1 3362
2 77046 1 3362
2 77047 1 3362
2 77048 1 3364
2 77049 1 3364
2 77050 1 3364
2 77051 1 3372
2 77052 1 3372
2 77053 1 3372
2 77054 1 3372
2 77055 1 3372
2 77056 1 3372
2 77057 1 3373
2 77058 1 3373
2 77059 1 3373
2 77060 1 3373
2 77061 1 3373
2 77062 1 3373
2 77063 1 3373
2 77064 1 3373
2 77065 1 3373
2 77066 1 3373
2 77067 1 3373
2 77068 1 3373
2 77069 1 3373
2 77070 1 3373
2 77071 1 3373
2 77072 1 3373
2 77073 1 3373
2 77074 1 3373
2 77075 1 3373
2 77076 1 3373
2 77077 1 3373
2 77078 1 3373
2 77079 1 3375
2 77080 1 3375
2 77081 1 3376
2 77082 1 3376
2 77083 1 3376
2 77084 1 3381
2 77085 1 3381
2 77086 1 3382
2 77087 1 3382
2 77088 1 3384
2 77089 1 3384
2 77090 1 3384
2 77091 1 3384
2 77092 1 3384
2 77093 1 3384
2 77094 1 3384
2 77095 1 3384
2 77096 1 3384
2 77097 1 3384
2 77098 1 3384
2 77099 1 3384
2 77100 1 3384
2 77101 1 3384
2 77102 1 3384
2 77103 1 3384
2 77104 1 3384
2 77105 1 3384
2 77106 1 3384
2 77107 1 3384
2 77108 1 3384
2 77109 1 3384
2 77110 1 3384
2 77111 1 3385
2 77112 1 3385
2 77113 1 3385
2 77114 1 3385
2 77115 1 3385
2 77116 1 3385
2 77117 1 3385
2 77118 1 3385
2 77119 1 3386
2 77120 1 3386
2 77121 1 3386
2 77122 1 3386
2 77123 1 3386
2 77124 1 3386
2 77125 1 3386
2 77126 1 3386
2 77127 1 3386
2 77128 1 3386
2 77129 1 3386
2 77130 1 3386
2 77131 1 3386
2 77132 1 3386
2 77133 1 3386
2 77134 1 3386
2 77135 1 3386
2 77136 1 3386
2 77137 1 3386
2 77138 1 3386
2 77139 1 3386
2 77140 1 3386
2 77141 1 3386
2 77142 1 3386
2 77143 1 3386
2 77144 1 3386
2 77145 1 3386
2 77146 1 3386
2 77147 1 3386
2 77148 1 3386
2 77149 1 3386
2 77150 1 3386
2 77151 1 3386
2 77152 1 3386
2 77153 1 3386
2 77154 1 3386
2 77155 1 3386
2 77156 1 3386
2 77157 1 3386
2 77158 1 3386
2 77159 1 3386
2 77160 1 3386
2 77161 1 3386
2 77162 1 3386
2 77163 1 3386
2 77164 1 3386
2 77165 1 3386
2 77166 1 3387
2 77167 1 3387
2 77168 1 3387
2 77169 1 3388
2 77170 1 3388
2 77171 1 3389
2 77172 1 3389
2 77173 1 3389
2 77174 1 3390
2 77175 1 3390
2 77176 1 3390
2 77177 1 3390
2 77178 1 3390
2 77179 1 3390
2 77180 1 3391
2 77181 1 3391
2 77182 1 3391
2 77183 1 3391
2 77184 1 3395
2 77185 1 3395
2 77186 1 3395
2 77187 1 3396
2 77188 1 3396
2 77189 1 3397
2 77190 1 3397
2 77191 1 3398
2 77192 1 3398
2 77193 1 3398
2 77194 1 3398
2 77195 1 3398
2 77196 1 3398
2 77197 1 3406
2 77198 1 3406
2 77199 1 3409
2 77200 1 3409
2 77201 1 3411
2 77202 1 3411
2 77203 1 3411
2 77204 1 3411
2 77205 1 3411
2 77206 1 3411
2 77207 1 3411
2 77208 1 3411
2 77209 1 3411
2 77210 1 3411
2 77211 1 3412
2 77212 1 3412
2 77213 1 3412
2 77214 1 3413
2 77215 1 3413
2 77216 1 3413
2 77217 1 3413
2 77218 1 3413
2 77219 1 3413
2 77220 1 3413
2 77221 1 3413
2 77222 1 3413
2 77223 1 3421
2 77224 1 3421
2 77225 1 3427
2 77226 1 3427
2 77227 1 3427
2 77228 1 3427
2 77229 1 3427
2 77230 1 3427
2 77231 1 3427
2 77232 1 3427
2 77233 1 3427
2 77234 1 3427
2 77235 1 3427
2 77236 1 3427
2 77237 1 3427
2 77238 1 3427
2 77239 1 3427
2 77240 1 3436
2 77241 1 3436
2 77242 1 3436
2 77243 1 3436
2 77244 1 3437
2 77245 1 3437
2 77246 1 3441
2 77247 1 3441
2 77248 1 3441
2 77249 1 3441
2 77250 1 3441
2 77251 1 3441
2 77252 1 3441
2 77253 1 3441
2 77254 1 3441
2 77255 1 3441
2 77256 1 3441
2 77257 1 3441
2 77258 1 3441
2 77259 1 3441
2 77260 1 3441
2 77261 1 3441
2 77262 1 3441
2 77263 1 3441
2 77264 1 3441
2 77265 1 3441
2 77266 1 3441
2 77267 1 3441
2 77268 1 3441
2 77269 1 3441
2 77270 1 3441
2 77271 1 3441
2 77272 1 3441
2 77273 1 3441
2 77274 1 3441
2 77275 1 3441
2 77276 1 3441
2 77277 1 3441
2 77278 1 3442
2 77279 1 3442
2 77280 1 3448
2 77281 1 3448
2 77282 1 3448
2 77283 1 3448
2 77284 1 3449
2 77285 1 3449
2 77286 1 3450
2 77287 1 3450
2 77288 1 3453
2 77289 1 3453
2 77290 1 3453
2 77291 1 3453
2 77292 1 3454
2 77293 1 3454
2 77294 1 3454
2 77295 1 3454
2 77296 1 3458
2 77297 1 3458
2 77298 1 3458
2 77299 1 3459
2 77300 1 3459
2 77301 1 3459
2 77302 1 3459
2 77303 1 3459
2 77304 1 3472
2 77305 1 3472
2 77306 1 3473
2 77307 1 3473
2 77308 1 3473
2 77309 1 3473
2 77310 1 3473
2 77311 1 3473
2 77312 1 3473
2 77313 1 3473
2 77314 1 3473
2 77315 1 3474
2 77316 1 3474
2 77317 1 3474
2 77318 1 3474
2 77319 1 3475
2 77320 1 3475
2 77321 1 3475
2 77322 1 3475
2 77323 1 3479
2 77324 1 3479
2 77325 1 3479
2 77326 1 3479
2 77327 1 3481
2 77328 1 3481
2 77329 1 3493
2 77330 1 3493
2 77331 1 3494
2 77332 1 3494
2 77333 1 3505
2 77334 1 3505
2 77335 1 3512
2 77336 1 3512
2 77337 1 3512
2 77338 1 3512
2 77339 1 3512
2 77340 1 3512
2 77341 1 3512
2 77342 1 3512
2 77343 1 3512
2 77344 1 3512
2 77345 1 3512
2 77346 1 3512
2 77347 1 3512
2 77348 1 3512
2 77349 1 3512
2 77350 1 3512
2 77351 1 3513
2 77352 1 3513
2 77353 1 3522
2 77354 1 3522
2 77355 1 3522
2 77356 1 3522
2 77357 1 3522
2 77358 1 3522
2 77359 1 3522
2 77360 1 3522
2 77361 1 3522
2 77362 1 3522
2 77363 1 3523
2 77364 1 3523
2 77365 1 3523
2 77366 1 3526
2 77367 1 3526
2 77368 1 3527
2 77369 1 3527
2 77370 1 3527
2 77371 1 3527
2 77372 1 3527
2 77373 1 3527
2 77374 1 3527
2 77375 1 3527
2 77376 1 3528
2 77377 1 3528
2 77378 1 3528
2 77379 1 3528
2 77380 1 3530
2 77381 1 3530
2 77382 1 3531
2 77383 1 3531
2 77384 1 3531
2 77385 1 3531
2 77386 1 3531
2 77387 1 3532
2 77388 1 3532
2 77389 1 3532
2 77390 1 3533
2 77391 1 3533
2 77392 1 3533
2 77393 1 3533
2 77394 1 3533
2 77395 1 3533
2 77396 1 3533
2 77397 1 3533
2 77398 1 3533
2 77399 1 3533
2 77400 1 3533
2 77401 1 3534
2 77402 1 3534
2 77403 1 3535
2 77404 1 3535
2 77405 1 3535
2 77406 1 3535
2 77407 1 3535
2 77408 1 3544
2 77409 1 3544
2 77410 1 3544
2 77411 1 3544
2 77412 1 3544
2 77413 1 3544
2 77414 1 3544
2 77415 1 3544
2 77416 1 3544
2 77417 1 3544
2 77418 1 3544
2 77419 1 3544
2 77420 1 3544
2 77421 1 3544
2 77422 1 3544
2 77423 1 3544
2 77424 1 3544
2 77425 1 3544
2 77426 1 3544
2 77427 1 3544
2 77428 1 3544
2 77429 1 3544
2 77430 1 3544
2 77431 1 3544
2 77432 1 3545
2 77433 1 3545
2 77434 1 3545
2 77435 1 3563
2 77436 1 3563
2 77437 1 3563
2 77438 1 3563
2 77439 1 3565
2 77440 1 3565
2 77441 1 3565
2 77442 1 3565
2 77443 1 3565
2 77444 1 3566
2 77445 1 3566
2 77446 1 3579
2 77447 1 3579
2 77448 1 3579
2 77449 1 3579
2 77450 1 3579
2 77451 1 3579
2 77452 1 3579
2 77453 1 3579
2 77454 1 3587
2 77455 1 3587
2 77456 1 3587
2 77457 1 3587
2 77458 1 3587
2 77459 1 3587
2 77460 1 3587
2 77461 1 3587
2 77462 1 3587
2 77463 1 3587
2 77464 1 3587
2 77465 1 3587
2 77466 1 3587
2 77467 1 3587
2 77468 1 3587
2 77469 1 3587
2 77470 1 3587
2 77471 1 3587
2 77472 1 3587
2 77473 1 3587
2 77474 1 3587
2 77475 1 3587
2 77476 1 3587
2 77477 1 3589
2 77478 1 3589
2 77479 1 3589
2 77480 1 3589
2 77481 1 3589
2 77482 1 3589
2 77483 1 3589
2 77484 1 3589
2 77485 1 3591
2 77486 1 3591
2 77487 1 3592
2 77488 1 3592
2 77489 1 3592
2 77490 1 3592
2 77491 1 3592
2 77492 1 3592
2 77493 1 3592
2 77494 1 3592
2 77495 1 3592
2 77496 1 3592
2 77497 1 3593
2 77498 1 3593
2 77499 1 3594
2 77500 1 3594
2 77501 1 3595
2 77502 1 3595
2 77503 1 3595
2 77504 1 3595
2 77505 1 3595
2 77506 1 3595
2 77507 1 3595
2 77508 1 3595
2 77509 1 3597
2 77510 1 3597
2 77511 1 3597
2 77512 1 3597
2 77513 1 3597
2 77514 1 3605
2 77515 1 3605
2 77516 1 3605
2 77517 1 3605
2 77518 1 3605
2 77519 1 3605
2 77520 1 3605
2 77521 1 3605
2 77522 1 3607
2 77523 1 3607
2 77524 1 3608
2 77525 1 3608
2 77526 1 3609
2 77527 1 3609
2 77528 1 3609
2 77529 1 3609
2 77530 1 3609
2 77531 1 3609
2 77532 1 3610
2 77533 1 3610
2 77534 1 3610
2 77535 1 3619
2 77536 1 3619
2 77537 1 3619
2 77538 1 3620
2 77539 1 3620
2 77540 1 3620
2 77541 1 3620
2 77542 1 3620
2 77543 1 3620
2 77544 1 3621
2 77545 1 3621
2 77546 1 3621
2 77547 1 3621
2 77548 1 3622
2 77549 1 3622
2 77550 1 3629
2 77551 1 3629
2 77552 1 3629
2 77553 1 3629
2 77554 1 3629
2 77555 1 3629
2 77556 1 3629
2 77557 1 3630
2 77558 1 3630
2 77559 1 3631
2 77560 1 3631
2 77561 1 3637
2 77562 1 3637
2 77563 1 3637
2 77564 1 3645
2 77565 1 3645
2 77566 1 3645
2 77567 1 3646
2 77568 1 3646
2 77569 1 3646
2 77570 1 3647
2 77571 1 3647
2 77572 1 3647
2 77573 1 3649
2 77574 1 3649
2 77575 1 3649
2 77576 1 3649
2 77577 1 3650
2 77578 1 3650
2 77579 1 3665
2 77580 1 3665
2 77581 1 3665
2 77582 1 3665
2 77583 1 3665
2 77584 1 3665
2 77585 1 3665
2 77586 1 3665
2 77587 1 3665
2 77588 1 3665
2 77589 1 3665
2 77590 1 3665
2 77591 1 3665
2 77592 1 3665
2 77593 1 3665
2 77594 1 3665
2 77595 1 3665
2 77596 1 3675
2 77597 1 3675
2 77598 1 3675
2 77599 1 3675
2 77600 1 3677
2 77601 1 3677
2 77602 1 3686
2 77603 1 3686
2 77604 1 3686
2 77605 1 3686
2 77606 1 3686
2 77607 1 3686
2 77608 1 3686
2 77609 1 3686
2 77610 1 3686
2 77611 1 3687
2 77612 1 3687
2 77613 1 3687
2 77614 1 3688
2 77615 1 3688
2 77616 1 3688
2 77617 1 3688
2 77618 1 3688
2 77619 1 3688
2 77620 1 3688
2 77621 1 3689
2 77622 1 3689
2 77623 1 3691
2 77624 1 3691
2 77625 1 3701
2 77626 1 3701
2 77627 1 3703
2 77628 1 3703
2 77629 1 3703
2 77630 1 3711
2 77631 1 3711
2 77632 1 3711
2 77633 1 3711
2 77634 1 3711
2 77635 1 3711
2 77636 1 3712
2 77637 1 3712
2 77638 1 3712
2 77639 1 3712
2 77640 1 3712
2 77641 1 3712
2 77642 1 3713
2 77643 1 3713
2 77644 1 3726
2 77645 1 3726
2 77646 1 3727
2 77647 1 3727
2 77648 1 3727
2 77649 1 3727
2 77650 1 3727
2 77651 1 3727
2 77652 1 3727
2 77653 1 3727
2 77654 1 3728
2 77655 1 3728
2 77656 1 3728
2 77657 1 3728
2 77658 1 3728
2 77659 1 3728
2 77660 1 3728
2 77661 1 3728
2 77662 1 3728
2 77663 1 3728
2 77664 1 3728
2 77665 1 3728
2 77666 1 3728
2 77667 1 3728
2 77668 1 3728
2 77669 1 3728
2 77670 1 3728
2 77671 1 3728
2 77672 1 3728
2 77673 1 3728
2 77674 1 3728
2 77675 1 3728
2 77676 1 3728
2 77677 1 3728
2 77678 1 3728
2 77679 1 3728
2 77680 1 3728
2 77681 1 3728
2 77682 1 3728
2 77683 1 3730
2 77684 1 3730
2 77685 1 3730
2 77686 1 3730
2 77687 1 3731
2 77688 1 3731
2 77689 1 3732
2 77690 1 3732
2 77691 1 3733
2 77692 1 3733
2 77693 1 3734
2 77694 1 3734
2 77695 1 3735
2 77696 1 3735
2 77697 1 3735
2 77698 1 3735
2 77699 1 3736
2 77700 1 3736
2 77701 1 3736
2 77702 1 3736
2 77703 1 3747
2 77704 1 3747
2 77705 1 3747
2 77706 1 3747
2 77707 1 3747
2 77708 1 3747
2 77709 1 3747
2 77710 1 3747
2 77711 1 3748
2 77712 1 3748
2 77713 1 3748
2 77714 1 3748
2 77715 1 3748
2 77716 1 3748
2 77717 1 3748
2 77718 1 3748
2 77719 1 3748
2 77720 1 3749
2 77721 1 3749
2 77722 1 3753
2 77723 1 3753
2 77724 1 3753
2 77725 1 3753
2 77726 1 3754
2 77727 1 3754
2 77728 1 3754
2 77729 1 3754
2 77730 1 3754
2 77731 1 3754
2 77732 1 3754
2 77733 1 3754
2 77734 1 3754
2 77735 1 3754
2 77736 1 3754
2 77737 1 3754
2 77738 1 3754
2 77739 1 3754
2 77740 1 3764
2 77741 1 3764
2 77742 1 3765
2 77743 1 3765
2 77744 1 3768
2 77745 1 3768
2 77746 1 3768
2 77747 1 3775
2 77748 1 3775
2 77749 1 3775
2 77750 1 3776
2 77751 1 3776
2 77752 1 3783
2 77753 1 3783
2 77754 1 3786
2 77755 1 3786
2 77756 1 3791
2 77757 1 3791
2 77758 1 3791
2 77759 1 3792
2 77760 1 3792
2 77761 1 3793
2 77762 1 3793
2 77763 1 3793
2 77764 1 3793
2 77765 1 3793
2 77766 1 3793
2 77767 1 3793
2 77768 1 3793
2 77769 1 3793
2 77770 1 3793
2 77771 1 3793
2 77772 1 3805
2 77773 1 3805
2 77774 1 3814
2 77775 1 3814
2 77776 1 3814
2 77777 1 3814
2 77778 1 3814
2 77779 1 3814
2 77780 1 3814
2 77781 1 3814
2 77782 1 3814
2 77783 1 3814
2 77784 1 3814
2 77785 1 3814
2 77786 1 3815
2 77787 1 3815
2 77788 1 3816
2 77789 1 3816
2 77790 1 3816
2 77791 1 3816
2 77792 1 3817
2 77793 1 3817
2 77794 1 3818
2 77795 1 3818
2 77796 1 3818
2 77797 1 3818
2 77798 1 3818
2 77799 1 3818
2 77800 1 3818
2 77801 1 3818
2 77802 1 3818
2 77803 1 3818
2 77804 1 3818
2 77805 1 3818
2 77806 1 3818
2 77807 1 3818
2 77808 1 3819
2 77809 1 3819
2 77810 1 3819
2 77811 1 3819
2 77812 1 3819
2 77813 1 3819
2 77814 1 3819
2 77815 1 3820
2 77816 1 3820
2 77817 1 3820
2 77818 1 3820
2 77819 1 3820
2 77820 1 3820
2 77821 1 3820
2 77822 1 3820
2 77823 1 3820
2 77824 1 3820
2 77825 1 3820
2 77826 1 3820
2 77827 1 3820
2 77828 1 3820
2 77829 1 3821
2 77830 1 3821
2 77831 1 3821
2 77832 1 3821
2 77833 1 3821
2 77834 1 3821
2 77835 1 3821
2 77836 1 3821
2 77837 1 3822
2 77838 1 3822
2 77839 1 3822
2 77840 1 3822
2 77841 1 3822
2 77842 1 3822
2 77843 1 3822
2 77844 1 3823
2 77845 1 3823
2 77846 1 3823
2 77847 1 3823
2 77848 1 3823
2 77849 1 3823
2 77850 1 3823
2 77851 1 3823
2 77852 1 3823
2 77853 1 3823
2 77854 1 3823
2 77855 1 3823
2 77856 1 3823
2 77857 1 3823
2 77858 1 3823
2 77859 1 3823
2 77860 1 3823
2 77861 1 3823
2 77862 1 3823
2 77863 1 3823
2 77864 1 3823
2 77865 1 3823
2 77866 1 3823
2 77867 1 3823
2 77868 1 3823
2 77869 1 3823
2 77870 1 3823
2 77871 1 3823
2 77872 1 3823
2 77873 1 3823
2 77874 1 3823
2 77875 1 3823
2 77876 1 3823
2 77877 1 3823
2 77878 1 3823
2 77879 1 3823
2 77880 1 3823
2 77881 1 3823
2 77882 1 3823
2 77883 1 3823
2 77884 1 3823
2 77885 1 3823
2 77886 1 3824
2 77887 1 3824
2 77888 1 3824
2 77889 1 3824
2 77890 1 3824
2 77891 1 3824
2 77892 1 3824
2 77893 1 3824
2 77894 1 3824
2 77895 1 3824
2 77896 1 3824
2 77897 1 3824
2 77898 1 3824
2 77899 1 3826
2 77900 1 3826
2 77901 1 3826
2 77902 1 3826
2 77903 1 3827
2 77904 1 3827
2 77905 1 3828
2 77906 1 3828
2 77907 1 3841
2 77908 1 3841
2 77909 1 3841
2 77910 1 3841
2 77911 1 3841
2 77912 1 3842
2 77913 1 3842
2 77914 1 3842
2 77915 1 3842
2 77916 1 3845
2 77917 1 3845
2 77918 1 3845
2 77919 1 3845
2 77920 1 3845
2 77921 1 3856
2 77922 1 3856
2 77923 1 3856
2 77924 1 3858
2 77925 1 3858
2 77926 1 3859
2 77927 1 3859
2 77928 1 3860
2 77929 1 3860
2 77930 1 3860
2 77931 1 3860
2 77932 1 3861
2 77933 1 3861
2 77934 1 3864
2 77935 1 3864
2 77936 1 3865
2 77937 1 3865
2 77938 1 3875
2 77939 1 3875
2 77940 1 3875
2 77941 1 3880
2 77942 1 3880
2 77943 1 3880
2 77944 1 3880
2 77945 1 3880
2 77946 1 3880
2 77947 1 3880
2 77948 1 3880
2 77949 1 3880
2 77950 1 3880
2 77951 1 3880
2 77952 1 3881
2 77953 1 3881
2 77954 1 3881
2 77955 1 3881
2 77956 1 3881
2 77957 1 3881
2 77958 1 3881
2 77959 1 3881
2 77960 1 3881
2 77961 1 3881
2 77962 1 3881
2 77963 1 3883
2 77964 1 3883
2 77965 1 3883
2 77966 1 3883
2 77967 1 3883
2 77968 1 3883
2 77969 1 3883
2 77970 1 3883
2 77971 1 3886
2 77972 1 3886
2 77973 1 3886
2 77974 1 3886
2 77975 1 3886
2 77976 1 3886
2 77977 1 3886
2 77978 1 3886
2 77979 1 3886
2 77980 1 3886
2 77981 1 3886
2 77982 1 3886
2 77983 1 3886
2 77984 1 3886
2 77985 1 3886
2 77986 1 3886
2 77987 1 3886
2 77988 1 3886
2 77989 1 3886
2 77990 1 3886
2 77991 1 3886
2 77992 1 3886
2 77993 1 3886
2 77994 1 3886
2 77995 1 3886
2 77996 1 3886
2 77997 1 3886
2 77998 1 3886
2 77999 1 3886
2 78000 1 3886
2 78001 1 3886
2 78002 1 3886
2 78003 1 3886
2 78004 1 3887
2 78005 1 3887
2 78006 1 3887
2 78007 1 3887
2 78008 1 3887
2 78009 1 3887
2 78010 1 3887
2 78011 1 3887
2 78012 1 3887
2 78013 1 3887
2 78014 1 3887
2 78015 1 3887
2 78016 1 3888
2 78017 1 3888
2 78018 1 3888
2 78019 1 3888
2 78020 1 3888
2 78021 1 3888
2 78022 1 3888
2 78023 1 3889
2 78024 1 3889
2 78025 1 3889
2 78026 1 3889
2 78027 1 3890
2 78028 1 3890
2 78029 1 3891
2 78030 1 3891
2 78031 1 3891
2 78032 1 3891
2 78033 1 3891
2 78034 1 3893
2 78035 1 3893
2 78036 1 3897
2 78037 1 3897
2 78038 1 3897
2 78039 1 3900
2 78040 1 3900
2 78041 1 3900
2 78042 1 3900
2 78043 1 3900
2 78044 1 3900
2 78045 1 3900
2 78046 1 3900
2 78047 1 3900
2 78048 1 3900
2 78049 1 3900
2 78050 1 3900
2 78051 1 3901
2 78052 1 3901
2 78053 1 3902
2 78054 1 3902
2 78055 1 3902
2 78056 1 3902
2 78057 1 3902
2 78058 1 3903
2 78059 1 3903
2 78060 1 3903
2 78061 1 3903
2 78062 1 3903
2 78063 1 3905
2 78064 1 3905
2 78065 1 3905
2 78066 1 3905
2 78067 1 3914
2 78068 1 3914
2 78069 1 3914
2 78070 1 3914
2 78071 1 3914
2 78072 1 3914
2 78073 1 3914
2 78074 1 3914
2 78075 1 3914
2 78076 1 3914
2 78077 1 3914
2 78078 1 3914
2 78079 1 3914
2 78080 1 3914
2 78081 1 3914
2 78082 1 3914
2 78083 1 3914
2 78084 1 3914
2 78085 1 3914
2 78086 1 3914
2 78087 1 3914
2 78088 1 3914
2 78089 1 3914
2 78090 1 3914
2 78091 1 3915
2 78092 1 3915
2 78093 1 3917
2 78094 1 3917
2 78095 1 3918
2 78096 1 3918
2 78097 1 3918
2 78098 1 3918
2 78099 1 3918
2 78100 1 3918
2 78101 1 3918
2 78102 1 3918
2 78103 1 3926
2 78104 1 3926
2 78105 1 3927
2 78106 1 3927
2 78107 1 3940
2 78108 1 3940
2 78109 1 3943
2 78110 1 3943
2 78111 1 3945
2 78112 1 3945
2 78113 1 3945
2 78114 1 3952
2 78115 1 3952
2 78116 1 3952
2 78117 1 3952
2 78118 1 3952
2 78119 1 3952
2 78120 1 3952
2 78121 1 3953
2 78122 1 3953
2 78123 1 3953
2 78124 1 3966
2 78125 1 3966
2 78126 1 3966
2 78127 1 3966
2 78128 1 3970
2 78129 1 3970
2 78130 1 3973
2 78131 1 3973
2 78132 1 3973
2 78133 1 3973
2 78134 1 3973
2 78135 1 3973
2 78136 1 3973
2 78137 1 3973
2 78138 1 3974
2 78139 1 3974
2 78140 1 3974
2 78141 1 3974
2 78142 1 3974
2 78143 1 3974
2 78144 1 3974
2 78145 1 3974
2 78146 1 3974
2 78147 1 3974
2 78148 1 3974
2 78149 1 3974
2 78150 1 3981
2 78151 1 3981
2 78152 1 3981
2 78153 1 3981
2 78154 1 3981
2 78155 1 3981
2 78156 1 3981
2 78157 1 3981
2 78158 1 3981
2 78159 1 3981
2 78160 1 3981
2 78161 1 3981
2 78162 1 3981
2 78163 1 3981
2 78164 1 3981
2 78165 1 3981
2 78166 1 3981
2 78167 1 3981
2 78168 1 3982
2 78169 1 3982
2 78170 1 3982
2 78171 1 3982
2 78172 1 3982
2 78173 1 3982
2 78174 1 3982
2 78175 1 3982
2 78176 1 3982
2 78177 1 3982
2 78178 1 3982
2 78179 1 3989
2 78180 1 3989
2 78181 1 3989
2 78182 1 3990
2 78183 1 3990
2 78184 1 3999
2 78185 1 3999
2 78186 1 3999
2 78187 1 4000
2 78188 1 4000
2 78189 1 4000
2 78190 1 4001
2 78191 1 4001
2 78192 1 4001
2 78193 1 4001
2 78194 1 4001
2 78195 1 4002
2 78196 1 4002
2 78197 1 4003
2 78198 1 4003
2 78199 1 4003
2 78200 1 4003
2 78201 1 4003
2 78202 1 4003
2 78203 1 4004
2 78204 1 4004
2 78205 1 4004
2 78206 1 4004
2 78207 1 4004
2 78208 1 4004
2 78209 1 4004
2 78210 1 4005
2 78211 1 4005
2 78212 1 4005
2 78213 1 4005
2 78214 1 4005
2 78215 1 4005
2 78216 1 4005
2 78217 1 4005
2 78218 1 4007
2 78219 1 4007
2 78220 1 4007
2 78221 1 4007
2 78222 1 4007
2 78223 1 4009
2 78224 1 4009
2 78225 1 4009
2 78226 1 4010
2 78227 1 4010
2 78228 1 4010
2 78229 1 4010
2 78230 1 4011
2 78231 1 4011
2 78232 1 4011
2 78233 1 4011
2 78234 1 4011
2 78235 1 4016
2 78236 1 4016
2 78237 1 4016
2 78238 1 4016
2 78239 1 4016
2 78240 1 4016
2 78241 1 4016
2 78242 1 4016
2 78243 1 4016
2 78244 1 4016
2 78245 1 4016
2 78246 1 4016
2 78247 1 4016
2 78248 1 4016
2 78249 1 4016
2 78250 1 4017
2 78251 1 4017
2 78252 1 4017
2 78253 1 4017
2 78254 1 4017
2 78255 1 4017
2 78256 1 4017
2 78257 1 4020
2 78258 1 4020
2 78259 1 4029
2 78260 1 4029
2 78261 1 4030
2 78262 1 4030
2 78263 1 4030
2 78264 1 4030
2 78265 1 4030
2 78266 1 4030
2 78267 1 4030
2 78268 1 4030
2 78269 1 4030
2 78270 1 4030
2 78271 1 4030
2 78272 1 4030
2 78273 1 4030
2 78274 1 4030
2 78275 1 4030
2 78276 1 4030
2 78277 1 4030
2 78278 1 4031
2 78279 1 4031
2 78280 1 4031
2 78281 1 4032
2 78282 1 4032
2 78283 1 4032
2 78284 1 4032
2 78285 1 4032
2 78286 1 4032
2 78287 1 4032
2 78288 1 4032
2 78289 1 4032
2 78290 1 4032
2 78291 1 4032
2 78292 1 4032
2 78293 1 4032
2 78294 1 4032
2 78295 1 4032
2 78296 1 4032
2 78297 1 4032
2 78298 1 4032
2 78299 1 4032
2 78300 1 4032
2 78301 1 4033
2 78302 1 4033
2 78303 1 4033
2 78304 1 4033
2 78305 1 4033
2 78306 1 4034
2 78307 1 4034
2 78308 1 4034
2 78309 1 4034
2 78310 1 4034
2 78311 1 4034
2 78312 1 4034
2 78313 1 4034
2 78314 1 4034
2 78315 1 4034
2 78316 1 4034
2 78317 1 4034
2 78318 1 4034
2 78319 1 4034
2 78320 1 4034
2 78321 1 4034
2 78322 1 4034
2 78323 1 4034
2 78324 1 4034
2 78325 1 4034
2 78326 1 4034
2 78327 1 4034
2 78328 1 4034
2 78329 1 4034
2 78330 1 4034
2 78331 1 4034
2 78332 1 4034
2 78333 1 4035
2 78334 1 4035
2 78335 1 4035
2 78336 1 4035
2 78337 1 4035
2 78338 1 4035
2 78339 1 4036
2 78340 1 4036
2 78341 1 4036
2 78342 1 4036
2 78343 1 4037
2 78344 1 4037
2 78345 1 4037
2 78346 1 4037
2 78347 1 4037
2 78348 1 4037
2 78349 1 4037
2 78350 1 4037
2 78351 1 4037
2 78352 1 4037
2 78353 1 4037
2 78354 1 4037
2 78355 1 4038
2 78356 1 4038
2 78357 1 4038
2 78358 1 4038
2 78359 1 4038
2 78360 1 4038
2 78361 1 4038
2 78362 1 4038
2 78363 1 4038
2 78364 1 4038
2 78365 1 4038
2 78366 1 4038
2 78367 1 4038
2 78368 1 4039
2 78369 1 4039
2 78370 1 4040
2 78371 1 4040
2 78372 1 4043
2 78373 1 4043
2 78374 1 4043
2 78375 1 4043
2 78376 1 4043
2 78377 1 4050
2 78378 1 4050
2 78379 1 4051
2 78380 1 4051
2 78381 1 4051
2 78382 1 4051
2 78383 1 4052
2 78384 1 4052
2 78385 1 4052
2 78386 1 4060
2 78387 1 4060
2 78388 1 4060
2 78389 1 4061
2 78390 1 4061
2 78391 1 4061
2 78392 1 4061
2 78393 1 4061
2 78394 1 4064
2 78395 1 4064
2 78396 1 4064
2 78397 1 4064
2 78398 1 4065
2 78399 1 4065
2 78400 1 4066
2 78401 1 4066
2 78402 1 4069
2 78403 1 4069
2 78404 1 4074
2 78405 1 4074
2 78406 1 4074
2 78407 1 4075
2 78408 1 4075
2 78409 1 4075
2 78410 1 4075
2 78411 1 4075
2 78412 1 4075
2 78413 1 4075
2 78414 1 4076
2 78415 1 4076
2 78416 1 4076
2 78417 1 4077
2 78418 1 4077
2 78419 1 4077
2 78420 1 4077
2 78421 1 4078
2 78422 1 4078
2 78423 1 4079
2 78424 1 4079
2 78425 1 4079
2 78426 1 4079
2 78427 1 4081
2 78428 1 4081
2 78429 1 4083
2 78430 1 4083
2 78431 1 4083
2 78432 1 4086
2 78433 1 4086
2 78434 1 4086
2 78435 1 4086
2 78436 1 4087
2 78437 1 4087
2 78438 1 4087
2 78439 1 4087
2 78440 1 4087
2 78441 1 4113
2 78442 1 4113
2 78443 1 4113
2 78444 1 4113
2 78445 1 4113
2 78446 1 4113
2 78447 1 4113
2 78448 1 4113
2 78449 1 4113
2 78450 1 4113
2 78451 1 4113
2 78452 1 4113
2 78453 1 4114
2 78454 1 4114
2 78455 1 4114
2 78456 1 4115
2 78457 1 4115
2 78458 1 4115
2 78459 1 4115
2 78460 1 4115
2 78461 1 4115
2 78462 1 4115
2 78463 1 4116
2 78464 1 4116
2 78465 1 4116
2 78466 1 4119
2 78467 1 4119
2 78468 1 4119
2 78469 1 4120
2 78470 1 4120
2 78471 1 4127
2 78472 1 4127
2 78473 1 4135
2 78474 1 4135
2 78475 1 4135
2 78476 1 4135
2 78477 1 4135
2 78478 1 4135
2 78479 1 4135
2 78480 1 4135
2 78481 1 4135
2 78482 1 4135
2 78483 1 4135
2 78484 1 4135
2 78485 1 4135
2 78486 1 4135
2 78487 1 4135
2 78488 1 4135
2 78489 1 4135
2 78490 1 4135
2 78491 1 4135
2 78492 1 4135
2 78493 1 4135
2 78494 1 4135
2 78495 1 4137
2 78496 1 4137
2 78497 1 4137
2 78498 1 4137
2 78499 1 4137
2 78500 1 4137
2 78501 1 4137
2 78502 1 4137
2 78503 1 4137
2 78504 1 4137
2 78505 1 4137
2 78506 1 4138
2 78507 1 4138
2 78508 1 4138
2 78509 1 4138
2 78510 1 4139
2 78511 1 4139
2 78512 1 4141
2 78513 1 4141
2 78514 1 4141
2 78515 1 4142
2 78516 1 4142
2 78517 1 4145
2 78518 1 4145
2 78519 1 4145
2 78520 1 4145
2 78521 1 4145
2 78522 1 4145
2 78523 1 4145
2 78524 1 4145
2 78525 1 4145
2 78526 1 4145
2 78527 1 4145
2 78528 1 4145
2 78529 1 4145
2 78530 1 4145
2 78531 1 4145
2 78532 1 4145
2 78533 1 4146
2 78534 1 4146
2 78535 1 4146
2 78536 1 4146
2 78537 1 4146
2 78538 1 4147
2 78539 1 4147
2 78540 1 4148
2 78541 1 4148
2 78542 1 4149
2 78543 1 4149
2 78544 1 4155
2 78545 1 4155
2 78546 1 4155
2 78547 1 4155
2 78548 1 4155
2 78549 1 4155
2 78550 1 4155
2 78551 1 4157
2 78552 1 4157
2 78553 1 4157
2 78554 1 4157
2 78555 1 4177
2 78556 1 4177
2 78557 1 4178
2 78558 1 4178
2 78559 1 4179
2 78560 1 4179
2 78561 1 4179
2 78562 1 4179
2 78563 1 4179
2 78564 1 4179
2 78565 1 4180
2 78566 1 4180
2 78567 1 4180
2 78568 1 4181
2 78569 1 4181
2 78570 1 4193
2 78571 1 4193
2 78572 1 4193
2 78573 1 4193
2 78574 1 4193
2 78575 1 4194
2 78576 1 4194
2 78577 1 4195
2 78578 1 4195
2 78579 1 4195
2 78580 1 4195
2 78581 1 4195
2 78582 1 4218
2 78583 1 4218
2 78584 1 4227
2 78585 1 4227
2 78586 1 4228
2 78587 1 4228
2 78588 1 4228
2 78589 1 4229
2 78590 1 4229
2 78591 1 4229
2 78592 1 4230
2 78593 1 4230
2 78594 1 4230
2 78595 1 4230
2 78596 1 4230
2 78597 1 4230
2 78598 1 4230
2 78599 1 4230
2 78600 1 4231
2 78601 1 4231
2 78602 1 4237
2 78603 1 4237
2 78604 1 4237
2 78605 1 4237
2 78606 1 4238
2 78607 1 4238
2 78608 1 4238
2 78609 1 4238
2 78610 1 4238
2 78611 1 4238
2 78612 1 4238
2 78613 1 4238
2 78614 1 4238
2 78615 1 4238
2 78616 1 4238
2 78617 1 4238
2 78618 1 4238
2 78619 1 4238
2 78620 1 4238
2 78621 1 4239
2 78622 1 4239
2 78623 1 4239
2 78624 1 4240
2 78625 1 4240
2 78626 1 4241
2 78627 1 4241
2 78628 1 4242
2 78629 1 4242
2 78630 1 4242
2 78631 1 4242
2 78632 1 4242
2 78633 1 4242
2 78634 1 4242
2 78635 1 4242
2 78636 1 4242
2 78637 1 4242
2 78638 1 4242
2 78639 1 4242
2 78640 1 4242
2 78641 1 4242
2 78642 1 4242
2 78643 1 4243
2 78644 1 4243
2 78645 1 4243
2 78646 1 4243
2 78647 1 4243
2 78648 1 4243
2 78649 1 4243
2 78650 1 4244
2 78651 1 4244
2 78652 1 4245
2 78653 1 4245
2 78654 1 4245
2 78655 1 4245
2 78656 1 4253
2 78657 1 4253
2 78658 1 4254
2 78659 1 4254
2 78660 1 4255
2 78661 1 4255
2 78662 1 4266
2 78663 1 4266
2 78664 1 4266
2 78665 1 4266
2 78666 1 4266
2 78667 1 4267
2 78668 1 4267
2 78669 1 4268
2 78670 1 4268
2 78671 1 4268
2 78672 1 4269
2 78673 1 4269
2 78674 1 4270
2 78675 1 4270
2 78676 1 4270
2 78677 1 4270
2 78678 1 4270
2 78679 1 4270
2 78680 1 4270
2 78681 1 4270
2 78682 1 4270
2 78683 1 4270
2 78684 1 4270
2 78685 1 4270
2 78686 1 4270
2 78687 1 4270
2 78688 1 4270
2 78689 1 4270
2 78690 1 4270
2 78691 1 4271
2 78692 1 4271
2 78693 1 4273
2 78694 1 4273
2 78695 1 4278
2 78696 1 4278
2 78697 1 4278
2 78698 1 4278
2 78699 1 4278
2 78700 1 4278
2 78701 1 4278
2 78702 1 4286
2 78703 1 4286
2 78704 1 4291
2 78705 1 4291
2 78706 1 4293
2 78707 1 4293
2 78708 1 4294
2 78709 1 4294
2 78710 1 4303
2 78711 1 4303
2 78712 1 4303
2 78713 1 4303
2 78714 1 4311
2 78715 1 4311
2 78716 1 4311
2 78717 1 4311
2 78718 1 4311
2 78719 1 4311
2 78720 1 4312
2 78721 1 4312
2 78722 1 4316
2 78723 1 4316
2 78724 1 4316
2 78725 1 4317
2 78726 1 4317
2 78727 1 4317
2 78728 1 4318
2 78729 1 4318
2 78730 1 4331
2 78731 1 4331
2 78732 1 4331
2 78733 1 4331
2 78734 1 4331
2 78735 1 4331
2 78736 1 4331
2 78737 1 4332
2 78738 1 4332
2 78739 1 4332
2 78740 1 4332
2 78741 1 4333
2 78742 1 4333
2 78743 1 4333
2 78744 1 4333
2 78745 1 4333
2 78746 1 4334
2 78747 1 4334
2 78748 1 4334
2 78749 1 4334
2 78750 1 4334
2 78751 1 4334
2 78752 1 4334
2 78753 1 4334
2 78754 1 4335
2 78755 1 4335
2 78756 1 4335
2 78757 1 4335
2 78758 1 4335
2 78759 1 4336
2 78760 1 4336
2 78761 1 4336
2 78762 1 4336
2 78763 1 4336
2 78764 1 4336
2 78765 1 4336
2 78766 1 4336
2 78767 1 4336
2 78768 1 4336
2 78769 1 4336
2 78770 1 4336
2 78771 1 4337
2 78772 1 4337
2 78773 1 4339
2 78774 1 4339
2 78775 1 4340
2 78776 1 4340
2 78777 1 4340
2 78778 1 4341
2 78779 1 4341
2 78780 1 4342
2 78781 1 4342
2 78782 1 4351
2 78783 1 4351
2 78784 1 4351
2 78785 1 4352
2 78786 1 4352
2 78787 1 4354
2 78788 1 4354
2 78789 1 4354
2 78790 1 4354
2 78791 1 4354
2 78792 1 4354
2 78793 1 4356
2 78794 1 4356
2 78795 1 4356
2 78796 1 4361
2 78797 1 4361
2 78798 1 4361
2 78799 1 4361
2 78800 1 4361
2 78801 1 4361
2 78802 1 4361
2 78803 1 4361
2 78804 1 4362
2 78805 1 4362
2 78806 1 4363
2 78807 1 4363
2 78808 1 4365
2 78809 1 4365
2 78810 1 4372
2 78811 1 4372
2 78812 1 4372
2 78813 1 4372
2 78814 1 4372
2 78815 1 4373
2 78816 1 4373
2 78817 1 4373
2 78818 1 4373
2 78819 1 4373
2 78820 1 4374
2 78821 1 4374
2 78822 1 4374
2 78823 1 4374
2 78824 1 4374
2 78825 1 4374
2 78826 1 4374
2 78827 1 4374
2 78828 1 4374
2 78829 1 4377
2 78830 1 4377
2 78831 1 4379
2 78832 1 4379
2 78833 1 4379
2 78834 1 4379
2 78835 1 4379
2 78836 1 4379
2 78837 1 4379
2 78838 1 4380
2 78839 1 4380
2 78840 1 4380
2 78841 1 4380
2 78842 1 4381
2 78843 1 4381
2 78844 1 4382
2 78845 1 4382
2 78846 1 4382
2 78847 1 4382
2 78848 1 4382
2 78849 1 4382
2 78850 1 4382
2 78851 1 4383
2 78852 1 4383
2 78853 1 4383
2 78854 1 4383
2 78855 1 4383
2 78856 1 4383
2 78857 1 4383
2 78858 1 4383
2 78859 1 4383
2 78860 1 4383
2 78861 1 4383
2 78862 1 4383
2 78863 1 4383
2 78864 1 4383
2 78865 1 4383
2 78866 1 4383
2 78867 1 4383
2 78868 1 4383
2 78869 1 4383
2 78870 1 4383
2 78871 1 4383
2 78872 1 4383
2 78873 1 4383
2 78874 1 4383
2 78875 1 4383
2 78876 1 4383
2 78877 1 4383
2 78878 1 4383
2 78879 1 4383
2 78880 1 4383
2 78881 1 4383
2 78882 1 4383
2 78883 1 4383
2 78884 1 4383
2 78885 1 4383
2 78886 1 4383
2 78887 1 4383
2 78888 1 4385
2 78889 1 4385
2 78890 1 4385
2 78891 1 4387
2 78892 1 4387
2 78893 1 4394
2 78894 1 4394
2 78895 1 4395
2 78896 1 4395
2 78897 1 4396
2 78898 1 4396
2 78899 1 4403
2 78900 1 4403
2 78901 1 4403
2 78902 1 4406
2 78903 1 4406
2 78904 1 4406
2 78905 1 4406
2 78906 1 4406
2 78907 1 4406
2 78908 1 4406
2 78909 1 4406
2 78910 1 4406
2 78911 1 4406
2 78912 1 4406
2 78913 1 4406
2 78914 1 4406
2 78915 1 4406
2 78916 1 4407
2 78917 1 4407
2 78918 1 4407
2 78919 1 4407
2 78920 1 4407
2 78921 1 4407
2 78922 1 4407
2 78923 1 4407
2 78924 1 4415
2 78925 1 4415
2 78926 1 4415
2 78927 1 4415
2 78928 1 4415
2 78929 1 4415
2 78930 1 4415
2 78931 1 4415
2 78932 1 4415
2 78933 1 4415
2 78934 1 4415
2 78935 1 4415
2 78936 1 4415
2 78937 1 4416
2 78938 1 4416
2 78939 1 4416
2 78940 1 4417
2 78941 1 4417
2 78942 1 4417
2 78943 1 4418
2 78944 1 4418
2 78945 1 4418
2 78946 1 4421
2 78947 1 4421
2 78948 1 4421
2 78949 1 4421
2 78950 1 4421
2 78951 1 4421
2 78952 1 4421
2 78953 1 4421
2 78954 1 4421
2 78955 1 4423
2 78956 1 4423
2 78957 1 4428
2 78958 1 4428
2 78959 1 4429
2 78960 1 4429
2 78961 1 4429
2 78962 1 4431
2 78963 1 4431
2 78964 1 4443
2 78965 1 4443
2 78966 1 4443
2 78967 1 4443
2 78968 1 4443
2 78969 1 4443
2 78970 1 4443
2 78971 1 4443
2 78972 1 4443
2 78973 1 4443
2 78974 1 4443
2 78975 1 4444
2 78976 1 4444
2 78977 1 4445
2 78978 1 4445
2 78979 1 4445
2 78980 1 4456
2 78981 1 4456
2 78982 1 4456
2 78983 1 4456
2 78984 1 4456
2 78985 1 4456
2 78986 1 4456
2 78987 1 4456
2 78988 1 4456
2 78989 1 4456
2 78990 1 4456
2 78991 1 4456
2 78992 1 4456
2 78993 1 4456
2 78994 1 4457
2 78995 1 4457
2 78996 1 4457
2 78997 1 4457
2 78998 1 4457
2 78999 1 4457
2 79000 1 4457
2 79001 1 4457
2 79002 1 4457
2 79003 1 4459
2 79004 1 4459
2 79005 1 4459
2 79006 1 4480
2 79007 1 4480
2 79008 1 4480
2 79009 1 4484
2 79010 1 4484
2 79011 1 4489
2 79012 1 4489
2 79013 1 4489
2 79014 1 4489
2 79015 1 4503
2 79016 1 4503
2 79017 1 4503
2 79018 1 4503
2 79019 1 4504
2 79020 1 4504
2 79021 1 4505
2 79022 1 4505
2 79023 1 4517
2 79024 1 4517
2 79025 1 4517
2 79026 1 4517
2 79027 1 4517
2 79028 1 4517
2 79029 1 4517
2 79030 1 4517
2 79031 1 4517
2 79032 1 4518
2 79033 1 4518
2 79034 1 4519
2 79035 1 4519
2 79036 1 4519
2 79037 1 4519
2 79038 1 4519
2 79039 1 4519
2 79040 1 4519
2 79041 1 4519
2 79042 1 4519
2 79043 1 4519
2 79044 1 4521
2 79045 1 4521
2 79046 1 4521
2 79047 1 4521
2 79048 1 4521
2 79049 1 4521
2 79050 1 4521
2 79051 1 4522
2 79052 1 4522
2 79053 1 4522
2 79054 1 4522
2 79055 1 4522
2 79056 1 4522
2 79057 1 4522
2 79058 1 4522
2 79059 1 4523
2 79060 1 4523
2 79061 1 4523
2 79062 1 4523
2 79063 1 4523
2 79064 1 4523
2 79065 1 4523
2 79066 1 4523
2 79067 1 4524
2 79068 1 4524
2 79069 1 4524
2 79070 1 4524
2 79071 1 4524
2 79072 1 4524
2 79073 1 4524
2 79074 1 4524
2 79075 1 4524
2 79076 1 4524
2 79077 1 4524
2 79078 1 4524
2 79079 1 4524
2 79080 1 4525
2 79081 1 4525
2 79082 1 4525
2 79083 1 4525
2 79084 1 4525
2 79085 1 4525
2 79086 1 4525
2 79087 1 4525
2 79088 1 4525
2 79089 1 4525
2 79090 1 4529
2 79091 1 4529
2 79092 1 4533
2 79093 1 4533
2 79094 1 4533
2 79095 1 4537
2 79096 1 4537
2 79097 1 4537
2 79098 1 4544
2 79099 1 4544
2 79100 1 4544
2 79101 1 4544
2 79102 1 4545
2 79103 1 4545
2 79104 1 4545
2 79105 1 4545
2 79106 1 4545
2 79107 1 4548
2 79108 1 4548
2 79109 1 4549
2 79110 1 4549
2 79111 1 4549
2 79112 1 4549
2 79113 1 4550
2 79114 1 4550
2 79115 1 4550
2 79116 1 4550
2 79117 1 4550
2 79118 1 4550
2 79119 1 4550
2 79120 1 4550
2 79121 1 4550
2 79122 1 4550
2 79123 1 4552
2 79124 1 4552
2 79125 1 4552
2 79126 1 4553
2 79127 1 4553
2 79128 1 4554
2 79129 1 4554
2 79130 1 4554
2 79131 1 4554
2 79132 1 4554
2 79133 1 4555
2 79134 1 4555
2 79135 1 4563
2 79136 1 4563
2 79137 1 4567
2 79138 1 4567
2 79139 1 4573
2 79140 1 4573
2 79141 1 4574
2 79142 1 4574
2 79143 1 4575
2 79144 1 4575
2 79145 1 4575
2 79146 1 4575
2 79147 1 4575
2 79148 1 4576
2 79149 1 4576
2 79150 1 4576
2 79151 1 4577
2 79152 1 4577
2 79153 1 4577
2 79154 1 4577
2 79155 1 4577
2 79156 1 4577
2 79157 1 4577
2 79158 1 4577
2 79159 1 4577
2 79160 1 4577
2 79161 1 4577
2 79162 1 4577
2 79163 1 4577
2 79164 1 4577
2 79165 1 4577
2 79166 1 4577
2 79167 1 4577
2 79168 1 4577
2 79169 1 4577
2 79170 1 4577
2 79171 1 4578
2 79172 1 4578
2 79173 1 4578
2 79174 1 4579
2 79175 1 4579
2 79176 1 4579
2 79177 1 4588
2 79178 1 4588
2 79179 1 4588
2 79180 1 4588
2 79181 1 4588
2 79182 1 4588
2 79183 1 4588
2 79184 1 4588
2 79185 1 4588
2 79186 1 4589
2 79187 1 4589
2 79188 1 4589
2 79189 1 4589
2 79190 1 4589
2 79191 1 4593
2 79192 1 4593
2 79193 1 4593
2 79194 1 4593
2 79195 1 4593
2 79196 1 4593
2 79197 1 4594
2 79198 1 4594
2 79199 1 4594
2 79200 1 4594
2 79201 1 4594
2 79202 1 4594
2 79203 1 4594
2 79204 1 4595
2 79205 1 4595
2 79206 1 4595
2 79207 1 4595
2 79208 1 4604
2 79209 1 4604
2 79210 1 4604
2 79211 1 4604
2 79212 1 4607
2 79213 1 4607
2 79214 1 4607
2 79215 1 4607
2 79216 1 4607
2 79217 1 4607
2 79218 1 4607
2 79219 1 4607
2 79220 1 4607
2 79221 1 4607
2 79222 1 4607
2 79223 1 4608
2 79224 1 4608
2 79225 1 4609
2 79226 1 4609
2 79227 1 4609
2 79228 1 4609
2 79229 1 4610
2 79230 1 4610
2 79231 1 4610
2 79232 1 4610
2 79233 1 4610
2 79234 1 4610
2 79235 1 4610
2 79236 1 4610
2 79237 1 4610
2 79238 1 4611
2 79239 1 4611
2 79240 1 4612
2 79241 1 4612
2 79242 1 4613
2 79243 1 4613
2 79244 1 4613
2 79245 1 4613
2 79246 1 4613
2 79247 1 4614
2 79248 1 4614
2 79249 1 4622
2 79250 1 4622
2 79251 1 4635
2 79252 1 4635
2 79253 1 4635
2 79254 1 4635
2 79255 1 4635
2 79256 1 4635
2 79257 1 4635
2 79258 1 4635
2 79259 1 4635
2 79260 1 4635
2 79261 1 4635
2 79262 1 4635
2 79263 1 4635
2 79264 1 4635
2 79265 1 4635
2 79266 1 4635
2 79267 1 4635
2 79268 1 4635
2 79269 1 4635
2 79270 1 4635
2 79271 1 4636
2 79272 1 4636
2 79273 1 4637
2 79274 1 4637
2 79275 1 4640
2 79276 1 4640
2 79277 1 4640
2 79278 1 4640
2 79279 1 4642
2 79280 1 4642
2 79281 1 4643
2 79282 1 4643
2 79283 1 4643
2 79284 1 4643
2 79285 1 4646
2 79286 1 4646
2 79287 1 4646
2 79288 1 4646
2 79289 1 4647
2 79290 1 4647
2 79291 1 4647
2 79292 1 4647
2 79293 1 4648
2 79294 1 4648
2 79295 1 4648
2 79296 1 4649
2 79297 1 4649
2 79298 1 4649
2 79299 1 4649
2 79300 1 4649
2 79301 1 4649
2 79302 1 4649
2 79303 1 4649
2 79304 1 4649
2 79305 1 4649
2 79306 1 4650
2 79307 1 4650
2 79308 1 4650
2 79309 1 4650
2 79310 1 4659
2 79311 1 4659
2 79312 1 4659
2 79313 1 4659
2 79314 1 4663
2 79315 1 4663
2 79316 1 4671
2 79317 1 4671
2 79318 1 4677
2 79319 1 4677
2 79320 1 4677
2 79321 1 4677
2 79322 1 4678
2 79323 1 4678
2 79324 1 4678
2 79325 1 4678
2 79326 1 4678
2 79327 1 4678
2 79328 1 4679
2 79329 1 4679
2 79330 1 4685
2 79331 1 4685
2 79332 1 4685
2 79333 1 4685
2 79334 1 4685
2 79335 1 4685
2 79336 1 4685
2 79337 1 4685
2 79338 1 4685
2 79339 1 4685
2 79340 1 4685
2 79341 1 4685
2 79342 1 4685
2 79343 1 4686
2 79344 1 4686
2 79345 1 4686
2 79346 1 4687
2 79347 1 4687
2 79348 1 4687
2 79349 1 4688
2 79350 1 4688
2 79351 1 4688
2 79352 1 4697
2 79353 1 4697
2 79354 1 4697
2 79355 1 4697
2 79356 1 4705
2 79357 1 4705
2 79358 1 4705
2 79359 1 4705
2 79360 1 4705
2 79361 1 4705
2 79362 1 4705
2 79363 1 4705
2 79364 1 4705
2 79365 1 4705
2 79366 1 4705
2 79367 1 4706
2 79368 1 4706
2 79369 1 4706
2 79370 1 4706
2 79371 1 4706
2 79372 1 4706
2 79373 1 4718
2 79374 1 4718
2 79375 1 4718
2 79376 1 4720
2 79377 1 4720
2 79378 1 4720
2 79379 1 4720
2 79380 1 4720
2 79381 1 4720
2 79382 1 4720
2 79383 1 4721
2 79384 1 4721
2 79385 1 4722
2 79386 1 4722
2 79387 1 4722
2 79388 1 4722
2 79389 1 4722
2 79390 1 4723
2 79391 1 4723
2 79392 1 4724
2 79393 1 4724
2 79394 1 4725
2 79395 1 4725
2 79396 1 4738
2 79397 1 4738
2 79398 1 4738
2 79399 1 4738
2 79400 1 4738
2 79401 1 4738
2 79402 1 4739
2 79403 1 4739
2 79404 1 4739
2 79405 1 4740
2 79406 1 4740
2 79407 1 4746
2 79408 1 4746
2 79409 1 4746
2 79410 1 4746
2 79411 1 4746
2 79412 1 4748
2 79413 1 4748
2 79414 1 4748
2 79415 1 4752
2 79416 1 4752
2 79417 1 4760
2 79418 1 4760
2 79419 1 4761
2 79420 1 4761
2 79421 1 4761
2 79422 1 4761
2 79423 1 4761
2 79424 1 4763
2 79425 1 4763
2 79426 1 4763
2 79427 1 4782
2 79428 1 4782
2 79429 1 4790
2 79430 1 4790
2 79431 1 4790
2 79432 1 4790
2 79433 1 4790
2 79434 1 4790
2 79435 1 4790
2 79436 1 4790
2 79437 1 4790
2 79438 1 4791
2 79439 1 4791
2 79440 1 4791
2 79441 1 4791
2 79442 1 4791
2 79443 1 4791
2 79444 1 4791
2 79445 1 4799
2 79446 1 4799
2 79447 1 4799
2 79448 1 4799
2 79449 1 4799
2 79450 1 4800
2 79451 1 4800
2 79452 1 4800
2 79453 1 4800
2 79454 1 4800
2 79455 1 4800
2 79456 1 4800
2 79457 1 4800
2 79458 1 4800
2 79459 1 4800
2 79460 1 4800
2 79461 1 4800
2 79462 1 4800
2 79463 1 4800
2 79464 1 4801
2 79465 1 4801
2 79466 1 4802
2 79467 1 4802
2 79468 1 4807
2 79469 1 4807
2 79470 1 4810
2 79471 1 4810
2 79472 1 4810
2 79473 1 4850
2 79474 1 4850
2 79475 1 4852
2 79476 1 4852
2 79477 1 4853
2 79478 1 4853
2 79479 1 4853
2 79480 1 4853
2 79481 1 4865
2 79482 1 4865
2 79483 1 4865
2 79484 1 4865
2 79485 1 4865
2 79486 1 4865
2 79487 1 4865
2 79488 1 4865
2 79489 1 4865
2 79490 1 4865
2 79491 1 4865
2 79492 1 4865
2 79493 1 4865
2 79494 1 4865
2 79495 1 4865
2 79496 1 4865
2 79497 1 4865
2 79498 1 4865
2 79499 1 4865
2 79500 1 4865
2 79501 1 4865
2 79502 1 4866
2 79503 1 4866
2 79504 1 4866
2 79505 1 4866
2 79506 1 4867
2 79507 1 4867
2 79508 1 4867
2 79509 1 4869
2 79510 1 4869
2 79511 1 4869
2 79512 1 4869
2 79513 1 4869
2 79514 1 4870
2 79515 1 4870
2 79516 1 4870
2 79517 1 4870
2 79518 1 4870
2 79519 1 4870
2 79520 1 4870
2 79521 1 4870
2 79522 1 4870
2 79523 1 4871
2 79524 1 4871
2 79525 1 4871
2 79526 1 4872
2 79527 1 4872
2 79528 1 4880
2 79529 1 4880
2 79530 1 4886
2 79531 1 4886
2 79532 1 4887
2 79533 1 4887
2 79534 1 4888
2 79535 1 4888
2 79536 1 4889
2 79537 1 4889
2 79538 1 4889
2 79539 1 4889
2 79540 1 4889
2 79541 1 4889
2 79542 1 4889
2 79543 1 4890
2 79544 1 4890
2 79545 1 4890
2 79546 1 4902
2 79547 1 4902
2 79548 1 4905
2 79549 1 4905
2 79550 1 4905
2 79551 1 4905
2 79552 1 4905
2 79553 1 4905
2 79554 1 4905
2 79555 1 4905
2 79556 1 4905
2 79557 1 4905
2 79558 1 4905
2 79559 1 4905
2 79560 1 4905
2 79561 1 4905
2 79562 1 4906
2 79563 1 4906
2 79564 1 4906
2 79565 1 4907
2 79566 1 4907
2 79567 1 4907
2 79568 1 4907
2 79569 1 4907
2 79570 1 4907
2 79571 1 4907
2 79572 1 4907
2 79573 1 4911
2 79574 1 4911
2 79575 1 4911
2 79576 1 4930
2 79577 1 4930
2 79578 1 4930
2 79579 1 4935
2 79580 1 4935
2 79581 1 4935
2 79582 1 4936
2 79583 1 4936
2 79584 1 4936
2 79585 1 4936
2 79586 1 4948
2 79587 1 4948
2 79588 1 4948
2 79589 1 4948
2 79590 1 4958
2 79591 1 4958
2 79592 1 4963
2 79593 1 4963
2 79594 1 4965
2 79595 1 4965
2 79596 1 4965
2 79597 1 4965
2 79598 1 4965
2 79599 1 4965
2 79600 1 4965
2 79601 1 4965
2 79602 1 4965
2 79603 1 4965
2 79604 1 4966
2 79605 1 4966
2 79606 1 4966
2 79607 1 4966
2 79608 1 4966
2 79609 1 4966
2 79610 1 4966
2 79611 1 4966
2 79612 1 4966
2 79613 1 4967
2 79614 1 4967
2 79615 1 4980
2 79616 1 4980
2 79617 1 4980
2 79618 1 4980
2 79619 1 4980
2 79620 1 4981
2 79621 1 4981
2 79622 1 4981
2 79623 1 4982
2 79624 1 4982
2 79625 1 4982
2 79626 1 4983
2 79627 1 4983
2 79628 1 4983
2 79629 1 4984
2 79630 1 4984
2 79631 1 4984
2 79632 1 4984
2 79633 1 4985
2 79634 1 4985
2 79635 1 4986
2 79636 1 4986
2 79637 1 4986
2 79638 1 4986
2 79639 1 4986
2 79640 1 4986
2 79641 1 4986
2 79642 1 4986
2 79643 1 4986
2 79644 1 4987
2 79645 1 4987
2 79646 1 5006
2 79647 1 5006
2 79648 1 5006
2 79649 1 5006
2 79650 1 5006
2 79651 1 5008
2 79652 1 5008
2 79653 1 5008
2 79654 1 5008
2 79655 1 5008
2 79656 1 5008
2 79657 1 5013
2 79658 1 5013
2 79659 1 5013
2 79660 1 5013
2 79661 1 5013
2 79662 1 5013
2 79663 1 5014
2 79664 1 5014
2 79665 1 5016
2 79666 1 5016
2 79667 1 5017
2 79668 1 5017
2 79669 1 5017
2 79670 1 5017
2 79671 1 5017
2 79672 1 5018
2 79673 1 5018
2 79674 1 5018
2 79675 1 5018
2 79676 1 5019
2 79677 1 5019
2 79678 1 5019
2 79679 1 5019
2 79680 1 5027
2 79681 1 5027
2 79682 1 5027
2 79683 1 5027
2 79684 1 5027
2 79685 1 5027
2 79686 1 5028
2 79687 1 5028
2 79688 1 5028
2 79689 1 5028
2 79690 1 5028
2 79691 1 5031
2 79692 1 5031
2 79693 1 5031
2 79694 1 5032
2 79695 1 5032
2 79696 1 5032
2 79697 1 5041
2 79698 1 5041
2 79699 1 5041
2 79700 1 5044
2 79701 1 5044
2 79702 1 5060
2 79703 1 5060
2 79704 1 5060
2 79705 1 5060
2 79706 1 5060
2 79707 1 5068
2 79708 1 5068
2 79709 1 5068
2 79710 1 5068
2 79711 1 5069
2 79712 1 5069
2 79713 1 5069
2 79714 1 5069
2 79715 1 5071
2 79716 1 5071
2 79717 1 5073
2 79718 1 5073
2 79719 1 5078
2 79720 1 5078
2 79721 1 5086
2 79722 1 5086
2 79723 1 5086
2 79724 1 5086
2 79725 1 5086
2 79726 1 5086
2 79727 1 5086
2 79728 1 5086
2 79729 1 5094
2 79730 1 5094
2 79731 1 5094
2 79732 1 5095
2 79733 1 5095
2 79734 1 5095
2 79735 1 5095
2 79736 1 5097
2 79737 1 5097
2 79738 1 5100
2 79739 1 5100
2 79740 1 5101
2 79741 1 5101
2 79742 1 5108
2 79743 1 5108
2 79744 1 5108
2 79745 1 5108
2 79746 1 5118
2 79747 1 5118
2 79748 1 5118
2 79749 1 5126
2 79750 1 5126
2 79751 1 5127
2 79752 1 5127
2 79753 1 5128
2 79754 1 5128
2 79755 1 5128
2 79756 1 5128
2 79757 1 5128
2 79758 1 5129
2 79759 1 5129
2 79760 1 5129
2 79761 1 5131
2 79762 1 5131
2 79763 1 5132
2 79764 1 5132
2 79765 1 5134
2 79766 1 5134
2 79767 1 5141
2 79768 1 5141
2 79769 1 5141
2 79770 1 5141
2 79771 1 5141
2 79772 1 5142
2 79773 1 5142
2 79774 1 5148
2 79775 1 5148
2 79776 1 5148
2 79777 1 5148
2 79778 1 5148
2 79779 1 5153
2 79780 1 5153
2 79781 1 5153
2 79782 1 5153
2 79783 1 5153
2 79784 1 5153
2 79785 1 5165
2 79786 1 5165
2 79787 1 5165
2 79788 1 5174
2 79789 1 5174
2 79790 1 5174
2 79791 1 5174
2 79792 1 5174
2 79793 1 5174
2 79794 1 5174
2 79795 1 5174
2 79796 1 5174
2 79797 1 5182
2 79798 1 5182
2 79799 1 5182
2 79800 1 5182
2 79801 1 5182
2 79802 1 5182
2 79803 1 5182
2 79804 1 5183
2 79805 1 5183
2 79806 1 5208
2 79807 1 5208
2 79808 1 5211
2 79809 1 5211
2 79810 1 5211
2 79811 1 5211
2 79812 1 5211
2 79813 1 5211
2 79814 1 5211
2 79815 1 5211
2 79816 1 5225
2 79817 1 5225
2 79818 1 5225
2 79819 1 5225
2 79820 1 5225
2 79821 1 5225
2 79822 1 5225
2 79823 1 5225
2 79824 1 5225
2 79825 1 5225
2 79826 1 5225
2 79827 1 5225
2 79828 1 5225
2 79829 1 5225
2 79830 1 5225
2 79831 1 5225
2 79832 1 5225
2 79833 1 5230
2 79834 1 5230
2 79835 1 5230
2 79836 1 5230
2 79837 1 5238
2 79838 1 5238
2 79839 1 5238
2 79840 1 5238
2 79841 1 5238
2 79842 1 5238
2 79843 1 5238
2 79844 1 5240
2 79845 1 5240
2 79846 1 5243
2 79847 1 5243
2 79848 1 5243
2 79849 1 5243
2 79850 1 5243
2 79851 1 5243
2 79852 1 5243
2 79853 1 5243
2 79854 1 5243
2 79855 1 5244
2 79856 1 5244
2 79857 1 5244
2 79858 1 5244
2 79859 1 5244
2 79860 1 5244
2 79861 1 5252
2 79862 1 5252
2 79863 1 5252
2 79864 1 5252
2 79865 1 5252
2 79866 1 5252
2 79867 1 5252
2 79868 1 5254
2 79869 1 5254
2 79870 1 5254
2 79871 1 5254
2 79872 1 5255
2 79873 1 5255
2 79874 1 5255
2 79875 1 5255
2 79876 1 5255
2 79877 1 5255
2 79878 1 5255
2 79879 1 5255
2 79880 1 5255
2 79881 1 5255
2 79882 1 5255
2 79883 1 5255
2 79884 1 5255
2 79885 1 5255
2 79886 1 5255
2 79887 1 5255
2 79888 1 5255
2 79889 1 5255
2 79890 1 5255
2 79891 1 5255
2 79892 1 5255
2 79893 1 5255
2 79894 1 5255
2 79895 1 5255
2 79896 1 5255
2 79897 1 5255
2 79898 1 5255
2 79899 1 5255
2 79900 1 5255
2 79901 1 5255
2 79902 1 5255
2 79903 1 5255
2 79904 1 5255
2 79905 1 5255
2 79906 1 5255
2 79907 1 5255
2 79908 1 5255
2 79909 1 5255
2 79910 1 5255
2 79911 1 5255
2 79912 1 5255
2 79913 1 5255
2 79914 1 5255
2 79915 1 5255
2 79916 1 5255
2 79917 1 5263
2 79918 1 5263
2 79919 1 5264
2 79920 1 5264
2 79921 1 5265
2 79922 1 5265
2 79923 1 5265
2 79924 1 5266
2 79925 1 5266
2 79926 1 5267
2 79927 1 5267
2 79928 1 5275
2 79929 1 5275
2 79930 1 5275
2 79931 1 5275
2 79932 1 5275
2 79933 1 5275
2 79934 1 5276
2 79935 1 5276
2 79936 1 5277
2 79937 1 5277
2 79938 1 5278
2 79939 1 5278
2 79940 1 5280
2 79941 1 5280
2 79942 1 5280
2 79943 1 5280
2 79944 1 5280
2 79945 1 5280
2 79946 1 5290
2 79947 1 5290
2 79948 1 5290
2 79949 1 5292
2 79950 1 5292
2 79951 1 5292
2 79952 1 5292
2 79953 1 5292
2 79954 1 5292
2 79955 1 5292
2 79956 1 5294
2 79957 1 5294
2 79958 1 5294
2 79959 1 5294
2 79960 1 5294
2 79961 1 5294
2 79962 1 5294
2 79963 1 5295
2 79964 1 5295
2 79965 1 5295
2 79966 1 5295
2 79967 1 5295
2 79968 1 5295
2 79969 1 5298
2 79970 1 5298
2 79971 1 5298
2 79972 1 5298
2 79973 1 5298
2 79974 1 5298
2 79975 1 5298
2 79976 1 5298
2 79977 1 5298
2 79978 1 5298
2 79979 1 5299
2 79980 1 5299
2 79981 1 5299
2 79982 1 5299
2 79983 1 5299
2 79984 1 5299
2 79985 1 5299
2 79986 1 5299
2 79987 1 5299
2 79988 1 5299
2 79989 1 5299
2 79990 1 5300
2 79991 1 5300
2 79992 1 5301
2 79993 1 5301
2 79994 1 5301
2 79995 1 5301
2 79996 1 5301
2 79997 1 5301
2 79998 1 5301
2 79999 1 5301
2 80000 1 5302
2 80001 1 5302
2 80002 1 5302
2 80003 1 5303
2 80004 1 5303
2 80005 1 5303
2 80006 1 5303
2 80007 1 5303
2 80008 1 5303
2 80009 1 5317
2 80010 1 5317
2 80011 1 5317
2 80012 1 5320
2 80013 1 5320
2 80014 1 5320
2 80015 1 5320
2 80016 1 5321
2 80017 1 5321
2 80018 1 5322
2 80019 1 5322
2 80020 1 5322
2 80021 1 5322
2 80022 1 5322
2 80023 1 5323
2 80024 1 5323
2 80025 1 5334
2 80026 1 5334
2 80027 1 5345
2 80028 1 5345
2 80029 1 5356
2 80030 1 5356
2 80031 1 5356
2 80032 1 5356
2 80033 1 5357
2 80034 1 5357
2 80035 1 5357
2 80036 1 5357
2 80037 1 5368
2 80038 1 5368
2 80039 1 5382
2 80040 1 5382
2 80041 1 5383
2 80042 1 5383
2 80043 1 5384
2 80044 1 5384
2 80045 1 5384
2 80046 1 5384
2 80047 1 5384
2 80048 1 5384
2 80049 1 5384
2 80050 1 5384
2 80051 1 5385
2 80052 1 5385
2 80053 1 5385
2 80054 1 5389
2 80055 1 5389
2 80056 1 5389
2 80057 1 5389
2 80058 1 5389
2 80059 1 5389
2 80060 1 5389
2 80061 1 5406
2 80062 1 5406
2 80063 1 5406
2 80064 1 5406
2 80065 1 5408
2 80066 1 5408
2 80067 1 5422
2 80068 1 5422
2 80069 1 5423
2 80070 1 5423
2 80071 1 5423
2 80072 1 5423
2 80073 1 5423
2 80074 1 5423
2 80075 1 5424
2 80076 1 5424
2 80077 1 5424
2 80078 1 5425
2 80079 1 5425
2 80080 1 5425
2 80081 1 5425
2 80082 1 5425
2 80083 1 5426
2 80084 1 5426
2 80085 1 5426
2 80086 1 5435
2 80087 1 5435
2 80088 1 5435
2 80089 1 5435
2 80090 1 5435
2 80091 1 5436
2 80092 1 5436
2 80093 1 5446
2 80094 1 5446
2 80095 1 5446
2 80096 1 5446
2 80097 1 5447
2 80098 1 5447
2 80099 1 5448
2 80100 1 5448
2 80101 1 5455
2 80102 1 5455
2 80103 1 5456
2 80104 1 5456
2 80105 1 5456
2 80106 1 5456
2 80107 1 5456
2 80108 1 5456
2 80109 1 5456
2 80110 1 5456
2 80111 1 5457
2 80112 1 5457
2 80113 1 5464
2 80114 1 5464
2 80115 1 5474
2 80116 1 5474
2 80117 1 5474
2 80118 1 5474
2 80119 1 5475
2 80120 1 5475
2 80121 1 5475
2 80122 1 5475
2 80123 1 5484
2 80124 1 5484
2 80125 1 5499
2 80126 1 5499
2 80127 1 5499
2 80128 1 5500
2 80129 1 5500
2 80130 1 5503
2 80131 1 5503
2 80132 1 5513
2 80133 1 5513
2 80134 1 5513
2 80135 1 5513
2 80136 1 5513
2 80137 1 5515
2 80138 1 5515
2 80139 1 5515
2 80140 1 5515
2 80141 1 5516
2 80142 1 5516
2 80143 1 5524
2 80144 1 5524
2 80145 1 5525
2 80146 1 5525
2 80147 1 5525
2 80148 1 5525
2 80149 1 5534
2 80150 1 5534
2 80151 1 5536
2 80152 1 5536
2 80153 1 5536
2 80154 1 5545
2 80155 1 5545
2 80156 1 5545
2 80157 1 5545
2 80158 1 5545
2 80159 1 5545
2 80160 1 5545
2 80161 1 5545
2 80162 1 5546
2 80163 1 5546
2 80164 1 5546
2 80165 1 5546
2 80166 1 5549
2 80167 1 5549
2 80168 1 5566
2 80169 1 5566
2 80170 1 5566
2 80171 1 5566
2 80172 1 5575
2 80173 1 5575
2 80174 1 5576
2 80175 1 5576
2 80176 1 5576
2 80177 1 5576
2 80178 1 5576
2 80179 1 5576
2 80180 1 5577
2 80181 1 5577
2 80182 1 5591
2 80183 1 5591
2 80184 1 5591
2 80185 1 5591
2 80186 1 5608
2 80187 1 5608
2 80188 1 5609
2 80189 1 5609
2 80190 1 5610
2 80191 1 5610
2 80192 1 5610
2 80193 1 5610
2 80194 1 5610
2 80195 1 5610
2 80196 1 5610
2 80197 1 5617
2 80198 1 5617
2 80199 1 5617
2 80200 1 5627
2 80201 1 5627
2 80202 1 5627
2 80203 1 5627
2 80204 1 5627
2 80205 1 5627
2 80206 1 5628
2 80207 1 5628
2 80208 1 5628
2 80209 1 5628
2 80210 1 5635
2 80211 1 5635
2 80212 1 5644
2 80213 1 5644
2 80214 1 5644
2 80215 1 5651
2 80216 1 5651
2 80217 1 5655
2 80218 1 5655
2 80219 1 5660
2 80220 1 5660
2 80221 1 5660
2 80222 1 5660
2 80223 1 5661
2 80224 1 5661
2 80225 1 5685
2 80226 1 5685
2 80227 1 5685
2 80228 1 5685
2 80229 1 5692
2 80230 1 5692
2 80231 1 5700
2 80232 1 5700
2 80233 1 5700
2 80234 1 5704
2 80235 1 5704
2 80236 1 5712
2 80237 1 5712
2 80238 1 5712
2 80239 1 5717
2 80240 1 5717
2 80241 1 5717
2 80242 1 5717
2 80243 1 5720
2 80244 1 5720
2 80245 1 5720
2 80246 1 5720
2 80247 1 5725
2 80248 1 5725
2 80249 1 5738
2 80250 1 5738
2 80251 1 5739
2 80252 1 5739
2 80253 1 5741
2 80254 1 5741
2 80255 1 5741
2 80256 1 5753
2 80257 1 5753
2 80258 1 5756
2 80259 1 5756
2 80260 1 5756
2 80261 1 5756
2 80262 1 5757
2 80263 1 5757
2 80264 1 5764
2 80265 1 5764
2 80266 1 5765
2 80267 1 5765
2 80268 1 5765
2 80269 1 5765
2 80270 1 5765
2 80271 1 5765
2 80272 1 5765
2 80273 1 5765
2 80274 1 5765
2 80275 1 5765
2 80276 1 5765
2 80277 1 5765
2 80278 1 5765
2 80279 1 5766
2 80280 1 5766
2 80281 1 5766
2 80282 1 5766
2 80283 1 5766
2 80284 1 5766
2 80285 1 5766
2 80286 1 5767
2 80287 1 5767
2 80288 1 5777
2 80289 1 5777
2 80290 1 5788
2 80291 1 5788
2 80292 1 5796
2 80293 1 5796
2 80294 1 5796
2 80295 1 5797
2 80296 1 5797
2 80297 1 5797
2 80298 1 5797
2 80299 1 5797
2 80300 1 5797
2 80301 1 5797
2 80302 1 5797
2 80303 1 5799
2 80304 1 5799
2 80305 1 5799
2 80306 1 5799
2 80307 1 5799
2 80308 1 5799
2 80309 1 5805
2 80310 1 5805
2 80311 1 5815
2 80312 1 5815
2 80313 1 5819
2 80314 1 5819
2 80315 1 5827
2 80316 1 5827
2 80317 1 5835
2 80318 1 5835
2 80319 1 5836
2 80320 1 5836
2 80321 1 5836
2 80322 1 5837
2 80323 1 5837
2 80324 1 5837
2 80325 1 5837
2 80326 1 5837
2 80327 1 5837
2 80328 1 5837
2 80329 1 5837
2 80330 1 5837
2 80331 1 5837
2 80332 1 5863
2 80333 1 5863
2 80334 1 5863
2 80335 1 5863
2 80336 1 5864
2 80337 1 5864
2 80338 1 5866
2 80339 1 5866
2 80340 1 5866
2 80341 1 5866
2 80342 1 5866
2 80343 1 5867
2 80344 1 5867
2 80345 1 5867
2 80346 1 5885
2 80347 1 5885
2 80348 1 5896
2 80349 1 5896
2 80350 1 5896
2 80351 1 5903
2 80352 1 5903
2 80353 1 5910
2 80354 1 5910
2 80355 1 5910
2 80356 1 5910
2 80357 1 5910
2 80358 1 5910
2 80359 1 5910
2 80360 1 5911
2 80361 1 5911
2 80362 1 5917
2 80363 1 5917
2 80364 1 5918
2 80365 1 5918
2 80366 1 5925
2 80367 1 5925
2 80368 1 5925
2 80369 1 5927
2 80370 1 5927
2 80371 1 5930
2 80372 1 5930
2 80373 1 5930
2 80374 1 5930
2 80375 1 5930
2 80376 1 5930
2 80377 1 5930
2 80378 1 5931
2 80379 1 5931
2 80380 1 5934
2 80381 1 5934
2 80382 1 5935
2 80383 1 5935
2 80384 1 5935
2 80385 1 5935
2 80386 1 5935
2 80387 1 5938
2 80388 1 5938
2 80389 1 5950
2 80390 1 5950
2 80391 1 5961
2 80392 1 5961
2 80393 1 5962
2 80394 1 5962
2 80395 1 5962
2 80396 1 5962
2 80397 1 5962
2 80398 1 5962
2 80399 1 5962
2 80400 1 5962
2 80401 1 5962
2 80402 1 5962
2 80403 1 5962
2 80404 1 5965
2 80405 1 5965
2 80406 1 5972
2 80407 1 5972
2 80408 1 5973
2 80409 1 5973
2 80410 1 5973
2 80411 1 5977
2 80412 1 5977
2 80413 1 5977
2 80414 1 5977
2 80415 1 5977
2 80416 1 5977
2 80417 1 5977
2 80418 1 5977
2 80419 1 5977
2 80420 1 5977
2 80421 1 5977
2 80422 1 5977
2 80423 1 5977
2 80424 1 5977
2 80425 1 5977
2 80426 1 5977
2 80427 1 5977
2 80428 1 5977
2 80429 1 5977
2 80430 1 5977
2 80431 1 5977
2 80432 1 5977
2 80433 1 5977
2 80434 1 5977
2 80435 1 5977
2 80436 1 5977
2 80437 1 5977
2 80438 1 5977
2 80439 1 5977
2 80440 1 5977
2 80441 1 5977
2 80442 1 5977
2 80443 1 5977
2 80444 1 5977
2 80445 1 5978
2 80446 1 5978
2 80447 1 5978
2 80448 1 5978
2 80449 1 5978
2 80450 1 5978
2 80451 1 5978
2 80452 1 5979
2 80453 1 5979
2 80454 1 5979
2 80455 1 5980
2 80456 1 5980
2 80457 1 5980
2 80458 1 5980
2 80459 1 5980
2 80460 1 5980
2 80461 1 5980
2 80462 1 5980
2 80463 1 5980
2 80464 1 5981
2 80465 1 5981
2 80466 1 5992
2 80467 1 5992
2 80468 1 5992
2 80469 1 5992
2 80470 1 5994
2 80471 1 5994
2 80472 1 5995
2 80473 1 5995
2 80474 1 6004
2 80475 1 6004
2 80476 1 6004
2 80477 1 6004
2 80478 1 6004
2 80479 1 6005
2 80480 1 6005
2 80481 1 6005
2 80482 1 6005
2 80483 1 6006
2 80484 1 6006
2 80485 1 6006
2 80486 1 6007
2 80487 1 6007
2 80488 1 6007
2 80489 1 6007
2 80490 1 6007
2 80491 1 6007
2 80492 1 6007
2 80493 1 6007
2 80494 1 6007
2 80495 1 6007
2 80496 1 6007
2 80497 1 6007
2 80498 1 6007
2 80499 1 6007
2 80500 1 6007
2 80501 1 6010
2 80502 1 6010
2 80503 1 6010
2 80504 1 6010
2 80505 1 6010
2 80506 1 6010
2 80507 1 6010
2 80508 1 6010
2 80509 1 6011
2 80510 1 6011
2 80511 1 6011
2 80512 1 6011
2 80513 1 6011
2 80514 1 6011
2 80515 1 6011
2 80516 1 6011
2 80517 1 6011
2 80518 1 6011
2 80519 1 6011
2 80520 1 6011
2 80521 1 6011
2 80522 1 6011
2 80523 1 6011
2 80524 1 6011
2 80525 1 6011
2 80526 1 6011
2 80527 1 6012
2 80528 1 6012
2 80529 1 6012
2 80530 1 6012
2 80531 1 6014
2 80532 1 6014
2 80533 1 6015
2 80534 1 6015
2 80535 1 6015
2 80536 1 6023
2 80537 1 6023
2 80538 1 6027
2 80539 1 6027
2 80540 1 6030
2 80541 1 6030
2 80542 1 6030
2 80543 1 6031
2 80544 1 6031
2 80545 1 6031
2 80546 1 6031
2 80547 1 6031
2 80548 1 6031
2 80549 1 6044
2 80550 1 6044
2 80551 1 6044
2 80552 1 6044
2 80553 1 6044
2 80554 1 6044
2 80555 1 6044
2 80556 1 6044
2 80557 1 6044
2 80558 1 6044
2 80559 1 6044
2 80560 1 6044
2 80561 1 6044
2 80562 1 6044
2 80563 1 6044
2 80564 1 6044
2 80565 1 6044
2 80566 1 6044
2 80567 1 6045
2 80568 1 6045
2 80569 1 6045
2 80570 1 6045
2 80571 1 6045
2 80572 1 6046
2 80573 1 6046
2 80574 1 6047
2 80575 1 6047
2 80576 1 6047
2 80577 1 6047
2 80578 1 6061
2 80579 1 6061
2 80580 1 6061
2 80581 1 6061
2 80582 1 6063
2 80583 1 6063
2 80584 1 6072
2 80585 1 6072
2 80586 1 6072
2 80587 1 6072
2 80588 1 6072
2 80589 1 6072
2 80590 1 6073
2 80591 1 6073
2 80592 1 6073
2 80593 1 6073
2 80594 1 6073
2 80595 1 6073
2 80596 1 6074
2 80597 1 6074
2 80598 1 6075
2 80599 1 6075
2 80600 1 6076
2 80601 1 6076
2 80602 1 6076
2 80603 1 6085
2 80604 1 6085
2 80605 1 6085
2 80606 1 6085
2 80607 1 6085
2 80608 1 6086
2 80609 1 6086
2 80610 1 6094
2 80611 1 6094
2 80612 1 6094
2 80613 1 6103
2 80614 1 6103
2 80615 1 6105
2 80616 1 6105
2 80617 1 6109
2 80618 1 6109
2 80619 1 6110
2 80620 1 6110
2 80621 1 6110
2 80622 1 6111
2 80623 1 6111
2 80624 1 6111
2 80625 1 6111
2 80626 1 6111
2 80627 1 6111
2 80628 1 6111
2 80629 1 6112
2 80630 1 6112
2 80631 1 6116
2 80632 1 6116
2 80633 1 6116
2 80634 1 6133
2 80635 1 6133
2 80636 1 6133
2 80637 1 6133
2 80638 1 6133
2 80639 1 6134
2 80640 1 6134
2 80641 1 6143
2 80642 1 6143
2 80643 1 6143
2 80644 1 6151
2 80645 1 6151
2 80646 1 6159
2 80647 1 6159
2 80648 1 6159
2 80649 1 6161
2 80650 1 6161
2 80651 1 6161
2 80652 1 6175
2 80653 1 6175
2 80654 1 6183
2 80655 1 6183
2 80656 1 6183
2 80657 1 6185
2 80658 1 6185
2 80659 1 6185
2 80660 1 6185
2 80661 1 6185
2 80662 1 6185
2 80663 1 6192
2 80664 1 6192
2 80665 1 6192
2 80666 1 6192
2 80667 1 6192
2 80668 1 6200
2 80669 1 6200
2 80670 1 6200
2 80671 1 6200
2 80672 1 6200
2 80673 1 6200
2 80674 1 6200
2 80675 1 6201
2 80676 1 6201
2 80677 1 6208
2 80678 1 6208
2 80679 1 6208
2 80680 1 6208
2 80681 1 6208
2 80682 1 6208
2 80683 1 6208
2 80684 1 6221
2 80685 1 6221
2 80686 1 6221
2 80687 1 6222
2 80688 1 6222
2 80689 1 6222
2 80690 1 6230
2 80691 1 6230
2 80692 1 6233
2 80693 1 6233
2 80694 1 6235
2 80695 1 6235
2 80696 1 6238
2 80697 1 6238
2 80698 1 6238
2 80699 1 6238
2 80700 1 6239
2 80701 1 6239
2 80702 1 6239
2 80703 1 6239
2 80704 1 6239
2 80705 1 6241
2 80706 1 6241
2 80707 1 6247
2 80708 1 6247
2 80709 1 6249
2 80710 1 6249
2 80711 1 6249
2 80712 1 6249
2 80713 1 6249
2 80714 1 6249
2 80715 1 6249
2 80716 1 6249
2 80717 1 6250
2 80718 1 6250
2 80719 1 6253
2 80720 1 6253
2 80721 1 6255
2 80722 1 6255
2 80723 1 6285
2 80724 1 6285
2 80725 1 6285
2 80726 1 6285
2 80727 1 6285
2 80728 1 6285
2 80729 1 6285
2 80730 1 6286
2 80731 1 6286
2 80732 1 6286
2 80733 1 6289
2 80734 1 6289
2 80735 1 6289
2 80736 1 6289
2 80737 1 6292
2 80738 1 6292
2 80739 1 6292
2 80740 1 6292
2 80741 1 6294
2 80742 1 6294
2 80743 1 6297
2 80744 1 6297
2 80745 1 6298
2 80746 1 6298
2 80747 1 6300
2 80748 1 6300
2 80749 1 6307
2 80750 1 6307
2 80751 1 6307
2 80752 1 6317
2 80753 1 6317
2 80754 1 6318
2 80755 1 6318
2 80756 1 6319
2 80757 1 6319
2 80758 1 6327
2 80759 1 6327
2 80760 1 6327
2 80761 1 6327
2 80762 1 6327
2 80763 1 6327
2 80764 1 6327
2 80765 1 6332
2 80766 1 6332
2 80767 1 6332
2 80768 1 6332
2 80769 1 6332
2 80770 1 6332
2 80771 1 6332
2 80772 1 6332
2 80773 1 6333
2 80774 1 6333
2 80775 1 6333
2 80776 1 6333
2 80777 1 6334
2 80778 1 6334
2 80779 1 6334
2 80780 1 6336
2 80781 1 6336
2 80782 1 6336
2 80783 1 6336
2 80784 1 6338
2 80785 1 6338
2 80786 1 6338
2 80787 1 6338
2 80788 1 6338
2 80789 1 6338
2 80790 1 6338
2 80791 1 6338
2 80792 1 6338
2 80793 1 6340
2 80794 1 6340
2 80795 1 6341
2 80796 1 6341
2 80797 1 6341
2 80798 1 6341
2 80799 1 6341
2 80800 1 6341
2 80801 1 6341
2 80802 1 6341
2 80803 1 6341
2 80804 1 6341
2 80805 1 6341
2 80806 1 6341
2 80807 1 6341
2 80808 1 6341
2 80809 1 6341
2 80810 1 6341
2 80811 1 6341
2 80812 1 6341
2 80813 1 6341
2 80814 1 6341
2 80815 1 6341
2 80816 1 6341
2 80817 1 6341
2 80818 1 6341
2 80819 1 6341
2 80820 1 6341
2 80821 1 6341
2 80822 1 6341
2 80823 1 6342
2 80824 1 6342
2 80825 1 6342
2 80826 1 6342
2 80827 1 6342
2 80828 1 6342
2 80829 1 6342
2 80830 1 6342
2 80831 1 6343
2 80832 1 6343
2 80833 1 6343
2 80834 1 6343
2 80835 1 6349
2 80836 1 6349
2 80837 1 6349
2 80838 1 6349
2 80839 1 6349
2 80840 1 6349
2 80841 1 6359
2 80842 1 6359
2 80843 1 6362
2 80844 1 6362
2 80845 1 6362
2 80846 1 6362
2 80847 1 6365
2 80848 1 6365
2 80849 1 6365
2 80850 1 6365
2 80851 1 6365
2 80852 1 6366
2 80853 1 6366
2 80854 1 6368
2 80855 1 6368
2 80856 1 6370
2 80857 1 6370
2 80858 1 6373
2 80859 1 6373
2 80860 1 6373
2 80861 1 6373
2 80862 1 6373
2 80863 1 6373
2 80864 1 6373
2 80865 1 6373
2 80866 1 6373
2 80867 1 6373
2 80868 1 6373
2 80869 1 6373
2 80870 1 6373
2 80871 1 6373
2 80872 1 6373
2 80873 1 6373
2 80874 1 6373
2 80875 1 6373
2 80876 1 6373
2 80877 1 6373
2 80878 1 6373
2 80879 1 6374
2 80880 1 6374
2 80881 1 6374
2 80882 1 6382
2 80883 1 6382
2 80884 1 6382
2 80885 1 6382
2 80886 1 6382
2 80887 1 6384
2 80888 1 6384
2 80889 1 6384
2 80890 1 6384
2 80891 1 6385
2 80892 1 6385
2 80893 1 6385
2 80894 1 6393
2 80895 1 6393
2 80896 1 6393
2 80897 1 6393
2 80898 1 6393
2 80899 1 6393
2 80900 1 6393
2 80901 1 6396
2 80902 1 6396
2 80903 1 6406
2 80904 1 6406
2 80905 1 6406
2 80906 1 6406
2 80907 1 6406
2 80908 1 6407
2 80909 1 6407
2 80910 1 6407
2 80911 1 6407
2 80912 1 6407
2 80913 1 6407
2 80914 1 6407
2 80915 1 6407
2 80916 1 6407
2 80917 1 6407
2 80918 1 6407
2 80919 1 6413
2 80920 1 6413
2 80921 1 6413
2 80922 1 6413
2 80923 1 6438
2 80924 1 6438
2 80925 1 6439
2 80926 1 6439
2 80927 1 6439
2 80928 1 6439
2 80929 1 6439
2 80930 1 6439
2 80931 1 6439
2 80932 1 6439
2 80933 1 6439
2 80934 1 6439
2 80935 1 6439
2 80936 1 6439
2 80937 1 6439
2 80938 1 6439
2 80939 1 6440
2 80940 1 6440
2 80941 1 6440
2 80942 1 6440
2 80943 1 6440
2 80944 1 6440
2 80945 1 6443
2 80946 1 6443
2 80947 1 6443
2 80948 1 6443
2 80949 1 6443
2 80950 1 6444
2 80951 1 6444
2 80952 1 6448
2 80953 1 6448
2 80954 1 6462
2 80955 1 6462
2 80956 1 6464
2 80957 1 6464
2 80958 1 6464
2 80959 1 6464
2 80960 1 6464
2 80961 1 6465
2 80962 1 6465
2 80963 1 6465
2 80964 1 6474
2 80965 1 6474
2 80966 1 6474
2 80967 1 6475
2 80968 1 6475
2 80969 1 6477
2 80970 1 6477
2 80971 1 6477
2 80972 1 6477
2 80973 1 6477
2 80974 1 6477
2 80975 1 6477
2 80976 1 6478
2 80977 1 6478
2 80978 1 6482
2 80979 1 6482
2 80980 1 6483
2 80981 1 6483
2 80982 1 6483
2 80983 1 6483
2 80984 1 6483
2 80985 1 6483
2 80986 1 6483
2 80987 1 6483
2 80988 1 6485
2 80989 1 6485
2 80990 1 6485
2 80991 1 6485
2 80992 1 6485
2 80993 1 6488
2 80994 1 6488
2 80995 1 6507
2 80996 1 6507
2 80997 1 6507
2 80998 1 6507
2 80999 1 6509
2 81000 1 6509
2 81001 1 6512
2 81002 1 6512
2 81003 1 6512
2 81004 1 6516
2 81005 1 6516
2 81006 1 6525
2 81007 1 6525
2 81008 1 6525
2 81009 1 6525
2 81010 1 6525
2 81011 1 6525
2 81012 1 6525
2 81013 1 6525
2 81014 1 6525
2 81015 1 6529
2 81016 1 6529
2 81017 1 6529
2 81018 1 6529
2 81019 1 6529
2 81020 1 6529
2 81021 1 6529
2 81022 1 6529
2 81023 1 6530
2 81024 1 6530
2 81025 1 6530
2 81026 1 6530
2 81027 1 6530
2 81028 1 6530
2 81029 1 6530
2 81030 1 6531
2 81031 1 6531
2 81032 1 6544
2 81033 1 6544
2 81034 1 6544
2 81035 1 6544
2 81036 1 6544
2 81037 1 6544
2 81038 1 6544
2 81039 1 6544
2 81040 1 6544
2 81041 1 6544
2 81042 1 6544
2 81043 1 6544
2 81044 1 6544
2 81045 1 6544
2 81046 1 6544
2 81047 1 6544
2 81048 1 6546
2 81049 1 6546
2 81050 1 6546
2 81051 1 6546
2 81052 1 6547
2 81053 1 6547
2 81054 1 6547
2 81055 1 6547
2 81056 1 6548
2 81057 1 6548
2 81058 1 6548
2 81059 1 6550
2 81060 1 6550
2 81061 1 6551
2 81062 1 6551
2 81063 1 6552
2 81064 1 6552
2 81065 1 6556
2 81066 1 6556
2 81067 1 6556
2 81068 1 6556
2 81069 1 6556
2 81070 1 6556
2 81071 1 6556
2 81072 1 6556
2 81073 1 6557
2 81074 1 6557
2 81075 1 6557
2 81076 1 6557
2 81077 1 6557
2 81078 1 6557
2 81079 1 6557
2 81080 1 6557
2 81081 1 6557
2 81082 1 6557
2 81083 1 6557
2 81084 1 6558
2 81085 1 6558
2 81086 1 6559
2 81087 1 6559
2 81088 1 6559
2 81089 1 6559
2 81090 1 6559
2 81091 1 6563
2 81092 1 6563
2 81093 1 6570
2 81094 1 6570
2 81095 1 6574
2 81096 1 6574
2 81097 1 6575
2 81098 1 6575
2 81099 1 6575
2 81100 1 6575
2 81101 1 6575
2 81102 1 6576
2 81103 1 6576
2 81104 1 6576
2 81105 1 6577
2 81106 1 6577
2 81107 1 6609
2 81108 1 6609
2 81109 1 6610
2 81110 1 6610
2 81111 1 6610
2 81112 1 6610
2 81113 1 6610
2 81114 1 6610
2 81115 1 6610
2 81116 1 6610
2 81117 1 6610
2 81118 1 6610
2 81119 1 6610
2 81120 1 6610
2 81121 1 6610
2 81122 1 6610
2 81123 1 6611
2 81124 1 6611
2 81125 1 6611
2 81126 1 6611
2 81127 1 6611
2 81128 1 6613
2 81129 1 6613
2 81130 1 6627
2 81131 1 6627
2 81132 1 6627
2 81133 1 6628
2 81134 1 6628
2 81135 1 6628
2 81136 1 6628
2 81137 1 6628
2 81138 1 6628
2 81139 1 6628
2 81140 1 6628
2 81141 1 6628
2 81142 1 6628
2 81143 1 6628
2 81144 1 6628
2 81145 1 6628
2 81146 1 6628
2 81147 1 6628
2 81148 1 6638
2 81149 1 6638
2 81150 1 6652
2 81151 1 6652
2 81152 1 6652
2 81153 1 6654
2 81154 1 6654
2 81155 1 6656
2 81156 1 6656
2 81157 1 6657
2 81158 1 6657
2 81159 1 6657
2 81160 1 6657
2 81161 1 6658
2 81162 1 6658
2 81163 1 6658
2 81164 1 6658
2 81165 1 6659
2 81166 1 6659
2 81167 1 6660
2 81168 1 6660
2 81169 1 6660
2 81170 1 6661
2 81171 1 6661
2 81172 1 6662
2 81173 1 6662
2 81174 1 6665
2 81175 1 6665
2 81176 1 6669
2 81177 1 6669
2 81178 1 6669
2 81179 1 6671
2 81180 1 6671
2 81181 1 6672
2 81182 1 6672
2 81183 1 6679
2 81184 1 6679
2 81185 1 6679
2 81186 1 6679
2 81187 1 6679
2 81188 1 6679
2 81189 1 6680
2 81190 1 6680
2 81191 1 6680
2 81192 1 6680
2 81193 1 6688
2 81194 1 6688
2 81195 1 6690
2 81196 1 6690
2 81197 1 6690
2 81198 1 6690
2 81199 1 6690
2 81200 1 6691
2 81201 1 6691
2 81202 1 6691
2 81203 1 6693
2 81204 1 6693
2 81205 1 6695
2 81206 1 6695
2 81207 1 6697
2 81208 1 6697
2 81209 1 6699
2 81210 1 6699
2 81211 1 6723
2 81212 1 6723
2 81213 1 6724
2 81214 1 6724
2 81215 1 6724
2 81216 1 6724
2 81217 1 6724
2 81218 1 6724
2 81219 1 6725
2 81220 1 6725
2 81221 1 6732
2 81222 1 6732
2 81223 1 6732
2 81224 1 6732
2 81225 1 6735
2 81226 1 6735
2 81227 1 6735
2 81228 1 6740
2 81229 1 6740
2 81230 1 6742
2 81231 1 6742
2 81232 1 6742
2 81233 1 6743
2 81234 1 6743
2 81235 1 6743
2 81236 1 6743
2 81237 1 6743
2 81238 1 6743
2 81239 1 6745
2 81240 1 6745
2 81241 1 6746
2 81242 1 6746
2 81243 1 6759
2 81244 1 6759
2 81245 1 6759
2 81246 1 6759
2 81247 1 6759
2 81248 1 6759
2 81249 1 6759
2 81250 1 6759
2 81251 1 6759
2 81252 1 6759
2 81253 1 6759
2 81254 1 6759
2 81255 1 6759
2 81256 1 6759
2 81257 1 6759
2 81258 1 6759
2 81259 1 6759
2 81260 1 6759
2 81261 1 6759
2 81262 1 6759
2 81263 1 6759
2 81264 1 6759
2 81265 1 6759
2 81266 1 6760
2 81267 1 6760
2 81268 1 6760
2 81269 1 6760
2 81270 1 6760
2 81271 1 6760
2 81272 1 6760
2 81273 1 6760
2 81274 1 6765
2 81275 1 6765
2 81276 1 6765
2 81277 1 6765
2 81278 1 6765
2 81279 1 6772
2 81280 1 6772
2 81281 1 6773
2 81282 1 6773
2 81283 1 6775
2 81284 1 6775
2 81285 1 6780
2 81286 1 6780
2 81287 1 6780
2 81288 1 6785
2 81289 1 6785
2 81290 1 6799
2 81291 1 6799
2 81292 1 6800
2 81293 1 6800
2 81294 1 6801
2 81295 1 6801
2 81296 1 6801
2 81297 1 6801
2 81298 1 6802
2 81299 1 6802
2 81300 1 6802
2 81301 1 6805
2 81302 1 6805
2 81303 1 6805
2 81304 1 6805
2 81305 1 6805
2 81306 1 6805
2 81307 1 6805
2 81308 1 6805
2 81309 1 6823
2 81310 1 6823
2 81311 1 6825
2 81312 1 6825
2 81313 1 6827
2 81314 1 6827
2 81315 1 6828
2 81316 1 6828
2 81317 1 6829
2 81318 1 6829
2 81319 1 6829
2 81320 1 6843
2 81321 1 6843
2 81322 1 6864
2 81323 1 6864
2 81324 1 6864
2 81325 1 6864
2 81326 1 6864
2 81327 1 6864
2 81328 1 6864
2 81329 1 6864
2 81330 1 6864
2 81331 1 6864
2 81332 1 6864
2 81333 1 6864
2 81334 1 6864
2 81335 1 6864
2 81336 1 6864
2 81337 1 6864
2 81338 1 6864
2 81339 1 6864
2 81340 1 6864
2 81341 1 6864
2 81342 1 6864
2 81343 1 6873
2 81344 1 6873
2 81345 1 6875
2 81346 1 6875
2 81347 1 6875
2 81348 1 6875
2 81349 1 6875
2 81350 1 6887
2 81351 1 6887
2 81352 1 6887
2 81353 1 6887
2 81354 1 6887
2 81355 1 6887
2 81356 1 6887
2 81357 1 6887
2 81358 1 6888
2 81359 1 6888
2 81360 1 6888
2 81361 1 6888
2 81362 1 6888
2 81363 1 6891
2 81364 1 6891
2 81365 1 6891
2 81366 1 6891
2 81367 1 6891
2 81368 1 6891
2 81369 1 6893
2 81370 1 6893
2 81371 1 6900
2 81372 1 6900
2 81373 1 6900
2 81374 1 6900
2 81375 1 6901
2 81376 1 6901
2 81377 1 6901
2 81378 1 6901
2 81379 1 6905
2 81380 1 6905
2 81381 1 6905
2 81382 1 6905
2 81383 1 6905
2 81384 1 6905
2 81385 1 6905
2 81386 1 6905
2 81387 1 6905
2 81388 1 6905
2 81389 1 6905
2 81390 1 6905
2 81391 1 6905
2 81392 1 6905
2 81393 1 6905
2 81394 1 6905
2 81395 1 6905
2 81396 1 6905
2 81397 1 6905
2 81398 1 6905
2 81399 1 6905
2 81400 1 6905
2 81401 1 6905
2 81402 1 6905
2 81403 1 6905
2 81404 1 6905
2 81405 1 6905
2 81406 1 6905
2 81407 1 6905
2 81408 1 6905
2 81409 1 6905
2 81410 1 6905
2 81411 1 6905
2 81412 1 6906
2 81413 1 6906
2 81414 1 6906
2 81415 1 6906
2 81416 1 6915
2 81417 1 6915
2 81418 1 6915
2 81419 1 6917
2 81420 1 6917
2 81421 1 6917
2 81422 1 6920
2 81423 1 6920
2 81424 1 6920
2 81425 1 6920
2 81426 1 6920
2 81427 1 6920
2 81428 1 6920
2 81429 1 6920
2 81430 1 6920
2 81431 1 6920
2 81432 1 6920
2 81433 1 6920
2 81434 1 6920
2 81435 1 6922
2 81436 1 6922
2 81437 1 6938
2 81438 1 6938
2 81439 1 6939
2 81440 1 6939
2 81441 1 6939
2 81442 1 6939
2 81443 1 6939
2 81444 1 6939
2 81445 1 6939
2 81446 1 6939
2 81447 1 6939
2 81448 1 6939
2 81449 1 6965
2 81450 1 6965
2 81451 1 6965
2 81452 1 6966
2 81453 1 6966
2 81454 1 6966
2 81455 1 6966
2 81456 1 6966
2 81457 1 6966
2 81458 1 6966
2 81459 1 6968
2 81460 1 6968
2 81461 1 6969
2 81462 1 6969
2 81463 1 6969
2 81464 1 6969
2 81465 1 6969
2 81466 1 6969
2 81467 1 6969
2 81468 1 6969
2 81469 1 6969
2 81470 1 6969
2 81471 1 6969
2 81472 1 6969
2 81473 1 6969
2 81474 1 6969
2 81475 1 6969
2 81476 1 6969
2 81477 1 6985
2 81478 1 6985
2 81479 1 6995
2 81480 1 6995
2 81481 1 6995
2 81482 1 6995
2 81483 1 6995
2 81484 1 6995
2 81485 1 7003
2 81486 1 7003
2 81487 1 7003
2 81488 1 7008
2 81489 1 7008
2 81490 1 7011
2 81491 1 7011
2 81492 1 7011
2 81493 1 7011
2 81494 1 7011
2 81495 1 7011
2 81496 1 7011
2 81497 1 7011
2 81498 1 7011
2 81499 1 7011
2 81500 1 7011
2 81501 1 7011
2 81502 1 7011
2 81503 1 7011
2 81504 1 7011
2 81505 1 7011
2 81506 1 7011
2 81507 1 7011
2 81508 1 7011
2 81509 1 7011
2 81510 1 7011
2 81511 1 7011
2 81512 1 7011
2 81513 1 7011
2 81514 1 7012
2 81515 1 7012
2 81516 1 7012
2 81517 1 7012
2 81518 1 7019
2 81519 1 7019
2 81520 1 7022
2 81521 1 7022
2 81522 1 7022
2 81523 1 7022
2 81524 1 7023
2 81525 1 7023
2 81526 1 7034
2 81527 1 7034
2 81528 1 7034
2 81529 1 7034
2 81530 1 7034
2 81531 1 7034
2 81532 1 7035
2 81533 1 7035
2 81534 1 7035
2 81535 1 7036
2 81536 1 7036
2 81537 1 7038
2 81538 1 7038
2 81539 1 7046
2 81540 1 7046
2 81541 1 7047
2 81542 1 7047
2 81543 1 7048
2 81544 1 7048
2 81545 1 7059
2 81546 1 7059
2 81547 1 7059
2 81548 1 7067
2 81549 1 7067
2 81550 1 7067
2 81551 1 7067
2 81552 1 7067
2 81553 1 7067
2 81554 1 7067
2 81555 1 7067
2 81556 1 7067
2 81557 1 7067
2 81558 1 7067
2 81559 1 7067
2 81560 1 7067
2 81561 1 7067
2 81562 1 7076
2 81563 1 7076
2 81564 1 7088
2 81565 1 7088
2 81566 1 7088
2 81567 1 7088
2 81568 1 7088
2 81569 1 7088
2 81570 1 7088
2 81571 1 7089
2 81572 1 7089
2 81573 1 7090
2 81574 1 7090
2 81575 1 7095
2 81576 1 7095
2 81577 1 7097
2 81578 1 7097
2 81579 1 7098
2 81580 1 7098
2 81581 1 7098
2 81582 1 7098
2 81583 1 7098
2 81584 1 7098
2 81585 1 7098
2 81586 1 7106
2 81587 1 7106
2 81588 1 7107
2 81589 1 7107
2 81590 1 7108
2 81591 1 7108
2 81592 1 7118
2 81593 1 7118
2 81594 1 7119
2 81595 1 7119
2 81596 1 7120
2 81597 1 7120
2 81598 1 7120
2 81599 1 7120
2 81600 1 7120
2 81601 1 7120
2 81602 1 7120
2 81603 1 7120
2 81604 1 7120
2 81605 1 7120
2 81606 1 7120
2 81607 1 7122
2 81608 1 7122
2 81609 1 7123
2 81610 1 7123
2 81611 1 7123
2 81612 1 7124
2 81613 1 7124
2 81614 1 7124
2 81615 1 7124
2 81616 1 7124
2 81617 1 7124
2 81618 1 7125
2 81619 1 7125
2 81620 1 7125
2 81621 1 7125
2 81622 1 7125
2 81623 1 7126
2 81624 1 7126
2 81625 1 7128
2 81626 1 7128
2 81627 1 7128
2 81628 1 7128
2 81629 1 7133
2 81630 1 7133
2 81631 1 7133
2 81632 1 7134
2 81633 1 7134
2 81634 1 7134
2 81635 1 7134
2 81636 1 7134
2 81637 1 7134
2 81638 1 7134
2 81639 1 7134
2 81640 1 7134
2 81641 1 7136
2 81642 1 7136
2 81643 1 7138
2 81644 1 7138
2 81645 1 7145
2 81646 1 7145
2 81647 1 7148
2 81648 1 7148
2 81649 1 7155
2 81650 1 7155
2 81651 1 7156
2 81652 1 7156
2 81653 1 7156
2 81654 1 7156
2 81655 1 7156
2 81656 1 7156
2 81657 1 7156
2 81658 1 7156
2 81659 1 7156
2 81660 1 7157
2 81661 1 7157
2 81662 1 7158
2 81663 1 7158
2 81664 1 7165
2 81665 1 7165
2 81666 1 7165
2 81667 1 7165
2 81668 1 7165
2 81669 1 7165
2 81670 1 7165
2 81671 1 7165
2 81672 1 7166
2 81673 1 7166
2 81674 1 7174
2 81675 1 7174
2 81676 1 7174
2 81677 1 7175
2 81678 1 7175
2 81679 1 7191
2 81680 1 7191
2 81681 1 7195
2 81682 1 7195
2 81683 1 7197
2 81684 1 7197
2 81685 1 7198
2 81686 1 7198
2 81687 1 7211
2 81688 1 7211
2 81689 1 7211
2 81690 1 7211
2 81691 1 7211
2 81692 1 7211
2 81693 1 7219
2 81694 1 7219
2 81695 1 7219
2 81696 1 7219
2 81697 1 7219
2 81698 1 7219
2 81699 1 7219
2 81700 1 7219
2 81701 1 7219
2 81702 1 7219
2 81703 1 7220
2 81704 1 7220
2 81705 1 7220
2 81706 1 7220
2 81707 1 7220
2 81708 1 7220
2 81709 1 7221
2 81710 1 7221
2 81711 1 7221
2 81712 1 7222
2 81713 1 7222
2 81714 1 7234
2 81715 1 7234
2 81716 1 7235
2 81717 1 7235
2 81718 1 7253
2 81719 1 7253
2 81720 1 7253
2 81721 1 7253
2 81722 1 7253
2 81723 1 7254
2 81724 1 7254
2 81725 1 7254
2 81726 1 7255
2 81727 1 7255
2 81728 1 7256
2 81729 1 7256
2 81730 1 7259
2 81731 1 7259
2 81732 1 7259
2 81733 1 7262
2 81734 1 7262
2 81735 1 7266
2 81736 1 7266
2 81737 1 7273
2 81738 1 7273
2 81739 1 7273
2 81740 1 7273
2 81741 1 7273
2 81742 1 7273
2 81743 1 7274
2 81744 1 7274
2 81745 1 7274
2 81746 1 7275
2 81747 1 7275
2 81748 1 7275
2 81749 1 7290
2 81750 1 7290
2 81751 1 7290
2 81752 1 7300
2 81753 1 7300
2 81754 1 7300
2 81755 1 7300
2 81756 1 7300
2 81757 1 7300
2 81758 1 7300
2 81759 1 7301
2 81760 1 7301
2 81761 1 7311
2 81762 1 7311
2 81763 1 7311
2 81764 1 7311
2 81765 1 7311
2 81766 1 7311
2 81767 1 7311
2 81768 1 7311
2 81769 1 7311
2 81770 1 7311
2 81771 1 7312
2 81772 1 7312
2 81773 1 7313
2 81774 1 7313
2 81775 1 7319
2 81776 1 7319
2 81777 1 7320
2 81778 1 7320
2 81779 1 7320
2 81780 1 7320
2 81781 1 7321
2 81782 1 7321
2 81783 1 7321
2 81784 1 7322
2 81785 1 7322
2 81786 1 7340
2 81787 1 7340
2 81788 1 7340
2 81789 1 7342
2 81790 1 7342
2 81791 1 7343
2 81792 1 7343
2 81793 1 7343
2 81794 1 7343
2 81795 1 7363
2 81796 1 7363
2 81797 1 7363
2 81798 1 7364
2 81799 1 7364
2 81800 1 7364
2 81801 1 7364
2 81802 1 7364
2 81803 1 7364
2 81804 1 7364
2 81805 1 7368
2 81806 1 7368
2 81807 1 7368
2 81808 1 7369
2 81809 1 7369
2 81810 1 7369
2 81811 1 7369
2 81812 1 7388
2 81813 1 7388
2 81814 1 7390
2 81815 1 7390
2 81816 1 7391
2 81817 1 7391
2 81818 1 7391
2 81819 1 7392
2 81820 1 7392
2 81821 1 7393
2 81822 1 7393
2 81823 1 7395
2 81824 1 7395
2 81825 1 7405
2 81826 1 7405
2 81827 1 7405
2 81828 1 7406
2 81829 1 7406
2 81830 1 7413
2 81831 1 7413
2 81832 1 7417
2 81833 1 7417
2 81834 1 7417
2 81835 1 7417
2 81836 1 7417
2 81837 1 7417
2 81838 1 7417
2 81839 1 7417
2 81840 1 7417
2 81841 1 7418
2 81842 1 7418
2 81843 1 7418
2 81844 1 7418
2 81845 1 7418
2 81846 1 7418
2 81847 1 7418
2 81848 1 7427
2 81849 1 7427
2 81850 1 7427
2 81851 1 7427
2 81852 1 7429
2 81853 1 7429
2 81854 1 7429
2 81855 1 7430
2 81856 1 7430
2 81857 1 7430
2 81858 1 7430
2 81859 1 7430
2 81860 1 7430
2 81861 1 7432
2 81862 1 7432
2 81863 1 7434
2 81864 1 7434
2 81865 1 7436
2 81866 1 7436
2 81867 1 7446
2 81868 1 7446
2 81869 1 7446
2 81870 1 7446
2 81871 1 7446
2 81872 1 7446
2 81873 1 7446
2 81874 1 7446
2 81875 1 7446
2 81876 1 7446
2 81877 1 7446
2 81878 1 7448
2 81879 1 7448
2 81880 1 7448
2 81881 1 7448
2 81882 1 7448
2 81883 1 7448
2 81884 1 7448
2 81885 1 7449
2 81886 1 7449
2 81887 1 7449
2 81888 1 7449
2 81889 1 7449
2 81890 1 7449
2 81891 1 7449
2 81892 1 7451
2 81893 1 7451
2 81894 1 7451
2 81895 1 7451
2 81896 1 7451
2 81897 1 7451
2 81898 1 7451
2 81899 1 7452
2 81900 1 7452
2 81901 1 7452
2 81902 1 7452
2 81903 1 7455
2 81904 1 7455
2 81905 1 7456
2 81906 1 7456
2 81907 1 7458
2 81908 1 7458
2 81909 1 7458
2 81910 1 7458
2 81911 1 7460
2 81912 1 7460
2 81913 1 7460
2 81914 1 7460
2 81915 1 7460
2 81916 1 7460
2 81917 1 7460
2 81918 1 7460
2 81919 1 7461
2 81920 1 7461
2 81921 1 7461
2 81922 1 7461
2 81923 1 7461
2 81924 1 7463
2 81925 1 7463
2 81926 1 7463
2 81927 1 7472
2 81928 1 7472
2 81929 1 7475
2 81930 1 7475
2 81931 1 7475
2 81932 1 7490
2 81933 1 7490
2 81934 1 7490
2 81935 1 7490
2 81936 1 7490
2 81937 1 7491
2 81938 1 7491
2 81939 1 7491
2 81940 1 7491
2 81941 1 7492
2 81942 1 7492
2 81943 1 7498
2 81944 1 7498
2 81945 1 7502
2 81946 1 7502
2 81947 1 7502
2 81948 1 7505
2 81949 1 7505
2 81950 1 7505
2 81951 1 7505
2 81952 1 7505
2 81953 1 7505
2 81954 1 7505
2 81955 1 7506
2 81956 1 7506
2 81957 1 7506
2 81958 1 7506
2 81959 1 7506
2 81960 1 7506
2 81961 1 7506
2 81962 1 7506
2 81963 1 7506
2 81964 1 7506
2 81965 1 7506
2 81966 1 7516
2 81967 1 7516
2 81968 1 7525
2 81969 1 7525
2 81970 1 7525
2 81971 1 7525
2 81972 1 7536
2 81973 1 7536
2 81974 1 7536
2 81975 1 7538
2 81976 1 7538
2 81977 1 7538
2 81978 1 7539
2 81979 1 7539
2 81980 1 7539
2 81981 1 7541
2 81982 1 7541
2 81983 1 7541
2 81984 1 7541
2 81985 1 7541
2 81986 1 7541
2 81987 1 7550
2 81988 1 7550
2 81989 1 7551
2 81990 1 7551
2 81991 1 7551
2 81992 1 7568
2 81993 1 7568
2 81994 1 7569
2 81995 1 7569
2 81996 1 7601
2 81997 1 7601
2 81998 1 7601
2 81999 1 7601
2 82000 1 7601
2 82001 1 7601
2 82002 1 7601
2 82003 1 7601
2 82004 1 7601
2 82005 1 7601
2 82006 1 7602
2 82007 1 7602
2 82008 1 7602
2 82009 1 7602
2 82010 1 7603
2 82011 1 7603
2 82012 1 7603
2 82013 1 7603
2 82014 1 7603
2 82015 1 7603
2 82016 1 7603
2 82017 1 7603
2 82018 1 7603
2 82019 1 7603
2 82020 1 7603
2 82021 1 7603
2 82022 1 7603
2 82023 1 7603
2 82024 1 7603
2 82025 1 7603
2 82026 1 7603
2 82027 1 7603
2 82028 1 7603
2 82029 1 7605
2 82030 1 7605
2 82031 1 7605
2 82032 1 7606
2 82033 1 7606
2 82034 1 7614
2 82035 1 7614
2 82036 1 7614
2 82037 1 7614
2 82038 1 7614
2 82039 1 7615
2 82040 1 7615
2 82041 1 7616
2 82042 1 7616
2 82043 1 7618
2 82044 1 7618
2 82045 1 7622
2 82046 1 7622
2 82047 1 7623
2 82048 1 7623
2 82049 1 7628
2 82050 1 7628
2 82051 1 7628
2 82052 1 7629
2 82053 1 7629
2 82054 1 7630
2 82055 1 7630
2 82056 1 7630
2 82057 1 7633
2 82058 1 7633
2 82059 1 7633
2 82060 1 7645
2 82061 1 7645
2 82062 1 7646
2 82063 1 7646
2 82064 1 7646
2 82065 1 7646
2 82066 1 7646
2 82067 1 7646
2 82068 1 7646
2 82069 1 7646
2 82070 1 7646
2 82071 1 7656
2 82072 1 7656
2 82073 1 7656
2 82074 1 7661
2 82075 1 7661
2 82076 1 7696
2 82077 1 7696
2 82078 1 7696
2 82079 1 7706
2 82080 1 7706
2 82081 1 7706
2 82082 1 7710
2 82083 1 7710
2 82084 1 7712
2 82085 1 7712
2 82086 1 7712
2 82087 1 7712
2 82088 1 7715
2 82089 1 7715
2 82090 1 7716
2 82091 1 7716
2 82092 1 7716
2 82093 1 7716
2 82094 1 7716
2 82095 1 7716
2 82096 1 7716
2 82097 1 7716
2 82098 1 7716
2 82099 1 7716
2 82100 1 7716
2 82101 1 7716
2 82102 1 7716
2 82103 1 7716
2 82104 1 7716
2 82105 1 7716
2 82106 1 7716
2 82107 1 7716
2 82108 1 7716
2 82109 1 7716
2 82110 1 7716
2 82111 1 7716
2 82112 1 7716
2 82113 1 7716
2 82114 1 7716
2 82115 1 7717
2 82116 1 7717
2 82117 1 7717
2 82118 1 7717
2 82119 1 7717
2 82120 1 7717
2 82121 1 7725
2 82122 1 7725
2 82123 1 7725
2 82124 1 7725
2 82125 1 7726
2 82126 1 7726
2 82127 1 7726
2 82128 1 7726
2 82129 1 7726
2 82130 1 7726
2 82131 1 7729
2 82132 1 7729
2 82133 1 7733
2 82134 1 7733
2 82135 1 7733
2 82136 1 7734
2 82137 1 7734
2 82138 1 7735
2 82139 1 7735
2 82140 1 7735
2 82141 1 7744
2 82142 1 7744
2 82143 1 7745
2 82144 1 7745
2 82145 1 7746
2 82146 1 7746
2 82147 1 7748
2 82148 1 7748
2 82149 1 7749
2 82150 1 7749
2 82151 1 7756
2 82152 1 7756
2 82153 1 7756
2 82154 1 7756
2 82155 1 7756
2 82156 1 7756
2 82157 1 7756
2 82158 1 7756
2 82159 1 7756
2 82160 1 7756
2 82161 1 7757
2 82162 1 7757
2 82163 1 7758
2 82164 1 7758
2 82165 1 7768
2 82166 1 7768
2 82167 1 7773
2 82168 1 7773
2 82169 1 7773
2 82170 1 7774
2 82171 1 7774
2 82172 1 7774
2 82173 1 7796
2 82174 1 7796
2 82175 1 7797
2 82176 1 7797
2 82177 1 7817
2 82178 1 7817
2 82179 1 7817
2 82180 1 7826
2 82181 1 7826
2 82182 1 7826
2 82183 1 7826
2 82184 1 7826
2 82185 1 7826
2 82186 1 7826
2 82187 1 7834
2 82188 1 7834
2 82189 1 7834
2 82190 1 7834
2 82191 1 7848
2 82192 1 7848
2 82193 1 7848
2 82194 1 7848
2 82195 1 7848
2 82196 1 7848
2 82197 1 7848
2 82198 1 7848
2 82199 1 7848
2 82200 1 7848
2 82201 1 7848
2 82202 1 7848
2 82203 1 7848
2 82204 1 7848
2 82205 1 7848
2 82206 1 7848
2 82207 1 7848
2 82208 1 7848
2 82209 1 7848
2 82210 1 7848
2 82211 1 7848
2 82212 1 7848
2 82213 1 7848
2 82214 1 7848
2 82215 1 7848
2 82216 1 7848
2 82217 1 7848
2 82218 1 7848
2 82219 1 7848
2 82220 1 7849
2 82221 1 7849
2 82222 1 7849
2 82223 1 7849
2 82224 1 7849
2 82225 1 7850
2 82226 1 7850
2 82227 1 7851
2 82228 1 7851
2 82229 1 7854
2 82230 1 7854
2 82231 1 7854
2 82232 1 7867
2 82233 1 7867
2 82234 1 7868
2 82235 1 7868
2 82236 1 7868
2 82237 1 7868
2 82238 1 7868
2 82239 1 7868
2 82240 1 7868
2 82241 1 7868
2 82242 1 7868
2 82243 1 7873
2 82244 1 7873
2 82245 1 7874
2 82246 1 7874
2 82247 1 7874
2 82248 1 7874
2 82249 1 7874
2 82250 1 7874
2 82251 1 7879
2 82252 1 7879
2 82253 1 7879
2 82254 1 7890
2 82255 1 7890
2 82256 1 7891
2 82257 1 7891
2 82258 1 7904
2 82259 1 7904
2 82260 1 7904
2 82261 1 7904
2 82262 1 7908
2 82263 1 7908
2 82264 1 7923
2 82265 1 7923
2 82266 1 7930
2 82267 1 7930
2 82268 1 7939
2 82269 1 7939
2 82270 1 7939
2 82271 1 7939
2 82272 1 7939
2 82273 1 7939
2 82274 1 7939
2 82275 1 7939
2 82276 1 7940
2 82277 1 7940
2 82278 1 7940
2 82279 1 7948
2 82280 1 7948
2 82281 1 7948
2 82282 1 7975
2 82283 1 7975
2 82284 1 7976
2 82285 1 7976
2 82286 1 7988
2 82287 1 7988
2 82288 1 7988
2 82289 1 7988
2 82290 1 8012
2 82291 1 8012
2 82292 1 8012
2 82293 1 8012
2 82294 1 8013
2 82295 1 8013
2 82296 1 8016
2 82297 1 8016
2 82298 1 8017
2 82299 1 8017
2 82300 1 8020
2 82301 1 8020
2 82302 1 8032
2 82303 1 8032
2 82304 1 8032
2 82305 1 8033
2 82306 1 8033
2 82307 1 8036
2 82308 1 8036
2 82309 1 8036
2 82310 1 8036
2 82311 1 8037
2 82312 1 8037
2 82313 1 8037
2 82314 1 8047
2 82315 1 8047
2 82316 1 8047
2 82317 1 8072
2 82318 1 8072
2 82319 1 8072
2 82320 1 8072
2 82321 1 8073
2 82322 1 8073
2 82323 1 8084
2 82324 1 8084
2 82325 1 8093
2 82326 1 8093
2 82327 1 8093
2 82328 1 8095
2 82329 1 8095
2 82330 1 8096
2 82331 1 8096
2 82332 1 8096
2 82333 1 8096
2 82334 1 8096
2 82335 1 8098
2 82336 1 8098
2 82337 1 8098
2 82338 1 8099
2 82339 1 8099
2 82340 1 8102
2 82341 1 8102
2 82342 1 8102
2 82343 1 8102
2 82344 1 8115
2 82345 1 8115
2 82346 1 8126
2 82347 1 8126
2 82348 1 8127
2 82349 1 8127
2 82350 1 8138
2 82351 1 8138
2 82352 1 8138
2 82353 1 8138
2 82354 1 8139
2 82355 1 8139
2 82356 1 8139
2 82357 1 8189
2 82358 1 8189
2 82359 1 8190
2 82360 1 8190
2 82361 1 8191
2 82362 1 8191
2 82363 1 8191
2 82364 1 8191
2 82365 1 8191
2 82366 1 8191
2 82367 1 8191
2 82368 1 8191
2 82369 1 8206
2 82370 1 8206
2 82371 1 8207
2 82372 1 8207
2 82373 1 8208
2 82374 1 8208
2 82375 1 8208
2 82376 1 8208
2 82377 1 8208
2 82378 1 8208
2 82379 1 8208
2 82380 1 8208
2 82381 1 8208
2 82382 1 8208
2 82383 1 8208
2 82384 1 8208
2 82385 1 8208
2 82386 1 8208
2 82387 1 8208
2 82388 1 8208
2 82389 1 8208
2 82390 1 8209
2 82391 1 8209
2 82392 1 8209
2 82393 1 8209
2 82394 1 8210
2 82395 1 8210
2 82396 1 8210
2 82397 1 8210
2 82398 1 8211
2 82399 1 8211
2 82400 1 8211
2 82401 1 8225
2 82402 1 8225
2 82403 1 8225
2 82404 1 8225
2 82405 1 8225
2 82406 1 8225
2 82407 1 8225
2 82408 1 8225
2 82409 1 8225
2 82410 1 8225
2 82411 1 8225
2 82412 1 8225
2 82413 1 8225
2 82414 1 8225
2 82415 1 8225
2 82416 1 8225
2 82417 1 8225
2 82418 1 8225
2 82419 1 8225
2 82420 1 8225
2 82421 1 8225
2 82422 1 8225
2 82423 1 8225
2 82424 1 8225
2 82425 1 8225
2 82426 1 8225
2 82427 1 8225
2 82428 1 8225
2 82429 1 8225
2 82430 1 8225
2 82431 1 8225
2 82432 1 8226
2 82433 1 8226
2 82434 1 8227
2 82435 1 8227
2 82436 1 8227
2 82437 1 8227
2 82438 1 8227
2 82439 1 8228
2 82440 1 8228
2 82441 1 8228
2 82442 1 8228
2 82443 1 8228
2 82444 1 8228
2 82445 1 8228
2 82446 1 8228
2 82447 1 8228
2 82448 1 8228
2 82449 1 8229
2 82450 1 8229
2 82451 1 8229
2 82452 1 8229
2 82453 1 8236
2 82454 1 8236
2 82455 1 8244
2 82456 1 8244
2 82457 1 8273
2 82458 1 8273
2 82459 1 8273
2 82460 1 8281
2 82461 1 8281
2 82462 1 8282
2 82463 1 8282
2 82464 1 8283
2 82465 1 8283
2 82466 1 8284
2 82467 1 8284
2 82468 1 8284
2 82469 1 8284
2 82470 1 8285
2 82471 1 8285
2 82472 1 8285
2 82473 1 8285
2 82474 1 8285
2 82475 1 8285
2 82476 1 8285
2 82477 1 8295
2 82478 1 8295
2 82479 1 8303
2 82480 1 8303
2 82481 1 8309
2 82482 1 8309
2 82483 1 8310
2 82484 1 8310
2 82485 1 8310
2 82486 1 8313
2 82487 1 8313
2 82488 1 8317
2 82489 1 8317
2 82490 1 8317
2 82491 1 8317
2 82492 1 8335
2 82493 1 8335
2 82494 1 8335
2 82495 1 8339
2 82496 1 8339
2 82497 1 8342
2 82498 1 8342
2 82499 1 8342
2 82500 1 8342
2 82501 1 8351
2 82502 1 8351
2 82503 1 8352
2 82504 1 8352
2 82505 1 8352
2 82506 1 8353
2 82507 1 8353
2 82508 1 8353
2 82509 1 8353
2 82510 1 8358
2 82511 1 8358
2 82512 1 8374
2 82513 1 8374
2 82514 1 8374
2 82515 1 8382
2 82516 1 8382
2 82517 1 8382
2 82518 1 8382
2 82519 1 8402
2 82520 1 8402
2 82521 1 8402
2 82522 1 8402
2 82523 1 8404
2 82524 1 8404
2 82525 1 8404
2 82526 1 8404
2 82527 1 8404
2 82528 1 8404
2 82529 1 8404
2 82530 1 8404
2 82531 1 8404
2 82532 1 8404
2 82533 1 8404
2 82534 1 8404
2 82535 1 8404
2 82536 1 8404
2 82537 1 8405
2 82538 1 8405
2 82539 1 8405
2 82540 1 8405
2 82541 1 8406
2 82542 1 8406
2 82543 1 8406
2 82544 1 8406
2 82545 1 8414
2 82546 1 8414
2 82547 1 8415
2 82548 1 8415
2 82549 1 8415
2 82550 1 8415
2 82551 1 8415
2 82552 1 8415
2 82553 1 8415
2 82554 1 8415
2 82555 1 8415
2 82556 1 8415
2 82557 1 8415
2 82558 1 8415
2 82559 1 8415
2 82560 1 8415
2 82561 1 8415
2 82562 1 8415
2 82563 1 8415
2 82564 1 8415
2 82565 1 8415
2 82566 1 8415
2 82567 1 8415
2 82568 1 8415
2 82569 1 8415
2 82570 1 8415
2 82571 1 8415
2 82572 1 8415
2 82573 1 8415
2 82574 1 8415
2 82575 1 8415
2 82576 1 8415
2 82577 1 8415
2 82578 1 8415
2 82579 1 8415
2 82580 1 8415
2 82581 1 8415
2 82582 1 8415
2 82583 1 8415
2 82584 1 8415
2 82585 1 8415
2 82586 1 8415
2 82587 1 8415
2 82588 1 8415
2 82589 1 8416
2 82590 1 8416
2 82591 1 8416
2 82592 1 8416
2 82593 1 8416
2 82594 1 8416
2 82595 1 8416
2 82596 1 8416
2 82597 1 8416
2 82598 1 8416
2 82599 1 8416
2 82600 1 8416
2 82601 1 8417
2 82602 1 8417
2 82603 1 8418
2 82604 1 8418
2 82605 1 8420
2 82606 1 8420
2 82607 1 8420
2 82608 1 8420
2 82609 1 8420
2 82610 1 8423
2 82611 1 8423
2 82612 1 8423
2 82613 1 8425
2 82614 1 8425
2 82615 1 8451
2 82616 1 8451
2 82617 1 8451
2 82618 1 8451
2 82619 1 8451
2 82620 1 8451
2 82621 1 8451
2 82622 1 8454
2 82623 1 8454
2 82624 1 8454
2 82625 1 8454
2 82626 1 8462
2 82627 1 8462
2 82628 1 8464
2 82629 1 8464
2 82630 1 8464
2 82631 1 8464
2 82632 1 8464
2 82633 1 8464
2 82634 1 8464
2 82635 1 8464
2 82636 1 8483
2 82637 1 8483
2 82638 1 8483
2 82639 1 8483
2 82640 1 8483
2 82641 1 8483
2 82642 1 8483
2 82643 1 8483
2 82644 1 8483
2 82645 1 8483
2 82646 1 8483
2 82647 1 8483
2 82648 1 8489
2 82649 1 8489
2 82650 1 8489
2 82651 1 8489
2 82652 1 8489
2 82653 1 8489
2 82654 1 8489
2 82655 1 8489
2 82656 1 8489
2 82657 1 8489
2 82658 1 8489
2 82659 1 8489
2 82660 1 8489
2 82661 1 8489
2 82662 1 8489
2 82663 1 8489
2 82664 1 8489
2 82665 1 8489
2 82666 1 8489
2 82667 1 8491
2 82668 1 8491
2 82669 1 8496
2 82670 1 8496
2 82671 1 8501
2 82672 1 8501
2 82673 1 8506
2 82674 1 8506
2 82675 1 8506
2 82676 1 8506
2 82677 1 8506
2 82678 1 8506
2 82679 1 8506
2 82680 1 8506
2 82681 1 8506
2 82682 1 8506
2 82683 1 8506
2 82684 1 8506
2 82685 1 8506
2 82686 1 8506
2 82687 1 8506
2 82688 1 8506
2 82689 1 8506
2 82690 1 8506
2 82691 1 8514
2 82692 1 8514
2 82693 1 8514
2 82694 1 8515
2 82695 1 8515
2 82696 1 8516
2 82697 1 8516
2 82698 1 8524
2 82699 1 8524
2 82700 1 8539
2 82701 1 8539
2 82702 1 8540
2 82703 1 8540
2 82704 1 8541
2 82705 1 8541
2 82706 1 8541
2 82707 1 8542
2 82708 1 8542
2 82709 1 8548
2 82710 1 8548
2 82711 1 8548
2 82712 1 8548
2 82713 1 8548
2 82714 1 8548
2 82715 1 8548
2 82716 1 8548
2 82717 1 8549
2 82718 1 8549
2 82719 1 8549
2 82720 1 8549
2 82721 1 8549
2 82722 1 8550
2 82723 1 8550
2 82724 1 8577
2 82725 1 8577
2 82726 1 8581
2 82727 1 8581
2 82728 1 8589
2 82729 1 8589
2 82730 1 8590
2 82731 1 8590
2 82732 1 8598
2 82733 1 8598
2 82734 1 8600
2 82735 1 8600
2 82736 1 8602
2 82737 1 8602
2 82738 1 8606
2 82739 1 8606
2 82740 1 8609
2 82741 1 8609
2 82742 1 8609
2 82743 1 8609
2 82744 1 8610
2 82745 1 8610
2 82746 1 8610
2 82747 1 8625
2 82748 1 8625
2 82749 1 8625
2 82750 1 8633
2 82751 1 8633
2 82752 1 8633
2 82753 1 8634
2 82754 1 8634
2 82755 1 8642
2 82756 1 8642
2 82757 1 8658
2 82758 1 8658
2 82759 1 8688
2 82760 1 8688
2 82761 1 8689
2 82762 1 8689
2 82763 1 8692
2 82764 1 8692
2 82765 1 8693
2 82766 1 8693
2 82767 1 8694
2 82768 1 8694
2 82769 1 8703
2 82770 1 8703
2 82771 1 8703
2 82772 1 8718
2 82773 1 8718
2 82774 1 8722
2 82775 1 8722
2 82776 1 8729
2 82777 1 8729
2 82778 1 8742
2 82779 1 8742
2 82780 1 8742
2 82781 1 8743
2 82782 1 8743
2 82783 1 8743
2 82784 1 8743
2 82785 1 8743
2 82786 1 8743
2 82787 1 8743
2 82788 1 8743
2 82789 1 8743
2 82790 1 8744
2 82791 1 8744
2 82792 1 8754
2 82793 1 8754
2 82794 1 8754
2 82795 1 8764
2 82796 1 8764
2 82797 1 8764
2 82798 1 8764
2 82799 1 8764
2 82800 1 8764
2 82801 1 8764
2 82802 1 8764
2 82803 1 8764
2 82804 1 8764
2 82805 1 8764
2 82806 1 8764
2 82807 1 8764
2 82808 1 8764
2 82809 1 8764
2 82810 1 8764
2 82811 1 8764
2 82812 1 8765
2 82813 1 8765
2 82814 1 8775
2 82815 1 8775
2 82816 1 8788
2 82817 1 8788
2 82818 1 8789
2 82819 1 8789
2 82820 1 8796
2 82821 1 8796
2 82822 1 8797
2 82823 1 8797
2 82824 1 8800
2 82825 1 8800
2 82826 1 8806
2 82827 1 8806
2 82828 1 8806
2 82829 1 8818
2 82830 1 8818
2 82831 1 8829
2 82832 1 8829
2 82833 1 8840
2 82834 1 8840
2 82835 1 8840
2 82836 1 8840
2 82837 1 8843
2 82838 1 8843
2 82839 1 8844
2 82840 1 8844
2 82841 1 8844
2 82842 1 8845
2 82843 1 8845
2 82844 1 8845
2 82845 1 8845
2 82846 1 8845
2 82847 1 8845
2 82848 1 8845
2 82849 1 8846
2 82850 1 8846
2 82851 1 8846
2 82852 1 8846
2 82853 1 8846
2 82854 1 8847
2 82855 1 8847
2 82856 1 8847
2 82857 1 8847
2 82858 1 8847
2 82859 1 8847
2 82860 1 8848
2 82861 1 8848
2 82862 1 8861
2 82863 1 8861
2 82864 1 8861
2 82865 1 8864
2 82866 1 8864
2 82867 1 8864
2 82868 1 8864
2 82869 1 8864
2 82870 1 8864
2 82871 1 8864
2 82872 1 8864
2 82873 1 8864
2 82874 1 8864
2 82875 1 8864
2 82876 1 8864
2 82877 1 8864
2 82878 1 8864
2 82879 1 8864
2 82880 1 8864
2 82881 1 8864
2 82882 1 8864
2 82883 1 8864
2 82884 1 8864
2 82885 1 8864
2 82886 1 8864
2 82887 1 8865
2 82888 1 8865
2 82889 1 8865
2 82890 1 8866
2 82891 1 8866
2 82892 1 8867
2 82893 1 8867
2 82894 1 8867
2 82895 1 8867
2 82896 1 8868
2 82897 1 8868
2 82898 1 8869
2 82899 1 8869
2 82900 1 8874
2 82901 1 8874
2 82902 1 8883
2 82903 1 8883
2 82904 1 8883
2 82905 1 8884
2 82906 1 8884
2 82907 1 8884
2 82908 1 8884
2 82909 1 8884
2 82910 1 8884
2 82911 1 8884
2 82912 1 8886
2 82913 1 8886
2 82914 1 8886
2 82915 1 8886
2 82916 1 8886
2 82917 1 8889
2 82918 1 8889
2 82919 1 8889
2 82920 1 8889
2 82921 1 8889
2 82922 1 8889
2 82923 1 8889
2 82924 1 8889
2 82925 1 8889
2 82926 1 8889
2 82927 1 8889
2 82928 1 8889
2 82929 1 8889
2 82930 1 8889
2 82931 1 8889
2 82932 1 8889
2 82933 1 8889
2 82934 1 8890
2 82935 1 8890
2 82936 1 8890
2 82937 1 8890
2 82938 1 8890
2 82939 1 8890
2 82940 1 8890
2 82941 1 8890
2 82942 1 8890
2 82943 1 8890
2 82944 1 8890
2 82945 1 8890
2 82946 1 8890
2 82947 1 8890
2 82948 1 8890
2 82949 1 8890
2 82950 1 8890
2 82951 1 8890
2 82952 1 8890
2 82953 1 8890
2 82954 1 8890
2 82955 1 8890
2 82956 1 8890
2 82957 1 8890
2 82958 1 8890
2 82959 1 8890
2 82960 1 8890
2 82961 1 8890
2 82962 1 8890
2 82963 1 8890
2 82964 1 8890
2 82965 1 8890
2 82966 1 8890
2 82967 1 8890
2 82968 1 8890
2 82969 1 8890
2 82970 1 8890
2 82971 1 8890
2 82972 1 8890
2 82973 1 8890
2 82974 1 8890
2 82975 1 8890
2 82976 1 8890
2 82977 1 8890
2 82978 1 8890
2 82979 1 8890
2 82980 1 8890
2 82981 1 8890
2 82982 1 8890
2 82983 1 8890
2 82984 1 8890
2 82985 1 8890
2 82986 1 8890
2 82987 1 8890
2 82988 1 8891
2 82989 1 8891
2 82990 1 8899
2 82991 1 8899
2 82992 1 8899
2 82993 1 8899
2 82994 1 8900
2 82995 1 8900
2 82996 1 8901
2 82997 1 8901
2 82998 1 8901
2 82999 1 8901
2 83000 1 8901
2 83001 1 8901
2 83002 1 8901
2 83003 1 8901
2 83004 1 8913
2 83005 1 8913
2 83006 1 8913
2 83007 1 8913
2 83008 1 8913
2 83009 1 8914
2 83010 1 8914
2 83011 1 8933
2 83012 1 8933
2 83013 1 8933
2 83014 1 8933
2 83015 1 8933
2 83016 1 8939
2 83017 1 8939
2 83018 1 8939
2 83019 1 8939
2 83020 1 8939
2 83021 1 8939
2 83022 1 8939
2 83023 1 8939
2 83024 1 8939
2 83025 1 8939
2 83026 1 8939
2 83027 1 8939
2 83028 1 8940
2 83029 1 8940
2 83030 1 8940
2 83031 1 8940
2 83032 1 8954
2 83033 1 8954
2 83034 1 8978
2 83035 1 8978
2 83036 1 8978
2 83037 1 8978
2 83038 1 8978
2 83039 1 8988
2 83040 1 8988
2 83041 1 8989
2 83042 1 8989
2 83043 1 8989
2 83044 1 9013
2 83045 1 9013
2 83046 1 9015
2 83047 1 9015
2 83048 1 9015
2 83049 1 9015
2 83050 1 9015
2 83051 1 9015
2 83052 1 9023
2 83053 1 9023
2 83054 1 9038
2 83055 1 9038
2 83056 1 9038
2 83057 1 9062
2 83058 1 9062
2 83059 1 9062
2 83060 1 9062
2 83061 1 9062
2 83062 1 9062
2 83063 1 9062
2 83064 1 9062
2 83065 1 9064
2 83066 1 9064
2 83067 1 9064
2 83068 1 9071
2 83069 1 9071
2 83070 1 9079
2 83071 1 9079
2 83072 1 9084
2 83073 1 9084
2 83074 1 9084
2 83075 1 9084
2 83076 1 9084
2 83077 1 9084
2 83078 1 9085
2 83079 1 9085
2 83080 1 9085
2 83081 1 9085
2 83082 1 9085
2 83083 1 9085
2 83084 1 9085
2 83085 1 9085
2 83086 1 9085
2 83087 1 9086
2 83088 1 9086
2 83089 1 9087
2 83090 1 9087
2 83091 1 9095
2 83092 1 9095
2 83093 1 9097
2 83094 1 9097
2 83095 1 9113
2 83096 1 9113
2 83097 1 9113
2 83098 1 9123
2 83099 1 9123
2 83100 1 9123
2 83101 1 9124
2 83102 1 9124
2 83103 1 9125
2 83104 1 9125
2 83105 1 9131
2 83106 1 9131
2 83107 1 9132
2 83108 1 9132
2 83109 1 9162
2 83110 1 9162
2 83111 1 9173
2 83112 1 9173
2 83113 1 9182
2 83114 1 9182
2 83115 1 9200
2 83116 1 9200
2 83117 1 9219
2 83118 1 9219
2 83119 1 9220
2 83120 1 9220
2 83121 1 9227
2 83122 1 9227
2 83123 1 9227
2 83124 1 9227
2 83125 1 9227
2 83126 1 9229
2 83127 1 9229
2 83128 1 9229
2 83129 1 9231
2 83130 1 9231
2 83131 1 9246
2 83132 1 9246
2 83133 1 9248
2 83134 1 9248
2 83135 1 9248
2 83136 1 9248
2 83137 1 9248
2 83138 1 9248
2 83139 1 9249
2 83140 1 9249
2 83141 1 9249
2 83142 1 9249
2 83143 1 9249
2 83144 1 9249
2 83145 1 9252
2 83146 1 9252
2 83147 1 9252
2 83148 1 9264
2 83149 1 9264
2 83150 1 9308
2 83151 1 9308
2 83152 1 9308
2 83153 1 9308
2 83154 1 9326
2 83155 1 9326
2 83156 1 9331
2 83157 1 9331
2 83158 1 9331
2 83159 1 9331
2 83160 1 9331
2 83161 1 9331
2 83162 1 9331
2 83163 1 9331
2 83164 1 9331
2 83165 1 9331
2 83166 1 9331
2 83167 1 9331
2 83168 1 9331
2 83169 1 9331
2 83170 1 9331
2 83171 1 9331
2 83172 1 9331
2 83173 1 9331
2 83174 1 9331
2 83175 1 9331
2 83176 1 9332
2 83177 1 9332
2 83178 1 9333
2 83179 1 9333
2 83180 1 9333
2 83181 1 9341
2 83182 1 9341
2 83183 1 9341
2 83184 1 9341
2 83185 1 9341
2 83186 1 9342
2 83187 1 9342
2 83188 1 9342
2 83189 1 9345
2 83190 1 9345
2 83191 1 9348
2 83192 1 9348
2 83193 1 9357
2 83194 1 9357
2 83195 1 9358
2 83196 1 9358
2 83197 1 9359
2 83198 1 9359
2 83199 1 9359
2 83200 1 9363
2 83201 1 9363
2 83202 1 9363
2 83203 1 9369
2 83204 1 9369
2 83205 1 9375
2 83206 1 9375
2 83207 1 9376
2 83208 1 9376
2 83209 1 9377
2 83210 1 9377
2 83211 1 9380
2 83212 1 9380
2 83213 1 9387
2 83214 1 9387
2 83215 1 9390
2 83216 1 9390
2 83217 1 9400
2 83218 1 9400
2 83219 1 9400
2 83220 1 9400
2 83221 1 9400
2 83222 1 9400
2 83223 1 9402
2 83224 1 9402
2 83225 1 9403
2 83226 1 9403
2 83227 1 9404
2 83228 1 9404
2 83229 1 9408
2 83230 1 9408
2 83231 1 9409
2 83232 1 9409
2 83233 1 9409
2 83234 1 9409
2 83235 1 9411
2 83236 1 9411
2 83237 1 9411
2 83238 1 9413
2 83239 1 9413
2 83240 1 9413
2 83241 1 9414
2 83242 1 9414
2 83243 1 9421
2 83244 1 9421
2 83245 1 9421
2 83246 1 9421
2 83247 1 9422
2 83248 1 9422
2 83249 1 9422
2 83250 1 9422
2 83251 1 9422
2 83252 1 9422
2 83253 1 9422
2 83254 1 9422
2 83255 1 9422
2 83256 1 9422
2 83257 1 9422
2 83258 1 9422
2 83259 1 9422
2 83260 1 9422
2 83261 1 9425
2 83262 1 9425
2 83263 1 9425
2 83264 1 9427
2 83265 1 9427
2 83266 1 9427
2 83267 1 9428
2 83268 1 9428
2 83269 1 9428
2 83270 1 9428
2 83271 1 9428
2 83272 1 9430
2 83273 1 9430
2 83274 1 9430
2 83275 1 9431
2 83276 1 9431
2 83277 1 9432
2 83278 1 9432
2 83279 1 9453
2 83280 1 9453
2 83281 1 9453
2 83282 1 9453
2 83283 1 9454
2 83284 1 9454
2 83285 1 9458
2 83286 1 9458
2 83287 1 9458
2 83288 1 9466
2 83289 1 9466
2 83290 1 9466
2 83291 1 9466
2 83292 1 9467
2 83293 1 9467
2 83294 1 9468
2 83295 1 9468
2 83296 1 9469
2 83297 1 9469
2 83298 1 9472
2 83299 1 9472
2 83300 1 9473
2 83301 1 9473
2 83302 1 9473
2 83303 1 9473
2 83304 1 9473
2 83305 1 9473
2 83306 1 9494
2 83307 1 9494
2 83308 1 9495
2 83309 1 9495
2 83310 1 9495
2 83311 1 9495
2 83312 1 9495
2 83313 1 9503
2 83314 1 9503
2 83315 1 9503
2 83316 1 9504
2 83317 1 9504
2 83318 1 9505
2 83319 1 9505
2 83320 1 9526
2 83321 1 9526
2 83322 1 9527
2 83323 1 9527
2 83324 1 9529
2 83325 1 9529
2 83326 1 9541
2 83327 1 9541
2 83328 1 9541
2 83329 1 9541
2 83330 1 9542
2 83331 1 9542
2 83332 1 9544
2 83333 1 9544
2 83334 1 9546
2 83335 1 9546
2 83336 1 9547
2 83337 1 9547
2 83338 1 9547
2 83339 1 9550
2 83340 1 9550
2 83341 1 9551
2 83342 1 9551
2 83343 1 9552
2 83344 1 9552
2 83345 1 9552
2 83346 1 9557
2 83347 1 9557
2 83348 1 9565
2 83349 1 9565
2 83350 1 9565
2 83351 1 9565
2 83352 1 9565
2 83353 1 9566
2 83354 1 9566
2 83355 1 9566
2 83356 1 9566
2 83357 1 9566
2 83358 1 9567
2 83359 1 9567
2 83360 1 9569
2 83361 1 9569
2 83362 1 9585
2 83363 1 9585
2 83364 1 9585
2 83365 1 9585
2 83366 1 9585
2 83367 1 9585
2 83368 1 9586
2 83369 1 9586
2 83370 1 9586
2 83371 1 9594
2 83372 1 9594
2 83373 1 9595
2 83374 1 9595
2 83375 1 9595
2 83376 1 9595
2 83377 1 9595
2 83378 1 9599
2 83379 1 9599
2 83380 1 9606
2 83381 1 9606
2 83382 1 9606
2 83383 1 9606
2 83384 1 9607
2 83385 1 9607
2 83386 1 9612
2 83387 1 9612
2 83388 1 9612
2 83389 1 9631
2 83390 1 9631
2 83391 1 9632
2 83392 1 9632
2 83393 1 9632
2 83394 1 9632
2 83395 1 9632
2 83396 1 9635
2 83397 1 9635
2 83398 1 9635
2 83399 1 9636
2 83400 1 9636
2 83401 1 9658
2 83402 1 9658
2 83403 1 9658
2 83404 1 9658
2 83405 1 9658
2 83406 1 9658
2 83407 1 9658
2 83408 1 9659
2 83409 1 9659
2 83410 1 9675
2 83411 1 9675
2 83412 1 9676
2 83413 1 9676
2 83414 1 9696
2 83415 1 9696
2 83416 1 9696
2 83417 1 9696
2 83418 1 9696
2 83419 1 9696
2 83420 1 9696
2 83421 1 9707
2 83422 1 9707
2 83423 1 9707
2 83424 1 9707
2 83425 1 9707
2 83426 1 9708
2 83427 1 9708
2 83428 1 9708
2 83429 1 9716
2 83430 1 9716
2 83431 1 9717
2 83432 1 9717
2 83433 1 9717
2 83434 1 9720
2 83435 1 9720
2 83436 1 9720
2 83437 1 9721
2 83438 1 9721
2 83439 1 9722
2 83440 1 9722
2 83441 1 9722
2 83442 1 9722
2 83443 1 9722
2 83444 1 9722
2 83445 1 9722
2 83446 1 9722
2 83447 1 9723
2 83448 1 9723
2 83449 1 9724
2 83450 1 9724
2 83451 1 9734
2 83452 1 9734
2 83453 1 9734
2 83454 1 9734
2 83455 1 9734
2 83456 1 9734
2 83457 1 9734
2 83458 1 9743
2 83459 1 9743
2 83460 1 9743
2 83461 1 9743
2 83462 1 9743
2 83463 1 9743
2 83464 1 9751
2 83465 1 9751
2 83466 1 9751
2 83467 1 9751
2 83468 1 9752
2 83469 1 9752
2 83470 1 9752
2 83471 1 9752
2 83472 1 9752
2 83473 1 9752
2 83474 1 9752
2 83475 1 9753
2 83476 1 9753
2 83477 1 9757
2 83478 1 9757
2 83479 1 9775
2 83480 1 9775
2 83481 1 9775
2 83482 1 9775
2 83483 1 9775
2 83484 1 9784
2 83485 1 9784
2 83486 1 9786
2 83487 1 9786
2 83488 1 9786
2 83489 1 9788
2 83490 1 9788
2 83491 1 9788
2 83492 1 9789
2 83493 1 9789
2 83494 1 9799
2 83495 1 9799
2 83496 1 9806
2 83497 1 9806
2 83498 1 9820
2 83499 1 9820
2 83500 1 9820
2 83501 1 9820
2 83502 1 9848
2 83503 1 9848
2 83504 1 9859
2 83505 1 9859
2 83506 1 9861
2 83507 1 9861
2 83508 1 9861
2 83509 1 9861
2 83510 1 9861
2 83511 1 9862
2 83512 1 9862
2 83513 1 9875
2 83514 1 9875
2 83515 1 9876
2 83516 1 9876
2 83517 1 9876
2 83518 1 9876
2 83519 1 9876
2 83520 1 9876
2 83521 1 9902
2 83522 1 9902
2 83523 1 9923
2 83524 1 9923
2 83525 1 9932
2 83526 1 9932
2 83527 1 9945
2 83528 1 9945
2 83529 1 9964
2 83530 1 9964
2 83531 1 9964
2 83532 1 9964
2 83533 1 9990
2 83534 1 9990
2 83535 1 9990
2 83536 1 9990
2 83537 1 9990
2 83538 1 9990
2 83539 1 10000
2 83540 1 10000
2 83541 1 10003
2 83542 1 10003
2 83543 1 10015
2 83544 1 10015
2 83545 1 10044
2 83546 1 10044
2 83547 1 10075
2 83548 1 10075
2 83549 1 10085
2 83550 1 10085
2 83551 1 10085
2 83552 1 10085
2 83553 1 10085
2 83554 1 10085
2 83555 1 10085
2 83556 1 10085
2 83557 1 10087
2 83558 1 10087
2 83559 1 10087
2 83560 1 10087
2 83561 1 10087
2 83562 1 10087
2 83563 1 10088
2 83564 1 10088
2 83565 1 10106
2 83566 1 10106
2 83567 1 10114
2 83568 1 10114
2 83569 1 10134
2 83570 1 10134
2 83571 1 10134
2 83572 1 10135
2 83573 1 10135
2 83574 1 10135
2 83575 1 10135
2 83576 1 10164
2 83577 1 10164
2 83578 1 10165
2 83579 1 10165
2 83580 1 10178
2 83581 1 10178
2 83582 1 10187
2 83583 1 10187
2 83584 1 10187
2 83585 1 10187
2 83586 1 10187
2 83587 1 10187
2 83588 1 10224
2 83589 1 10224
2 83590 1 10224
2 83591 1 10225
2 83592 1 10225
2 83593 1 10240
2 83594 1 10240
2 83595 1 10254
2 83596 1 10254
2 83597 1 10254
2 83598 1 10255
2 83599 1 10255
2 83600 1 10263
2 83601 1 10263
2 83602 1 10263
2 83603 1 10263
2 83604 1 10287
2 83605 1 10287
2 83606 1 10287
2 83607 1 10288
2 83608 1 10288
2 83609 1 10328
2 83610 1 10328
2 83611 1 10328
2 83612 1 10360
2 83613 1 10360
2 83614 1 10362
2 83615 1 10362
2 83616 1 10362
2 83617 1 10362
2 83618 1 10376
2 83619 1 10376
2 83620 1 10384
2 83621 1 10384
2 83622 1 10384
2 83623 1 10384
2 83624 1 10385
2 83625 1 10385
2 83626 1 10385
2 83627 1 10386
2 83628 1 10386
2 83629 1 10415
2 83630 1 10415
2 83631 1 10419
2 83632 1 10419
2 83633 1 10438
2 83634 1 10438
2 83635 1 10438
2 83636 1 10438
2 83637 1 10438
2 83638 1 10438
2 83639 1 10438
2 83640 1 10445
2 83641 1 10445
2 83642 1 10445
2 83643 1 10445
2 83644 1 10445
2 83645 1 10445
2 83646 1 10445
2 83647 1 10446
2 83648 1 10446
2 83649 1 10457
2 83650 1 10457
2 83651 1 10457
2 83652 1 10457
2 83653 1 10458
2 83654 1 10458
2 83655 1 10458
2 83656 1 10458
2 83657 1 10458
2 83658 1 10461
2 83659 1 10461
2 83660 1 10461
2 83661 1 10461
2 83662 1 10461
2 83663 1 10461
2 83664 1 10461
2 83665 1 10461
2 83666 1 10461
2 83667 1 10461
2 83668 1 10461
2 83669 1 10461
2 83670 1 10461
2 83671 1 10463
2 83672 1 10463
2 83673 1 10492
2 83674 1 10492
2 83675 1 10492
2 83676 1 10493
2 83677 1 10493
2 83678 1 10511
2 83679 1 10511
2 83680 1 10511
2 83681 1 10511
2 83682 1 10511
2 83683 1 10511
2 83684 1 10511
2 83685 1 10512
2 83686 1 10512
2 83687 1 10512
2 83688 1 10512
2 83689 1 10513
2 83690 1 10513
2 83691 1 10521
2 83692 1 10521
2 83693 1 10527
2 83694 1 10527
2 83695 1 10565
2 83696 1 10565
2 83697 1 10565
2 83698 1 10598
2 83699 1 10598
2 83700 1 10599
2 83701 1 10599
2 83702 1 10601
2 83703 1 10601
2 83704 1 10617
2 83705 1 10617
2 83706 1 10620
2 83707 1 10620
2 83708 1 10623
2 83709 1 10623
2 83710 1 10631
2 83711 1 10631
2 83712 1 10638
2 83713 1 10638
2 83714 1 10650
2 83715 1 10650
2 83716 1 10651
2 83717 1 10651
2 83718 1 10652
2 83719 1 10652
2 83720 1 10652
2 83721 1 10661
2 83722 1 10661
2 83723 1 10661
2 83724 1 10661
2 83725 1 10662
2 83726 1 10662
2 83727 1 10662
2 83728 1 10662
2 83729 1 10679
2 83730 1 10679
2 83731 1 10690
2 83732 1 10690
2 83733 1 10691
2 83734 1 10691
2 83735 1 10692
2 83736 1 10692
2 83737 1 10697
2 83738 1 10697
2 83739 1 10698
2 83740 1 10698
2 83741 1 10700
2 83742 1 10700
2 83743 1 10735
2 83744 1 10735
2 83745 1 10736
2 83746 1 10736
2 83747 1 10736
2 83748 1 10742
2 83749 1 10742
2 83750 1 10742
2 83751 1 10744
2 83752 1 10744
2 83753 1 10745
2 83754 1 10745
2 83755 1 10750
2 83756 1 10750
2 83757 1 10753
2 83758 1 10753
2 83759 1 10755
2 83760 1 10755
2 83761 1 10770
2 83762 1 10770
2 83763 1 10770
2 83764 1 10772
2 83765 1 10772
2 83766 1 10782
2 83767 1 10782
2 83768 1 10793
2 83769 1 10793
2 83770 1 10803
2 83771 1 10803
2 83772 1 10803
2 83773 1 10807
2 83774 1 10807
2 83775 1 10807
2 83776 1 10812
2 83777 1 10812
2 83778 1 10812
2 83779 1 10812
2 83780 1 10812
2 83781 1 10812
2 83782 1 10822
2 83783 1 10822
2 83784 1 10829
2 83785 1 10829
2 83786 1 10830
2 83787 1 10830
2 83788 1 10830
2 83789 1 10833
2 83790 1 10833
2 83791 1 10834
2 83792 1 10834
2 83793 1 10834
2 83794 1 10834
2 83795 1 10835
2 83796 1 10835
2 83797 1 10837
2 83798 1 10837
2 83799 1 10843
2 83800 1 10843
2 83801 1 10848
2 83802 1 10848
2 83803 1 10854
2 83804 1 10854
2 83805 1 10854
2 83806 1 10859
2 83807 1 10859
2 83808 1 10872
2 83809 1 10872
2 83810 1 10882
2 83811 1 10882
2 83812 1 10883
2 83813 1 10883
2 83814 1 10883
2 83815 1 10883
2 83816 1 10883
2 83817 1 10883
2 83818 1 10884
2 83819 1 10884
2 83820 1 10885
2 83821 1 10885
2 83822 1 10885
2 83823 1 10886
2 83824 1 10886
2 83825 1 10912
2 83826 1 10912
2 83827 1 10912
2 83828 1 10912
2 83829 1 10912
2 83830 1 10912
2 83831 1 10951
2 83832 1 10951
2 83833 1 10951
2 83834 1 10967
2 83835 1 10967
2 83836 1 10977
2 83837 1 10977
2 83838 1 10977
2 83839 1 10977
2 83840 1 10977
2 83841 1 10978
2 83842 1 10978
2 83843 1 10986
2 83844 1 10986
2 83845 1 10986
2 83846 1 10987
2 83847 1 10987
2 83848 1 10987
2 83849 1 10995
2 83850 1 10995
2 83851 1 11004
2 83852 1 11004
2 83853 1 11016
2 83854 1 11016
2 83855 1 11016
2 83856 1 11046
2 83857 1 11046
2 83858 1 11065
2 83859 1 11065
2 83860 1 11069
2 83861 1 11069
2 83862 1 11070
2 83863 1 11070
2 83864 1 11070
2 83865 1 11075
2 83866 1 11075
2 83867 1 11075
2 83868 1 11075
2 83869 1 11077
2 83870 1 11077
2 83871 1 11077
2 83872 1 11081
2 83873 1 11081
2 83874 1 11081
2 83875 1 11081
2 83876 1 11089
2 83877 1 11089
2 83878 1 11099
2 83879 1 11099
2 83880 1 11112
2 83881 1 11112
2 83882 1 11122
2 83883 1 11122
2 83884 1 11123
2 83885 1 11123
2 83886 1 11131
2 83887 1 11131
2 83888 1 11134
2 83889 1 11134
2 83890 1 11140
2 83891 1 11140
2 83892 1 11141
2 83893 1 11141
2 83894 1 11142
2 83895 1 11142
2 83896 1 11142
2 83897 1 11143
2 83898 1 11143
2 83899 1 11170
2 83900 1 11170
2 83901 1 11206
2 83902 1 11206
2 83903 1 11206
2 83904 1 11206
2 83905 1 11206
2 83906 1 11206
2 83907 1 11207
2 83908 1 11207
2 83909 1 11207
2 83910 1 11208
2 83911 1 11208
2 83912 1 11208
2 83913 1 11208
2 83914 1 11211
2 83915 1 11211
2 83916 1 11222
2 83917 1 11222
2 83918 1 11222
2 83919 1 11222
2 83920 1 11222
2 83921 1 11231
2 83922 1 11231
2 83923 1 11231
2 83924 1 11231
2 83925 1 11231
2 83926 1 11231
2 83927 1 11232
2 83928 1 11232
2 83929 1 11248
2 83930 1 11248
2 83931 1 11248
2 83932 1 11249
2 83933 1 11249
2 83934 1 11249
2 83935 1 11249
2 83936 1 11249
2 83937 1 11250
2 83938 1 11250
2 83939 1 11251
2 83940 1 11251
2 83941 1 11251
2 83942 1 11275
2 83943 1 11275
2 83944 1 11275
2 83945 1 11275
2 83946 1 11275
2 83947 1 11275
2 83948 1 11276
2 83949 1 11276
2 83950 1 11276
2 83951 1 11276
2 83952 1 11276
2 83953 1 11276
2 83954 1 11276
2 83955 1 11276
2 83956 1 11276
2 83957 1 11276
2 83958 1 11276
2 83959 1 11276
2 83960 1 11276
2 83961 1 11276
2 83962 1 11276
2 83963 1 11276
2 83964 1 11276
2 83965 1 11276
2 83966 1 11276
2 83967 1 11276
2 83968 1 11276
2 83969 1 11277
2 83970 1 11277
2 83971 1 11292
2 83972 1 11292
2 83973 1 11292
2 83974 1 11292
2 83975 1 11292
2 83976 1 11292
2 83977 1 11292
2 83978 1 11300
2 83979 1 11300
2 83980 1 11301
2 83981 1 11301
2 83982 1 11315
2 83983 1 11315
2 83984 1 11316
2 83985 1 11316
2 83986 1 11321
2 83987 1 11321
2 83988 1 11344
2 83989 1 11344
2 83990 1 11353
2 83991 1 11353
2 83992 1 11365
2 83993 1 11365
2 83994 1 11380
2 83995 1 11380
2 83996 1 11381
2 83997 1 11381
2 83998 1 11381
2 83999 1 11381
2 84000 1 11381
2 84001 1 11381
2 84002 1 11381
2 84003 1 11381
2 84004 1 11381
2 84005 1 11381
2 84006 1 11381
2 84007 1 11381
2 84008 1 11381
2 84009 1 11381
2 84010 1 11381
2 84011 1 11381
2 84012 1 11381
2 84013 1 11381
2 84014 1 11381
2 84015 1 11381
2 84016 1 11381
2 84017 1 11381
2 84018 1 11381
2 84019 1 11381
2 84020 1 11381
2 84021 1 11383
2 84022 1 11383
2 84023 1 11383
2 84024 1 11386
2 84025 1 11386
2 84026 1 11386
2 84027 1 11386
2 84028 1 11386
2 84029 1 11386
2 84030 1 11387
2 84031 1 11387
2 84032 1 11387
2 84033 1 11392
2 84034 1 11392
2 84035 1 11393
2 84036 1 11393
2 84037 1 11393
2 84038 1 11394
2 84039 1 11394
2 84040 1 11401
2 84041 1 11401
2 84042 1 11404
2 84043 1 11404
2 84044 1 11404
2 84045 1 11404
2 84046 1 11404
2 84047 1 11404
2 84048 1 11404
2 84049 1 11411
2 84050 1 11411
2 84051 1 11412
2 84052 1 11412
2 84053 1 11428
2 84054 1 11428
2 84055 1 11428
2 84056 1 11428
2 84057 1 11428
2 84058 1 11428
2 84059 1 11428
2 84060 1 11428
2 84061 1 11428
2 84062 1 11428
2 84063 1 11428
2 84064 1 11428
2 84065 1 11428
2 84066 1 11428
2 84067 1 11428
2 84068 1 11428
2 84069 1 11428
2 84070 1 11428
2 84071 1 11428
2 84072 1 11429
2 84073 1 11429
2 84074 1 11453
2 84075 1 11453
2 84076 1 11453
2 84077 1 11454
2 84078 1 11454
2 84079 1 11454
2 84080 1 11454
2 84081 1 11454
2 84082 1 11454
2 84083 1 11454
2 84084 1 11454
2 84085 1 11454
2 84086 1 11454
2 84087 1 11454
2 84088 1 11454
2 84089 1 11455
2 84090 1 11455
2 84091 1 11458
2 84092 1 11458
2 84093 1 11475
2 84094 1 11475
2 84095 1 11475
2 84096 1 11476
2 84097 1 11476
2 84098 1 11497
2 84099 1 11497
2 84100 1 11498
2 84101 1 11498
2 84102 1 11498
2 84103 1 11506
2 84104 1 11506
2 84105 1 11516
2 84106 1 11516
2 84107 1 11533
2 84108 1 11533
2 84109 1 11533
2 84110 1 11547
2 84111 1 11547
2 84112 1 11567
2 84113 1 11567
2 84114 1 11567
2 84115 1 11582
2 84116 1 11582
2 84117 1 11582
2 84118 1 11582
2 84119 1 11591
2 84120 1 11591
2 84121 1 11591
2 84122 1 11591
2 84123 1 11603
2 84124 1 11603
2 84125 1 11603
2 84126 1 11603
2 84127 1 11603
2 84128 1 11603
2 84129 1 11603
2 84130 1 11603
2 84131 1 11604
2 84132 1 11604
2 84133 1 11604
2 84134 1 11611
2 84135 1 11611
2 84136 1 11629
2 84137 1 11629
2 84138 1 11629
2 84139 1 11649
2 84140 1 11649
2 84141 1 11651
2 84142 1 11651
2 84143 1 11665
2 84144 1 11665
2 84145 1 11667
2 84146 1 11667
2 84147 1 11687
2 84148 1 11687
2 84149 1 11691
2 84150 1 11691
2 84151 1 11691
2 84152 1 11692
2 84153 1 11692
2 84154 1 11692
2 84155 1 11692
2 84156 1 11692
2 84157 1 11693
2 84158 1 11693
2 84159 1 11701
2 84160 1 11701
2 84161 1 11702
2 84162 1 11702
2 84163 1 11702
2 84164 1 11702
2 84165 1 11702
2 84166 1 11702
2 84167 1 11702
2 84168 1 11704
2 84169 1 11704
2 84170 1 11709
2 84171 1 11709
2 84172 1 11709
2 84173 1 11709
2 84174 1 11709
2 84175 1 11709
2 84176 1 11709
2 84177 1 11709
2 84178 1 11709
2 84179 1 11709
2 84180 1 11709
2 84181 1 11709
2 84182 1 11709
2 84183 1 11709
2 84184 1 11709
2 84185 1 11725
2 84186 1 11725
2 84187 1 11725
2 84188 1 11725
2 84189 1 11725
2 84190 1 11725
2 84191 1 11725
2 84192 1 11725
2 84193 1 11725
2 84194 1 11725
2 84195 1 11725
2 84196 1 11725
2 84197 1 11725
2 84198 1 11725
2 84199 1 11725
2 84200 1 11726
2 84201 1 11726
2 84202 1 11726
2 84203 1 11726
2 84204 1 11726
2 84205 1 11726
2 84206 1 11726
2 84207 1 11726
2 84208 1 11727
2 84209 1 11727
2 84210 1 11738
2 84211 1 11738
2 84212 1 11778
2 84213 1 11778
2 84214 1 11778
2 84215 1 11778
2 84216 1 11791
2 84217 1 11791
2 84218 1 11808
2 84219 1 11808
2 84220 1 11808
2 84221 1 11808
2 84222 1 11808
2 84223 1 11808
2 84224 1 11808
2 84225 1 11808
2 84226 1 11809
2 84227 1 11809
2 84228 1 11826
2 84229 1 11826
2 84230 1 11873
2 84231 1 11873
2 84232 1 11874
2 84233 1 11874
2 84234 1 11875
2 84235 1 11875
2 84236 1 11875
2 84237 1 11875
2 84238 1 11875
2 84239 1 11875
2 84240 1 11875
2 84241 1 11875
2 84242 1 11875
2 84243 1 11875
2 84244 1 11875
2 84245 1 11875
2 84246 1 11876
2 84247 1 11876
2 84248 1 11876
2 84249 1 11876
2 84250 1 11876
2 84251 1 11876
2 84252 1 11878
2 84253 1 11878
2 84254 1 11890
2 84255 1 11890
2 84256 1 11891
2 84257 1 11891
2 84258 1 11893
2 84259 1 11893
2 84260 1 11924
2 84261 1 11924
2 84262 1 11924
2 84263 1 11924
2 84264 1 11924
2 84265 1 11924
2 84266 1 11924
2 84267 1 11924
2 84268 1 11924
2 84269 1 11927
2 84270 1 11927
2 84271 1 11937
2 84272 1 11937
2 84273 1 11937
2 84274 1 11937
2 84275 1 11941
2 84276 1 11941
2 84277 1 11941
2 84278 1 11941
2 84279 1 11941
2 84280 1 11942
2 84281 1 11942
2 84282 1 11942
2 84283 1 11944
2 84284 1 11944
2 84285 1 11944
2 84286 1 11944
2 84287 1 11961
2 84288 1 11961
2 84289 1 11962
2 84290 1 11962
2 84291 1 11963
2 84292 1 11963
2 84293 1 11963
2 84294 1 11966
2 84295 1 11966
2 84296 1 11966
2 84297 1 11966
2 84298 1 11966
2 84299 1 11966
2 84300 1 11966
2 84301 1 11966
2 84302 1 11966
2 84303 1 11966
2 84304 1 11966
2 84305 1 11976
2 84306 1 11976
2 84307 1 11982
2 84308 1 11982
2 84309 1 11994
2 84310 1 11994
2 84311 1 11994
2 84312 1 11994
2 84313 1 11994
2 84314 1 11994
2 84315 1 11994
2 84316 1 11994
2 84317 1 11994
2 84318 1 11994
2 84319 1 11995
2 84320 1 11995
2 84321 1 11996
2 84322 1 11996
2 84323 1 11996
2 84324 1 12019
2 84325 1 12019
2 84326 1 12020
2 84327 1 12020
2 84328 1 12020
2 84329 1 12020
2 84330 1 12020
2 84331 1 12020
2 84332 1 12021
2 84333 1 12021
2 84334 1 12021
2 84335 1 12039
2 84336 1 12039
2 84337 1 12039
2 84338 1 12039
2 84339 1 12039
2 84340 1 12039
2 84341 1 12039
2 84342 1 12040
2 84343 1 12040
2 84344 1 12040
2 84345 1 12040
2 84346 1 12040
2 84347 1 12040
2 84348 1 12040
2 84349 1 12040
2 84350 1 12040
2 84351 1 12040
2 84352 1 12040
2 84353 1 12040
2 84354 1 12042
2 84355 1 12042
2 84356 1 12044
2 84357 1 12044
2 84358 1 12046
2 84359 1 12046
2 84360 1 12083
2 84361 1 12083
2 84362 1 12084
2 84363 1 12084
2 84364 1 12084
2 84365 1 12084
2 84366 1 12084
2 84367 1 12084
2 84368 1 12084
2 84369 1 12084
2 84370 1 12084
2 84371 1 12084
2 84372 1 12084
2 84373 1 12084
2 84374 1 12084
2 84375 1 12084
2 84376 1 12084
2 84377 1 12084
2 84378 1 12084
2 84379 1 12084
2 84380 1 12085
2 84381 1 12085
2 84382 1 12085
2 84383 1 12086
2 84384 1 12086
2 84385 1 12086
2 84386 1 12087
2 84387 1 12087
2 84388 1 12090
2 84389 1 12090
2 84390 1 12090
2 84391 1 12091
2 84392 1 12091
2 84393 1 12091
2 84394 1 12108
2 84395 1 12108
2 84396 1 12117
2 84397 1 12117
2 84398 1 12117
2 84399 1 12138
2 84400 1 12138
2 84401 1 12138
2 84402 1 12139
2 84403 1 12139
2 84404 1 12139
2 84405 1 12140
2 84406 1 12140
2 84407 1 12141
2 84408 1 12141
2 84409 1 12141
2 84410 1 12141
2 84411 1 12141
2 84412 1 12141
2 84413 1 12141
2 84414 1 12141
2 84415 1 12141
2 84416 1 12141
2 84417 1 12142
2 84418 1 12142
2 84419 1 12143
2 84420 1 12143
2 84421 1 12145
2 84422 1 12145
2 84423 1 12145
2 84424 1 12146
2 84425 1 12146
2 84426 1 12150
2 84427 1 12150
2 84428 1 12151
2 84429 1 12151
2 84430 1 12152
2 84431 1 12152
2 84432 1 12171
2 84433 1 12171
2 84434 1 12172
2 84435 1 12172
2 84436 1 12172
2 84437 1 12183
2 84438 1 12183
2 84439 1 12183
2 84440 1 12185
2 84441 1 12185
2 84442 1 12196
2 84443 1 12196
2 84444 1 12197
2 84445 1 12197
2 84446 1 12197
2 84447 1 12197
2 84448 1 12197
2 84449 1 12200
2 84450 1 12200
2 84451 1 12201
2 84452 1 12201
2 84453 1 12201
2 84454 1 12201
2 84455 1 12201
2 84456 1 12201
2 84457 1 12201
2 84458 1 12201
2 84459 1 12201
2 84460 1 12201
2 84461 1 12202
2 84462 1 12202
2 84463 1 12203
2 84464 1 12203
2 84465 1 12218
2 84466 1 12218
2 84467 1 12218
2 84468 1 12219
2 84469 1 12219
2 84470 1 12219
2 84471 1 12219
2 84472 1 12219
2 84473 1 12219
2 84474 1 12219
2 84475 1 12219
2 84476 1 12220
2 84477 1 12220
2 84478 1 12221
2 84479 1 12221
2 84480 1 12221
2 84481 1 12221
2 84482 1 12221
2 84483 1 12221
2 84484 1 12222
2 84485 1 12222
2 84486 1 12222
2 84487 1 12222
2 84488 1 12222
2 84489 1 12222
2 84490 1 12223
2 84491 1 12223
2 84492 1 12230
2 84493 1 12230
2 84494 1 12238
2 84495 1 12238
2 84496 1 12241
2 84497 1 12241
2 84498 1 12242
2 84499 1 12242
2 84500 1 12242
2 84501 1 12242
2 84502 1 12242
2 84503 1 12242
2 84504 1 12242
2 84505 1 12242
2 84506 1 12244
2 84507 1 12244
2 84508 1 12250
2 84509 1 12250
2 84510 1 12255
2 84511 1 12255
2 84512 1 12255
2 84513 1 12255
2 84514 1 12256
2 84515 1 12256
2 84516 1 12258
2 84517 1 12258
2 84518 1 12259
2 84519 1 12259
2 84520 1 12259
2 84521 1 12259
2 84522 1 12260
2 84523 1 12260
2 84524 1 12275
2 84525 1 12275
2 84526 1 12275
2 84527 1 12276
2 84528 1 12276
2 84529 1 12277
2 84530 1 12277
2 84531 1 12277
2 84532 1 12277
2 84533 1 12281
2 84534 1 12281
2 84535 1 12283
2 84536 1 12283
2 84537 1 12283
2 84538 1 12291
2 84539 1 12291
2 84540 1 12291
2 84541 1 12291
2 84542 1 12298
2 84543 1 12298
2 84544 1 12299
2 84545 1 12299
2 84546 1 12299
2 84547 1 12311
2 84548 1 12311
2 84549 1 12311
2 84550 1 12311
2 84551 1 12311
2 84552 1 12312
2 84553 1 12312
2 84554 1 12312
2 84555 1 12324
2 84556 1 12324
2 84557 1 12324
2 84558 1 12324
2 84559 1 12324
2 84560 1 12325
2 84561 1 12325
2 84562 1 12344
2 84563 1 12344
2 84564 1 12344
2 84565 1 12344
2 84566 1 12345
2 84567 1 12345
2 84568 1 12345
2 84569 1 12345
2 84570 1 12345
2 84571 1 12346
2 84572 1 12346
2 84573 1 12346
2 84574 1 12346
2 84575 1 12346
2 84576 1 12346
2 84577 1 12346
2 84578 1 12346
2 84579 1 12346
2 84580 1 12346
2 84581 1 12349
2 84582 1 12349
2 84583 1 12349
2 84584 1 12353
2 84585 1 12353
2 84586 1 12361
2 84587 1 12361
2 84588 1 12361
2 84589 1 12361
2 84590 1 12361
2 84591 1 12361
2 84592 1 12361
2 84593 1 12361
2 84594 1 12361
2 84595 1 12361
2 84596 1 12361
2 84597 1 12361
2 84598 1 12361
2 84599 1 12363
2 84600 1 12363
2 84601 1 12376
2 84602 1 12376
2 84603 1 12376
2 84604 1 12376
2 84605 1 12387
2 84606 1 12387
2 84607 1 12387
2 84608 1 12423
2 84609 1 12423
2 84610 1 12423
2 84611 1 12423
2 84612 1 12423
2 84613 1 12423
2 84614 1 12423
2 84615 1 12426
2 84616 1 12426
2 84617 1 12426
2 84618 1 12426
2 84619 1 12428
2 84620 1 12428
2 84621 1 12429
2 84622 1 12429
2 84623 1 12432
2 84624 1 12432
2 84625 1 12434
2 84626 1 12434
2 84627 1 12434
2 84628 1 12438
2 84629 1 12438
2 84630 1 12498
2 84631 1 12498
2 84632 1 12498
2 84633 1 12499
2 84634 1 12499
2 84635 1 12499
2 84636 1 12499
2 84637 1 12499
2 84638 1 12499
2 84639 1 12499
2 84640 1 12509
2 84641 1 12509
2 84642 1 12509
2 84643 1 12516
2 84644 1 12516
2 84645 1 12525
2 84646 1 12525
2 84647 1 12525
2 84648 1 12525
2 84649 1 12525
2 84650 1 12525
2 84651 1 12525
2 84652 1 12525
2 84653 1 12525
2 84654 1 12525
2 84655 1 12525
2 84656 1 12525
2 84657 1 12525
2 84658 1 12525
2 84659 1 12525
2 84660 1 12525
2 84661 1 12525
2 84662 1 12525
2 84663 1 12525
2 84664 1 12525
2 84665 1 12525
2 84666 1 12525
2 84667 1 12525
2 84668 1 12525
2 84669 1 12525
2 84670 1 12525
2 84671 1 12525
2 84672 1 12525
2 84673 1 12525
2 84674 1 12525
2 84675 1 12525
2 84676 1 12525
2 84677 1 12525
2 84678 1 12525
2 84679 1 12525
2 84680 1 12525
2 84681 1 12525
2 84682 1 12525
2 84683 1 12525
2 84684 1 12525
2 84685 1 12525
2 84686 1 12525
2 84687 1 12525
2 84688 1 12525
2 84689 1 12525
2 84690 1 12525
2 84691 1 12525
2 84692 1 12525
2 84693 1 12525
2 84694 1 12525
2 84695 1 12525
2 84696 1 12525
2 84697 1 12525
2 84698 1 12525
2 84699 1 12525
2 84700 1 12525
2 84701 1 12525
2 84702 1 12525
2 84703 1 12525
2 84704 1 12525
2 84705 1 12525
2 84706 1 12526
2 84707 1 12526
2 84708 1 12526
2 84709 1 12526
2 84710 1 12542
2 84711 1 12542
2 84712 1 12552
2 84713 1 12552
2 84714 1 12578
2 84715 1 12578
2 84716 1 12579
2 84717 1 12579
2 84718 1 12588
2 84719 1 12588
2 84720 1 12588
2 84721 1 12598
2 84722 1 12598
2 84723 1 12598
2 84724 1 12598
2 84725 1 12598
2 84726 1 12599
2 84727 1 12599
2 84728 1 12599
2 84729 1 12605
2 84730 1 12605
2 84731 1 12605
2 84732 1 12605
2 84733 1 12617
2 84734 1 12617
2 84735 1 12619
2 84736 1 12619
2 84737 1 12622
2 84738 1 12622
2 84739 1 12637
2 84740 1 12637
2 84741 1 12637
2 84742 1 12637
2 84743 1 12637
2 84744 1 12637
2 84745 1 12637
2 84746 1 12654
2 84747 1 12654
2 84748 1 12654
2 84749 1 12655
2 84750 1 12655
2 84751 1 12656
2 84752 1 12656
2 84753 1 12672
2 84754 1 12672
2 84755 1 12672
2 84756 1 12672
2 84757 1 12672
2 84758 1 12672
2 84759 1 12683
2 84760 1 12683
2 84761 1 12691
2 84762 1 12691
2 84763 1 12691
2 84764 1 12692
2 84765 1 12692
2 84766 1 12697
2 84767 1 12697
2 84768 1 12697
2 84769 1 12698
2 84770 1 12698
2 84771 1 12698
2 84772 1 12698
2 84773 1 12706
2 84774 1 12706
2 84775 1 12706
2 84776 1 12706
2 84777 1 12706
2 84778 1 12706
2 84779 1 12706
2 84780 1 12706
2 84781 1 12706
2 84782 1 12706
2 84783 1 12706
2 84784 1 12706
2 84785 1 12706
2 84786 1 12706
2 84787 1 12706
2 84788 1 12706
2 84789 1 12706
2 84790 1 12706
2 84791 1 12706
2 84792 1 12706
2 84793 1 12708
2 84794 1 12708
2 84795 1 12708
2 84796 1 12708
2 84797 1 12708
2 84798 1 12708
2 84799 1 12708
2 84800 1 12708
2 84801 1 12708
2 84802 1 12709
2 84803 1 12709
2 84804 1 12709
2 84805 1 12733
2 84806 1 12733
2 84807 1 12734
2 84808 1 12734
2 84809 1 12734
2 84810 1 12735
2 84811 1 12735
2 84812 1 12737
2 84813 1 12737
2 84814 1 12739
2 84815 1 12739
2 84816 1 12748
2 84817 1 12748
2 84818 1 12753
2 84819 1 12753
2 84820 1 12756
2 84821 1 12756
2 84822 1 12766
2 84823 1 12766
2 84824 1 12767
2 84825 1 12767
2 84826 1 12770
2 84827 1 12770
2 84828 1 12771
2 84829 1 12771
2 84830 1 12781
2 84831 1 12781
2 84832 1 12788
2 84833 1 12788
2 84834 1 12801
2 84835 1 12801
2 84836 1 12802
2 84837 1 12802
2 84838 1 12804
2 84839 1 12804
2 84840 1 12806
2 84841 1 12806
2 84842 1 12806
2 84843 1 12807
2 84844 1 12807
2 84845 1 12808
2 84846 1 12808
2 84847 1 12808
2 84848 1 12820
2 84849 1 12820
2 84850 1 12838
2 84851 1 12838
2 84852 1 12839
2 84853 1 12839
2 84854 1 12841
2 84855 1 12841
2 84856 1 12841
2 84857 1 12845
2 84858 1 12845
2 84859 1 12848
2 84860 1 12848
2 84861 1 12848
2 84862 1 12848
2 84863 1 12848
2 84864 1 12851
2 84865 1 12851
2 84866 1 12851
2 84867 1 12851
2 84868 1 12861
2 84869 1 12861
2 84870 1 12867
2 84871 1 12867
2 84872 1 12867
2 84873 1 12867
2 84874 1 12867
2 84875 1 12867
2 84876 1 12867
2 84877 1 12867
2 84878 1 12867
2 84879 1 12868
2 84880 1 12868
2 84881 1 12869
2 84882 1 12869
2 84883 1 12869
2 84884 1 12869
2 84885 1 12869
2 84886 1 12869
2 84887 1 12869
2 84888 1 12869
2 84889 1 12869
2 84890 1 12871
2 84891 1 12871
2 84892 1 12872
2 84893 1 12872
2 84894 1 12873
2 84895 1 12873
2 84896 1 12873
2 84897 1 12883
2 84898 1 12883
2 84899 1 12883
2 84900 1 12883
2 84901 1 12886
2 84902 1 12886
2 84903 1 12887
2 84904 1 12887
2 84905 1 12888
2 84906 1 12888
2 84907 1 12889
2 84908 1 12889
2 84909 1 12890
2 84910 1 12890
2 84911 1 12890
2 84912 1 12890
2 84913 1 12891
2 84914 1 12891
2 84915 1 12899
2 84916 1 12899
2 84917 1 12899
2 84918 1 12899
2 84919 1 12899
2 84920 1 12899
2 84921 1 12899
2 84922 1 12900
2 84923 1 12900
2 84924 1 12900
2 84925 1 12900
2 84926 1 12900
2 84927 1 12900
2 84928 1 12900
2 84929 1 12900
2 84930 1 12900
2 84931 1 12900
2 84932 1 12900
2 84933 1 12903
2 84934 1 12903
2 84935 1 12903
2 84936 1 12909
2 84937 1 12909
2 84938 1 12909
2 84939 1 12909
2 84940 1 12918
2 84941 1 12918
2 84942 1 12918
2 84943 1 12918
2 84944 1 12921
2 84945 1 12921
2 84946 1 12921
2 84947 1 12923
2 84948 1 12923
2 84949 1 12935
2 84950 1 12935
2 84951 1 12937
2 84952 1 12937
2 84953 1 12937
2 84954 1 12937
2 84955 1 12937
2 84956 1 12942
2 84957 1 12942
2 84958 1 12946
2 84959 1 12946
2 84960 1 12947
2 84961 1 12947
2 84962 1 12947
2 84963 1 12947
2 84964 1 12949
2 84965 1 12949
2 84966 1 12951
2 84967 1 12951
2 84968 1 12952
2 84969 1 12952
2 84970 1 12952
2 84971 1 12960
2 84972 1 12960
2 84973 1 12964
2 84974 1 12964
2 84975 1 12964
2 84976 1 12965
2 84977 1 12965
2 84978 1 12965
2 84979 1 12965
2 84980 1 12965
2 84981 1 12965
2 84982 1 12965
2 84983 1 12965
2 84984 1 12965
2 84985 1 12965
2 84986 1 12965
2 84987 1 12965
2 84988 1 12965
2 84989 1 12965
2 84990 1 12965
2 84991 1 12965
2 84992 1 12965
2 84993 1 12965
2 84994 1 12965
2 84995 1 12965
2 84996 1 12965
2 84997 1 12968
2 84998 1 12968
2 84999 1 12968
2 85000 1 12968
2 85001 1 12983
2 85002 1 12983
2 85003 1 12983
2 85004 1 12983
2 85005 1 12983
2 85006 1 12992
2 85007 1 12992
2 85008 1 13010
2 85009 1 13010
2 85010 1 13037
2 85011 1 13037
2 85012 1 13053
2 85013 1 13053
2 85014 1 13055
2 85015 1 13055
2 85016 1 13057
2 85017 1 13057
2 85018 1 13057
2 85019 1 13057
2 85020 1 13057
2 85021 1 13057
2 85022 1 13057
2 85023 1 13058
2 85024 1 13058
2 85025 1 13058
2 85026 1 13061
2 85027 1 13061
2 85028 1 13063
2 85029 1 13063
2 85030 1 13083
2 85031 1 13083
2 85032 1 13099
2 85033 1 13099
2 85034 1 13099
2 85035 1 13100
2 85036 1 13100
2 85037 1 13106
2 85038 1 13106
2 85039 1 13111
2 85040 1 13111
2 85041 1 13111
2 85042 1 13111
2 85043 1 13112
2 85044 1 13112
2 85045 1 13112
2 85046 1 13112
2 85047 1 13114
2 85048 1 13114
2 85049 1 13123
2 85050 1 13123
2 85051 1 13124
2 85052 1 13124
2 85053 1 13126
2 85054 1 13126
2 85055 1 13139
2 85056 1 13139
2 85057 1 13163
2 85058 1 13163
2 85059 1 13164
2 85060 1 13164
2 85061 1 13164
2 85062 1 13164
2 85063 1 13164
2 85064 1 13167
2 85065 1 13167
2 85066 1 13168
2 85067 1 13168
2 85068 1 13168
2 85069 1 13170
2 85070 1 13170
2 85071 1 13171
2 85072 1 13171
2 85073 1 13175
2 85074 1 13175
2 85075 1 13175
2 85076 1 13175
2 85077 1 13175
2 85078 1 13175
2 85079 1 13176
2 85080 1 13176
2 85081 1 13184
2 85082 1 13184
2 85083 1 13184
2 85084 1 13184
2 85085 1 13184
2 85086 1 13184
2 85087 1 13184
2 85088 1 13184
2 85089 1 13184
2 85090 1 13184
2 85091 1 13184
2 85092 1 13193
2 85093 1 13193
2 85094 1 13193
2 85095 1 13193
2 85096 1 13193
2 85097 1 13194
2 85098 1 13194
2 85099 1 13194
2 85100 1 13194
2 85101 1 13194
2 85102 1 13195
2 85103 1 13195
2 85104 1 13196
2 85105 1 13196
2 85106 1 13204
2 85107 1 13204
2 85108 1 13204
2 85109 1 13204
2 85110 1 13204
2 85111 1 13205
2 85112 1 13205
2 85113 1 13207
2 85114 1 13207
2 85115 1 13220
2 85116 1 13220
2 85117 1 13220
2 85118 1 13229
2 85119 1 13229
2 85120 1 13229
2 85121 1 13230
2 85122 1 13230
2 85123 1 13231
2 85124 1 13231
2 85125 1 13231
2 85126 1 13235
2 85127 1 13235
2 85128 1 13235
2 85129 1 13235
2 85130 1 13235
2 85131 1 13235
2 85132 1 13235
2 85133 1 13235
2 85134 1 13235
2 85135 1 13235
2 85136 1 13235
2 85137 1 13235
2 85138 1 13235
2 85139 1 13235
2 85140 1 13235
2 85141 1 13235
2 85142 1 13235
2 85143 1 13235
2 85144 1 13235
2 85145 1 13236
2 85146 1 13236
2 85147 1 13236
2 85148 1 13236
2 85149 1 13236
2 85150 1 13236
2 85151 1 13236
2 85152 1 13236
2 85153 1 13236
2 85154 1 13236
2 85155 1 13236
2 85156 1 13236
2 85157 1 13236
2 85158 1 13236
2 85159 1 13236
2 85160 1 13236
2 85161 1 13236
2 85162 1 13236
2 85163 1 13236
2 85164 1 13236
2 85165 1 13236
2 85166 1 13236
2 85167 1 13236
2 85168 1 13236
2 85169 1 13236
2 85170 1 13236
2 85171 1 13236
2 85172 1 13236
2 85173 1 13236
2 85174 1 13236
2 85175 1 13236
2 85176 1 13236
2 85177 1 13236
2 85178 1 13236
2 85179 1 13236
2 85180 1 13236
2 85181 1 13236
2 85182 1 13236
2 85183 1 13236
2 85184 1 13236
2 85185 1 13236
2 85186 1 13236
2 85187 1 13236
2 85188 1 13236
2 85189 1 13236
2 85190 1 13238
2 85191 1 13238
2 85192 1 13263
2 85193 1 13263
2 85194 1 13263
2 85195 1 13264
2 85196 1 13264
2 85197 1 13264
2 85198 1 13265
2 85199 1 13265
2 85200 1 13265
2 85201 1 13265
2 85202 1 13269
2 85203 1 13269
2 85204 1 13269
2 85205 1 13269
2 85206 1 13269
2 85207 1 13271
2 85208 1 13271
2 85209 1 13271
2 85210 1 13271
2 85211 1 13272
2 85212 1 13272
2 85213 1 13273
2 85214 1 13273
2 85215 1 13273
2 85216 1 13274
2 85217 1 13274
2 85218 1 13274
2 85219 1 13275
2 85220 1 13275
2 85221 1 13275
2 85222 1 13275
2 85223 1 13275
2 85224 1 13277
2 85225 1 13277
2 85226 1 13280
2 85227 1 13280
2 85228 1 13281
2 85229 1 13281
2 85230 1 13290
2 85231 1 13290
2 85232 1 13290
2 85233 1 13291
2 85234 1 13291
2 85235 1 13293
2 85236 1 13293
2 85237 1 13302
2 85238 1 13302
2 85239 1 13302
2 85240 1 13305
2 85241 1 13305
2 85242 1 13305
2 85243 1 13308
2 85244 1 13308
2 85245 1 13309
2 85246 1 13309
2 85247 1 13309
2 85248 1 13318
2 85249 1 13318
2 85250 1 13326
2 85251 1 13326
2 85252 1 13326
2 85253 1 13327
2 85254 1 13327
2 85255 1 13327
2 85256 1 13334
2 85257 1 13334
2 85258 1 13334
2 85259 1 13335
2 85260 1 13335
2 85261 1 13336
2 85262 1 13336
2 85263 1 13336
2 85264 1 13336
2 85265 1 13336
2 85266 1 13339
2 85267 1 13339
2 85268 1 13339
2 85269 1 13360
2 85270 1 13360
2 85271 1 13362
2 85272 1 13362
2 85273 1 13378
2 85274 1 13378
2 85275 1 13386
2 85276 1 13386
2 85277 1 13397
2 85278 1 13397
2 85279 1 13397
2 85280 1 13397
2 85281 1 13397
2 85282 1 13397
2 85283 1 13397
2 85284 1 13403
2 85285 1 13403
2 85286 1 13413
2 85287 1 13413
2 85288 1 13413
2 85289 1 13413
2 85290 1 13413
2 85291 1 13413
2 85292 1 13413
2 85293 1 13413
2 85294 1 13413
2 85295 1 13413
2 85296 1 13413
2 85297 1 13413
2 85298 1 13413
2 85299 1 13413
2 85300 1 13413
2 85301 1 13413
2 85302 1 13413
2 85303 1 13413
2 85304 1 13413
2 85305 1 13413
2 85306 1 13413
2 85307 1 13413
2 85308 1 13413
2 85309 1 13432
2 85310 1 13432
2 85311 1 13432
2 85312 1 13432
2 85313 1 13432
2 85314 1 13432
2 85315 1 13441
2 85316 1 13441
2 85317 1 13455
2 85318 1 13455
2 85319 1 13455
2 85320 1 13458
2 85321 1 13458
2 85322 1 13476
2 85323 1 13476
2 85324 1 13476
2 85325 1 13476
2 85326 1 13479
2 85327 1 13479
2 85328 1 13479
2 85329 1 13482
2 85330 1 13482
2 85331 1 13482
2 85332 1 13494
2 85333 1 13494
2 85334 1 13501
2 85335 1 13501
2 85336 1 13501
2 85337 1 13501
2 85338 1 13501
2 85339 1 13501
2 85340 1 13501
2 85341 1 13502
2 85342 1 13502
2 85343 1 13502
2 85344 1 13503
2 85345 1 13503
2 85346 1 13508
2 85347 1 13508
2 85348 1 13508
2 85349 1 13508
2 85350 1 13508
2 85351 1 13508
2 85352 1 13508
2 85353 1 13508
2 85354 1 13508
2 85355 1 13509
2 85356 1 13509
2 85357 1 13510
2 85358 1 13510
2 85359 1 13510
2 85360 1 13510
2 85361 1 13510
2 85362 1 13516
2 85363 1 13516
2 85364 1 13516
2 85365 1 13516
2 85366 1 13516
2 85367 1 13517
2 85368 1 13517
2 85369 1 13529
2 85370 1 13529
2 85371 1 13533
2 85372 1 13533
2 85373 1 13549
2 85374 1 13549
2 85375 1 13550
2 85376 1 13550
2 85377 1 13551
2 85378 1 13551
2 85379 1 13551
2 85380 1 13551
2 85381 1 13551
2 85382 1 13551
2 85383 1 13551
2 85384 1 13551
2 85385 1 13551
2 85386 1 13551
2 85387 1 13552
2 85388 1 13552
2 85389 1 13564
2 85390 1 13564
2 85391 1 13566
2 85392 1 13566
2 85393 1 13567
2 85394 1 13567
2 85395 1 13567
2 85396 1 13567
2 85397 1 13567
2 85398 1 13567
2 85399 1 13567
2 85400 1 13570
2 85401 1 13570
2 85402 1 13571
2 85403 1 13571
2 85404 1 13571
2 85405 1 13571
2 85406 1 13572
2 85407 1 13572
2 85408 1 13572
2 85409 1 13572
2 85410 1 13572
2 85411 1 13572
2 85412 1 13576
2 85413 1 13576
2 85414 1 13577
2 85415 1 13577
2 85416 1 13577
2 85417 1 13587
2 85418 1 13587
2 85419 1 13589
2 85420 1 13589
2 85421 1 13594
2 85422 1 13594
2 85423 1 13595
2 85424 1 13595
2 85425 1 13595
2 85426 1 13595
2 85427 1 13595
2 85428 1 13595
2 85429 1 13596
2 85430 1 13596
2 85431 1 13606
2 85432 1 13606
2 85433 1 13607
2 85434 1 13607
2 85435 1 13607
2 85436 1 13607
2 85437 1 13607
2 85438 1 13614
2 85439 1 13614
2 85440 1 13626
2 85441 1 13626
2 85442 1 13630
2 85443 1 13630
2 85444 1 13630
2 85445 1 13638
2 85446 1 13638
2 85447 1 13639
2 85448 1 13639
2 85449 1 13640
2 85450 1 13640
2 85451 1 13640
2 85452 1 13660
2 85453 1 13660
2 85454 1 13660
2 85455 1 13668
2 85456 1 13668
2 85457 1 13668
2 85458 1 13668
2 85459 1 13668
2 85460 1 13668
2 85461 1 13668
2 85462 1 13668
2 85463 1 13668
2 85464 1 13668
2 85465 1 13668
2 85466 1 13668
2 85467 1 13681
2 85468 1 13681
2 85469 1 13681
2 85470 1 13681
2 85471 1 13681
2 85472 1 13681
2 85473 1 13681
2 85474 1 13682
2 85475 1 13682
2 85476 1 13682
2 85477 1 13682
2 85478 1 13683
2 85479 1 13683
2 85480 1 13684
2 85481 1 13684
2 85482 1 13684
2 85483 1 13684
2 85484 1 13684
2 85485 1 13684
2 85486 1 13684
2 85487 1 13684
2 85488 1 13684
2 85489 1 13684
2 85490 1 13684
2 85491 1 13687
2 85492 1 13687
2 85493 1 13693
2 85494 1 13693
2 85495 1 13693
2 85496 1 13693
2 85497 1 13693
2 85498 1 13694
2 85499 1 13694
2 85500 1 13713
2 85501 1 13713
2 85502 1 13758
2 85503 1 13758
2 85504 1 13774
2 85505 1 13774
2 85506 1 13774
2 85507 1 13774
2 85508 1 13774
2 85509 1 13774
2 85510 1 13775
2 85511 1 13775
2 85512 1 13775
2 85513 1 13775
2 85514 1 13778
2 85515 1 13778
2 85516 1 13782
2 85517 1 13782
2 85518 1 13798
2 85519 1 13798
2 85520 1 13798
2 85521 1 13798
2 85522 1 13798
2 85523 1 13813
2 85524 1 13813
2 85525 1 13813
2 85526 1 13824
2 85527 1 13824
2 85528 1 13824
2 85529 1 13824
2 85530 1 13824
2 85531 1 13824
2 85532 1 13828
2 85533 1 13828
2 85534 1 13828
2 85535 1 13829
2 85536 1 13829
2 85537 1 13829
2 85538 1 13829
2 85539 1 13829
2 85540 1 13829
2 85541 1 13829
2 85542 1 13830
2 85543 1 13830
2 85544 1 13830
2 85545 1 13830
2 85546 1 13830
2 85547 1 13830
2 85548 1 13830
2 85549 1 13830
2 85550 1 13830
2 85551 1 13830
2 85552 1 13830
2 85553 1 13830
2 85554 1 13831
2 85555 1 13831
2 85556 1 13831
2 85557 1 13831
2 85558 1 13831
2 85559 1 13831
2 85560 1 13839
2 85561 1 13839
2 85562 1 13849
2 85563 1 13849
2 85564 1 13850
2 85565 1 13850
2 85566 1 13850
2 85567 1 13851
2 85568 1 13851
2 85569 1 13851
2 85570 1 13851
2 85571 1 13851
2 85572 1 13851
2 85573 1 13851
2 85574 1 13851
2 85575 1 13851
2 85576 1 13851
2 85577 1 13856
2 85578 1 13856
2 85579 1 13868
2 85580 1 13868
2 85581 1 13886
2 85582 1 13886
2 85583 1 13912
2 85584 1 13912
2 85585 1 13916
2 85586 1 13916
2 85587 1 13916
2 85588 1 13916
2 85589 1 13918
2 85590 1 13918
2 85591 1 13918
2 85592 1 13918
2 85593 1 13919
2 85594 1 13919
2 85595 1 13919
2 85596 1 13919
2 85597 1 13920
2 85598 1 13920
2 85599 1 13921
2 85600 1 13921
2 85601 1 13927
2 85602 1 13927
2 85603 1 13927
2 85604 1 13932
2 85605 1 13932
2 85606 1 13936
2 85607 1 13936
2 85608 1 13939
2 85609 1 13939
2 85610 1 13939
2 85611 1 13939
2 85612 1 13965
2 85613 1 13965
2 85614 1 13965
2 85615 1 13968
2 85616 1 13968
2 85617 1 13968
2 85618 1 13969
2 85619 1 13969
2 85620 1 13988
2 85621 1 13988
2 85622 1 13988
2 85623 1 13988
2 85624 1 13988
2 85625 1 13988
2 85626 1 13988
2 85627 1 13988
2 85628 1 13989
2 85629 1 13989
2 85630 1 13989
2 85631 1 14001
2 85632 1 14001
2 85633 1 14001
2 85634 1 14011
2 85635 1 14011
2 85636 1 14011
2 85637 1 14012
2 85638 1 14012
2 85639 1 14012
2 85640 1 14012
2 85641 1 14012
2 85642 1 14026
2 85643 1 14026
2 85644 1 14026
2 85645 1 14026
2 85646 1 14026
2 85647 1 14026
2 85648 1 14026
2 85649 1 14026
2 85650 1 14026
2 85651 1 14027
2 85652 1 14027
2 85653 1 14027
2 85654 1 14027
2 85655 1 14027
2 85656 1 14027
2 85657 1 14027
2 85658 1 14027
2 85659 1 14028
2 85660 1 14028
2 85661 1 14028
2 85662 1 14030
2 85663 1 14030
2 85664 1 14031
2 85665 1 14031
2 85666 1 14032
2 85667 1 14032
2 85668 1 14032
2 85669 1 14033
2 85670 1 14033
2 85671 1 14033
2 85672 1 14035
2 85673 1 14035
2 85674 1 14040
2 85675 1 14040
2 85676 1 14049
2 85677 1 14049
2 85678 1 14049
2 85679 1 14050
2 85680 1 14050
2 85681 1 14051
2 85682 1 14051
2 85683 1 14051
2 85684 1 14051
2 85685 1 14051
2 85686 1 14051
2 85687 1 14051
2 85688 1 14051
2 85689 1 14051
2 85690 1 14051
2 85691 1 14051
2 85692 1 14051
2 85693 1 14051
2 85694 1 14051
2 85695 1 14051
2 85696 1 14051
2 85697 1 14051
2 85698 1 14051
2 85699 1 14051
2 85700 1 14051
2 85701 1 14051
2 85702 1 14051
2 85703 1 14051
2 85704 1 14051
2 85705 1 14051
2 85706 1 14051
2 85707 1 14052
2 85708 1 14052
2 85709 1 14053
2 85710 1 14053
2 85711 1 14056
2 85712 1 14056
2 85713 1 14056
2 85714 1 14077
2 85715 1 14077
2 85716 1 14098
2 85717 1 14098
2 85718 1 14101
2 85719 1 14101
2 85720 1 14102
2 85721 1 14102
2 85722 1 14102
2 85723 1 14102
2 85724 1 14102
2 85725 1 14102
2 85726 1 14102
2 85727 1 14102
2 85728 1 14102
2 85729 1 14102
2 85730 1 14102
2 85731 1 14103
2 85732 1 14103
2 85733 1 14113
2 85734 1 14113
2 85735 1 14113
2 85736 1 14114
2 85737 1 14114
2 85738 1 14139
2 85739 1 14139
2 85740 1 14139
2 85741 1 14139
2 85742 1 14139
2 85743 1 14139
2 85744 1 14143
2 85745 1 14143
2 85746 1 14156
2 85747 1 14156
2 85748 1 14169
2 85749 1 14169
2 85750 1 14177
2 85751 1 14177
2 85752 1 14177
2 85753 1 14190
2 85754 1 14190
2 85755 1 14198
2 85756 1 14198
2 85757 1 14198
2 85758 1 14198
2 85759 1 14199
2 85760 1 14199
2 85761 1 14199
2 85762 1 14199
2 85763 1 14199
2 85764 1 14199
2 85765 1 14200
2 85766 1 14200
2 85767 1 14210
2 85768 1 14210
2 85769 1 14211
2 85770 1 14211
2 85771 1 14225
2 85772 1 14225
2 85773 1 14225
2 85774 1 14225
2 85775 1 14225
2 85776 1 14225
2 85777 1 14225
2 85778 1 14225
2 85779 1 14225
2 85780 1 14225
2 85781 1 14226
2 85782 1 14226
2 85783 1 14226
2 85784 1 14226
2 85785 1 14226
2 85786 1 14226
2 85787 1 14226
2 85788 1 14230
2 85789 1 14230
2 85790 1 14230
2 85791 1 14233
2 85792 1 14233
2 85793 1 14233
2 85794 1 14233
2 85795 1 14233
2 85796 1 14233
2 85797 1 14233
2 85798 1 14233
2 85799 1 14233
2 85800 1 14233
2 85801 1 14233
2 85802 1 14233
2 85803 1 14233
2 85804 1 14233
2 85805 1 14233
2 85806 1 14233
2 85807 1 14233
2 85808 1 14233
2 85809 1 14233
2 85810 1 14233
2 85811 1 14233
2 85812 1 14234
2 85813 1 14234
2 85814 1 14234
2 85815 1 14234
2 85816 1 14234
2 85817 1 14234
2 85818 1 14250
2 85819 1 14250
2 85820 1 14258
2 85821 1 14258
2 85822 1 14258
2 85823 1 14258
2 85824 1 14258
2 85825 1 14259
2 85826 1 14259
2 85827 1 14268
2 85828 1 14268
2 85829 1 14268
2 85830 1 14268
2 85831 1 14269
2 85832 1 14269
2 85833 1 14285
2 85834 1 14285
2 85835 1 14285
2 85836 1 14285
2 85837 1 14285
2 85838 1 14285
2 85839 1 14285
2 85840 1 14286
2 85841 1 14286
2 85842 1 14286
2 85843 1 14286
2 85844 1 14286
2 85845 1 14286
2 85846 1 14287
2 85847 1 14287
2 85848 1 14293
2 85849 1 14293
2 85850 1 14308
2 85851 1 14308
2 85852 1 14308
2 85853 1 14308
2 85854 1 14308
2 85855 1 14308
2 85856 1 14334
2 85857 1 14334
2 85858 1 14335
2 85859 1 14335
2 85860 1 14335
2 85861 1 14335
2 85862 1 14346
2 85863 1 14346
2 85864 1 14353
2 85865 1 14353
2 85866 1 14380
2 85867 1 14380
2 85868 1 14381
2 85869 1 14381
2 85870 1 14383
2 85871 1 14383
2 85872 1 14390
2 85873 1 14390
2 85874 1 14396
2 85875 1 14396
2 85876 1 14396
2 85877 1 14397
2 85878 1 14397
2 85879 1 14397
2 85880 1 14397
2 85881 1 14397
2 85882 1 14397
2 85883 1 14397
2 85884 1 14397
2 85885 1 14397
2 85886 1 14410
2 85887 1 14410
2 85888 1 14411
2 85889 1 14411
2 85890 1 14412
2 85891 1 14412
2 85892 1 14412
2 85893 1 14412
2 85894 1 14412
2 85895 1 14412
2 85896 1 14414
2 85897 1 14414
2 85898 1 14414
2 85899 1 14414
2 85900 1 14414
2 85901 1 14415
2 85902 1 14415
2 85903 1 14415
2 85904 1 14431
2 85905 1 14431
2 85906 1 14438
2 85907 1 14438
2 85908 1 14438
2 85909 1 14438
2 85910 1 14453
2 85911 1 14453
2 85912 1 14455
2 85913 1 14455
2 85914 1 14467
2 85915 1 14467
2 85916 1 14477
2 85917 1 14477
2 85918 1 14478
2 85919 1 14478
2 85920 1 14478
2 85921 1 14478
2 85922 1 14495
2 85923 1 14495
2 85924 1 14497
2 85925 1 14497
2 85926 1 14497
2 85927 1 14498
2 85928 1 14498
2 85929 1 14504
2 85930 1 14504
2 85931 1 14504
2 85932 1 14504
2 85933 1 14513
2 85934 1 14513
2 85935 1 14513
2 85936 1 14515
2 85937 1 14515
2 85938 1 14533
2 85939 1 14533
2 85940 1 14534
2 85941 1 14534
2 85942 1 14534
2 85943 1 14534
2 85944 1 14537
2 85945 1 14537
2 85946 1 14545
2 85947 1 14545
2 85948 1 14546
2 85949 1 14546
2 85950 1 14552
2 85951 1 14552
2 85952 1 14553
2 85953 1 14553
2 85954 1 14557
2 85955 1 14557
2 85956 1 14557
2 85957 1 14558
2 85958 1 14558
2 85959 1 14558
2 85960 1 14558
2 85961 1 14558
2 85962 1 14558
2 85963 1 14558
2 85964 1 14568
2 85965 1 14568
2 85966 1 14570
2 85967 1 14570
2 85968 1 14572
2 85969 1 14572
2 85970 1 14573
2 85971 1 14573
2 85972 1 14573
2 85973 1 14573
2 85974 1 14573
2 85975 1 14581
2 85976 1 14581
2 85977 1 14587
2 85978 1 14587
2 85979 1 14587
2 85980 1 14588
2 85981 1 14588
2 85982 1 14593
2 85983 1 14593
2 85984 1 14593
2 85985 1 14593
2 85986 1 14593
2 85987 1 14594
2 85988 1 14594
2 85989 1 14594
2 85990 1 14594
2 85991 1 14595
2 85992 1 14595
2 85993 1 14597
2 85994 1 14597
2 85995 1 14602
2 85996 1 14602
2 85997 1 14605
2 85998 1 14605
2 85999 1 14605
2 86000 1 14656
2 86001 1 14656
2 86002 1 14656
2 86003 1 14657
2 86004 1 14657
2 86005 1 14658
2 86006 1 14658
2 86007 1 14658
2 86008 1 14670
2 86009 1 14670
2 86010 1 14677
2 86011 1 14677
2 86012 1 14682
2 86013 1 14682
2 86014 1 14682
2 86015 1 14682
2 86016 1 14682
2 86017 1 14682
2 86018 1 14682
2 86019 1 14682
2 86020 1 14683
2 86021 1 14683
2 86022 1 14684
2 86023 1 14684
2 86024 1 14702
2 86025 1 14702
2 86026 1 14702
2 86027 1 14702
2 86028 1 14702
2 86029 1 14702
2 86030 1 14702
2 86031 1 14702
2 86032 1 14715
2 86033 1 14715
2 86034 1 14716
2 86035 1 14716
2 86036 1 14718
2 86037 1 14718
2 86038 1 14718
2 86039 1 14734
2 86040 1 14734
2 86041 1 14734
2 86042 1 14734
2 86043 1 14734
2 86044 1 14734
2 86045 1 14734
2 86046 1 14734
2 86047 1 14735
2 86048 1 14735
2 86049 1 14743
2 86050 1 14743
2 86051 1 14743
2 86052 1 14753
2 86053 1 14753
2 86054 1 14753
2 86055 1 14753
2 86056 1 14753
2 86057 1 14753
2 86058 1 14753
2 86059 1 14756
2 86060 1 14756
2 86061 1 14756
2 86062 1 14756
2 86063 1 14756
2 86064 1 14756
2 86065 1 14756
2 86066 1 14756
2 86067 1 14756
2 86068 1 14756
2 86069 1 14756
2 86070 1 14756
2 86071 1 14756
2 86072 1 14756
2 86073 1 14756
2 86074 1 14757
2 86075 1 14757
2 86076 1 14758
2 86077 1 14758
2 86078 1 14761
2 86079 1 14761
2 86080 1 14761
2 86081 1 14768
2 86082 1 14768
2 86083 1 14768
2 86084 1 14768
2 86085 1 14770
2 86086 1 14770
2 86087 1 14770
2 86088 1 14770
2 86089 1 14770
2 86090 1 14770
2 86091 1 14784
2 86092 1 14784
2 86093 1 14784
2 86094 1 14784
2 86095 1 14784
2 86096 1 14786
2 86097 1 14786
2 86098 1 14788
2 86099 1 14788
2 86100 1 14790
2 86101 1 14790
2 86102 1 14802
2 86103 1 14802
2 86104 1 14802
2 86105 1 14802
2 86106 1 14802
2 86107 1 14802
2 86108 1 14802
2 86109 1 14802
2 86110 1 14802
2 86111 1 14802
2 86112 1 14802
2 86113 1 14802
2 86114 1 14805
2 86115 1 14805
2 86116 1 14805
2 86117 1 14805
2 86118 1 14805
2 86119 1 14805
2 86120 1 14805
2 86121 1 14805
2 86122 1 14805
2 86123 1 14805
2 86124 1 14805
2 86125 1 14805
2 86126 1 14805
2 86127 1 14805
2 86128 1 14805
2 86129 1 14805
2 86130 1 14806
2 86131 1 14806
2 86132 1 14806
2 86133 1 14806
2 86134 1 14834
2 86135 1 14834
2 86136 1 14835
2 86137 1 14835
2 86138 1 14836
2 86139 1 14836
2 86140 1 14836
2 86141 1 14838
2 86142 1 14838
2 86143 1 14838
2 86144 1 14838
2 86145 1 14840
2 86146 1 14840
2 86147 1 14842
2 86148 1 14842
2 86149 1 14843
2 86150 1 14843
2 86151 1 14854
2 86152 1 14854
2 86153 1 14855
2 86154 1 14855
2 86155 1 14866
2 86156 1 14866
2 86157 1 14870
2 86158 1 14870
2 86159 1 14870
2 86160 1 14870
2 86161 1 14872
2 86162 1 14872
2 86163 1 14872
2 86164 1 14900
2 86165 1 14900
2 86166 1 14900
2 86167 1 14938
2 86168 1 14938
2 86169 1 14938
2 86170 1 14941
2 86171 1 14941
2 86172 1 14941
2 86173 1 14945
2 86174 1 14945
2 86175 1 14946
2 86176 1 14946
2 86177 1 14946
2 86178 1 14946
2 86179 1 14962
2 86180 1 14962
2 86181 1 14966
2 86182 1 14966
2 86183 1 14966
2 86184 1 14970
2 86185 1 14970
2 86186 1 14972
2 86187 1 14972
2 86188 1 14989
2 86189 1 14989
2 86190 1 14991
2 86191 1 14991
2 86192 1 14991
2 86193 1 14992
2 86194 1 14992
2 86195 1 14995
2 86196 1 14995
2 86197 1 14995
2 86198 1 14996
2 86199 1 14996
2 86200 1 14996
2 86201 1 14996
2 86202 1 14996
2 86203 1 14998
2 86204 1 14998
2 86205 1 15002
2 86206 1 15002
2 86207 1 15002
2 86208 1 15002
2 86209 1 15002
2 86210 1 15002
2 86211 1 15003
2 86212 1 15003
2 86213 1 15003
2 86214 1 15003
2 86215 1 15003
2 86216 1 15011
2 86217 1 15011
2 86218 1 15068
2 86219 1 15068
2 86220 1 15069
2 86221 1 15069
2 86222 1 15093
2 86223 1 15093
2 86224 1 15121
2 86225 1 15121
2 86226 1 15129
2 86227 1 15129
2 86228 1 15148
2 86229 1 15148
2 86230 1 15167
2 86231 1 15167
2 86232 1 15177
2 86233 1 15177
2 86234 1 15177
2 86235 1 15177
2 86236 1 15177
2 86237 1 15177
2 86238 1 15177
2 86239 1 15177
2 86240 1 15177
2 86241 1 15177
2 86242 1 15177
2 86243 1 15178
2 86244 1 15178
2 86245 1 15178
2 86246 1 15178
2 86247 1 15178
2 86248 1 15179
2 86249 1 15179
2 86250 1 15210
2 86251 1 15210
2 86252 1 15211
2 86253 1 15211
2 86254 1 15211
2 86255 1 15223
2 86256 1 15223
2 86257 1 15231
2 86258 1 15231
2 86259 1 15231
2 86260 1 15255
2 86261 1 15255
2 86262 1 15255
2 86263 1 15255
2 86264 1 15255
2 86265 1 15255
2 86266 1 15256
2 86267 1 15256
2 86268 1 15256
2 86269 1 15256
2 86270 1 15256
2 86271 1 15256
2 86272 1 15256
2 86273 1 15257
2 86274 1 15257
2 86275 1 15264
2 86276 1 15264
2 86277 1 15264
2 86278 1 15264
2 86279 1 15283
2 86280 1 15283
2 86281 1 15284
2 86282 1 15284
2 86283 1 15284
2 86284 1 15284
2 86285 1 15284
2 86286 1 15300
2 86287 1 15300
2 86288 1 15300
2 86289 1 15300
2 86290 1 15300
2 86291 1 15300
2 86292 1 15300
2 86293 1 15300
2 86294 1 15300
2 86295 1 15300
2 86296 1 15300
2 86297 1 15300
2 86298 1 15300
2 86299 1 15300
2 86300 1 15306
2 86301 1 15306
2 86302 1 15306
2 86303 1 15306
2 86304 1 15306
2 86305 1 15306
2 86306 1 15306
2 86307 1 15306
2 86308 1 15314
2 86309 1 15314
2 86310 1 15314
2 86311 1 15316
2 86312 1 15316
2 86313 1 15316
2 86314 1 15316
2 86315 1 15316
2 86316 1 15316
2 86317 1 15316
2 86318 1 15316
2 86319 1 15316
2 86320 1 15316
2 86321 1 15317
2 86322 1 15317
2 86323 1 15317
2 86324 1 15317
2 86325 1 15318
2 86326 1 15318
2 86327 1 15318
2 86328 1 15318
2 86329 1 15318
2 86330 1 15318
2 86331 1 15318
2 86332 1 15318
2 86333 1 15318
2 86334 1 15318
2 86335 1 15318
2 86336 1 15331
2 86337 1 15331
2 86338 1 15344
2 86339 1 15344
2 86340 1 15344
2 86341 1 15344
2 86342 1 15344
2 86343 1 15368
2 86344 1 15368
2 86345 1 15368
2 86346 1 15369
2 86347 1 15369
2 86348 1 15369
2 86349 1 15385
2 86350 1 15385
2 86351 1 15386
2 86352 1 15386
2 86353 1 15386
2 86354 1 15386
2 86355 1 15426
2 86356 1 15426
2 86357 1 15426
2 86358 1 15457
2 86359 1 15457
2 86360 1 15461
2 86361 1 15461
2 86362 1 15466
2 86363 1 15466
2 86364 1 15466
2 86365 1 15468
2 86366 1 15468
2 86367 1 15478
2 86368 1 15478
2 86369 1 15478
2 86370 1 15478
2 86371 1 15479
2 86372 1 15479
2 86373 1 15479
2 86374 1 15479
2 86375 1 15484
2 86376 1 15484
2 86377 1 15517
2 86378 1 15517
2 86379 1 15555
2 86380 1 15555
2 86381 1 15555
2 86382 1 15555
2 86383 1 15570
2 86384 1 15570
2 86385 1 15570
2 86386 1 15574
2 86387 1 15574
2 86388 1 15579
2 86389 1 15579
2 86390 1 15582
2 86391 1 15582
2 86392 1 15589
2 86393 1 15589
2 86394 1 15589
2 86395 1 15600
2 86396 1 15600
2 86397 1 15617
2 86398 1 15617
2 86399 1 15620
2 86400 1 15620
2 86401 1 15627
2 86402 1 15627
2 86403 1 15627
2 86404 1 15627
2 86405 1 15647
2 86406 1 15647
2 86407 1 15647
2 86408 1 15647
2 86409 1 15647
2 86410 1 15695
2 86411 1 15695
2 86412 1 15695
2 86413 1 15695
2 86414 1 15748
2 86415 1 15748
2 86416 1 15756
2 86417 1 15756
2 86418 1 15757
2 86419 1 15757
2 86420 1 15762
2 86421 1 15762
2 86422 1 15762
2 86423 1 15762
2 86424 1 15762
2 86425 1 15774
2 86426 1 15774
2 86427 1 15786
2 86428 1 15786
2 86429 1 15786
2 86430 1 15793
2 86431 1 15793
2 86432 1 15794
2 86433 1 15794
2 86434 1 15794
2 86435 1 15819
2 86436 1 15819
2 86437 1 15820
2 86438 1 15820
2 86439 1 15820
2 86440 1 15820
2 86441 1 15820
2 86442 1 15821
2 86443 1 15821
2 86444 1 15821
2 86445 1 15822
2 86446 1 15822
2 86447 1 15823
2 86448 1 15823
2 86449 1 15856
2 86450 1 15856
2 86451 1 15858
2 86452 1 15858
2 86453 1 15858
2 86454 1 15858
2 86455 1 15858
2 86456 1 15858
2 86457 1 15858
2 86458 1 15858
2 86459 1 15858
2 86460 1 15858
2 86461 1 15858
2 86462 1 15858
2 86463 1 15858
2 86464 1 15858
2 86465 1 15858
2 86466 1 15858
2 86467 1 15858
2 86468 1 15858
2 86469 1 15858
2 86470 1 15858
2 86471 1 15858
2 86472 1 15858
2 86473 1 15858
2 86474 1 15858
2 86475 1 15858
2 86476 1 15858
2 86477 1 15858
2 86478 1 15858
2 86479 1 15858
2 86480 1 15858
2 86481 1 15858
2 86482 1 15858
2 86483 1 15858
2 86484 1 15858
2 86485 1 15858
2 86486 1 15858
2 86487 1 15858
2 86488 1 15858
2 86489 1 15858
2 86490 1 15858
2 86491 1 15858
2 86492 1 15858
2 86493 1 15858
2 86494 1 15858
2 86495 1 15858
2 86496 1 15858
2 86497 1 15858
2 86498 1 15858
2 86499 1 15858
2 86500 1 15858
2 86501 1 15858
2 86502 1 15858
2 86503 1 15858
2 86504 1 15858
2 86505 1 15858
2 86506 1 15858
2 86507 1 15858
2 86508 1 15858
2 86509 1 15858
2 86510 1 15858
2 86511 1 15859
2 86512 1 15859
2 86513 1 15859
2 86514 1 15859
2 86515 1 15859
2 86516 1 15859
2 86517 1 15860
2 86518 1 15860
2 86519 1 15861
2 86520 1 15861
2 86521 1 15864
2 86522 1 15864
2 86523 1 15864
2 86524 1 15864
2 86525 1 15864
2 86526 1 15865
2 86527 1 15865
2 86528 1 15874
2 86529 1 15874
2 86530 1 15874
2 86531 1 15874
2 86532 1 15874
2 86533 1 15874
2 86534 1 15875
2 86535 1 15875
2 86536 1 15875
2 86537 1 15887
2 86538 1 15887
2 86539 1 15887
2 86540 1 15888
2 86541 1 15888
2 86542 1 15888
2 86543 1 15898
2 86544 1 15898
2 86545 1 15898
2 86546 1 15898
2 86547 1 15898
2 86548 1 15898
2 86549 1 15899
2 86550 1 15899
2 86551 1 15900
2 86552 1 15900
2 86553 1 15900
2 86554 1 15900
2 86555 1 15900
2 86556 1 15900
2 86557 1 15900
2 86558 1 15900
2 86559 1 15900
2 86560 1 15900
2 86561 1 15900
2 86562 1 15900
2 86563 1 15900
2 86564 1 15900
2 86565 1 15900
2 86566 1 15900
2 86567 1 15900
2 86568 1 15900
2 86569 1 15900
2 86570 1 15900
2 86571 1 15900
2 86572 1 15900
2 86573 1 15900
2 86574 1 15900
2 86575 1 15900
2 86576 1 15910
2 86577 1 15910
2 86578 1 15910
2 86579 1 15910
2 86580 1 15910
2 86581 1 15910
2 86582 1 15910
2 86583 1 15910
2 86584 1 15910
2 86585 1 15910
2 86586 1 15911
2 86587 1 15911
2 86588 1 15916
2 86589 1 15916
2 86590 1 15916
2 86591 1 15917
2 86592 1 15917
2 86593 1 15917
2 86594 1 15917
2 86595 1 15918
2 86596 1 15918
2 86597 1 15918
2 86598 1 15918
2 86599 1 15931
2 86600 1 15931
2 86601 1 15931
2 86602 1 15931
2 86603 1 15932
2 86604 1 15932
2 86605 1 15932
2 86606 1 15933
2 86607 1 15933
2 86608 1 15934
2 86609 1 15934
2 86610 1 15937
2 86611 1 15937
2 86612 1 15937
2 86613 1 15937
2 86614 1 15937
2 86615 1 15937
2 86616 1 15938
2 86617 1 15938
2 86618 1 15940
2 86619 1 15940
2 86620 1 15940
2 86621 1 15940
2 86622 1 15948
2 86623 1 15948
2 86624 1 15948
2 86625 1 15951
2 86626 1 15951
2 86627 1 15951
2 86628 1 15953
2 86629 1 15953
2 86630 1 15954
2 86631 1 15954
2 86632 1 15963
2 86633 1 15963
2 86634 1 15963
2 86635 1 15963
2 86636 1 15967
2 86637 1 15967
2 86638 1 15968
2 86639 1 15968
2 86640 1 15968
2 86641 1 15968
2 86642 1 15968
2 86643 1 15968
2 86644 1 15969
2 86645 1 15969
2 86646 1 15969
2 86647 1 15982
2 86648 1 15982
2 86649 1 15982
2 86650 1 15982
2 86651 1 15982
2 86652 1 15982
2 86653 1 15982
2 86654 1 15982
2 86655 1 15983
2 86656 1 15983
2 86657 1 15983
2 86658 1 15984
2 86659 1 15984
2 86660 1 15984
2 86661 1 15986
2 86662 1 15986
2 86663 1 15987
2 86664 1 15987
2 86665 1 15987
2 86666 1 15987
2 86667 1 15987
2 86668 1 15987
2 86669 1 15987
2 86670 1 15987
2 86671 1 15987
2 86672 1 15987
2 86673 1 15987
2 86674 1 15987
2 86675 1 15987
2 86676 1 15987
2 86677 1 15987
2 86678 1 15987
2 86679 1 15987
2 86680 1 15988
2 86681 1 15988
2 86682 1 15988
2 86683 1 15989
2 86684 1 15989
2 86685 1 15989
2 86686 1 16026
2 86687 1 16026
2 86688 1 16026
2 86689 1 16026
2 86690 1 16027
2 86691 1 16027
2 86692 1 16027
2 86693 1 16028
2 86694 1 16028
2 86695 1 16028
2 86696 1 16028
2 86697 1 16029
2 86698 1 16029
2 86699 1 16029
2 86700 1 16029
2 86701 1 16029
2 86702 1 16029
2 86703 1 16029
2 86704 1 16029
2 86705 1 16029
2 86706 1 16031
2 86707 1 16031
2 86708 1 16031
2 86709 1 16031
2 86710 1 16031
2 86711 1 16031
2 86712 1 16031
2 86713 1 16031
2 86714 1 16031
2 86715 1 16034
2 86716 1 16034
2 86717 1 16034
2 86718 1 16034
2 86719 1 16034
2 86720 1 16034
2 86721 1 16034
2 86722 1 16034
2 86723 1 16034
2 86724 1 16034
2 86725 1 16034
2 86726 1 16034
2 86727 1 16034
2 86728 1 16034
2 86729 1 16034
2 86730 1 16034
2 86731 1 16034
2 86732 1 16034
2 86733 1 16034
2 86734 1 16034
2 86735 1 16034
2 86736 1 16035
2 86737 1 16035
2 86738 1 16035
2 86739 1 16035
2 86740 1 16035
2 86741 1 16035
2 86742 1 16035
2 86743 1 16035
2 86744 1 16035
2 86745 1 16035
2 86746 1 16035
2 86747 1 16042
2 86748 1 16042
2 86749 1 16049
2 86750 1 16049
2 86751 1 16049
2 86752 1 16064
2 86753 1 16064
2 86754 1 16064
2 86755 1 16084
2 86756 1 16084
2 86757 1 16084
2 86758 1 16086
2 86759 1 16086
2 86760 1 16086
2 86761 1 16101
2 86762 1 16101
2 86763 1 16102
2 86764 1 16102
2 86765 1 16107
2 86766 1 16107
2 86767 1 16108
2 86768 1 16108
2 86769 1 16117
2 86770 1 16117
2 86771 1 16118
2 86772 1 16118
2 86773 1 16119
2 86774 1 16119
2 86775 1 16121
2 86776 1 16121
2 86777 1 16121
2 86778 1 16131
2 86779 1 16131
2 86780 1 16131
2 86781 1 16142
2 86782 1 16142
2 86783 1 16154
2 86784 1 16154
2 86785 1 16158
2 86786 1 16158
2 86787 1 16182
2 86788 1 16182
2 86789 1 16185
2 86790 1 16185
2 86791 1 16185
2 86792 1 16185
2 86793 1 16185
2 86794 1 16187
2 86795 1 16187
2 86796 1 16188
2 86797 1 16188
2 86798 1 16192
2 86799 1 16192
2 86800 1 16192
2 86801 1 16192
2 86802 1 16192
2 86803 1 16192
2 86804 1 16192
2 86805 1 16192
2 86806 1 16193
2 86807 1 16193
2 86808 1 16193
2 86809 1 16198
2 86810 1 16198
2 86811 1 16198
2 86812 1 16203
2 86813 1 16203
2 86814 1 16206
2 86815 1 16206
2 86816 1 16232
2 86817 1 16232
2 86818 1 16233
2 86819 1 16233
2 86820 1 16233
2 86821 1 16241
2 86822 1 16241
2 86823 1 16242
2 86824 1 16242
2 86825 1 16242
2 86826 1 16249
2 86827 1 16249
2 86828 1 16249
2 86829 1 16250
2 86830 1 16250
2 86831 1 16250
2 86832 1 16250
2 86833 1 16250
2 86834 1 16251
2 86835 1 16251
2 86836 1 16259
2 86837 1 16259
2 86838 1 16259
2 86839 1 16259
2 86840 1 16259
2 86841 1 16259
2 86842 1 16259
2 86843 1 16260
2 86844 1 16260
2 86845 1 16267
2 86846 1 16267
2 86847 1 16267
2 86848 1 16267
2 86849 1 16267
2 86850 1 16267
2 86851 1 16267
2 86852 1 16268
2 86853 1 16268
2 86854 1 16268
2 86855 1 16268
2 86856 1 16278
2 86857 1 16278
2 86858 1 16287
2 86859 1 16287
2 86860 1 16293
2 86861 1 16293
2 86862 1 16293
2 86863 1 16293
2 86864 1 16313
2 86865 1 16313
2 86866 1 16331
2 86867 1 16331
2 86868 1 16331
2 86869 1 16337
2 86870 1 16337
2 86871 1 16337
2 86872 1 16338
2 86873 1 16338
2 86874 1 16338
2 86875 1 16338
2 86876 1 16346
2 86877 1 16346
2 86878 1 16346
2 86879 1 16347
2 86880 1 16347
2 86881 1 16347
2 86882 1 16347
2 86883 1 16347
2 86884 1 16347
2 86885 1 16347
2 86886 1 16352
2 86887 1 16352
2 86888 1 16369
2 86889 1 16369
2 86890 1 16369
2 86891 1 16369
2 86892 1 16369
2 86893 1 16375
2 86894 1 16375
2 86895 1 16386
2 86896 1 16386
2 86897 1 16386
2 86898 1 16386
2 86899 1 16386
2 86900 1 16387
2 86901 1 16387
2 86902 1 16400
2 86903 1 16400
2 86904 1 16400
2 86905 1 16400
2 86906 1 16401
2 86907 1 16401
2 86908 1 16412
2 86909 1 16412
2 86910 1 16412
2 86911 1 16412
2 86912 1 16412
2 86913 1 16413
2 86914 1 16413
2 86915 1 16414
2 86916 1 16414
2 86917 1 16414
2 86918 1 16414
2 86919 1 16417
2 86920 1 16417
2 86921 1 16417
2 86922 1 16417
2 86923 1 16417
2 86924 1 16417
2 86925 1 16417
2 86926 1 16417
2 86927 1 16417
2 86928 1 16418
2 86929 1 16418
2 86930 1 16418
2 86931 1 16437
2 86932 1 16437
2 86933 1 16437
2 86934 1 16437
2 86935 1 16437
2 86936 1 16437
2 86937 1 16437
2 86938 1 16437
2 86939 1 16437
2 86940 1 16437
2 86941 1 16437
2 86942 1 16438
2 86943 1 16438
2 86944 1 16439
2 86945 1 16439
2 86946 1 16439
2 86947 1 16439
2 86948 1 16439
2 86949 1 16439
2 86950 1 16439
2 86951 1 16439
2 86952 1 16446
2 86953 1 16446
2 86954 1 16446
2 86955 1 16447
2 86956 1 16447
2 86957 1 16467
2 86958 1 16467
2 86959 1 16467
2 86960 1 16467
2 86961 1 16492
2 86962 1 16492
2 86963 1 16492
2 86964 1 16501
2 86965 1 16501
2 86966 1 16501
2 86967 1 16506
2 86968 1 16506
2 86969 1 16506
2 86970 1 16512
2 86971 1 16512
2 86972 1 16512
2 86973 1 16513
2 86974 1 16513
2 86975 1 16520
2 86976 1 16520
2 86977 1 16520
2 86978 1 16520
2 86979 1 16521
2 86980 1 16521
2 86981 1 16521
2 86982 1 16523
2 86983 1 16523
2 86984 1 16540
2 86985 1 16540
2 86986 1 16540
2 86987 1 16540
2 86988 1 16541
2 86989 1 16541
2 86990 1 16541
2 86991 1 16541
2 86992 1 16542
2 86993 1 16542
2 86994 1 16542
2 86995 1 16542
2 86996 1 16542
2 86997 1 16542
2 86998 1 16542
2 86999 1 16542
2 87000 1 16542
2 87001 1 16542
2 87002 1 16542
2 87003 1 16559
2 87004 1 16559
2 87005 1 16559
2 87006 1 16559
2 87007 1 16565
2 87008 1 16565
2 87009 1 16565
2 87010 1 16565
2 87011 1 16597
2 87012 1 16597
2 87013 1 16597
2 87014 1 16597
2 87015 1 16597
2 87016 1 16597
2 87017 1 16597
2 87018 1 16597
2 87019 1 16597
2 87020 1 16597
2 87021 1 16598
2 87022 1 16598
2 87023 1 16599
2 87024 1 16599
2 87025 1 16599
2 87026 1 16599
2 87027 1 16600
2 87028 1 16600
2 87029 1 16604
2 87030 1 16604
2 87031 1 16604
2 87032 1 16606
2 87033 1 16606
2 87034 1 16616
2 87035 1 16616
2 87036 1 16617
2 87037 1 16617
2 87038 1 16649
2 87039 1 16649
2 87040 1 16651
2 87041 1 16651
2 87042 1 16678
2 87043 1 16678
2 87044 1 16678
2 87045 1 16685
2 87046 1 16685
2 87047 1 16685
2 87048 1 16695
2 87049 1 16695
2 87050 1 16695
2 87051 1 16713
2 87052 1 16713
2 87053 1 16714
2 87054 1 16714
2 87055 1 16724
2 87056 1 16724
2 87057 1 16724
2 87058 1 16734
2 87059 1 16734
2 87060 1 16734
2 87061 1 16735
2 87062 1 16735
2 87063 1 16736
2 87064 1 16736
2 87065 1 16762
2 87066 1 16762
2 87067 1 16769
2 87068 1 16769
2 87069 1 16769
2 87070 1 16769
2 87071 1 16770
2 87072 1 16770
2 87073 1 16778
2 87074 1 16778
2 87075 1 16779
2 87076 1 16779
2 87077 1 16832
2 87078 1 16832
2 87079 1 16840
2 87080 1 16840
2 87081 1 16847
2 87082 1 16847
2 87083 1 16859
2 87084 1 16859
2 87085 1 16859
2 87086 1 16859
2 87087 1 16861
2 87088 1 16861
2 87089 1 16867
2 87090 1 16867
2 87091 1 16867
2 87092 1 16880
2 87093 1 16880
2 87094 1 16880
2 87095 1 16880
2 87096 1 16881
2 87097 1 16881
2 87098 1 16881
2 87099 1 16881
2 87100 1 16881
2 87101 1 16911
2 87102 1 16911
2 87103 1 16920
2 87104 1 16920
2 87105 1 16949
2 87106 1 16949
2 87107 1 16949
2 87108 1 16949
2 87109 1 16950
2 87110 1 16950
2 87111 1 16976
2 87112 1 16976
2 87113 1 16981
2 87114 1 16981
2 87115 1 16981
2 87116 1 16981
2 87117 1 16981
2 87118 1 16981
2 87119 1 16981
2 87120 1 16981
2 87121 1 16993
2 87122 1 16993
2 87123 1 16993
2 87124 1 17034
2 87125 1 17034
2 87126 1 17034
2 87127 1 17035
2 87128 1 17035
2 87129 1 17037
2 87130 1 17037
2 87131 1 17037
2 87132 1 17040
2 87133 1 17040
2 87134 1 17045
2 87135 1 17045
2 87136 1 17045
2 87137 1 17045
2 87138 1 17045
2 87139 1 17045
2 87140 1 17045
2 87141 1 17045
2 87142 1 17046
2 87143 1 17046
2 87144 1 17046
2 87145 1 17047
2 87146 1 17047
2 87147 1 17047
2 87148 1 17069
2 87149 1 17069
2 87150 1 17069
2 87151 1 17069
2 87152 1 17069
2 87153 1 17069
2 87154 1 17069
2 87155 1 17091
2 87156 1 17091
2 87157 1 17093
2 87158 1 17093
2 87159 1 17110
2 87160 1 17110
2 87161 1 17110
2 87162 1 17112
2 87163 1 17112
2 87164 1 17112
2 87165 1 17113
2 87166 1 17113
2 87167 1 17113
2 87168 1 17113
2 87169 1 17113
2 87170 1 17115
2 87171 1 17115
2 87172 1 17115
2 87173 1 17115
2 87174 1 17115
2 87175 1 17118
2 87176 1 17118
2 87177 1 17124
2 87178 1 17124
2 87179 1 17124
2 87180 1 17124
2 87181 1 17124
2 87182 1 17124
2 87183 1 17124
2 87184 1 17124
2 87185 1 17124
2 87186 1 17124
2 87187 1 17124
2 87188 1 17125
2 87189 1 17125
2 87190 1 17125
2 87191 1 17133
2 87192 1 17133
2 87193 1 17134
2 87194 1 17134
2 87195 1 17143
2 87196 1 17143
2 87197 1 17143
2 87198 1 17143
2 87199 1 17143
2 87200 1 17143
2 87201 1 17143
2 87202 1 17143
2 87203 1 17143
2 87204 1 17143
2 87205 1 17143
2 87206 1 17143
2 87207 1 17143
2 87208 1 17143
2 87209 1 17143
2 87210 1 17143
2 87211 1 17143
2 87212 1 17143
2 87213 1 17144
2 87214 1 17144
2 87215 1 17144
2 87216 1 17144
2 87217 1 17144
2 87218 1 17144
2 87219 1 17145
2 87220 1 17145
2 87221 1 17146
2 87222 1 17146
2 87223 1 17146
2 87224 1 17146
2 87225 1 17147
2 87226 1 17147
2 87227 1 17147
2 87228 1 17147
2 87229 1 17148
2 87230 1 17148
2 87231 1 17154
2 87232 1 17154
2 87233 1 17154
2 87234 1 17154
2 87235 1 17154
2 87236 1 17154
2 87237 1 17154
2 87238 1 17154
2 87239 1 17154
2 87240 1 17154
2 87241 1 17155
2 87242 1 17155
2 87243 1 17167
2 87244 1 17167
2 87245 1 17183
2 87246 1 17183
2 87247 1 17183
2 87248 1 17183
2 87249 1 17184
2 87250 1 17184
2 87251 1 17195
2 87252 1 17195
2 87253 1 17214
2 87254 1 17214
2 87255 1 17214
2 87256 1 17214
2 87257 1 17214
2 87258 1 17214
2 87259 1 17214
2 87260 1 17214
2 87261 1 17214
2 87262 1 17214
2 87263 1 17214
2 87264 1 17214
2 87265 1 17214
2 87266 1 17214
2 87267 1 17214
2 87268 1 17214
2 87269 1 17214
2 87270 1 17214
2 87271 1 17214
2 87272 1 17214
2 87273 1 17214
2 87274 1 17214
2 87275 1 17215
2 87276 1 17215
2 87277 1 17220
2 87278 1 17220
2 87279 1 17220
2 87280 1 17225
2 87281 1 17225
2 87282 1 17242
2 87283 1 17242
2 87284 1 17245
2 87285 1 17245
2 87286 1 17245
2 87287 1 17245
2 87288 1 17245
2 87289 1 17269
2 87290 1 17269
2 87291 1 17270
2 87292 1 17270
2 87293 1 17278
2 87294 1 17278
2 87295 1 17300
2 87296 1 17300
2 87297 1 17301
2 87298 1 17301
2 87299 1 17302
2 87300 1 17302
2 87301 1 17303
2 87302 1 17303
2 87303 1 17303
2 87304 1 17308
2 87305 1 17308
2 87306 1 17322
2 87307 1 17322
2 87308 1 17322
2 87309 1 17326
2 87310 1 17326
2 87311 1 17333
2 87312 1 17333
2 87313 1 17334
2 87314 1 17334
2 87315 1 17334
2 87316 1 17334
2 87317 1 17335
2 87318 1 17335
2 87319 1 17341
2 87320 1 17341
2 87321 1 17341
2 87322 1 17341
2 87323 1 17352
2 87324 1 17352
2 87325 1 17352
2 87326 1 17354
2 87327 1 17354
2 87328 1 17360
2 87329 1 17360
2 87330 1 17361
2 87331 1 17361
2 87332 1 17361
2 87333 1 17361
2 87334 1 17376
2 87335 1 17376
2 87336 1 17376
2 87337 1 17376
2 87338 1 17376
2 87339 1 17376
2 87340 1 17376
2 87341 1 17376
2 87342 1 17376
2 87343 1 17376
2 87344 1 17376
2 87345 1 17376
2 87346 1 17376
2 87347 1 17376
2 87348 1 17377
2 87349 1 17377
2 87350 1 17379
2 87351 1 17379
2 87352 1 17379
2 87353 1 17380
2 87354 1 17380
2 87355 1 17383
2 87356 1 17383
2 87357 1 17384
2 87358 1 17384
2 87359 1 17395
2 87360 1 17395
2 87361 1 17424
2 87362 1 17424
2 87363 1 17446
2 87364 1 17446
2 87365 1 17449
2 87366 1 17449
2 87367 1 17449
2 87368 1 17452
2 87369 1 17452
2 87370 1 17452
2 87371 1 17453
2 87372 1 17453
2 87373 1 17453
2 87374 1 17461
2 87375 1 17461
2 87376 1 17461
2 87377 1 17462
2 87378 1 17462
2 87379 1 17469
2 87380 1 17469
2 87381 1 17475
2 87382 1 17475
2 87383 1 17475
2 87384 1 17475
2 87385 1 17476
2 87386 1 17476
2 87387 1 17476
2 87388 1 17495
2 87389 1 17495
2 87390 1 17508
2 87391 1 17508
2 87392 1 17508
2 87393 1 17509
2 87394 1 17509
2 87395 1 17510
2 87396 1 17510
2 87397 1 17511
2 87398 1 17511
2 87399 1 17547
2 87400 1 17547
2 87401 1 17560
2 87402 1 17560
2 87403 1 17571
2 87404 1 17571
2 87405 1 17584
2 87406 1 17584
2 87407 1 17585
2 87408 1 17585
2 87409 1 17586
2 87410 1 17586
2 87411 1 17587
2 87412 1 17587
2 87413 1 17590
2 87414 1 17590
2 87415 1 17609
2 87416 1 17609
2 87417 1 17623
2 87418 1 17623
2 87419 1 17623
2 87420 1 17623
2 87421 1 17624
2 87422 1 17624
2 87423 1 17653
2 87424 1 17653
2 87425 1 17665
2 87426 1 17665
2 87427 1 17665
2 87428 1 17665
2 87429 1 17665
2 87430 1 17666
2 87431 1 17666
2 87432 1 17666
2 87433 1 17666
2 87434 1 17666
2 87435 1 17682
2 87436 1 17682
2 87437 1 17683
2 87438 1 17683
2 87439 1 17685
2 87440 1 17685
2 87441 1 17688
2 87442 1 17688
2 87443 1 17688
2 87444 1 17688
2 87445 1 17688
2 87446 1 17688
2 87447 1 17688
2 87448 1 17688
2 87449 1 17689
2 87450 1 17689
2 87451 1 17696
2 87452 1 17696
2 87453 1 17696
2 87454 1 17696
2 87455 1 17696
2 87456 1 17696
2 87457 1 17697
2 87458 1 17697
2 87459 1 17697
2 87460 1 17704
2 87461 1 17704
2 87462 1 17704
2 87463 1 17704
2 87464 1 17704
2 87465 1 17704
2 87466 1 17704
2 87467 1 17704
2 87468 1 17705
2 87469 1 17705
2 87470 1 17713
2 87471 1 17713
2 87472 1 17715
2 87473 1 17715
2 87474 1 17719
2 87475 1 17719
2 87476 1 17719
2 87477 1 17719
2 87478 1 17719
2 87479 1 17719
2 87480 1 17719
2 87481 1 17724
2 87482 1 17724
2 87483 1 17728
2 87484 1 17728
2 87485 1 17728
2 87486 1 17728
2 87487 1 17728
2 87488 1 17728
2 87489 1 17728
2 87490 1 17740
2 87491 1 17740
2 87492 1 17751
2 87493 1 17751
2 87494 1 17755
2 87495 1 17755
2 87496 1 17755
2 87497 1 17755
2 87498 1 17755
2 87499 1 17755
2 87500 1 17755
2 87501 1 17755
2 87502 1 17755
2 87503 1 17755
2 87504 1 17755
2 87505 1 17755
2 87506 1 17755
2 87507 1 17755
2 87508 1 17779
2 87509 1 17779
2 87510 1 17781
2 87511 1 17781
2 87512 1 17787
2 87513 1 17787
2 87514 1 17787
2 87515 1 17787
2 87516 1 17788
2 87517 1 17788
2 87518 1 17802
2 87519 1 17802
2 87520 1 17810
2 87521 1 17810
2 87522 1 17810
2 87523 1 17821
2 87524 1 17821
2 87525 1 17830
2 87526 1 17830
2 87527 1 17849
2 87528 1 17849
2 87529 1 17849
2 87530 1 17849
2 87531 1 17849
2 87532 1 17849
2 87533 1 17849
2 87534 1 17849
2 87535 1 17849
2 87536 1 17849
2 87537 1 17849
2 87538 1 17849
2 87539 1 17849
2 87540 1 17849
2 87541 1 17849
2 87542 1 17849
2 87543 1 17850
2 87544 1 17850
2 87545 1 17850
2 87546 1 17859
2 87547 1 17859
2 87548 1 17859
2 87549 1 17859
2 87550 1 17859
2 87551 1 17859
2 87552 1 17859
2 87553 1 17859
2 87554 1 17859
2 87555 1 17859
2 87556 1 17859
2 87557 1 17859
2 87558 1 17859
2 87559 1 17860
2 87560 1 17860
2 87561 1 17860
2 87562 1 17860
2 87563 1 17860
2 87564 1 17860
2 87565 1 17860
2 87566 1 17860
2 87567 1 17861
2 87568 1 17861
2 87569 1 17866
2 87570 1 17866
2 87571 1 17888
2 87572 1 17888
2 87573 1 17891
2 87574 1 17891
2 87575 1 17901
2 87576 1 17901
2 87577 1 17901
2 87578 1 17901
2 87579 1 17901
2 87580 1 17901
2 87581 1 17901
2 87582 1 17901
2 87583 1 17901
2 87584 1 17922
2 87585 1 17922
2 87586 1 17929
2 87587 1 17929
2 87588 1 17937
2 87589 1 17937
2 87590 1 17941
2 87591 1 17941
2 87592 1 17961
2 87593 1 17961
2 87594 1 17961
2 87595 1 17961
2 87596 1 17962
2 87597 1 17962
2 87598 1 17986
2 87599 1 17986
2 87600 1 17987
2 87601 1 17987
2 87602 1 18026
2 87603 1 18026
2 87604 1 18026
2 87605 1 18026
2 87606 1 18027
2 87607 1 18027
2 87608 1 18027
2 87609 1 18027
2 87610 1 18027
2 87611 1 18027
2 87612 1 18028
2 87613 1 18028
2 87614 1 18030
2 87615 1 18030
2 87616 1 18030
2 87617 1 18030
2 87618 1 18038
2 87619 1 18038
2 87620 1 18040
2 87621 1 18040
2 87622 1 18046
2 87623 1 18046
2 87624 1 18046
2 87625 1 18046
2 87626 1 18046
2 87627 1 18046
2 87628 1 18046
2 87629 1 18046
2 87630 1 18046
2 87631 1 18046
2 87632 1 18047
2 87633 1 18047
2 87634 1 18047
2 87635 1 18047
2 87636 1 18048
2 87637 1 18048
2 87638 1 18048
2 87639 1 18048
2 87640 1 18048
2 87641 1 18048
2 87642 1 18048
2 87643 1 18049
2 87644 1 18049
2 87645 1 18051
2 87646 1 18051
2 87647 1 18051
2 87648 1 18051
2 87649 1 18051
2 87650 1 18052
2 87651 1 18052
2 87652 1 18053
2 87653 1 18053
2 87654 1 18060
2 87655 1 18060
2 87656 1 18060
2 87657 1 18073
2 87658 1 18073
2 87659 1 18073
2 87660 1 18073
2 87661 1 18073
2 87662 1 18073
2 87663 1 18073
2 87664 1 18081
2 87665 1 18081
2 87666 1 18081
2 87667 1 18081
2 87668 1 18081
2 87669 1 18089
2 87670 1 18089
2 87671 1 18089
2 87672 1 18089
2 87673 1 18098
2 87674 1 18098
2 87675 1 18098
2 87676 1 18098
2 87677 1 18098
2 87678 1 18099
2 87679 1 18099
2 87680 1 18099
2 87681 1 18113
2 87682 1 18113
2 87683 1 18113
2 87684 1 18121
2 87685 1 18121
2 87686 1 18121
2 87687 1 18121
2 87688 1 18121
2 87689 1 18121
2 87690 1 18147
2 87691 1 18147
2 87692 1 18147
2 87693 1 18148
2 87694 1 18148
2 87695 1 18148
2 87696 1 18194
2 87697 1 18194
2 87698 1 18194
2 87699 1 18195
2 87700 1 18195
2 87701 1 18195
2 87702 1 18196
2 87703 1 18196
2 87704 1 18197
2 87705 1 18197
2 87706 1 18197
2 87707 1 18198
2 87708 1 18198
2 87709 1 18208
2 87710 1 18208
2 87711 1 18208
2 87712 1 18208
2 87713 1 18208
2 87714 1 18210
2 87715 1 18210
2 87716 1 18224
2 87717 1 18224
2 87718 1 18260
2 87719 1 18260
2 87720 1 18276
2 87721 1 18276
2 87722 1 18276
2 87723 1 18277
2 87724 1 18277
2 87725 1 18277
2 87726 1 18281
2 87727 1 18281
2 87728 1 18281
2 87729 1 18281
2 87730 1 18281
2 87731 1 18281
2 87732 1 18281
2 87733 1 18281
2 87734 1 18282
2 87735 1 18282
2 87736 1 18282
2 87737 1 18284
2 87738 1 18284
2 87739 1 18284
2 87740 1 18292
2 87741 1 18292
2 87742 1 18308
2 87743 1 18308
2 87744 1 18308
2 87745 1 18309
2 87746 1 18309
2 87747 1 18312
2 87748 1 18312
2 87749 1 18335
2 87750 1 18335
2 87751 1 18335
2 87752 1 18386
2 87753 1 18386
2 87754 1 18386
2 87755 1 18386
2 87756 1 18387
2 87757 1 18387
2 87758 1 18388
2 87759 1 18388
2 87760 1 18388
2 87761 1 18388
2 87762 1 18388
2 87763 1 18412
2 87764 1 18412
2 87765 1 18413
2 87766 1 18413
2 87767 1 18446
2 87768 1 18446
2 87769 1 18446
2 87770 1 18446
2 87771 1 18446
2 87772 1 18448
2 87773 1 18448
2 87774 1 18454
2 87775 1 18454
2 87776 1 18454
2 87777 1 18462
2 87778 1 18462
2 87779 1 18466
2 87780 1 18466
2 87781 1 18466
2 87782 1 18466
2 87783 1 18469
2 87784 1 18469
2 87785 1 18469
2 87786 1 18469
2 87787 1 18469
2 87788 1 18470
2 87789 1 18470
2 87790 1 18470
2 87791 1 18507
2 87792 1 18507
2 87793 1 18507
2 87794 1 18507
2 87795 1 18507
2 87796 1 18507
2 87797 1 18508
2 87798 1 18508
2 87799 1 18508
2 87800 1 18508
2 87801 1 18515
2 87802 1 18515
2 87803 1 18523
2 87804 1 18523
2 87805 1 18523
2 87806 1 18524
2 87807 1 18524
2 87808 1 18524
2 87809 1 18538
2 87810 1 18538
2 87811 1 18538
2 87812 1 18538
2 87813 1 18538
2 87814 1 18538
2 87815 1 18538
2 87816 1 18542
2 87817 1 18542
2 87818 1 18555
2 87819 1 18555
2 87820 1 18556
2 87821 1 18556
2 87822 1 18556
2 87823 1 18556
2 87824 1 18561
2 87825 1 18561
2 87826 1 18561
2 87827 1 18561
2 87828 1 18561
2 87829 1 18561
2 87830 1 18561
2 87831 1 18564
2 87832 1 18564
2 87833 1 18572
2 87834 1 18572
2 87835 1 18572
2 87836 1 18572
2 87837 1 18572
2 87838 1 18572
2 87839 1 18573
2 87840 1 18573
2 87841 1 18575
2 87842 1 18575
2 87843 1 18582
2 87844 1 18582
2 87845 1 18582
2 87846 1 18582
2 87847 1 18582
2 87848 1 18582
2 87849 1 18583
2 87850 1 18583
2 87851 1 18583
2 87852 1 18585
2 87853 1 18585
2 87854 1 18586
2 87855 1 18586
2 87856 1 18586
2 87857 1 18586
2 87858 1 18586
2 87859 1 18587
2 87860 1 18587
2 87861 1 18587
2 87862 1 18587
2 87863 1 18587
2 87864 1 18587
2 87865 1 18589
2 87866 1 18589
2 87867 1 18596
2 87868 1 18596
2 87869 1 18596
2 87870 1 18597
2 87871 1 18597
2 87872 1 18598
2 87873 1 18598
2 87874 1 18598
2 87875 1 18598
2 87876 1 18598
2 87877 1 18598
2 87878 1 18615
2 87879 1 18615
2 87880 1 18615
2 87881 1 18615
2 87882 1 18620
2 87883 1 18620
2 87884 1 18620
2 87885 1 18620
2 87886 1 18620
2 87887 1 18625
2 87888 1 18625
2 87889 1 18625
2 87890 1 18625
2 87891 1 18625
2 87892 1 18630
2 87893 1 18630
2 87894 1 18630
2 87895 1 18641
2 87896 1 18641
2 87897 1 18641
2 87898 1 18641
2 87899 1 18649
2 87900 1 18649
2 87901 1 18649
2 87902 1 18649
2 87903 1 18649
2 87904 1 18649
2 87905 1 18650
2 87906 1 18650
2 87907 1 18659
2 87908 1 18659
2 87909 1 18660
2 87910 1 18660
2 87911 1 18660
2 87912 1 18660
2 87913 1 18660
2 87914 1 18660
2 87915 1 18660
2 87916 1 18660
2 87917 1 18661
2 87918 1 18661
2 87919 1 18662
2 87920 1 18662
2 87921 1 18662
2 87922 1 18662
2 87923 1 18662
2 87924 1 18663
2 87925 1 18663
2 87926 1 18664
2 87927 1 18664
2 87928 1 18664
2 87929 1 18677
2 87930 1 18677
2 87931 1 18677
2 87932 1 18678
2 87933 1 18678
2 87934 1 18678
2 87935 1 18678
2 87936 1 18678
2 87937 1 18678
2 87938 1 18678
2 87939 1 18678
2 87940 1 18678
2 87941 1 18678
2 87942 1 18678
2 87943 1 18678
2 87944 1 18678
2 87945 1 18678
2 87946 1 18679
2 87947 1 18679
2 87948 1 18680
2 87949 1 18680
2 87950 1 18681
2 87951 1 18681
2 87952 1 18681
2 87953 1 18683
2 87954 1 18683
2 87955 1 18683
2 87956 1 18708
2 87957 1 18708
2 87958 1 18716
2 87959 1 18716
2 87960 1 18716
2 87961 1 18716
2 87962 1 18726
2 87963 1 18726
2 87964 1 18726
2 87965 1 18726
2 87966 1 18726
2 87967 1 18745
2 87968 1 18745
2 87969 1 18745
2 87970 1 18745
2 87971 1 18746
2 87972 1 18746
2 87973 1 18768
2 87974 1 18768
2 87975 1 18768
2 87976 1 18776
2 87977 1 18776
2 87978 1 18779
2 87979 1 18779
2 87980 1 18779
2 87981 1 18780
2 87982 1 18780
2 87983 1 18780
2 87984 1 18780
2 87985 1 18781
2 87986 1 18781
2 87987 1 18788
2 87988 1 18788
2 87989 1 18789
2 87990 1 18789
2 87991 1 18789
2 87992 1 18789
2 87993 1 18789
2 87994 1 18789
2 87995 1 18789
2 87996 1 18789
2 87997 1 18789
2 87998 1 18789
2 87999 1 18789
2 88000 1 18791
2 88001 1 18791
2 88002 1 18832
2 88003 1 18832
2 88004 1 18832
2 88005 1 18832
2 88006 1 18832
2 88007 1 18832
2 88008 1 18832
2 88009 1 18832
2 88010 1 18832
2 88011 1 18832
2 88012 1 18832
2 88013 1 18832
2 88014 1 18832
2 88015 1 18832
2 88016 1 18832
2 88017 1 18832
2 88018 1 18832
2 88019 1 18833
2 88020 1 18833
2 88021 1 18833
2 88022 1 18834
2 88023 1 18834
2 88024 1 18834
2 88025 1 18834
2 88026 1 18835
2 88027 1 18835
2 88028 1 18835
2 88029 1 18836
2 88030 1 18836
2 88031 1 18836
2 88032 1 18837
2 88033 1 18837
2 88034 1 18848
2 88035 1 18848
2 88036 1 18848
2 88037 1 18848
2 88038 1 18849
2 88039 1 18849
2 88040 1 18849
2 88041 1 18851
2 88042 1 18851
2 88043 1 18851
2 88044 1 18851
2 88045 1 18851
2 88046 1 18851
2 88047 1 18851
2 88048 1 18851
2 88049 1 18851
2 88050 1 18851
2 88051 1 18853
2 88052 1 18853
2 88053 1 18854
2 88054 1 18854
2 88055 1 18855
2 88056 1 18855
2 88057 1 18857
2 88058 1 18857
2 88059 1 18859
2 88060 1 18859
2 88061 1 18859
2 88062 1 18873
2 88063 1 18873
2 88064 1 18874
2 88065 1 18874
2 88066 1 18876
2 88067 1 18876
2 88068 1 18883
2 88069 1 18883
2 88070 1 18884
2 88071 1 18884
2 88072 1 18884
2 88073 1 18884
2 88074 1 18888
2 88075 1 18888
2 88076 1 18898
2 88077 1 18898
2 88078 1 18899
2 88079 1 18899
2 88080 1 18899
2 88081 1 18899
2 88082 1 18899
2 88083 1 18901
2 88084 1 18901
2 88085 1 18901
2 88086 1 18909
2 88087 1 18909
2 88088 1 18909
2 88089 1 18909
2 88090 1 18909
2 88091 1 18910
2 88092 1 18910
2 88093 1 18910
2 88094 1 18910
2 88095 1 18910
2 88096 1 18910
2 88097 1 18912
2 88098 1 18912
2 88099 1 18912
2 88100 1 18920
2 88101 1 18920
2 88102 1 18920
2 88103 1 18920
2 88104 1 18936
2 88105 1 18936
2 88106 1 18936
2 88107 1 18940
2 88108 1 18940
2 88109 1 18940
2 88110 1 18940
2 88111 1 18940
2 88112 1 18940
2 88113 1 18941
2 88114 1 18941
2 88115 1 18965
2 88116 1 18965
2 88117 1 18981
2 88118 1 18981
2 88119 1 18981
2 88120 1 18981
2 88121 1 18981
2 88122 1 18981
2 88123 1 18981
2 88124 1 18981
2 88125 1 18981
2 88126 1 18981
2 88127 1 18981
2 88128 1 18981
2 88129 1 18981
2 88130 1 18981
2 88131 1 18981
2 88132 1 18981
2 88133 1 18981
2 88134 1 18981
2 88135 1 18981
2 88136 1 18981
2 88137 1 18982
2 88138 1 18982
2 88139 1 18982
2 88140 1 18982
2 88141 1 18983
2 88142 1 18983
2 88143 1 18983
2 88144 1 18983
2 88145 1 18983
2 88146 1 18983
2 88147 1 18983
2 88148 1 18983
2 88149 1 18983
2 88150 1 18983
2 88151 1 18983
2 88152 1 18983
2 88153 1 18983
2 88154 1 18983
2 88155 1 18991
2 88156 1 18991
2 88157 1 18997
2 88158 1 18997
2 88159 1 19000
2 88160 1 19000
2 88161 1 19000
2 88162 1 19004
2 88163 1 19004
2 88164 1 19005
2 88165 1 19005
2 88166 1 19005
2 88167 1 19005
2 88168 1 19012
2 88169 1 19012
2 88170 1 19013
2 88171 1 19013
2 88172 1 19028
2 88173 1 19028
2 88174 1 19029
2 88175 1 19029
2 88176 1 19032
2 88177 1 19032
2 88178 1 19032
2 88179 1 19032
2 88180 1 19032
2 88181 1 19037
2 88182 1 19037
2 88183 1 19039
2 88184 1 19039
2 88185 1 19039
2 88186 1 19039
2 88187 1 19039
2 88188 1 19039
2 88189 1 19039
2 88190 1 19043
2 88191 1 19043
2 88192 1 19044
2 88193 1 19044
2 88194 1 19044
2 88195 1 19044
2 88196 1 19054
2 88197 1 19054
2 88198 1 19073
2 88199 1 19073
2 88200 1 19073
2 88201 1 19073
2 88202 1 19074
2 88203 1 19074
2 88204 1 19082
2 88205 1 19082
2 88206 1 19083
2 88207 1 19083
2 88208 1 19083
2 88209 1 19083
2 88210 1 19085
2 88211 1 19085
2 88212 1 19085
2 88213 1 19097
2 88214 1 19097
2 88215 1 19097
2 88216 1 19097
2 88217 1 19111
2 88218 1 19111
2 88219 1 19119
2 88220 1 19119
2 88221 1 19119
2 88222 1 19119
2 88223 1 19119
2 88224 1 19123
2 88225 1 19123
2 88226 1 19123
2 88227 1 19123
2 88228 1 19135
2 88229 1 19135
2 88230 1 19142
2 88231 1 19142
2 88232 1 19148
2 88233 1 19148
2 88234 1 19149
2 88235 1 19149
2 88236 1 19151
2 88237 1 19151
2 88238 1 19151
2 88239 1 19151
2 88240 1 19151
2 88241 1 19151
2 88242 1 19151
2 88243 1 19151
2 88244 1 19151
2 88245 1 19151
2 88246 1 19151
2 88247 1 19151
2 88248 1 19151
2 88249 1 19151
2 88250 1 19151
2 88251 1 19151
2 88252 1 19151
2 88253 1 19152
2 88254 1 19152
2 88255 1 19166
2 88256 1 19166
2 88257 1 19166
2 88258 1 19166
2 88259 1 19166
2 88260 1 19167
2 88261 1 19167
2 88262 1 19177
2 88263 1 19177
2 88264 1 19177
2 88265 1 19177
2 88266 1 19177
2 88267 1 19177
2 88268 1 19177
2 88269 1 19177
2 88270 1 19177
2 88271 1 19177
2 88272 1 19177
2 88273 1 19177
2 88274 1 19177
2 88275 1 19177
2 88276 1 19177
2 88277 1 19178
2 88278 1 19178
2 88279 1 19178
2 88280 1 19178
2 88281 1 19178
2 88282 1 19191
2 88283 1 19191
2 88284 1 19191
2 88285 1 19191
2 88286 1 19191
2 88287 1 19204
2 88288 1 19204
2 88289 1 19204
2 88290 1 19204
2 88291 1 19209
2 88292 1 19209
2 88293 1 19216
2 88294 1 19216
2 88295 1 19223
2 88296 1 19223
2 88297 1 19223
2 88298 1 19223
2 88299 1 19223
2 88300 1 19223
2 88301 1 19223
2 88302 1 19223
2 88303 1 19223
2 88304 1 19223
2 88305 1 19223
2 88306 1 19223
2 88307 1 19223
2 88308 1 19223
2 88309 1 19223
2 88310 1 19223
2 88311 1 19223
2 88312 1 19223
2 88313 1 19223
2 88314 1 19223
2 88315 1 19224
2 88316 1 19224
2 88317 1 19224
2 88318 1 19224
2 88319 1 19225
2 88320 1 19225
2 88321 1 19225
2 88322 1 19225
2 88323 1 19225
2 88324 1 19225
2 88325 1 19225
2 88326 1 19225
2 88327 1 19225
2 88328 1 19225
2 88329 1 19225
2 88330 1 19225
2 88331 1 19225
2 88332 1 19225
2 88333 1 19225
2 88334 1 19225
2 88335 1 19225
2 88336 1 19225
2 88337 1 19225
2 88338 1 19225
2 88339 1 19225
2 88340 1 19225
2 88341 1 19225
2 88342 1 19225
2 88343 1 19225
2 88344 1 19225
2 88345 1 19227
2 88346 1 19227
2 88347 1 19230
2 88348 1 19230
2 88349 1 19230
2 88350 1 19230
2 88351 1 19230
2 88352 1 19230
2 88353 1 19230
2 88354 1 19230
2 88355 1 19230
2 88356 1 19230
2 88357 1 19230
2 88358 1 19230
2 88359 1 19230
2 88360 1 19230
2 88361 1 19230
2 88362 1 19230
2 88363 1 19230
2 88364 1 19230
2 88365 1 19230
2 88366 1 19230
2 88367 1 19230
2 88368 1 19230
2 88369 1 19231
2 88370 1 19231
2 88371 1 19231
2 88372 1 19231
2 88373 1 19231
2 88374 1 19231
2 88375 1 19231
2 88376 1 19231
2 88377 1 19231
2 88378 1 19231
2 88379 1 19231
2 88380 1 19231
2 88381 1 19267
2 88382 1 19267
2 88383 1 19267
2 88384 1 19267
2 88385 1 19267
2 88386 1 19267
2 88387 1 19267
2 88388 1 19267
2 88389 1 19267
2 88390 1 19267
2 88391 1 19267
2 88392 1 19267
2 88393 1 19281
2 88394 1 19281
2 88395 1 19281
2 88396 1 19281
2 88397 1 19281
2 88398 1 19281
2 88399 1 19281
2 88400 1 19281
2 88401 1 19281
2 88402 1 19282
2 88403 1 19282
2 88404 1 19282
2 88405 1 19282
2 88406 1 19282
2 88407 1 19282
2 88408 1 19282
2 88409 1 19290
2 88410 1 19290
2 88411 1 19291
2 88412 1 19291
2 88413 1 19295
2 88414 1 19295
2 88415 1 19295
2 88416 1 19295
2 88417 1 19312
2 88418 1 19312
2 88419 1 19316
2 88420 1 19316
2 88421 1 19317
2 88422 1 19317
2 88423 1 19319
2 88424 1 19319
2 88425 1 19336
2 88426 1 19336
2 88427 1 19340
2 88428 1 19340
2 88429 1 19340
2 88430 1 19340
2 88431 1 19340
2 88432 1 19340
2 88433 1 19342
2 88434 1 19342
2 88435 1 19343
2 88436 1 19343
2 88437 1 19353
2 88438 1 19353
2 88439 1 19353
2 88440 1 19360
2 88441 1 19360
2 88442 1 19368
2 88443 1 19368
2 88444 1 19370
2 88445 1 19370
2 88446 1 19384
2 88447 1 19384
2 88448 1 19384
2 88449 1 19413
2 88450 1 19413
2 88451 1 19413
2 88452 1 19421
2 88453 1 19421
2 88454 1 19425
2 88455 1 19425
2 88456 1 19425
2 88457 1 19425
2 88458 1 19439
2 88459 1 19439
2 88460 1 19473
2 88461 1 19473
2 88462 1 19473
2 88463 1 19473
2 88464 1 19473
2 88465 1 19473
2 88466 1 19473
2 88467 1 19473
2 88468 1 19473
2 88469 1 19480
2 88470 1 19480
2 88471 1 19503
2 88472 1 19503
2 88473 1 19504
2 88474 1 19504
2 88475 1 19504
2 88476 1 19514
2 88477 1 19514
2 88478 1 19525
2 88479 1 19525
2 88480 1 19525
2 88481 1 19525
2 88482 1 19525
2 88483 1 19540
2 88484 1 19540
2 88485 1 19540
2 88486 1 19541
2 88487 1 19541
2 88488 1 19541
2 88489 1 19543
2 88490 1 19543
2 88491 1 19551
2 88492 1 19551
2 88493 1 19551
2 88494 1 19562
2 88495 1 19562
2 88496 1 19564
2 88497 1 19564
2 88498 1 19565
2 88499 1 19565
2 88500 1 19570
2 88501 1 19570
2 88502 1 19571
2 88503 1 19571
2 88504 1 19571
2 88505 1 19571
2 88506 1 19574
2 88507 1 19574
2 88508 1 19600
2 88509 1 19600
2 88510 1 19600
2 88511 1 19601
2 88512 1 19601
2 88513 1 19601
2 88514 1 19606
2 88515 1 19606
2 88516 1 19606
2 88517 1 19606
2 88518 1 19606
2 88519 1 19606
2 88520 1 19607
2 88521 1 19607
2 88522 1 19609
2 88523 1 19609
2 88524 1 19609
2 88525 1 19609
2 88526 1 19609
2 88527 1 19609
2 88528 1 19609
2 88529 1 19609
2 88530 1 19609
2 88531 1 19609
2 88532 1 19609
2 88533 1 19609
2 88534 1 19609
2 88535 1 19609
2 88536 1 19609
2 88537 1 19609
2 88538 1 19609
2 88539 1 19609
2 88540 1 19610
2 88541 1 19610
2 88542 1 19610
2 88543 1 19610
2 88544 1 19610
2 88545 1 19610
2 88546 1 19610
2 88547 1 19610
2 88548 1 19610
2 88549 1 19610
2 88550 1 19618
2 88551 1 19618
2 88552 1 19618
2 88553 1 19618
2 88554 1 19618
2 88555 1 19618
2 88556 1 19618
2 88557 1 19618
2 88558 1 19618
2 88559 1 19618
2 88560 1 19618
2 88561 1 19618
2 88562 1 19618
2 88563 1 19621
2 88564 1 19621
2 88565 1 19625
2 88566 1 19625
2 88567 1 19628
2 88568 1 19628
2 88569 1 19629
2 88570 1 19629
2 88571 1 19629
2 88572 1 19629
2 88573 1 19633
2 88574 1 19633
2 88575 1 19647
2 88576 1 19647
2 88577 1 19647
2 88578 1 19647
2 88579 1 19648
2 88580 1 19648
2 88581 1 19648
2 88582 1 19649
2 88583 1 19649
2 88584 1 19649
2 88585 1 19649
2 88586 1 19657
2 88587 1 19657
2 88588 1 19657
2 88589 1 19658
2 88590 1 19658
2 88591 1 19676
2 88592 1 19676
2 88593 1 19676
2 88594 1 19676
2 88595 1 19676
2 88596 1 19676
2 88597 1 19676
2 88598 1 19676
2 88599 1 19676
2 88600 1 19676
2 88601 1 19676
2 88602 1 19676
2 88603 1 19676
2 88604 1 19676
2 88605 1 19676
2 88606 1 19676
2 88607 1 19676
2 88608 1 19676
2 88609 1 19676
2 88610 1 19677
2 88611 1 19677
2 88612 1 19677
2 88613 1 19678
2 88614 1 19678
2 88615 1 19678
2 88616 1 19678
2 88617 1 19679
2 88618 1 19679
2 88619 1 19680
2 88620 1 19680
2 88621 1 19680
2 88622 1 19680
2 88623 1 19683
2 88624 1 19683
2 88625 1 19687
2 88626 1 19687
2 88627 1 19692
2 88628 1 19692
2 88629 1 19692
2 88630 1 19692
2 88631 1 19710
2 88632 1 19710
2 88633 1 19718
2 88634 1 19718
2 88635 1 19719
2 88636 1 19719
2 88637 1 19740
2 88638 1 19740
2 88639 1 19740
2 88640 1 19745
2 88641 1 19745
2 88642 1 19747
2 88643 1 19747
2 88644 1 19770
2 88645 1 19770
2 88646 1 19770
2 88647 1 19770
2 88648 1 19770
2 88649 1 19770
2 88650 1 19770
2 88651 1 19770
2 88652 1 19770
2 88653 1 19771
2 88654 1 19771
2 88655 1 19771
2 88656 1 19772
2 88657 1 19772
2 88658 1 19772
2 88659 1 19772
2 88660 1 19772
2 88661 1 19772
2 88662 1 19772
2 88663 1 19772
2 88664 1 19772
2 88665 1 19772
2 88666 1 19772
2 88667 1 19772
2 88668 1 19772
2 88669 1 19772
2 88670 1 19772
2 88671 1 19775
2 88672 1 19775
2 88673 1 19780
2 88674 1 19780
2 88675 1 19780
2 88676 1 19782
2 88677 1 19782
2 88678 1 19784
2 88679 1 19784
2 88680 1 19784
2 88681 1 19788
2 88682 1 19788
2 88683 1 19789
2 88684 1 19789
2 88685 1 19789
2 88686 1 19789
2 88687 1 19789
2 88688 1 19789
2 88689 1 19789
2 88690 1 19789
2 88691 1 19789
2 88692 1 19789
2 88693 1 19789
2 88694 1 19789
2 88695 1 19789
2 88696 1 19789
2 88697 1 19789
2 88698 1 19789
2 88699 1 19789
2 88700 1 19789
2 88701 1 19789
2 88702 1 19789
2 88703 1 19789
2 88704 1 19789
2 88705 1 19789
2 88706 1 19789
2 88707 1 19789
2 88708 1 19789
2 88709 1 19789
2 88710 1 19789
2 88711 1 19789
2 88712 1 19790
2 88713 1 19790
2 88714 1 19797
2 88715 1 19797
2 88716 1 19797
2 88717 1 19797
2 88718 1 19797
2 88719 1 19797
2 88720 1 19797
2 88721 1 19797
2 88722 1 19797
2 88723 1 19797
2 88724 1 19797
2 88725 1 19798
2 88726 1 19798
2 88727 1 19804
2 88728 1 19804
2 88729 1 19810
2 88730 1 19810
2 88731 1 19810
2 88732 1 19810
2 88733 1 19810
2 88734 1 19810
2 88735 1 19811
2 88736 1 19811
2 88737 1 19811
2 88738 1 19811
2 88739 1 19812
2 88740 1 19812
2 88741 1 19812
2 88742 1 19812
2 88743 1 19812
2 88744 1 19828
2 88745 1 19828
2 88746 1 19828
2 88747 1 19828
2 88748 1 19828
2 88749 1 19828
2 88750 1 19828
2 88751 1 19828
2 88752 1 19832
2 88753 1 19832
2 88754 1 19832
2 88755 1 19832
2 88756 1 19832
2 88757 1 19832
2 88758 1 19832
2 88759 1 19832
2 88760 1 19832
2 88761 1 19832
2 88762 1 19833
2 88763 1 19833
2 88764 1 19833
2 88765 1 19833
2 88766 1 19842
2 88767 1 19842
2 88768 1 19842
2 88769 1 19842
2 88770 1 19842
2 88771 1 19842
2 88772 1 19872
2 88773 1 19872
2 88774 1 19872
2 88775 1 19872
2 88776 1 19872
2 88777 1 19872
2 88778 1 19873
2 88779 1 19873
2 88780 1 19873
2 88781 1 19880
2 88782 1 19880
2 88783 1 19901
2 88784 1 19901
2 88785 1 19901
2 88786 1 19928
2 88787 1 19928
2 88788 1 19946
2 88789 1 19946
2 88790 1 19946
2 88791 1 19946
2 88792 1 19946
2 88793 1 19946
2 88794 1 19970
2 88795 1 19970
2 88796 1 19989
2 88797 1 19989
2 88798 1 19989
2 88799 1 19989
2 88800 1 19989
2 88801 1 19990
2 88802 1 19990
2 88803 1 19990
2 88804 1 20006
2 88805 1 20006
2 88806 1 20007
2 88807 1 20007
2 88808 1 20010
2 88809 1 20010
2 88810 1 20010
2 88811 1 20010
2 88812 1 20010
2 88813 1 20010
2 88814 1 20010
2 88815 1 20011
2 88816 1 20011
2 88817 1 20011
2 88818 1 20011
2 88819 1 20016
2 88820 1 20016
2 88821 1 20028
2 88822 1 20028
2 88823 1 20028
2 88824 1 20028
2 88825 1 20028
2 88826 1 20029
2 88827 1 20029
2 88828 1 20045
2 88829 1 20045
2 88830 1 20045
2 88831 1 20053
2 88832 1 20053
2 88833 1 20054
2 88834 1 20054
2 88835 1 20054
2 88836 1 20054
2 88837 1 20071
2 88838 1 20071
2 88839 1 20093
2 88840 1 20093
2 88841 1 20103
2 88842 1 20103
2 88843 1 20121
2 88844 1 20121
2 88845 1 20121
2 88846 1 20121
2 88847 1 20122
2 88848 1 20122
2 88849 1 20122
2 88850 1 20122
2 88851 1 20122
2 88852 1 20132
2 88853 1 20132
2 88854 1 20132
2 88855 1 20132
2 88856 1 20132
2 88857 1 20132
2 88858 1 20132
2 88859 1 20133
2 88860 1 20133
2 88861 1 20134
2 88862 1 20134
2 88863 1 20143
2 88864 1 20143
2 88865 1 20143
2 88866 1 20143
2 88867 1 20154
2 88868 1 20154
2 88869 1 20154
2 88870 1 20154
2 88871 1 20154
2 88872 1 20154
2 88873 1 20154
2 88874 1 20154
2 88875 1 20154
2 88876 1 20154
2 88877 1 20154
2 88878 1 20154
2 88879 1 20156
2 88880 1 20156
2 88881 1 20157
2 88882 1 20157
2 88883 1 20157
2 88884 1 20184
2 88885 1 20184
2 88886 1 20188
2 88887 1 20188
2 88888 1 20188
2 88889 1 20189
2 88890 1 20189
2 88891 1 20194
2 88892 1 20194
2 88893 1 20194
2 88894 1 20194
2 88895 1 20202
2 88896 1 20202
2 88897 1 20202
2 88898 1 20202
2 88899 1 20202
2 88900 1 20202
2 88901 1 20202
2 88902 1 20202
2 88903 1 20202
2 88904 1 20202
2 88905 1 20202
2 88906 1 20202
2 88907 1 20202
2 88908 1 20202
2 88909 1 20202
2 88910 1 20202
2 88911 1 20202
2 88912 1 20202
2 88913 1 20202
2 88914 1 20202
2 88915 1 20202
2 88916 1 20202
2 88917 1 20202
2 88918 1 20202
2 88919 1 20209
2 88920 1 20209
2 88921 1 20209
2 88922 1 20209
2 88923 1 20209
2 88924 1 20209
2 88925 1 20209
2 88926 1 20209
2 88927 1 20209
2 88928 1 20220
2 88929 1 20220
2 88930 1 20220
2 88931 1 20222
2 88932 1 20222
2 88933 1 20222
2 88934 1 20228
2 88935 1 20228
2 88936 1 20228
2 88937 1 20229
2 88938 1 20229
2 88939 1 20232
2 88940 1 20232
2 88941 1 20232
2 88942 1 20244
2 88943 1 20244
2 88944 1 20247
2 88945 1 20247
2 88946 1 20247
2 88947 1 20248
2 88948 1 20248
2 88949 1 20248
2 88950 1 20248
2 88951 1 20248
2 88952 1 20248
2 88953 1 20248
2 88954 1 20265
2 88955 1 20265
2 88956 1 20265
2 88957 1 20265
2 88958 1 20265
2 88959 1 20280
2 88960 1 20280
2 88961 1 20300
2 88962 1 20300
2 88963 1 20300
2 88964 1 20300
2 88965 1 20300
2 88966 1 20300
2 88967 1 20339
2 88968 1 20339
2 88969 1 20339
2 88970 1 20339
2 88971 1 20339
2 88972 1 20345
2 88973 1 20345
2 88974 1 20353
2 88975 1 20353
2 88976 1 20364
2 88977 1 20364
2 88978 1 20364
2 88979 1 20365
2 88980 1 20365
2 88981 1 20365
2 88982 1 20366
2 88983 1 20366
2 88984 1 20366
2 88985 1 20377
2 88986 1 20377
2 88987 1 20378
2 88988 1 20378
2 88989 1 20379
2 88990 1 20379
2 88991 1 20379
2 88992 1 20379
2 88993 1 20380
2 88994 1 20380
2 88995 1 20387
2 88996 1 20387
2 88997 1 20387
2 88998 1 20388
2 88999 1 20388
2 89000 1 20391
2 89001 1 20391
2 89002 1 20391
2 89003 1 20391
2 89004 1 20399
2 89005 1 20399
2 89006 1 20399
2 89007 1 20399
2 89008 1 20399
2 89009 1 20399
2 89010 1 20400
2 89011 1 20400
2 89012 1 20407
2 89013 1 20407
2 89014 1 20407
2 89015 1 20408
2 89016 1 20408
2 89017 1 20408
2 89018 1 20408
2 89019 1 20409
2 89020 1 20409
2 89021 1 20410
2 89022 1 20410
2 89023 1 20410
2 89024 1 20410
2 89025 1 20410
2 89026 1 20411
2 89027 1 20411
2 89028 1 20426
2 89029 1 20426
2 89030 1 20427
2 89031 1 20427
2 89032 1 20427
2 89033 1 20461
2 89034 1 20461
2 89035 1 20490
2 89036 1 20490
2 89037 1 20504
2 89038 1 20504
2 89039 1 20504
2 89040 1 20504
2 89041 1 20504
2 89042 1 20505
2 89043 1 20505
2 89044 1 20505
2 89045 1 20505
2 89046 1 20514
2 89047 1 20514
2 89048 1 20514
2 89049 1 20514
2 89050 1 20514
2 89051 1 20514
2 89052 1 20514
2 89053 1 20514
2 89054 1 20514
2 89055 1 20514
2 89056 1 20514
2 89057 1 20514
2 89058 1 20514
2 89059 1 20514
2 89060 1 20514
2 89061 1 20514
2 89062 1 20514
2 89063 1 20514
2 89064 1 20515
2 89065 1 20515
2 89066 1 20518
2 89067 1 20518
2 89068 1 20531
2 89069 1 20531
2 89070 1 20545
2 89071 1 20545
2 89072 1 20546
2 89073 1 20546
2 89074 1 20549
2 89075 1 20549
2 89076 1 20549
2 89077 1 20549
2 89078 1 20584
2 89079 1 20584
2 89080 1 20584
2 89081 1 20584
2 89082 1 20584
2 89083 1 20584
2 89084 1 20584
2 89085 1 20584
2 89086 1 20584
2 89087 1 20584
2 89088 1 20584
2 89089 1 20584
2 89090 1 20584
2 89091 1 20584
2 89092 1 20584
2 89093 1 20584
2 89094 1 20584
2 89095 1 20584
2 89096 1 20594
2 89097 1 20594
2 89098 1 20594
2 89099 1 20594
2 89100 1 20594
2 89101 1 20594
2 89102 1 20594
2 89103 1 20594
2 89104 1 20594
2 89105 1 20594
2 89106 1 20594
2 89107 1 20594
2 89108 1 20594
2 89109 1 20594
2 89110 1 20594
2 89111 1 20595
2 89112 1 20595
2 89113 1 20596
2 89114 1 20596
2 89115 1 20596
2 89116 1 20596
2 89117 1 20596
2 89118 1 20596
2 89119 1 20596
2 89120 1 20596
2 89121 1 20596
2 89122 1 20596
2 89123 1 20596
2 89124 1 20596
2 89125 1 20596
2 89126 1 20596
2 89127 1 20596
2 89128 1 20596
2 89129 1 20596
2 89130 1 20596
2 89131 1 20596
2 89132 1 20596
2 89133 1 20596
2 89134 1 20596
2 89135 1 20596
2 89136 1 20596
2 89137 1 20596
2 89138 1 20596
2 89139 1 20596
2 89140 1 20596
2 89141 1 20596
2 89142 1 20596
2 89143 1 20596
2 89144 1 20617
2 89145 1 20617
2 89146 1 20623
2 89147 1 20623
2 89148 1 20631
2 89149 1 20631
2 89150 1 20631
2 89151 1 20631
2 89152 1 20631
2 89153 1 20631
2 89154 1 20632
2 89155 1 20632
2 89156 1 20632
2 89157 1 20632
2 89158 1 20643
2 89159 1 20643
2 89160 1 20643
2 89161 1 20643
2 89162 1 20643
2 89163 1 20643
2 89164 1 20643
2 89165 1 20644
2 89166 1 20644
2 89167 1 20644
2 89168 1 20644
2 89169 1 20644
2 89170 1 20654
2 89171 1 20654
2 89172 1 20654
2 89173 1 20654
2 89174 1 20654
2 89175 1 20655
2 89176 1 20655
2 89177 1 20655
2 89178 1 20658
2 89179 1 20658
2 89180 1 20658
2 89181 1 20659
2 89182 1 20659
2 89183 1 20660
2 89184 1 20660
2 89185 1 20660
2 89186 1 20660
2 89187 1 20660
2 89188 1 20660
2 89189 1 20675
2 89190 1 20675
2 89191 1 20675
2 89192 1 20675
2 89193 1 20678
2 89194 1 20678
2 89195 1 20678
2 89196 1 20694
2 89197 1 20694
2 89198 1 20694
2 89199 1 20694
2 89200 1 20696
2 89201 1 20696
2 89202 1 20699
2 89203 1 20699
2 89204 1 20699
2 89205 1 20699
2 89206 1 20699
2 89207 1 20699
2 89208 1 20701
2 89209 1 20701
2 89210 1 20715
2 89211 1 20715
2 89212 1 20726
2 89213 1 20726
2 89214 1 20727
2 89215 1 20727
2 89216 1 20760
2 89217 1 20760
2 89218 1 20760
2 89219 1 20773
2 89220 1 20773
2 89221 1 20773
2 89222 1 20773
2 89223 1 20773
2 89224 1 20773
2 89225 1 20773
2 89226 1 20773
2 89227 1 20773
2 89228 1 20773
2 89229 1 20773
2 89230 1 20773
2 89231 1 20773
2 89232 1 20773
2 89233 1 20773
2 89234 1 20773
2 89235 1 20773
2 89236 1 20773
2 89237 1 20773
2 89238 1 20773
2 89239 1 20773
2 89240 1 20774
2 89241 1 20774
2 89242 1 20774
2 89243 1 20774
2 89244 1 20775
2 89245 1 20775
2 89246 1 20775
2 89247 1 20775
2 89248 1 20775
2 89249 1 20775
2 89250 1 20775
2 89251 1 20776
2 89252 1 20776
2 89253 1 20776
2 89254 1 20776
2 89255 1 20776
2 89256 1 20776
2 89257 1 20776
2 89258 1 20776
2 89259 1 20776
2 89260 1 20776
2 89261 1 20776
2 89262 1 20776
2 89263 1 20776
2 89264 1 20776
2 89265 1 20776
2 89266 1 20776
2 89267 1 20776
2 89268 1 20776
2 89269 1 20776
2 89270 1 20776
2 89271 1 20776
2 89272 1 20777
2 89273 1 20777
2 89274 1 20784
2 89275 1 20784
2 89276 1 20788
2 89277 1 20788
2 89278 1 20788
2 89279 1 20800
2 89280 1 20800
2 89281 1 20801
2 89282 1 20801
2 89283 1 20824
2 89284 1 20824
2 89285 1 20824
2 89286 1 20824
2 89287 1 20833
2 89288 1 20833
2 89289 1 20834
2 89290 1 20834
2 89291 1 20834
2 89292 1 20834
2 89293 1 20835
2 89294 1 20835
2 89295 1 20835
2 89296 1 20835
2 89297 1 20835
2 89298 1 20835
2 89299 1 20847
2 89300 1 20847
2 89301 1 20847
2 89302 1 20848
2 89303 1 20848
2 89304 1 20848
2 89305 1 20858
2 89306 1 20858
2 89307 1 20859
2 89308 1 20859
2 89309 1 20869
2 89310 1 20869
2 89311 1 20869
2 89312 1 20869
2 89313 1 20869
2 89314 1 20870
2 89315 1 20870
2 89316 1 20870
2 89317 1 20870
2 89318 1 20870
2 89319 1 20870
2 89320 1 20870
2 89321 1 20871
2 89322 1 20871
2 89323 1 20871
2 89324 1 20871
2 89325 1 20871
2 89326 1 20871
2 89327 1 20875
2 89328 1 20875
2 89329 1 20875
2 89330 1 20878
2 89331 1 20878
2 89332 1 20888
2 89333 1 20888
2 89334 1 20888
2 89335 1 20888
2 89336 1 20889
2 89337 1 20889
2 89338 1 20889
2 89339 1 20890
2 89340 1 20890
2 89341 1 20890
2 89342 1 20890
2 89343 1 20898
2 89344 1 20898
2 89345 1 20899
2 89346 1 20899
2 89347 1 20899
2 89348 1 20900
2 89349 1 20900
2 89350 1 20913
2 89351 1 20913
2 89352 1 20915
2 89353 1 20915
2 89354 1 20915
2 89355 1 20915
2 89356 1 20915
2 89357 1 20915
2 89358 1 20915
2 89359 1 20915
2 89360 1 20915
2 89361 1 20915
2 89362 1 20915
2 89363 1 20916
2 89364 1 20916
2 89365 1 20916
2 89366 1 20927
2 89367 1 20927
2 89368 1 20941
2 89369 1 20941
2 89370 1 20941
2 89371 1 20941
2 89372 1 20942
2 89373 1 20942
2 89374 1 20943
2 89375 1 20943
2 89376 1 20943
2 89377 1 20957
2 89378 1 20957
2 89379 1 20957
2 89380 1 20958
2 89381 1 20958
2 89382 1 20958
2 89383 1 20961
2 89384 1 20961
2 89385 1 20961
2 89386 1 20961
2 89387 1 20961
2 89388 1 20961
2 89389 1 20961
2 89390 1 20961
2 89391 1 20961
2 89392 1 20962
2 89393 1 20962
2 89394 1 20962
2 89395 1 20962
2 89396 1 20993
2 89397 1 20993
2 89398 1 20998
2 89399 1 20998
2 89400 1 20998
2 89401 1 21007
2 89402 1 21007
2 89403 1 21007
2 89404 1 21007
2 89405 1 21007
2 89406 1 21008
2 89407 1 21008
2 89408 1 21008
2 89409 1 21008
2 89410 1 21008
2 89411 1 21010
2 89412 1 21010
2 89413 1 21011
2 89414 1 21011
2 89415 1 21013
2 89416 1 21013
2 89417 1 21013
2 89418 1 21013
2 89419 1 21014
2 89420 1 21014
2 89421 1 21017
2 89422 1 21017
2 89423 1 21027
2 89424 1 21027
2 89425 1 21027
2 89426 1 21027
2 89427 1 21027
2 89428 1 21027
2 89429 1 21027
2 89430 1 21035
2 89431 1 21035
2 89432 1 21035
2 89433 1 21035
2 89434 1 21035
2 89435 1 21048
2 89436 1 21048
2 89437 1 21048
2 89438 1 21049
2 89439 1 21049
2 89440 1 21057
2 89441 1 21057
2 89442 1 21061
2 89443 1 21061
2 89444 1 21068
2 89445 1 21068
2 89446 1 21068
2 89447 1 21068
2 89448 1 21068
2 89449 1 21068
2 89450 1 21068
2 89451 1 21068
2 89452 1 21069
2 89453 1 21069
2 89454 1 21072
2 89455 1 21072
2 89456 1 21072
2 89457 1 21072
2 89458 1 21072
2 89459 1 21072
2 89460 1 21084
2 89461 1 21084
2 89462 1 21115
2 89463 1 21115
2 89464 1 21115
2 89465 1 21115
2 89466 1 21115
2 89467 1 21115
2 89468 1 21115
2 89469 1 21116
2 89470 1 21116
2 89471 1 21116
2 89472 1 21118
2 89473 1 21118
2 89474 1 21119
2 89475 1 21119
2 89476 1 21119
2 89477 1 21119
2 89478 1 21119
2 89479 1 21119
2 89480 1 21120
2 89481 1 21120
2 89482 1 21127
2 89483 1 21127
2 89484 1 21136
2 89485 1 21136
2 89486 1 21165
2 89487 1 21165
2 89488 1 21165
2 89489 1 21171
2 89490 1 21171
2 89491 1 21171
2 89492 1 21180
2 89493 1 21180
2 89494 1 21181
2 89495 1 21181
2 89496 1 21181
2 89497 1 21181
2 89498 1 21181
2 89499 1 21196
2 89500 1 21196
2 89501 1 21196
2 89502 1 21196
2 89503 1 21196
2 89504 1 21196
2 89505 1 21196
2 89506 1 21196
2 89507 1 21196
2 89508 1 21196
2 89509 1 21196
2 89510 1 21196
2 89511 1 21196
2 89512 1 21210
2 89513 1 21210
2 89514 1 21210
2 89515 1 21210
2 89516 1 21215
2 89517 1 21215
2 89518 1 21215
2 89519 1 21218
2 89520 1 21218
2 89521 1 21218
2 89522 1 21223
2 89523 1 21223
2 89524 1 21223
2 89525 1 21224
2 89526 1 21224
2 89527 1 21224
2 89528 1 21226
2 89529 1 21226
2 89530 1 21226
2 89531 1 21227
2 89532 1 21227
2 89533 1 21228
2 89534 1 21228
2 89535 1 21228
2 89536 1 21233
2 89537 1 21233
2 89538 1 21247
2 89539 1 21247
2 89540 1 21247
2 89541 1 21247
2 89542 1 21252
2 89543 1 21252
2 89544 1 21255
2 89545 1 21255
2 89546 1 21255
2 89547 1 21260
2 89548 1 21260
2 89549 1 21264
2 89550 1 21264
2 89551 1 21265
2 89552 1 21265
2 89553 1 21288
2 89554 1 21288
2 89555 1 21288
2 89556 1 21288
2 89557 1 21289
2 89558 1 21289
2 89559 1 21290
2 89560 1 21290
2 89561 1 21297
2 89562 1 21297
2 89563 1 21316
2 89564 1 21316
2 89565 1 21316
2 89566 1 21328
2 89567 1 21328
2 89568 1 21328
2 89569 1 21328
2 89570 1 21328
2 89571 1 21328
2 89572 1 21328
2 89573 1 21329
2 89574 1 21329
2 89575 1 21332
2 89576 1 21332
2 89577 1 21332
2 89578 1 21332
2 89579 1 21332
2 89580 1 21332
2 89581 1 21332
2 89582 1 21332
2 89583 1 21332
2 89584 1 21332
2 89585 1 21332
2 89586 1 21332
2 89587 1 21332
2 89588 1 21332
2 89589 1 21332
2 89590 1 21332
2 89591 1 21332
2 89592 1 21332
2 89593 1 21332
2 89594 1 21332
2 89595 1 21332
2 89596 1 21332
2 89597 1 21332
2 89598 1 21332
2 89599 1 21332
2 89600 1 21333
2 89601 1 21333
2 89602 1 21333
2 89603 1 21333
2 89604 1 21347
2 89605 1 21347
2 89606 1 21347
2 89607 1 21347
2 89608 1 21347
2 89609 1 21347
2 89610 1 21347
2 89611 1 21347
2 89612 1 21347
2 89613 1 21356
2 89614 1 21356
2 89615 1 21356
2 89616 1 21356
2 89617 1 21357
2 89618 1 21357
2 89619 1 21357
2 89620 1 21370
2 89621 1 21370
2 89622 1 21371
2 89623 1 21371
2 89624 1 21372
2 89625 1 21372
2 89626 1 21372
2 89627 1 21372
2 89628 1 21372
2 89629 1 21372
2 89630 1 21372
2 89631 1 21372
2 89632 1 21372
2 89633 1 21373
2 89634 1 21373
2 89635 1 21374
2 89636 1 21374
2 89637 1 21374
2 89638 1 21374
2 89639 1 21374
2 89640 1 21374
2 89641 1 21374
2 89642 1 21374
2 89643 1 21374
2 89644 1 21374
2 89645 1 21374
2 89646 1 21374
2 89647 1 21374
2 89648 1 21374
2 89649 1 21374
2 89650 1 21374
2 89651 1 21374
2 89652 1 21374
2 89653 1 21374
2 89654 1 21374
2 89655 1 21374
2 89656 1 21374
2 89657 1 21374
2 89658 1 21374
2 89659 1 21374
2 89660 1 21374
2 89661 1 21374
2 89662 1 21375
2 89663 1 21375
2 89664 1 21378
2 89665 1 21378
2 89666 1 21378
2 89667 1 21378
2 89668 1 21379
2 89669 1 21379
2 89670 1 21386
2 89671 1 21386
2 89672 1 21386
2 89673 1 21387
2 89674 1 21387
2 89675 1 21395
2 89676 1 21395
2 89677 1 21395
2 89678 1 21395
2 89679 1 21396
2 89680 1 21396
2 89681 1 21396
2 89682 1 21396
2 89683 1 21397
2 89684 1 21397
2 89685 1 21398
2 89686 1 21398
2 89687 1 21398
2 89688 1 21398
2 89689 1 21402
2 89690 1 21402
2 89691 1 21402
2 89692 1 21410
2 89693 1 21410
2 89694 1 21410
2 89695 1 21410
2 89696 1 21410
2 89697 1 21410
2 89698 1 21410
2 89699 1 21410
2 89700 1 21410
2 89701 1 21411
2 89702 1 21411
2 89703 1 21413
2 89704 1 21413
2 89705 1 21414
2 89706 1 21414
2 89707 1 21414
2 89708 1 21422
2 89709 1 21422
2 89710 1 21424
2 89711 1 21424
2 89712 1 21442
2 89713 1 21442
2 89714 1 21442
2 89715 1 21442
2 89716 1 21442
2 89717 1 21442
2 89718 1 21456
2 89719 1 21456
2 89720 1 21467
2 89721 1 21467
2 89722 1 21467
2 89723 1 21467
2 89724 1 21477
2 89725 1 21477
2 89726 1 21487
2 89727 1 21487
2 89728 1 21487
2 89729 1 21493
2 89730 1 21493
2 89731 1 21493
2 89732 1 21502
2 89733 1 21502
2 89734 1 21502
2 89735 1 21502
2 89736 1 21502
2 89737 1 21502
2 89738 1 21510
2 89739 1 21510
2 89740 1 21510
2 89741 1 21510
2 89742 1 21510
2 89743 1 21511
2 89744 1 21511
2 89745 1 21511
2 89746 1 21511
2 89747 1 21511
2 89748 1 21511
2 89749 1 21513
2 89750 1 21513
2 89751 1 21513
2 89752 1 21528
2 89753 1 21528
2 89754 1 21528
2 89755 1 21528
2 89756 1 21528
2 89757 1 21546
2 89758 1 21546
2 89759 1 21549
2 89760 1 21549
2 89761 1 21550
2 89762 1 21550
2 89763 1 21553
2 89764 1 21553
2 89765 1 21554
2 89766 1 21554
2 89767 1 21554
2 89768 1 21569
2 89769 1 21569
2 89770 1 21569
2 89771 1 21569
2 89772 1 21569
2 89773 1 21570
2 89774 1 21570
2 89775 1 21573
2 89776 1 21573
2 89777 1 21573
2 89778 1 21594
2 89779 1 21594
2 89780 1 21621
2 89781 1 21621
2 89782 1 21624
2 89783 1 21624
2 89784 1 21624
2 89785 1 21626
2 89786 1 21626
2 89787 1 21630
2 89788 1 21630
2 89789 1 21630
2 89790 1 21630
2 89791 1 21630
2 89792 1 21631
2 89793 1 21631
2 89794 1 21639
2 89795 1 21639
2 89796 1 21644
2 89797 1 21644
2 89798 1 21653
2 89799 1 21653
2 89800 1 21656
2 89801 1 21656
2 89802 1 21656
2 89803 1 21656
2 89804 1 21666
2 89805 1 21666
2 89806 1 21670
2 89807 1 21670
2 89808 1 21670
2 89809 1 21670
2 89810 1 21670
2 89811 1 21670
2 89812 1 21671
2 89813 1 21671
2 89814 1 21673
2 89815 1 21673
2 89816 1 21673
2 89817 1 21673
2 89818 1 21673
2 89819 1 21679
2 89820 1 21679
2 89821 1 21694
2 89822 1 21694
2 89823 1 21694
2 89824 1 21694
2 89825 1 21695
2 89826 1 21695
2 89827 1 21695
2 89828 1 21695
2 89829 1 21695
2 89830 1 21701
2 89831 1 21701
2 89832 1 21701
2 89833 1 21701
2 89834 1 21701
2 89835 1 21701
2 89836 1 21701
2 89837 1 21701
2 89838 1 21721
2 89839 1 21721
2 89840 1 21745
2 89841 1 21745
2 89842 1 21749
2 89843 1 21749
2 89844 1 21749
2 89845 1 21759
2 89846 1 21759
2 89847 1 21759
2 89848 1 21759
2 89849 1 21760
2 89850 1 21760
2 89851 1 21760
2 89852 1 21762
2 89853 1 21762
2 89854 1 21762
2 89855 1 21771
2 89856 1 21771
2 89857 1 21771
2 89858 1 21771
2 89859 1 21771
2 89860 1 21771
2 89861 1 21772
2 89862 1 21772
2 89863 1 21773
2 89864 1 21773
2 89865 1 21773
2 89866 1 21780
2 89867 1 21780
2 89868 1 21780
2 89869 1 21780
2 89870 1 21780
2 89871 1 21780
2 89872 1 21781
2 89873 1 21781
2 89874 1 21781
2 89875 1 21781
2 89876 1 21781
2 89877 1 21790
2 89878 1 21790
2 89879 1 21790
2 89880 1 21790
2 89881 1 21790
2 89882 1 21790
2 89883 1 21790
2 89884 1 21790
2 89885 1 21790
2 89886 1 21790
2 89887 1 21791
2 89888 1 21791
2 89889 1 21798
2 89890 1 21798
2 89891 1 21799
2 89892 1 21799
2 89893 1 21810
2 89894 1 21810
2 89895 1 21810
2 89896 1 21810
2 89897 1 21810
2 89898 1 21810
2 89899 1 21810
2 89900 1 21810
2 89901 1 21810
2 89902 1 21810
2 89903 1 21810
2 89904 1 21810
2 89905 1 21810
2 89906 1 21810
2 89907 1 21810
2 89908 1 21810
2 89909 1 21810
2 89910 1 21810
2 89911 1 21810
2 89912 1 21810
2 89913 1 21818
2 89914 1 21818
2 89915 1 21818
2 89916 1 21818
2 89917 1 21818
2 89918 1 21818
2 89919 1 21820
2 89920 1 21820
2 89921 1 21824
2 89922 1 21824
2 89923 1 21824
2 89924 1 21824
2 89925 1 21825
2 89926 1 21825
2 89927 1 21825
2 89928 1 21825
2 89929 1 21825
2 89930 1 21825
2 89931 1 21826
2 89932 1 21826
2 89933 1 21826
2 89934 1 21839
2 89935 1 21839
2 89936 1 21839
2 89937 1 21843
2 89938 1 21843
2 89939 1 21843
2 89940 1 21847
2 89941 1 21847
2 89942 1 21848
2 89943 1 21848
2 89944 1 21850
2 89945 1 21850
2 89946 1 21854
2 89947 1 21854
2 89948 1 21854
2 89949 1 21860
2 89950 1 21860
2 89951 1 21861
2 89952 1 21861
2 89953 1 21861
2 89954 1 21864
2 89955 1 21864
2 89956 1 21865
2 89957 1 21865
2 89958 1 21870
2 89959 1 21870
2 89960 1 21883
2 89961 1 21883
2 89962 1 21883
2 89963 1 21893
2 89964 1 21893
2 89965 1 21893
2 89966 1 21895
2 89967 1 21895
2 89968 1 21903
2 89969 1 21903
2 89970 1 21903
2 89971 1 21903
2 89972 1 21903
2 89973 1 21903
2 89974 1 21903
2 89975 1 21904
2 89976 1 21904
2 89977 1 21912
2 89978 1 21912
2 89979 1 21918
2 89980 1 21918
2 89981 1 21918
2 89982 1 21930
2 89983 1 21930
2 89984 1 21931
2 89985 1 21931
2 89986 1 21931
2 89987 1 21931
2 89988 1 21931
2 89989 1 21941
2 89990 1 21941
2 89991 1 21959
2 89992 1 21959
2 89993 1 21961
2 89994 1 21961
2 89995 1 21961
2 89996 1 21961
2 89997 1 21961
2 89998 1 21961
2 89999 1 21961
2 90000 1 21961
2 90001 1 21965
2 90002 1 21965
2 90003 1 21965
2 90004 1 21965
2 90005 1 21966
2 90006 1 21966
2 90007 1 21967
2 90008 1 21967
2 90009 1 21967
2 90010 1 21967
2 90011 1 21967
2 90012 1 21968
2 90013 1 21968
2 90014 1 21968
2 90015 1 21968
2 90016 1 21968
2 90017 1 21968
2 90018 1 21976
2 90019 1 21976
2 90020 1 21979
2 90021 1 21979
2 90022 1 21979
2 90023 1 21979
2 90024 1 21980
2 90025 1 21980
2 90026 1 21980
2 90027 1 21980
2 90028 1 21980
2 90029 1 21980
2 90030 1 21980
2 90031 1 21980
2 90032 1 21980
2 90033 1 21980
2 90034 1 21982
2 90035 1 21982
2 90036 1 21989
2 90037 1 21989
2 90038 1 21997
2 90039 1 21997
2 90040 1 21997
2 90041 1 21998
2 90042 1 21998
2 90043 1 21998
2 90044 1 21998
2 90045 1 22000
2 90046 1 22000
2 90047 1 22000
2 90048 1 22013
2 90049 1 22013
2 90050 1 22014
2 90051 1 22014
2 90052 1 22034
2 90053 1 22034
2 90054 1 22034
2 90055 1 22034
2 90056 1 22034
2 90057 1 22034
2 90058 1 22034
2 90059 1 22034
2 90060 1 22034
2 90061 1 22034
2 90062 1 22055
2 90063 1 22055
2 90064 1 22056
2 90065 1 22056
2 90066 1 22056
2 90067 1 22056
2 90068 1 22090
2 90069 1 22090
2 90070 1 22090
2 90071 1 22090
2 90072 1 22090
2 90073 1 22090
2 90074 1 22090
2 90075 1 22090
2 90076 1 22090
2 90077 1 22090
2 90078 1 22090
2 90079 1 22125
2 90080 1 22125
2 90081 1 22128
2 90082 1 22128
2 90083 1 22129
2 90084 1 22129
2 90085 1 22129
2 90086 1 22129
2 90087 1 22129
2 90088 1 22131
2 90089 1 22131
2 90090 1 22131
2 90091 1 22164
2 90092 1 22164
2 90093 1 22175
2 90094 1 22175
2 90095 1 22175
2 90096 1 22175
2 90097 1 22175
2 90098 1 22175
2 90099 1 22184
2 90100 1 22184
2 90101 1 22184
2 90102 1 22203
2 90103 1 22203
2 90104 1 22203
2 90105 1 22203
2 90106 1 22203
2 90107 1 22203
2 90108 1 22203
2 90109 1 22203
2 90110 1 22204
2 90111 1 22204
2 90112 1 22205
2 90113 1 22205
2 90114 1 22205
2 90115 1 22205
2 90116 1 22205
2 90117 1 22205
2 90118 1 22228
2 90119 1 22228
2 90120 1 22232
2 90121 1 22232
2 90122 1 22235
2 90123 1 22235
2 90124 1 22242
2 90125 1 22242
2 90126 1 22252
2 90127 1 22252
2 90128 1 22269
2 90129 1 22269
2 90130 1 22269
2 90131 1 22269
2 90132 1 22269
2 90133 1 22269
2 90134 1 22269
2 90135 1 22269
2 90136 1 22281
2 90137 1 22281
2 90138 1 22281
2 90139 1 22281
2 90140 1 22281
2 90141 1 22281
2 90142 1 22282
2 90143 1 22282
2 90144 1 22282
2 90145 1 22323
2 90146 1 22323
2 90147 1 22323
2 90148 1 22323
2 90149 1 22324
2 90150 1 22324
2 90151 1 22335
2 90152 1 22335
2 90153 1 22335
2 90154 1 22335
2 90155 1 22335
2 90156 1 22335
2 90157 1 22335
2 90158 1 22336
2 90159 1 22336
2 90160 1 22336
2 90161 1 22336
2 90162 1 22336
2 90163 1 22337
2 90164 1 22337
2 90165 1 22337
2 90166 1 22337
2 90167 1 22348
2 90168 1 22348
2 90169 1 22362
2 90170 1 22362
2 90171 1 22379
2 90172 1 22379
2 90173 1 22379
2 90174 1 22379
2 90175 1 22379
2 90176 1 22379
2 90177 1 22379
2 90178 1 22379
2 90179 1 22379
2 90180 1 22379
2 90181 1 22379
2 90182 1 22379
2 90183 1 22379
2 90184 1 22379
2 90185 1 22381
2 90186 1 22381
2 90187 1 22384
2 90188 1 22384
2 90189 1 22384
2 90190 1 22384
2 90191 1 22384
2 90192 1 22384
2 90193 1 22394
2 90194 1 22394
2 90195 1 22394
2 90196 1 22395
2 90197 1 22395
2 90198 1 22395
2 90199 1 22400
2 90200 1 22400
2 90201 1 22407
2 90202 1 22407
2 90203 1 22416
2 90204 1 22416
2 90205 1 22423
2 90206 1 22423
2 90207 1 22424
2 90208 1 22424
2 90209 1 22425
2 90210 1 22425
2 90211 1 22425
2 90212 1 22425
2 90213 1 22425
2 90214 1 22441
2 90215 1 22441
2 90216 1 22441
2 90217 1 22441
2 90218 1 22441
2 90219 1 22443
2 90220 1 22443
2 90221 1 22447
2 90222 1 22447
2 90223 1 22447
2 90224 1 22447
2 90225 1 22448
2 90226 1 22448
2 90227 1 22448
2 90228 1 22448
2 90229 1 22448
2 90230 1 22449
2 90231 1 22449
2 90232 1 22449
2 90233 1 22449
2 90234 1 22449
2 90235 1 22449
2 90236 1 22449
2 90237 1 22449
2 90238 1 22451
2 90239 1 22451
2 90240 1 22458
2 90241 1 22458
2 90242 1 22458
2 90243 1 22459
2 90244 1 22459
2 90245 1 22459
2 90246 1 22462
2 90247 1 22462
2 90248 1 22462
2 90249 1 22462
2 90250 1 22462
2 90251 1 22462
2 90252 1 22463
2 90253 1 22463
2 90254 1 22463
2 90255 1 22463
2 90256 1 22480
2 90257 1 22480
2 90258 1 22480
2 90259 1 22480
2 90260 1 22480
2 90261 1 22480
2 90262 1 22480
2 90263 1 22480
2 90264 1 22480
2 90265 1 22480
2 90266 1 22494
2 90267 1 22494
2 90268 1 22494
2 90269 1 22495
2 90270 1 22495
2 90271 1 22502
2 90272 1 22502
2 90273 1 22505
2 90274 1 22505
2 90275 1 22514
2 90276 1 22514
2 90277 1 22522
2 90278 1 22522
2 90279 1 22543
2 90280 1 22543
2 90281 1 22543
2 90282 1 22548
2 90283 1 22548
2 90284 1 22548
2 90285 1 22549
2 90286 1 22549
2 90287 1 22549
2 90288 1 22549
2 90289 1 22557
2 90290 1 22557
2 90291 1 22557
2 90292 1 22578
2 90293 1 22578
2 90294 1 22587
2 90295 1 22587
2 90296 1 22616
2 90297 1 22616
2 90298 1 22617
2 90299 1 22617
2 90300 1 22640
2 90301 1 22640
2 90302 1 22640
2 90303 1 22640
2 90304 1 22640
2 90305 1 22641
2 90306 1 22641
2 90307 1 22641
2 90308 1 22641
2 90309 1 22641
2 90310 1 22644
2 90311 1 22644
2 90312 1 22644
2 90313 1 22644
2 90314 1 22645
2 90315 1 22645
2 90316 1 22645
2 90317 1 22649
2 90318 1 22649
2 90319 1 22650
2 90320 1 22650
2 90321 1 22650
2 90322 1 22650
2 90323 1 22650
2 90324 1 22650
2 90325 1 22650
2 90326 1 22650
2 90327 1 22670
2 90328 1 22670
2 90329 1 22678
2 90330 1 22678
2 90331 1 22678
2 90332 1 22686
2 90333 1 22686
2 90334 1 22686
2 90335 1 22686
2 90336 1 22687
2 90337 1 22687
2 90338 1 22688
2 90339 1 22688
2 90340 1 22689
2 90341 1 22689
2 90342 1 22690
2 90343 1 22690
2 90344 1 22690
2 90345 1 22698
2 90346 1 22698
2 90347 1 22698
2 90348 1 22698
2 90349 1 22698
2 90350 1 22698
2 90351 1 22698
2 90352 1 22698
2 90353 1 22698
2 90354 1 22698
2 90355 1 22699
2 90356 1 22699
2 90357 1 22699
2 90358 1 22700
2 90359 1 22700
2 90360 1 22701
2 90361 1 22701
2 90362 1 22702
2 90363 1 22702
2 90364 1 22720
2 90365 1 22720
2 90366 1 22721
2 90367 1 22721
2 90368 1 22721
2 90369 1 22721
2 90370 1 22725
2 90371 1 22725
2 90372 1 22728
2 90373 1 22728
2 90374 1 22728
2 90375 1 22728
2 90376 1 22729
2 90377 1 22729
2 90378 1 22729
2 90379 1 22729
2 90380 1 22730
2 90381 1 22730
2 90382 1 22737
2 90383 1 22737
2 90384 1 22737
2 90385 1 22737
2 90386 1 22749
2 90387 1 22749
2 90388 1 22749
2 90389 1 22749
2 90390 1 22749
2 90391 1 22760
2 90392 1 22760
2 90393 1 22772
2 90394 1 22772
2 90395 1 22797
2 90396 1 22797
2 90397 1 22817
2 90398 1 22817
2 90399 1 22823
2 90400 1 22823
2 90401 1 22829
2 90402 1 22829
2 90403 1 22829
2 90404 1 22843
2 90405 1 22843
2 90406 1 22843
2 90407 1 22843
2 90408 1 22843
2 90409 1 22843
2 90410 1 22843
2 90411 1 22864
2 90412 1 22864
2 90413 1 22864
2 90414 1 22899
2 90415 1 22899
2 90416 1 22899
2 90417 1 22912
2 90418 1 22912
2 90419 1 22914
2 90420 1 22914
2 90421 1 22914
2 90422 1 22922
2 90423 1 22922
2 90424 1 22922
2 90425 1 22922
2 90426 1 22922
2 90427 1 22922
2 90428 1 22923
2 90429 1 22923
2 90430 1 22924
2 90431 1 22924
2 90432 1 22933
2 90433 1 22933
2 90434 1 22943
2 90435 1 22943
2 90436 1 22944
2 90437 1 22944
2 90438 1 22959
2 90439 1 22959
2 90440 1 22970
2 90441 1 22970
2 90442 1 22970
2 90443 1 22970
2 90444 1 22970
2 90445 1 22971
2 90446 1 22971
2 90447 1 23000
2 90448 1 23000
2 90449 1 23000
2 90450 1 23000
2 90451 1 23001
2 90452 1 23001
2 90453 1 23004
2 90454 1 23004
2 90455 1 23004
2 90456 1 23011
2 90457 1 23011
2 90458 1 23022
2 90459 1 23022
2 90460 1 23022
2 90461 1 23022
2 90462 1 23022
2 90463 1 23022
2 90464 1 23022
2 90465 1 23043
2 90466 1 23043
2 90467 1 23043
2 90468 1 23072
2 90469 1 23072
2 90470 1 23072
2 90471 1 23073
2 90472 1 23073
2 90473 1 23073
2 90474 1 23075
2 90475 1 23075
2 90476 1 23079
2 90477 1 23079
2 90478 1 23087
2 90479 1 23087
2 90480 1 23111
2 90481 1 23111
2 90482 1 23111
2 90483 1 23111
2 90484 1 23152
2 90485 1 23152
2 90486 1 23161
2 90487 1 23161
2 90488 1 23162
2 90489 1 23162
2 90490 1 23162
2 90491 1 23164
2 90492 1 23164
2 90493 1 23169
2 90494 1 23169
2 90495 1 23169
2 90496 1 23204
2 90497 1 23204
2 90498 1 23207
2 90499 1 23207
2 90500 1 23219
2 90501 1 23219
2 90502 1 23226
2 90503 1 23226
2 90504 1 23226
2 90505 1 23226
2 90506 1 23226
2 90507 1 23226
2 90508 1 23227
2 90509 1 23227
2 90510 1 23231
2 90511 1 23231
2 90512 1 23240
2 90513 1 23240
2 90514 1 23243
2 90515 1 23243
2 90516 1 23243
2 90517 1 23259
2 90518 1 23259
2 90519 1 23260
2 90520 1 23260
2 90521 1 23269
2 90522 1 23269
2 90523 1 23269
2 90524 1 23269
2 90525 1 23286
2 90526 1 23286
2 90527 1 23286
2 90528 1 23286
2 90529 1 23289
2 90530 1 23289
2 90531 1 23289
2 90532 1 23297
2 90533 1 23297
2 90534 1 23297
2 90535 1 23307
2 90536 1 23307
2 90537 1 23307
2 90538 1 23308
2 90539 1 23308
2 90540 1 23308
2 90541 1 23308
2 90542 1 23319
2 90543 1 23319
2 90544 1 23319
2 90545 1 23319
2 90546 1 23319
2 90547 1 23319
2 90548 1 23319
2 90549 1 23319
2 90550 1 23319
2 90551 1 23320
2 90552 1 23320
2 90553 1 23321
2 90554 1 23321
2 90555 1 23321
2 90556 1 23321
2 90557 1 23322
2 90558 1 23322
2 90559 1 23322
2 90560 1 23322
2 90561 1 23322
2 90562 1 23322
2 90563 1 23331
2 90564 1 23331
2 90565 1 23331
2 90566 1 23332
2 90567 1 23332
2 90568 1 23333
2 90569 1 23333
2 90570 1 23333
2 90571 1 23342
2 90572 1 23342
2 90573 1 23343
2 90574 1 23343
2 90575 1 23343
2 90576 1 23343
2 90577 1 23343
2 90578 1 23351
2 90579 1 23351
2 90580 1 23352
2 90581 1 23352
2 90582 1 23352
2 90583 1 23367
2 90584 1 23367
2 90585 1 23372
2 90586 1 23372
2 90587 1 23372
2 90588 1 23372
2 90589 1 23372
2 90590 1 23372
2 90591 1 23382
2 90592 1 23382
2 90593 1 23382
2 90594 1 23382
2 90595 1 23382
2 90596 1 23382
2 90597 1 23382
2 90598 1 23382
2 90599 1 23382
2 90600 1 23382
2 90601 1 23395
2 90602 1 23395
2 90603 1 23395
2 90604 1 23396
2 90605 1 23396
2 90606 1 23396
2 90607 1 23406
2 90608 1 23406
2 90609 1 23425
2 90610 1 23425
2 90611 1 23425
2 90612 1 23425
2 90613 1 23436
2 90614 1 23436
2 90615 1 23451
2 90616 1 23451
2 90617 1 23451
2 90618 1 23451
2 90619 1 23451
2 90620 1 23453
2 90621 1 23453
2 90622 1 23454
2 90623 1 23454
2 90624 1 23454
2 90625 1 23454
2 90626 1 23457
2 90627 1 23457
2 90628 1 23460
2 90629 1 23460
2 90630 1 23460
2 90631 1 23460
2 90632 1 23460
2 90633 1 23461
2 90634 1 23461
2 90635 1 23461
2 90636 1 23461
2 90637 1 23461
2 90638 1 23461
2 90639 1 23462
2 90640 1 23462
2 90641 1 23475
2 90642 1 23475
2 90643 1 23482
2 90644 1 23482
2 90645 1 23498
2 90646 1 23498
2 90647 1 23517
2 90648 1 23517
2 90649 1 23517
2 90650 1 23518
2 90651 1 23518
2 90652 1 23526
2 90653 1 23526
2 90654 1 23526
2 90655 1 23539
2 90656 1 23539
2 90657 1 23548
2 90658 1 23548
2 90659 1 23555
2 90660 1 23555
2 90661 1 23555
2 90662 1 23555
2 90663 1 23556
2 90664 1 23556
2 90665 1 23557
2 90666 1 23557
2 90667 1 23557
2 90668 1 23560
2 90669 1 23560
2 90670 1 23560
2 90671 1 23560
2 90672 1 23560
2 90673 1 23560
2 90674 1 23560
2 90675 1 23560
2 90676 1 23561
2 90677 1 23561
2 90678 1 23561
2 90679 1 23562
2 90680 1 23562
2 90681 1 23565
2 90682 1 23565
2 90683 1 23568
2 90684 1 23568
2 90685 1 23573
2 90686 1 23573
2 90687 1 23573
2 90688 1 23573
2 90689 1 23573
2 90690 1 23573
2 90691 1 23573
2 90692 1 23574
2 90693 1 23574
2 90694 1 23575
2 90695 1 23575
2 90696 1 23586
2 90697 1 23586
2 90698 1 23595
2 90699 1 23595
2 90700 1 23596
2 90701 1 23596
2 90702 1 23596
2 90703 1 23596
2 90704 1 23599
2 90705 1 23599
2 90706 1 23599
2 90707 1 23599
2 90708 1 23599
2 90709 1 23622
2 90710 1 23622
2 90711 1 23624
2 90712 1 23624
2 90713 1 23624
2 90714 1 23625
2 90715 1 23625
2 90716 1 23625
2 90717 1 23625
2 90718 1 23625
2 90719 1 23649
2 90720 1 23649
2 90721 1 23649
2 90722 1 23649
2 90723 1 23652
2 90724 1 23652
2 90725 1 23652
2 90726 1 23652
2 90727 1 23652
2 90728 1 23652
2 90729 1 23652
2 90730 1 23652
2 90731 1 23669
2 90732 1 23669
2 90733 1 23715
2 90734 1 23715
2 90735 1 23759
2 90736 1 23759
2 90737 1 23767
2 90738 1 23767
2 90739 1 23767
2 90740 1 23767
2 90741 1 23768
2 90742 1 23768
2 90743 1 23774
2 90744 1 23774
2 90745 1 23778
2 90746 1 23778
2 90747 1 23815
2 90748 1 23815
2 90749 1 23817
2 90750 1 23817
2 90751 1 23817
2 90752 1 23817
2 90753 1 23818
2 90754 1 23818
2 90755 1 23818
2 90756 1 23818
2 90757 1 23818
2 90758 1 23846
2 90759 1 23846
2 90760 1 23874
2 90761 1 23874
2 90762 1 23882
2 90763 1 23882
2 90764 1 23882
2 90765 1 23882
2 90766 1 23882
2 90767 1 23890
2 90768 1 23890
2 90769 1 23890
2 90770 1 23890
2 90771 1 23890
2 90772 1 23891
2 90773 1 23891
2 90774 1 23902
2 90775 1 23902
2 90776 1 23931
2 90777 1 23931
2 90778 1 23931
2 90779 1 23934
2 90780 1 23934
2 90781 1 23935
2 90782 1 23935
2 90783 1 23945
2 90784 1 23945
2 90785 1 23945
2 90786 1 23946
2 90787 1 23946
2 90788 1 23947
2 90789 1 23947
2 90790 1 23947
2 90791 1 23947
2 90792 1 23947
2 90793 1 23947
2 90794 1 23947
2 90795 1 23947
2 90796 1 23947
2 90797 1 23950
2 90798 1 23950
2 90799 1 23961
2 90800 1 23961
2 90801 1 23961
2 90802 1 23961
2 90803 1 23961
2 90804 1 23963
2 90805 1 23963
2 90806 1 23963
2 90807 1 23963
2 90808 1 23963
2 90809 1 23963
2 90810 1 23963
2 90811 1 23964
2 90812 1 23964
2 90813 1 23964
2 90814 1 23964
2 90815 1 23976
2 90816 1 23976
2 90817 1 23976
2 90818 1 23979
2 90819 1 23979
2 90820 1 23979
2 90821 1 23997
2 90822 1 23997
2 90823 1 23997
2 90824 1 23997
2 90825 1 23997
2 90826 1 23998
2 90827 1 23998
2 90828 1 23999
2 90829 1 23999
2 90830 1 23999
2 90831 1 23999
2 90832 1 24001
2 90833 1 24001
2 90834 1 24005
2 90835 1 24005
2 90836 1 24005
2 90837 1 24005
2 90838 1 24005
2 90839 1 24006
2 90840 1 24006
2 90841 1 24006
2 90842 1 24011
2 90843 1 24011
2 90844 1 24015
2 90845 1 24015
2 90846 1 24015
2 90847 1 24015
2 90848 1 24016
2 90849 1 24016
2 90850 1 24016
2 90851 1 24016
2 90852 1 24016
2 90853 1 24027
2 90854 1 24027
2 90855 1 24028
2 90856 1 24028
2 90857 1 24028
2 90858 1 24028
2 90859 1 24029
2 90860 1 24029
2 90861 1 24030
2 90862 1 24030
2 90863 1 24038
2 90864 1 24038
2 90865 1 24038
2 90866 1 24038
2 90867 1 24047
2 90868 1 24047
2 90869 1 24047
2 90870 1 24055
2 90871 1 24055
2 90872 1 24069
2 90873 1 24069
2 90874 1 24084
2 90875 1 24084
2 90876 1 24092
2 90877 1 24092
2 90878 1 24107
2 90879 1 24107
2 90880 1 24109
2 90881 1 24109
2 90882 1 24109
2 90883 1 24109
2 90884 1 24116
2 90885 1 24116
2 90886 1 24116
2 90887 1 24120
2 90888 1 24120
2 90889 1 24120
2 90890 1 24122
2 90891 1 24122
2 90892 1 24141
2 90893 1 24141
2 90894 1 24164
2 90895 1 24164
2 90896 1 24164
2 90897 1 24164
2 90898 1 24164
2 90899 1 24164
2 90900 1 24165
2 90901 1 24165
2 90902 1 24165
2 90903 1 24166
2 90904 1 24166
2 90905 1 24169
2 90906 1 24169
2 90907 1 24174
2 90908 1 24174
2 90909 1 24186
2 90910 1 24186
2 90911 1 24187
2 90912 1 24187
2 90913 1 24188
2 90914 1 24188
2 90915 1 24188
2 90916 1 24188
2 90917 1 24188
2 90918 1 24188
2 90919 1 24190
2 90920 1 24190
2 90921 1 24197
2 90922 1 24197
2 90923 1 24217
2 90924 1 24217
2 90925 1 24229
2 90926 1 24229
2 90927 1 24231
2 90928 1 24231
2 90929 1 24232
2 90930 1 24232
2 90931 1 24232
2 90932 1 24232
2 90933 1 24232
2 90934 1 24232
2 90935 1 24232
2 90936 1 24232
2 90937 1 24239
2 90938 1 24239
2 90939 1 24241
2 90940 1 24241
2 90941 1 24244
2 90942 1 24244
2 90943 1 24245
2 90944 1 24245
2 90945 1 24245
2 90946 1 24253
2 90947 1 24253
2 90948 1 24254
2 90949 1 24254
2 90950 1 24255
2 90951 1 24255
2 90952 1 24255
2 90953 1 24255
2 90954 1 24266
2 90955 1 24266
2 90956 1 24272
2 90957 1 24272
2 90958 1 24291
2 90959 1 24291
2 90960 1 24293
2 90961 1 24293
2 90962 1 24293
2 90963 1 24293
2 90964 1 24306
2 90965 1 24306
2 90966 1 24342
2 90967 1 24342
2 90968 1 24344
2 90969 1 24344
2 90970 1 24344
2 90971 1 24344
2 90972 1 24344
2 90973 1 24344
2 90974 1 24349
2 90975 1 24349
2 90976 1 24350
2 90977 1 24350
2 90978 1 24350
2 90979 1 24350
2 90980 1 24351
2 90981 1 24351
2 90982 1 24351
2 90983 1 24351
2 90984 1 24352
2 90985 1 24352
2 90986 1 24353
2 90987 1 24353
2 90988 1 24368
2 90989 1 24368
2 90990 1 24368
2 90991 1 24368
2 90992 1 24368
2 90993 1 24368
2 90994 1 24368
2 90995 1 24369
2 90996 1 24369
2 90997 1 24369
2 90998 1 24369
2 90999 1 24377
2 91000 1 24377
2 91001 1 24377
2 91002 1 24377
2 91003 1 24377
2 91004 1 24388
2 91005 1 24388
2 91006 1 24388
2 91007 1 24388
2 91008 1 24411
2 91009 1 24411
2 91010 1 24411
2 91011 1 24414
2 91012 1 24414
2 91013 1 24415
2 91014 1 24415
2 91015 1 24415
2 91016 1 24423
2 91017 1 24423
2 91018 1 24428
2 91019 1 24428
2 91020 1 24445
2 91021 1 24445
2 91022 1 24446
2 91023 1 24446
2 91024 1 24446
2 91025 1 24447
2 91026 1 24447
2 91027 1 24464
2 91028 1 24464
2 91029 1 24473
2 91030 1 24473
2 91031 1 24473
2 91032 1 24473
2 91033 1 24475
2 91034 1 24475
2 91035 1 24486
2 91036 1 24486
2 91037 1 24505
2 91038 1 24505
2 91039 1 24505
2 91040 1 24509
2 91041 1 24509
2 91042 1 24519
2 91043 1 24519
2 91044 1 24538
2 91045 1 24538
2 91046 1 24546
2 91047 1 24546
2 91048 1 24546
2 91049 1 24551
2 91050 1 24551
2 91051 1 24572
2 91052 1 24572
2 91053 1 24580
2 91054 1 24580
2 91055 1 24581
2 91056 1 24581
2 91057 1 24581
2 91058 1 24586
2 91059 1 24586
2 91060 1 24586
2 91061 1 24600
2 91062 1 24600
2 91063 1 24601
2 91064 1 24601
2 91065 1 24603
2 91066 1 24603
2 91067 1 24620
2 91068 1 24620
2 91069 1 24621
2 91070 1 24621
2 91071 1 24637
2 91072 1 24637
2 91073 1 24637
2 91074 1 24638
2 91075 1 24638
2 91076 1 24645
2 91077 1 24645
2 91078 1 24649
2 91079 1 24649
2 91080 1 24649
2 91081 1 24649
2 91082 1 24657
2 91083 1 24657
2 91084 1 24670
2 91085 1 24670
2 91086 1 24707
2 91087 1 24707
2 91088 1 24707
2 91089 1 24711
2 91090 1 24711
2 91091 1 24711
2 91092 1 24719
2 91093 1 24719
2 91094 1 24738
2 91095 1 24738
2 91096 1 24739
2 91097 1 24739
2 91098 1 24740
2 91099 1 24740
2 91100 1 24740
2 91101 1 24777
2 91102 1 24777
2 91103 1 24778
2 91104 1 24778
2 91105 1 24803
2 91106 1 24803
2 91107 1 24803
2 91108 1 24803
2 91109 1 24803
2 91110 1 24805
2 91111 1 24805
2 91112 1 24806
2 91113 1 24806
2 91114 1 24806
2 91115 1 24806
2 91116 1 24806
2 91117 1 24819
2 91118 1 24819
2 91119 1 24819
2 91120 1 24819
2 91121 1 24819
2 91122 1 24819
2 91123 1 24820
2 91124 1 24820
2 91125 1 24836
2 91126 1 24836
2 91127 1 24855
2 91128 1 24855
2 91129 1 24873
2 91130 1 24873
2 91131 1 24873
2 91132 1 24873
2 91133 1 24873
2 91134 1 24873
2 91135 1 24882
2 91136 1 24882
2 91137 1 24882
2 91138 1 24882
2 91139 1 24882
2 91140 1 24882
2 91141 1 24882
2 91142 1 24882
2 91143 1 24897
2 91144 1 24897
2 91145 1 24897
2 91146 1 24900
2 91147 1 24900
2 91148 1 24900
2 91149 1 24900
2 91150 1 24900
2 91151 1 24901
2 91152 1 24901
2 91153 1 24901
2 91154 1 24901
2 91155 1 24903
2 91156 1 24903
2 91157 1 24903
2 91158 1 24910
2 91159 1 24910
2 91160 1 24918
2 91161 1 24918
2 91162 1 24918
2 91163 1 24930
2 91164 1 24930
2 91165 1 24947
2 91166 1 24947
2 91167 1 24962
2 91168 1 24962
2 91169 1 24975
2 91170 1 24975
2 91171 1 24986
2 91172 1 24986
2 91173 1 24995
2 91174 1 24995
2 91175 1 24995
2 91176 1 25021
2 91177 1 25021
2 91178 1 25021
2 91179 1 25022
2 91180 1 25022
2 91181 1 25022
2 91182 1 25022
2 91183 1 25022
2 91184 1 25022
2 91185 1 25022
2 91186 1 25051
2 91187 1 25051
2 91188 1 25070
2 91189 1 25070
2 91190 1 25080
2 91191 1 25080
2 91192 1 25085
2 91193 1 25085
2 91194 1 25086
2 91195 1 25086
2 91196 1 25087
2 91197 1 25087
2 91198 1 25112
2 91199 1 25112
2 91200 1 25143
2 91201 1 25143
2 91202 1 25150
2 91203 1 25150
2 91204 1 25151
2 91205 1 25151
2 91206 1 25151
2 91207 1 25152
2 91208 1 25152
2 91209 1 25152
2 91210 1 25153
2 91211 1 25153
2 91212 1 25162
2 91213 1 25162
2 91214 1 25165
2 91215 1 25165
2 91216 1 25165
2 91217 1 25165
2 91218 1 25165
2 91219 1 25169
2 91220 1 25169
2 91221 1 25170
2 91222 1 25170
2 91223 1 25170
2 91224 1 25196
2 91225 1 25196
2 91226 1 25202
2 91227 1 25202
2 91228 1 25216
2 91229 1 25216
2 91230 1 25216
2 91231 1 25216
2 91232 1 25216
2 91233 1 25217
2 91234 1 25217
2 91235 1 25217
2 91236 1 25217
2 91237 1 25218
2 91238 1 25218
2 91239 1 25219
2 91240 1 25219
2 91241 1 25235
2 91242 1 25235
2 91243 1 25264
2 91244 1 25264
2 91245 1 25264
2 91246 1 25264
2 91247 1 25264
2 91248 1 25264
2 91249 1 25264
2 91250 1 25264
2 91251 1 25264
2 91252 1 25265
2 91253 1 25265
2 91254 1 25278
2 91255 1 25278
2 91256 1 25278
2 91257 1 25278
2 91258 1 25292
2 91259 1 25292
2 91260 1 25293
2 91261 1 25293
2 91262 1 25295
2 91263 1 25295
2 91264 1 25298
2 91265 1 25298
2 91266 1 25319
2 91267 1 25319
2 91268 1 25319
2 91269 1 25333
2 91270 1 25333
2 91271 1 25333
2 91272 1 25336
2 91273 1 25336
2 91274 1 25336
2 91275 1 25336
2 91276 1 25339
2 91277 1 25339
2 91278 1 25339
2 91279 1 25344
2 91280 1 25344
2 91281 1 25344
2 91282 1 25345
2 91283 1 25345
2 91284 1 25345
2 91285 1 25357
2 91286 1 25357
2 91287 1 25358
2 91288 1 25358
2 91289 1 25358
2 91290 1 25358
2 91291 1 25368
2 91292 1 25368
2 91293 1 25369
2 91294 1 25369
2 91295 1 25370
2 91296 1 25370
2 91297 1 25370
2 91298 1 25370
2 91299 1 25374
2 91300 1 25374
2 91301 1 25374
2 91302 1 25375
2 91303 1 25375
2 91304 1 25375
2 91305 1 25383
2 91306 1 25383
2 91307 1 25384
2 91308 1 25384
2 91309 1 25388
2 91310 1 25388
2 91311 1 25388
2 91312 1 25389
2 91313 1 25389
2 91314 1 25389
2 91315 1 25390
2 91316 1 25390
2 91317 1 25407
2 91318 1 25407
2 91319 1 25407
2 91320 1 25407
2 91321 1 25407
2 91322 1 25407
2 91323 1 25426
2 91324 1 25426
2 91325 1 25431
2 91326 1 25431
2 91327 1 25437
2 91328 1 25437
2 91329 1 25437
2 91330 1 25437
2 91331 1 25447
2 91332 1 25447
2 91333 1 25486
2 91334 1 25486
2 91335 1 25496
2 91336 1 25496
2 91337 1 25499
2 91338 1 25499
2 91339 1 25499
2 91340 1 25500
2 91341 1 25500
2 91342 1 25526
2 91343 1 25526
2 91344 1 25530
2 91345 1 25530
2 91346 1 25532
2 91347 1 25532
2 91348 1 25569
2 91349 1 25569
2 91350 1 25590
2 91351 1 25590
2 91352 1 25590
2 91353 1 25590
2 91354 1 25599
2 91355 1 25599
2 91356 1 25613
2 91357 1 25613
2 91358 1 25613
2 91359 1 25629
2 91360 1 25629
2 91361 1 25629
2 91362 1 25629
2 91363 1 25645
2 91364 1 25645
2 91365 1 25645
2 91366 1 25649
2 91367 1 25649
2 91368 1 25650
2 91369 1 25650
2 91370 1 25650
2 91371 1 25650
2 91372 1 25650
2 91373 1 25652
2 91374 1 25652
2 91375 1 25652
2 91376 1 25652
2 91377 1 25652
2 91378 1 25652
2 91379 1 25667
2 91380 1 25667
2 91381 1 25668
2 91382 1 25668
2 91383 1 25668
2 91384 1 25679
2 91385 1 25679
2 91386 1 25692
2 91387 1 25692
2 91388 1 25693
2 91389 1 25693
2 91390 1 25697
2 91391 1 25697
2 91392 1 25697
2 91393 1 25716
2 91394 1 25716
2 91395 1 25717
2 91396 1 25717
2 91397 1 25724
2 91398 1 25724
2 91399 1 25724
2 91400 1 25732
2 91401 1 25732
2 91402 1 25732
2 91403 1 25759
2 91404 1 25759
2 91405 1 25767
2 91406 1 25767
2 91407 1 25768
2 91408 1 25768
2 91409 1 25769
2 91410 1 25769
2 91411 1 25769
2 91412 1 25769
2 91413 1 25769
2 91414 1 25769
2 91415 1 25781
2 91416 1 25781
2 91417 1 25781
2 91418 1 25781
2 91419 1 25781
2 91420 1 25782
2 91421 1 25782
2 91422 1 25782
2 91423 1 25794
2 91424 1 25794
2 91425 1 25794
2 91426 1 25819
2 91427 1 25819
2 91428 1 25819
2 91429 1 25840
2 91430 1 25840
2 91431 1 25840
2 91432 1 25841
2 91433 1 25841
2 91434 1 25849
2 91435 1 25849
2 91436 1 25865
2 91437 1 25865
2 91438 1 25874
2 91439 1 25874
2 91440 1 25875
2 91441 1 25875
2 91442 1 25877
2 91443 1 25877
2 91444 1 25889
2 91445 1 25889
2 91446 1 25902
2 91447 1 25902
2 91448 1 25915
2 91449 1 25915
2 91450 1 25915
2 91451 1 25915
2 91452 1 25924
2 91453 1 25924
2 91454 1 25924
2 91455 1 25924
2 91456 1 25932
2 91457 1 25932
2 91458 1 25932
2 91459 1 25932
2 91460 1 25933
2 91461 1 25933
2 91462 1 25933
2 91463 1 25947
2 91464 1 25947
2 91465 1 25947
2 91466 1 25954
2 91467 1 25954
2 91468 1 25954
2 91469 1 25969
2 91470 1 25969
2 91471 1 25970
2 91472 1 25970
2 91473 1 25970
2 91474 1 25970
2 91475 1 25970
2 91476 1 25988
2 91477 1 25988
2 91478 1 25993
2 91479 1 25993
2 91480 1 25994
2 91481 1 25994
2 91482 1 26000
2 91483 1 26000
2 91484 1 26000
2 91485 1 26000
2 91486 1 26000
2 91487 1 26000
2 91488 1 26010
2 91489 1 26010
2 91490 1 26027
2 91491 1 26027
2 91492 1 26027
2 91493 1 26030
2 91494 1 26030
2 91495 1 26030
2 91496 1 26038
2 91497 1 26038
2 91498 1 26038
2 91499 1 26106
2 91500 1 26106
2 91501 1 26109
2 91502 1 26109
2 91503 1 26112
2 91504 1 26112
2 91505 1 26129
2 91506 1 26129
2 91507 1 26144
2 91508 1 26144
2 91509 1 26147
2 91510 1 26147
2 91511 1 26147
2 91512 1 26147
2 91513 1 26148
2 91514 1 26148
2 91515 1 26151
2 91516 1 26151
2 91517 1 26155
2 91518 1 26155
2 91519 1 26155
2 91520 1 26163
2 91521 1 26163
2 91522 1 26176
2 91523 1 26176
2 91524 1 26184
2 91525 1 26184
2 91526 1 26184
2 91527 1 26195
2 91528 1 26195
2 91529 1 26195
2 91530 1 26196
2 91531 1 26196
2 91532 1 26204
2 91533 1 26204
2 91534 1 26221
2 91535 1 26221
2 91536 1 26232
2 91537 1 26232
2 91538 1 26240
2 91539 1 26240
2 91540 1 26241
2 91541 1 26241
2 91542 1 26241
2 91543 1 26287
2 91544 1 26287
2 91545 1 26301
2 91546 1 26301
2 91547 1 26301
2 91548 1 26331
2 91549 1 26331
2 91550 1 26331
2 91551 1 26337
2 91552 1 26337
2 91553 1 26365
2 91554 1 26365
2 91555 1 26367
2 91556 1 26367
2 91557 1 26379
2 91558 1 26379
2 91559 1 26379
2 91560 1 26400
2 91561 1 26400
2 91562 1 26400
2 91563 1 26402
2 91564 1 26402
2 91565 1 26463
2 91566 1 26463
2 91567 1 26468
2 91568 1 26468
2 91569 1 26489
2 91570 1 26489
2 91571 1 26502
2 91572 1 26502
2 91573 1 26502
2 91574 1 26503
2 91575 1 26503
2 91576 1 26511
2 91577 1 26511
2 91578 1 26517
2 91579 1 26517
2 91580 1 26525
2 91581 1 26525
2 91582 1 26541
2 91583 1 26541
2 91584 1 26541
2 91585 1 26544
2 91586 1 26544
2 91587 1 26547
2 91588 1 26547
2 91589 1 26547
2 91590 1 26547
2 91591 1 26547
2 91592 1 26554
2 91593 1 26554
2 91594 1 26554
2 91595 1 26554
2 91596 1 26554
2 91597 1 26574
2 91598 1 26574
2 91599 1 26575
2 91600 1 26575
2 91601 1 26584
2 91602 1 26584
2 91603 1 26585
2 91604 1 26585
2 91605 1 26585
2 91606 1 26599
2 91607 1 26599
2 91608 1 26614
2 91609 1 26614
2 91610 1 26649
2 91611 1 26649
2 91612 1 26649
2 91613 1 26656
2 91614 1 26656
2 91615 1 26665
2 91616 1 26665
2 91617 1 26692
2 91618 1 26692
2 91619 1 26696
2 91620 1 26696
2 91621 1 26698
2 91622 1 26698
2 91623 1 26706
2 91624 1 26706
2 91625 1 26727
2 91626 1 26727
2 91627 1 26729
2 91628 1 26729
2 91629 1 26729
2 91630 1 26808
2 91631 1 26808
2 91632 1 26866
2 91633 1 26866
2 91634 1 26866
2 91635 1 26869
2 91636 1 26869
2 91637 1 26870
2 91638 1 26870
2 91639 1 26905
2 91640 1 26905
2 91641 1 26905
2 91642 1 26905
2 91643 1 26906
2 91644 1 26906
2 91645 1 26906
2 91646 1 26907
2 91647 1 26907
2 91648 1 26922
2 91649 1 26922
2 91650 1 26936
2 91651 1 26936
2 91652 1 26967
2 91653 1 26967
2 91654 1 26967
2 91655 1 26967
2 91656 1 26967
2 91657 1 26967
2 91658 1 26967
2 91659 1 26967
2 91660 1 26967
2 91661 1 26976
2 91662 1 26976
2 91663 1 26976
2 91664 1 26976
2 91665 1 26976
2 91666 1 26980
2 91667 1 26980
2 91668 1 26982
2 91669 1 26982
2 91670 1 26982
2 91671 1 26982
2 91672 1 26998
2 91673 1 26998
2 91674 1 27005
2 91675 1 27005
2 91676 1 27005
2 91677 1 27024
2 91678 1 27024
2 91679 1 27024
2 91680 1 27024
2 91681 1 27038
2 91682 1 27038
2 91683 1 27046
2 91684 1 27046
2 91685 1 27046
2 91686 1 27057
2 91687 1 27057
2 91688 1 27071
2 91689 1 27071
2 91690 1 27078
2 91691 1 27078
2 91692 1 27084
2 91693 1 27084
2 91694 1 27112
2 91695 1 27112
2 91696 1 27131
2 91697 1 27131
2 91698 1 27148
2 91699 1 27148
2 91700 1 27148
2 91701 1 27149
2 91702 1 27149
2 91703 1 27149
2 91704 1 27153
2 91705 1 27153
2 91706 1 27168
2 91707 1 27168
2 91708 1 27171
2 91709 1 27171
2 91710 1 27187
2 91711 1 27187
2 91712 1 27193
2 91713 1 27193
2 91714 1 27200
2 91715 1 27200
2 91716 1 27200
2 91717 1 27200
2 91718 1 27200
2 91719 1 27201
2 91720 1 27201
2 91721 1 27204
2 91722 1 27204
2 91723 1 27204
2 91724 1 27232
2 91725 1 27232
2 91726 1 27239
2 91727 1 27239
2 91728 1 27239
2 91729 1 27240
2 91730 1 27240
2 91731 1 27269
2 91732 1 27269
2 91733 1 27286
2 91734 1 27286
2 91735 1 27300
2 91736 1 27300
2 91737 1 27301
2 91738 1 27301
2 91739 1 27301
2 91740 1 27311
2 91741 1 27311
2 91742 1 27311
2 91743 1 27312
2 91744 1 27312
2 91745 1 27312
2 91746 1 27312
2 91747 1 27328
2 91748 1 27328
2 91749 1 27328
2 91750 1 27336
2 91751 1 27336
2 91752 1 27336
2 91753 1 27364
2 91754 1 27364
2 91755 1 27364
2 91756 1 27364
2 91757 1 27364
2 91758 1 27364
2 91759 1 27364
2 91760 1 27365
2 91761 1 27365
2 91762 1 27365
2 91763 1 27370
2 91764 1 27370
2 91765 1 27398
2 91766 1 27398
2 91767 1 27398
2 91768 1 27399
2 91769 1 27399
2 91770 1 27412
2 91771 1 27412
2 91772 1 27412
2 91773 1 27412
2 91774 1 27413
2 91775 1 27413
2 91776 1 27413
2 91777 1 27413
2 91778 1 27413
2 91779 1 27413
2 91780 1 27413
2 91781 1 27423
2 91782 1 27423
2 91783 1 27423
2 91784 1 27423
2 91785 1 27423
2 91786 1 27423
2 91787 1 27423
2 91788 1 27423
2 91789 1 27424
2 91790 1 27424
2 91791 1 27445
2 91792 1 27445
2 91793 1 27452
2 91794 1 27452
2 91795 1 27452
2 91796 1 27452
2 91797 1 27452
2 91798 1 27452
2 91799 1 27452
2 91800 1 27452
2 91801 1 27464
2 91802 1 27464
2 91803 1 27464
2 91804 1 27478
2 91805 1 27478
2 91806 1 27489
2 91807 1 27489
2 91808 1 27562
2 91809 1 27562
2 91810 1 27582
2 91811 1 27582
2 91812 1 27589
2 91813 1 27589
2 91814 1 27599
2 91815 1 27599
2 91816 1 27611
2 91817 1 27611
2 91818 1 27616
2 91819 1 27616
2 91820 1 27632
2 91821 1 27632
2 91822 1 27650
2 91823 1 27650
2 91824 1 27650
2 91825 1 27650
2 91826 1 27650
2 91827 1 27650
2 91828 1 27650
2 91829 1 27650
2 91830 1 27650
2 91831 1 27650
2 91832 1 27650
2 91833 1 27650
2 91834 1 27676
2 91835 1 27676
2 91836 1 27676
2 91837 1 27689
2 91838 1 27689
2 91839 1 27703
2 91840 1 27703
2 91841 1 27703
2 91842 1 27703
2 91843 1 27703
2 91844 1 27717
2 91845 1 27717
2 91846 1 27725
2 91847 1 27725
2 91848 1 27727
2 91849 1 27727
2 91850 1 27727
2 91851 1 27727
2 91852 1 27727
2 91853 1 27770
2 91854 1 27770
2 91855 1 27776
2 91856 1 27776
2 91857 1 27776
2 91858 1 27783
2 91859 1 27783
2 91860 1 27789
2 91861 1 27789
2 91862 1 27797
2 91863 1 27797
2 91864 1 27798
2 91865 1 27798
2 91866 1 27811
2 91867 1 27811
2 91868 1 27848
2 91869 1 27848
2 91870 1 27849
2 91871 1 27849
2 91872 1 27852
2 91873 1 27852
2 91874 1 27853
2 91875 1 27853
2 91876 1 27853
2 91877 1 27853
2 91878 1 27853
2 91879 1 27866
2 91880 1 27866
2 91881 1 27866
2 91882 1 27866
2 91883 1 27875
2 91884 1 27875
2 91885 1 27875
2 91886 1 27877
2 91887 1 27877
2 91888 1 27879
2 91889 1 27879
2 91890 1 27883
2 91891 1 27883
2 91892 1 27895
2 91893 1 27895
2 91894 1 27900
2 91895 1 27900
2 91896 1 27912
2 91897 1 27912
2 91898 1 27912
2 91899 1 27916
2 91900 1 27916
2 91901 1 27916
2 91902 1 27917
2 91903 1 27917
2 91904 1 27937
2 91905 1 27937
2 91906 1 27937
2 91907 1 27937
2 91908 1 27944
2 91909 1 27944
2 91910 1 27955
2 91911 1 27955
2 91912 1 27956
2 91913 1 27956
2 91914 1 27963
2 91915 1 27963
2 91916 1 27974
2 91917 1 27974
2 91918 1 27982
2 91919 1 27982
2 91920 1 28004
2 91921 1 28004
2 91922 1 28016
2 91923 1 28016
2 91924 1 28035
2 91925 1 28035
2 91926 1 28036
2 91927 1 28036
2 91928 1 28036
2 91929 1 28037
2 91930 1 28037
2 91931 1 28040
2 91932 1 28040
2 91933 1 28050
2 91934 1 28050
2 91935 1 28072
2 91936 1 28072
2 91937 1 28092
2 91938 1 28092
2 91939 1 28095
2 91940 1 28095
2 91941 1 28105
2 91942 1 28105
2 91943 1 28105
2 91944 1 28105
2 91945 1 28106
2 91946 1 28106
2 91947 1 28111
2 91948 1 28111
2 91949 1 28119
2 91950 1 28119
2 91951 1 28122
2 91952 1 28122
2 91953 1 28122
2 91954 1 28130
2 91955 1 28130
2 91956 1 28135
2 91957 1 28135
2 91958 1 28153
2 91959 1 28153
2 91960 1 28156
2 91961 1 28156
2 91962 1 28185
2 91963 1 28185
2 91964 1 28185
2 91965 1 28185
2 91966 1 28185
2 91967 1 28192
2 91968 1 28192
2 91969 1 28192
2 91970 1 28192
2 91971 1 28192
2 91972 1 28192
2 91973 1 28193
2 91974 1 28193
2 91975 1 28193
2 91976 1 28206
2 91977 1 28206
2 91978 1 28206
2 91979 1 28210
2 91980 1 28210
2 91981 1 28265
2 91982 1 28265
2 91983 1 28280
2 91984 1 28280
2 91985 1 28288
2 91986 1 28288
2 91987 1 28295
2 91988 1 28295
2 91989 1 28328
2 91990 1 28328
2 91991 1 28332
2 91992 1 28332
2 91993 1 28332
2 91994 1 28332
2 91995 1 28332
2 91996 1 28333
2 91997 1 28333
2 91998 1 28344
2 91999 1 28344
2 92000 1 28344
2 92001 1 28344
2 92002 1 28361
2 92003 1 28361
2 92004 1 28378
2 92005 1 28378
2 92006 1 28399
2 92007 1 28399
2 92008 1 28419
2 92009 1 28419
2 92010 1 28458
2 92011 1 28458
2 92012 1 28489
2 92013 1 28489
2 92014 1 28489
2 92015 1 28489
2 92016 1 28490
2 92017 1 28490
2 92018 1 28490
2 92019 1 28491
2 92020 1 28491
2 92021 1 28492
2 92022 1 28492
2 92023 1 28511
2 92024 1 28511
2 92025 1 28526
2 92026 1 28526
2 92027 1 28534
2 92028 1 28534
2 92029 1 28535
2 92030 1 28535
2 92031 1 28535
2 92032 1 28537
2 92033 1 28537
2 92034 1 28537
2 92035 1 28537
2 92036 1 28537
2 92037 1 28538
2 92038 1 28538
2 92039 1 28541
2 92040 1 28541
2 92041 1 28541
2 92042 1 28541
2 92043 1 28557
2 92044 1 28557
2 92045 1 28557
2 92046 1 28570
2 92047 1 28570
2 92048 1 28570
2 92049 1 28570
2 92050 1 28570
2 92051 1 28572
2 92052 1 28572
2 92053 1 28572
2 92054 1 28572
2 92055 1 28573
2 92056 1 28573
2 92057 1 28584
2 92058 1 28584
2 92059 1 28584
2 92060 1 28584
2 92061 1 28593
2 92062 1 28593
2 92063 1 28594
2 92064 1 28594
2 92065 1 28608
2 92066 1 28608
2 92067 1 28608
2 92068 1 28608
2 92069 1 28612
2 92070 1 28612
2 92071 1 28632
2 92072 1 28632
2 92073 1 28632
2 92074 1 28632
2 92075 1 28650
2 92076 1 28650
2 92077 1 28683
2 92078 1 28683
2 92079 1 28684
2 92080 1 28684
2 92081 1 28686
2 92082 1 28686
2 92083 1 28686
2 92084 1 28697
2 92085 1 28697
2 92086 1 28714
2 92087 1 28714
2 92088 1 28714
2 92089 1 28722
2 92090 1 28722
2 92091 1 28723
2 92092 1 28723
2 92093 1 28733
2 92094 1 28733
2 92095 1 28740
2 92096 1 28740
2 92097 1 28756
2 92098 1 28756
2 92099 1 28756
2 92100 1 28769
2 92101 1 28769
2 92102 1 28769
2 92103 1 28769
2 92104 1 28769
2 92105 1 28769
2 92106 1 28806
2 92107 1 28806
2 92108 1 28896
2 92109 1 28896
2 92110 1 28927
2 92111 1 28927
2 92112 1 28933
2 92113 1 28933
2 92114 1 28969
2 92115 1 28969
2 92116 1 29015
2 92117 1 29015
2 92118 1 29026
2 92119 1 29026
2 92120 1 29039
2 92121 1 29039
2 92122 1 29061
2 92123 1 29061
2 92124 1 29066
2 92125 1 29066
2 92126 1 29079
2 92127 1 29079
2 92128 1 29086
2 92129 1 29086
2 92130 1 29105
2 92131 1 29105
2 92132 1 29114
2 92133 1 29114
2 92134 1 29121
2 92135 1 29121
2 92136 1 29159
2 92137 1 29159
2 92138 1 29161
2 92139 1 29161
2 92140 1 29161
2 92141 1 29171
2 92142 1 29171
2 92143 1 29171
2 92144 1 29171
2 92145 1 29217
2 92146 1 29217
2 92147 1 29222
2 92148 1 29222
2 92149 1 29222
2 92150 1 29222
2 92151 1 29222
2 92152 1 29243
2 92153 1 29243
2 92154 1 29243
2 92155 1 29243
2 92156 1 29243
2 92157 1 29243
2 92158 1 29243
2 92159 1 29243
2 92160 1 29243
2 92161 1 29244
2 92162 1 29244
2 92163 1 29244
2 92164 1 29245
2 92165 1 29245
2 92166 1 29245
2 92167 1 29246
2 92168 1 29246
2 92169 1 29246
2 92170 1 29254
2 92171 1 29254
2 92172 1 29255
2 92173 1 29255
2 92174 1 29279
2 92175 1 29279
2 92176 1 29298
2 92177 1 29298
2 92178 1 29298
2 92179 1 29298
2 92180 1 29298
2 92181 1 29300
2 92182 1 29300
2 92183 1 29300
2 92184 1 29300
2 92185 1 29301
2 92186 1 29301
2 92187 1 29308
2 92188 1 29308
2 92189 1 29322
2 92190 1 29322
2 92191 1 29330
2 92192 1 29330
2 92193 1 29378
2 92194 1 29378
2 92195 1 29378
2 92196 1 29378
2 92197 1 29384
2 92198 1 29384
2 92199 1 29419
2 92200 1 29419
2 92201 1 29420
2 92202 1 29420
2 92203 1 29420
2 92204 1 29420
2 92205 1 29420
2 92206 1 29420
2 92207 1 29421
2 92208 1 29421
2 92209 1 29440
2 92210 1 29440
2 92211 1 29452
2 92212 1 29452
2 92213 1 29452
2 92214 1 29456
2 92215 1 29456
2 92216 1 29456
2 92217 1 29456
2 92218 1 29456
2 92219 1 29470
2 92220 1 29470
2 92221 1 29471
2 92222 1 29471
2 92223 1 29474
2 92224 1 29474
2 92225 1 29474
2 92226 1 29474
2 92227 1 29482
2 92228 1 29482
2 92229 1 29483
2 92230 1 29483
2 92231 1 29483
2 92232 1 29486
2 92233 1 29486
2 92234 1 29499
2 92235 1 29499
2 92236 1 29500
2 92237 1 29500
2 92238 1 29500
2 92239 1 29508
2 92240 1 29508
2 92241 1 29516
2 92242 1 29516
2 92243 1 29524
2 92244 1 29524
2 92245 1 29524
2 92246 1 29564
2 92247 1 29564
2 92248 1 29575
2 92249 1 29575
2 92250 1 29593
2 92251 1 29593
2 92252 1 29600
2 92253 1 29600
2 92254 1 29612
2 92255 1 29612
2 92256 1 29620
2 92257 1 29620
2 92258 1 29620
2 92259 1 29620
2 92260 1 29622
2 92261 1 29622
2 92262 1 29634
2 92263 1 29634
2 92264 1 29634
2 92265 1 29634
2 92266 1 29634
2 92267 1 29634
2 92268 1 29634
2 92269 1 29634
2 92270 1 29634
2 92271 1 29636
2 92272 1 29636
2 92273 1 29636
2 92274 1 29636
2 92275 1 29636
2 92276 1 29688
2 92277 1 29688
2 92278 1 29688
2 92279 1 29709
2 92280 1 29709
2 92281 1 29718
2 92282 1 29718
2 92283 1 29731
2 92284 1 29731
2 92285 1 29731
2 92286 1 29738
2 92287 1 29738
2 92288 1 29746
2 92289 1 29746
2 92290 1 29746
2 92291 1 29761
2 92292 1 29761
2 92293 1 29829
2 92294 1 29829
2 92295 1 29838
2 92296 1 29838
2 92297 1 29839
2 92298 1 29839
2 92299 1 29839
2 92300 1 29873
2 92301 1 29873
2 92302 1 29902
2 92303 1 29902
2 92304 1 29902
2 92305 1 29902
2 92306 1 29902
2 92307 1 29902
2 92308 1 29902
2 92309 1 29902
2 92310 1 29904
2 92311 1 29904
2 92312 1 29914
2 92313 1 29914
2 92314 1 29924
2 92315 1 29924
2 92316 1 29942
2 92317 1 29942
2 92318 1 29951
2 92319 1 29951
2 92320 1 29966
2 92321 1 29966
2 92322 1 29969
2 92323 1 29969
2 92324 1 29969
2 92325 1 29970
2 92326 1 29970
2 92327 1 29970
2 92328 1 29974
2 92329 1 29974
2 92330 1 29974
2 92331 1 29999
2 92332 1 29999
2 92333 1 30016
2 92334 1 30016
2 92335 1 30029
2 92336 1 30029
2 92337 1 30029
2 92338 1 30043
2 92339 1 30043
2 92340 1 30051
2 92341 1 30051
2 92342 1 30061
2 92343 1 30061
2 92344 1 30083
2 92345 1 30083
2 92346 1 30084
2 92347 1 30084
2 92348 1 30090
2 92349 1 30090
2 92350 1 30109
2 92351 1 30109
2 92352 1 30109
2 92353 1 30109
2 92354 1 30109
2 92355 1 30110
2 92356 1 30110
2 92357 1 30110
2 92358 1 30114
2 92359 1 30114
2 92360 1 30118
2 92361 1 30118
2 92362 1 30118
2 92363 1 30136
2 92364 1 30136
2 92365 1 30136
2 92366 1 30190
2 92367 1 30190
2 92368 1 30190
2 92369 1 30190
2 92370 1 30192
2 92371 1 30192
2 92372 1 30192
2 92373 1 30201
2 92374 1 30201
2 92375 1 30237
2 92376 1 30237
2 92377 1 30239
2 92378 1 30239
2 92379 1 30259
2 92380 1 30259
2 92381 1 30262
2 92382 1 30262
2 92383 1 30262
2 92384 1 30262
2 92385 1 30268
2 92386 1 30268
2 92387 1 30279
2 92388 1 30279
2 92389 1 30280
2 92390 1 30280
2 92391 1 30280
2 92392 1 30280
2 92393 1 30283
2 92394 1 30283
2 92395 1 30311
2 92396 1 30311
2 92397 1 30314
2 92398 1 30314
2 92399 1 30321
2 92400 1 30321
2 92401 1 30321
2 92402 1 30322
2 92403 1 30322
2 92404 1 30362
2 92405 1 30362
2 92406 1 30376
2 92407 1 30376
2 92408 1 30376
2 92409 1 30376
2 92410 1 30376
2 92411 1 30382
2 92412 1 30382
2 92413 1 30382
2 92414 1 30382
2 92415 1 30406
2 92416 1 30406
2 92417 1 30407
2 92418 1 30407
2 92419 1 30412
2 92420 1 30412
2 92421 1 30444
2 92422 1 30444
2 92423 1 30453
2 92424 1 30453
2 92425 1 30454
2 92426 1 30454
2 92427 1 30505
2 92428 1 30505
2 92429 1 30514
2 92430 1 30514
2 92431 1 30515
2 92432 1 30515
2 92433 1 30570
2 92434 1 30570
2 92435 1 30572
2 92436 1 30572
2 92437 1 30582
2 92438 1 30582
2 92439 1 30585
2 92440 1 30585
2 92441 1 30585
2 92442 1 30585
2 92443 1 30593
2 92444 1 30593
2 92445 1 30595
2 92446 1 30595
2 92447 1 30607
2 92448 1 30607
2 92449 1 30607
2 92450 1 30607
2 92451 1 30611
2 92452 1 30611
2 92453 1 30611
2 92454 1 30611
2 92455 1 30611
2 92456 1 30648
2 92457 1 30648
2 92458 1 30657
2 92459 1 30657
2 92460 1 30658
2 92461 1 30658
2 92462 1 30661
2 92463 1 30661
2 92464 1 30674
2 92465 1 30674
2 92466 1 30677
2 92467 1 30677
2 92468 1 30686
2 92469 1 30686
2 92470 1 30697
2 92471 1 30697
2 92472 1 30698
2 92473 1 30698
2 92474 1 30700
2 92475 1 30700
2 92476 1 30725
2 92477 1 30725
2 92478 1 30725
2 92479 1 30725
2 92480 1 30757
2 92481 1 30757
2 92482 1 30780
2 92483 1 30780
2 92484 1 30819
2 92485 1 30819
2 92486 1 30846
2 92487 1 30846
2 92488 1 30860
2 92489 1 30860
2 92490 1 30867
2 92491 1 30867
2 92492 1 30882
2 92493 1 30882
2 92494 1 30971
2 92495 1 30971
2 92496 1 31006
2 92497 1 31006
2 92498 1 31020
2 92499 1 31020
2 92500 1 31023
2 92501 1 31023
2 92502 1 31095
2 92503 1 31095
2 92504 1 31098
2 92505 1 31098
2 92506 1 31138
2 92507 1 31138
2 92508 1 31157
2 92509 1 31157
2 92510 1 31157
2 92511 1 31160
2 92512 1 31160
2 92513 1 31194
2 92514 1 31194
2 92515 1 31198
2 92516 1 31198
2 92517 1 31198
2 92518 1 31198
2 92519 1 31198
2 92520 1 31198
2 92521 1 31199
2 92522 1 31199
2 92523 1 31215
2 92524 1 31215
2 92525 1 31226
2 92526 1 31226
2 92527 1 31253
2 92528 1 31253
2 92529 1 31254
2 92530 1 31254
2 92531 1 31267
2 92532 1 31267
2 92533 1 31267
2 92534 1 31274
2 92535 1 31274
2 92536 1 31289
2 92537 1 31289
2 92538 1 31319
2 92539 1 31319
2 92540 1 31319
2 92541 1 31319
2 92542 1 31323
2 92543 1 31323
2 92544 1 31323
2 92545 1 31323
2 92546 1 31323
2 92547 1 31342
2 92548 1 31342
2 92549 1 31349
2 92550 1 31349
2 92551 1 31356
2 92552 1 31356
2 92553 1 31356
2 92554 1 31366
2 92555 1 31366
2 92556 1 31366
2 92557 1 31396
2 92558 1 31396
2 92559 1 31396
2 92560 1 31406
2 92561 1 31406
2 92562 1 31431
2 92563 1 31431
2 92564 1 31437
2 92565 1 31437
2 92566 1 31444
2 92567 1 31444
2 92568 1 31444
2 92569 1 31444
2 92570 1 31445
2 92571 1 31445
2 92572 1 31458
2 92573 1 31458
2 92574 1 31467
2 92575 1 31467
2 92576 1 31497
2 92577 1 31497
2 92578 1 31497
2 92579 1 31497
2 92580 1 31498
2 92581 1 31498
2 92582 1 31498
2 92583 1 31499
2 92584 1 31499
2 92585 1 31506
2 92586 1 31506
2 92587 1 31522
2 92588 1 31522
2 92589 1 31522
2 92590 1 31523
2 92591 1 31523
2 92592 1 31538
2 92593 1 31538
2 92594 1 31538
2 92595 1 31589
2 92596 1 31589
2 92597 1 31589
2 92598 1 31590
2 92599 1 31590
2 92600 1 31615
2 92601 1 31615
2 92602 1 31644
2 92603 1 31644
2 92604 1 31649
2 92605 1 31649
2 92606 1 31665
2 92607 1 31665
2 92608 1 31744
2 92609 1 31744
2 92610 1 31744
2 92611 1 31744
2 92612 1 31751
2 92613 1 31751
2 92614 1 31754
2 92615 1 31754
2 92616 1 31754
2 92617 1 31761
2 92618 1 31761
2 92619 1 31786
2 92620 1 31786
2 92621 1 31787
2 92622 1 31787
2 92623 1 31788
2 92624 1 31788
2 92625 1 31788
2 92626 1 31804
2 92627 1 31804
2 92628 1 31808
2 92629 1 31808
2 92630 1 31808
2 92631 1 31808
2 92632 1 31829
2 92633 1 31829
2 92634 1 31829
2 92635 1 31864
2 92636 1 31864
2 92637 1 31907
2 92638 1 31907
2 92639 1 31950
2 92640 1 31950
2 92641 1 31975
2 92642 1 31975
2 92643 1 31989
2 92644 1 31989
2 92645 1 31992
2 92646 1 31992
2 92647 1 31994
2 92648 1 31994
2 92649 1 32011
2 92650 1 32011
2 92651 1 32012
2 92652 1 32012
2 92653 1 32076
2 92654 1 32076
2 92655 1 32076
2 92656 1 32076
2 92657 1 32082
2 92658 1 32082
2 92659 1 32092
2 92660 1 32092
2 92661 1 32109
2 92662 1 32109
2 92663 1 32121
2 92664 1 32121
2 92665 1 32160
2 92666 1 32160
2 92667 1 32166
2 92668 1 32166
2 92669 1 32177
2 92670 1 32177
2 92671 1 32186
2 92672 1 32186
2 92673 1 32214
2 92674 1 32214
2 92675 1 32214
2 92676 1 32246
2 92677 1 32246
2 92678 1 32266
2 92679 1 32266
2 92680 1 32303
2 92681 1 32303
2 92682 1 32334
2 92683 1 32334
2 92684 1 32336
2 92685 1 32336
2 92686 1 32337
2 92687 1 32337
2 92688 1 32345
2 92689 1 32345
2 92690 1 32348
2 92691 1 32348
2 92692 1 32374
2 92693 1 32374
2 92694 1 32374
2 92695 1 32444
2 92696 1 32444
2 92697 1 32447
2 92698 1 32447
2 92699 1 32454
2 92700 1 32454
2 92701 1 32465
2 92702 1 32465
2 92703 1 32493
2 92704 1 32493
2 92705 1 32521
2 92706 1 32521
2 92707 1 32521
2 92708 1 32521
2 92709 1 32554
2 92710 1 32554
2 92711 1 32554
2 92712 1 32555
2 92713 1 32555
2 92714 1 32557
2 92715 1 32557
2 92716 1 32557
2 92717 1 32558
2 92718 1 32558
2 92719 1 32559
2 92720 1 32559
2 92721 1 32559
2 92722 1 32559
2 92723 1 32571
2 92724 1 32571
2 92725 1 32572
2 92726 1 32572
2 92727 1 32572
2 92728 1 32592
2 92729 1 32592
2 92730 1 32601
2 92731 1 32601
2 92732 1 32601
2 92733 1 32601
2 92734 1 32601
2 92735 1 32601
2 92736 1 32630
2 92737 1 32630
2 92738 1 32687
2 92739 1 32687
2 92740 1 32688
2 92741 1 32688
2 92742 1 32692
2 92743 1 32692
2 92744 1 32699
2 92745 1 32699
2 92746 1 32702
2 92747 1 32702
2 92748 1 32704
2 92749 1 32704
2 92750 1 32707
2 92751 1 32707
2 92752 1 32708
2 92753 1 32708
2 92754 1 32708
2 92755 1 32708
2 92756 1 32708
2 92757 1 32711
2 92758 1 32711
2 92759 1 32714
2 92760 1 32714
2 92761 1 32714
2 92762 1 32716
2 92763 1 32716
2 92764 1 32721
2 92765 1 32721
2 92766 1 32721
2 92767 1 32721
2 92768 1 32721
2 92769 1 32721
2 92770 1 32721
2 92771 1 32724
2 92772 1 32724
2 92773 1 32725
2 92774 1 32725
2 92775 1 32725
2 92776 1 32726
2 92777 1 32726
2 92778 1 32728
2 92779 1 32728
2 92780 1 32737
2 92781 1 32737
2 92782 1 32737
2 92783 1 32747
2 92784 1 32747
2 92785 1 32747
2 92786 1 32748
2 92787 1 32748
2 92788 1 32752
2 92789 1 32752
2 92790 1 32752
2 92791 1 32752
2 92792 1 32753
2 92793 1 32753
2 92794 1 32776
2 92795 1 32776
2 92796 1 32776
2 92797 1 32776
2 92798 1 32777
2 92799 1 32777
2 92800 1 32782
2 92801 1 32782
2 92802 1 32782
2 92803 1 32782
2 92804 1 32782
2 92805 1 32795
2 92806 1 32795
2 92807 1 32795
2 92808 1 32800
2 92809 1 32800
2 92810 1 32803
2 92811 1 32803
2 92812 1 32804
2 92813 1 32804
2 92814 1 32806
2 92815 1 32806
2 92816 1 32806
2 92817 1 32815
2 92818 1 32815
2 92819 1 32816
2 92820 1 32816
2 92821 1 32817
2 92822 1 32817
2 92823 1 32817
2 92824 1 32817
2 92825 1 32817
2 92826 1 32820
2 92827 1 32820
2 92828 1 32821
2 92829 1 32821
2 92830 1 32823
2 92831 1 32823
2 92832 1 32824
2 92833 1 32824
2 92834 1 32852
2 92835 1 32852
2 92836 1 32869
2 92837 1 32869
2 92838 1 32891
2 92839 1 32891
2 92840 1 32899
2 92841 1 32899
2 92842 1 32903
2 92843 1 32903
2 92844 1 32903
2 92845 1 32903
2 92846 1 32903
2 92847 1 32914
2 92848 1 32914
2 92849 1 32928
2 92850 1 32928
2 92851 1 32937
2 92852 1 32937
2 92853 1 32945
2 92854 1 32945
2 92855 1 32945
2 92856 1 32945
2 92857 1 32948
2 92858 1 32948
2 92859 1 32965
2 92860 1 32965
2 92861 1 32988
2 92862 1 32988
2 92863 1 33024
2 92864 1 33024
2 92865 1 33034
2 92866 1 33034
2 92867 1 33048
2 92868 1 33048
2 92869 1 33067
2 92870 1 33067
2 92871 1 33083
2 92872 1 33083
2 92873 1 33083
2 92874 1 33083
2 92875 1 33084
2 92876 1 33084
2 92877 1 33089
2 92878 1 33089
2 92879 1 33089
2 92880 1 33089
2 92881 1 33089
2 92882 1 33089
2 92883 1 33089
2 92884 1 33089
2 92885 1 33089
2 92886 1 33089
2 92887 1 33089
2 92888 1 33089
2 92889 1 33090
2 92890 1 33090
2 92891 1 33090
2 92892 1 33102
2 92893 1 33102
2 92894 1 33102
2 92895 1 33103
2 92896 1 33103
2 92897 1 33114
2 92898 1 33114
2 92899 1 33114
2 92900 1 33122
2 92901 1 33122
2 92902 1 33122
2 92903 1 33122
2 92904 1 33122
2 92905 1 33123
2 92906 1 33123
2 92907 1 33143
2 92908 1 33143
2 92909 1 33144
2 92910 1 33144
2 92911 1 33144
2 92912 1 33144
2 92913 1 33147
2 92914 1 33147
2 92915 1 33170
2 92916 1 33170
2 92917 1 33179
2 92918 1 33179
2 92919 1 33180
2 92920 1 33180
2 92921 1 33181
2 92922 1 33181
2 92923 1 33181
2 92924 1 33182
2 92925 1 33182
2 92926 1 33187
2 92927 1 33187
2 92928 1 33209
2 92929 1 33209
2 92930 1 33218
2 92931 1 33218
2 92932 1 33258
2 92933 1 33258
2 92934 1 33275
2 92935 1 33275
2 92936 1 33278
2 92937 1 33278
2 92938 1 33284
2 92939 1 33284
2 92940 1 33284
2 92941 1 33291
2 92942 1 33291
2 92943 1 33291
2 92944 1 33291
2 92945 1 33291
2 92946 1 33291
2 92947 1 33291
2 92948 1 33291
2 92949 1 33291
2 92950 1 33291
2 92951 1 33291
2 92952 1 33291
2 92953 1 33291
2 92954 1 33291
2 92955 1 33291
2 92956 1 33291
2 92957 1 33317
2 92958 1 33317
2 92959 1 33351
2 92960 1 33351
2 92961 1 33353
2 92962 1 33353
2 92963 1 33358
2 92964 1 33358
2 92965 1 33359
2 92966 1 33359
2 92967 1 33359
2 92968 1 33359
2 92969 1 33375
2 92970 1 33375
2 92971 1 33377
2 92972 1 33377
2 92973 1 33382
2 92974 1 33382
2 92975 1 33382
2 92976 1 33382
2 92977 1 33382
2 92978 1 33382
2 92979 1 33382
2 92980 1 33382
2 92981 1 33382
2 92982 1 33382
2 92983 1 33382
2 92984 1 33382
2 92985 1 33382
2 92986 1 33382
2 92987 1 33383
2 92988 1 33383
2 92989 1 33383
2 92990 1 33383
2 92991 1 33387
2 92992 1 33387
2 92993 1 33418
2 92994 1 33418
2 92995 1 33421
2 92996 1 33421
2 92997 1 33425
2 92998 1 33425
2 92999 1 33436
2 93000 1 33436
2 93001 1 33458
2 93002 1 33458
2 93003 1 33458
2 93004 1 33458
2 93005 1 33469
2 93006 1 33469
2 93007 1 33479
2 93008 1 33479
2 93009 1 33480
2 93010 1 33480
2 93011 1 33484
2 93012 1 33484
2 93013 1 33493
2 93014 1 33493
2 93015 1 33503
2 93016 1 33503
2 93017 1 33531
2 93018 1 33531
2 93019 1 33532
2 93020 1 33532
2 93021 1 33532
2 93022 1 33537
2 93023 1 33537
2 93024 1 33559
2 93025 1 33559
2 93026 1 33583
2 93027 1 33583
2 93028 1 33584
2 93029 1 33584
2 93030 1 33595
2 93031 1 33595
2 93032 1 33595
2 93033 1 33595
2 93034 1 33596
2 93035 1 33596
2 93036 1 33628
2 93037 1 33628
2 93038 1 33637
2 93039 1 33637
2 93040 1 33658
2 93041 1 33658
2 93042 1 33658
2 93043 1 33658
2 93044 1 33658
2 93045 1 33658
2 93046 1 33658
2 93047 1 33698
2 93048 1 33698
2 93049 1 33739
2 93050 1 33739
2 93051 1 33744
2 93052 1 33744
2 93053 1 33744
2 93054 1 33771
2 93055 1 33771
2 93056 1 33772
2 93057 1 33772
2 93058 1 33772
2 93059 1 33773
2 93060 1 33773
2 93061 1 33773
2 93062 1 33779
2 93063 1 33779
2 93064 1 33790
2 93065 1 33790
2 93066 1 33805
2 93067 1 33805
2 93068 1 33812
2 93069 1 33812
2 93070 1 33812
2 93071 1 33813
2 93072 1 33813
2 93073 1 33814
2 93074 1 33814
2 93075 1 33814
2 93076 1 33829
2 93077 1 33829
2 93078 1 33829
2 93079 1 33830
2 93080 1 33830
2 93081 1 33830
2 93082 1 33831
2 93083 1 33831
2 93084 1 33855
2 93085 1 33855
2 93086 1 33858
2 93087 1 33858
2 93088 1 33872
2 93089 1 33872
2 93090 1 33902
2 93091 1 33902
2 93092 1 33902
2 93093 1 33902
2 93094 1 33902
2 93095 1 33904
2 93096 1 33904
2 93097 1 33917
2 93098 1 33917
2 93099 1 33921
2 93100 1 33921
2 93101 1 33929
2 93102 1 33929
2 93103 1 33955
2 93104 1 33955
2 93105 1 33955
2 93106 1 33955
2 93107 1 33987
2 93108 1 33987
2 93109 1 34001
2 93110 1 34001
2 93111 1 34016
2 93112 1 34016
2 93113 1 34045
2 93114 1 34045
2 93115 1 34046
2 93116 1 34046
2 93117 1 34054
2 93118 1 34054
2 93119 1 34056
2 93120 1 34056
2 93121 1 34057
2 93122 1 34057
2 93123 1 34057
2 93124 1 34067
2 93125 1 34067
2 93126 1 34068
2 93127 1 34068
2 93128 1 34074
2 93129 1 34074
2 93130 1 34097
2 93131 1 34097
2 93132 1 34099
2 93133 1 34099
2 93134 1 34103
2 93135 1 34103
2 93136 1 34107
2 93137 1 34107
2 93138 1 34119
2 93139 1 34119
2 93140 1 34119
2 93141 1 34119
2 93142 1 34120
2 93143 1 34120
2 93144 1 34120
2 93145 1 34135
2 93146 1 34135
2 93147 1 34135
2 93148 1 34135
2 93149 1 34136
2 93150 1 34136
2 93151 1 34143
2 93152 1 34143
2 93153 1 34150
2 93154 1 34150
2 93155 1 34152
2 93156 1 34152
2 93157 1 34161
2 93158 1 34161
2 93159 1 34164
2 93160 1 34164
2 93161 1 34173
2 93162 1 34173
2 93163 1 34173
2 93164 1 34177
2 93165 1 34177
2 93166 1 34198
2 93167 1 34198
2 93168 1 34199
2 93169 1 34199
2 93170 1 34199
2 93171 1 34215
2 93172 1 34215
2 93173 1 34226
2 93174 1 34226
2 93175 1 34233
2 93176 1 34233
2 93177 1 34238
2 93178 1 34238
2 93179 1 34238
2 93180 1 34246
2 93181 1 34246
2 93182 1 34253
2 93183 1 34253
2 93184 1 34253
2 93185 1 34253
2 93186 1 34267
2 93187 1 34267
2 93188 1 34274
2 93189 1 34274
2 93190 1 34292
2 93191 1 34292
2 93192 1 34304
2 93193 1 34304
2 93194 1 34305
2 93195 1 34305
2 93196 1 34305
2 93197 1 34312
2 93198 1 34312
2 93199 1 34315
2 93200 1 34315
2 93201 1 34319
2 93202 1 34319
2 93203 1 34334
2 93204 1 34334
2 93205 1 34342
2 93206 1 34342
2 93207 1 34351
2 93208 1 34351
2 93209 1 34352
2 93210 1 34352
2 93211 1 34353
2 93212 1 34353
2 93213 1 34363
2 93214 1 34363
2 93215 1 34364
2 93216 1 34364
2 93217 1 34373
2 93218 1 34373
2 93219 1 34378
2 93220 1 34378
2 93221 1 34378
2 93222 1 34383
2 93223 1 34383
2 93224 1 34393
2 93225 1 34393
2 93226 1 34410
2 93227 1 34410
2 93228 1 34410
2 93229 1 34410
2 93230 1 34424
2 93231 1 34424
2 93232 1 34434
2 93233 1 34434
2 93234 1 34457
2 93235 1 34457
2 93236 1 34462
2 93237 1 34462
2 93238 1 34478
2 93239 1 34478
2 93240 1 34487
2 93241 1 34487
2 93242 1 34499
2 93243 1 34499
2 93244 1 34502
2 93245 1 34502
2 93246 1 34502
2 93247 1 34502
2 93248 1 34510
2 93249 1 34510
2 93250 1 34519
2 93251 1 34519
2 93252 1 34519
2 93253 1 34528
2 93254 1 34528
2 93255 1 34534
2 93256 1 34534
2 93257 1 34538
2 93258 1 34538
2 93259 1 34539
2 93260 1 34539
2 93261 1 34539
2 93262 1 34546
2 93263 1 34546
2 93264 1 34546
2 93265 1 34546
2 93266 1 34546
2 93267 1 34547
2 93268 1 34547
2 93269 1 34564
2 93270 1 34564
2 93271 1 34579
2 93272 1 34579
2 93273 1 34579
2 93274 1 34579
2 93275 1 34579
2 93276 1 34589
2 93277 1 34589
2 93278 1 34591
2 93279 1 34591
2 93280 1 34606
2 93281 1 34606
2 93282 1 34638
2 93283 1 34638
2 93284 1 34638
2 93285 1 34641
2 93286 1 34641
2 93287 1 34642
2 93288 1 34642
2 93289 1 34642
2 93290 1 34642
2 93291 1 34653
2 93292 1 34653
2 93293 1 34661
2 93294 1 34661
2 93295 1 34663
2 93296 1 34663
2 93297 1 34667
2 93298 1 34667
2 93299 1 34668
2 93300 1 34668
2 93301 1 34669
2 93302 1 34669
2 93303 1 34674
2 93304 1 34674
2 93305 1 34674
2 93306 1 34674
2 93307 1 34674
2 93308 1 34674
2 93309 1 34675
2 93310 1 34675
2 93311 1 34684
2 93312 1 34684
2 93313 1 34688
2 93314 1 34688
2 93315 1 34701
2 93316 1 34701
2 93317 1 34701
2 93318 1 34702
2 93319 1 34702
2 93320 1 34702
2 93321 1 34712
2 93322 1 34712
2 93323 1 34731
2 93324 1 34731
2 93325 1 34733
2 93326 1 34733
2 93327 1 34745
2 93328 1 34745
2 93329 1 34752
2 93330 1 34752
2 93331 1 34771
2 93332 1 34771
2 93333 1 34775
2 93334 1 34775
2 93335 1 34775
2 93336 1 34782
2 93337 1 34782
2 93338 1 34792
2 93339 1 34792
2 93340 1 34793
2 93341 1 34793
2 93342 1 34793
2 93343 1 34793
2 93344 1 34806
2 93345 1 34806
2 93346 1 34817
2 93347 1 34817
2 93348 1 34839
2 93349 1 34839
2 93350 1 34856
2 93351 1 34856
2 93352 1 34863
2 93353 1 34863
2 93354 1 34863
2 93355 1 34863
2 93356 1 34863
2 93357 1 34863
2 93358 1 34863
2 93359 1 34863
2 93360 1 34863
2 93361 1 34872
2 93362 1 34872
2 93363 1 34872
2 93364 1 34872
2 93365 1 34872
2 93366 1 34882
2 93367 1 34882
2 93368 1 34884
2 93369 1 34884
2 93370 1 34886
2 93371 1 34886
2 93372 1 34899
2 93373 1 34899
2 93374 1 34901
2 93375 1 34901
2 93376 1 34909
2 93377 1 34909
2 93378 1 34938
2 93379 1 34938
2 93380 1 34938
2 93381 1 34938
2 93382 1 34950
2 93383 1 34950
2 93384 1 34952
2 93385 1 34952
2 93386 1 34952
2 93387 1 34955
2 93388 1 34955
2 93389 1 34956
2 93390 1 34956
2 93391 1 34959
2 93392 1 34959
2 93393 1 34974
2 93394 1 34974
2 93395 1 34980
2 93396 1 34980
2 93397 1 34980
2 93398 1 34982
2 93399 1 34982
2 93400 1 34983
2 93401 1 34983
2 93402 1 34984
2 93403 1 34984
2 93404 1 34994
2 93405 1 34994
2 93406 1 34996
2 93407 1 34996
2 93408 1 34996
2 93409 1 35002
2 93410 1 35002
2 93411 1 35017
2 93412 1 35017
2 93413 1 35018
2 93414 1 35018
2 93415 1 35018
2 93416 1 35018
2 93417 1 35020
2 93418 1 35020
2 93419 1 35020
2 93420 1 35022
2 93421 1 35022
2 93422 1 35022
2 93423 1 35024
2 93424 1 35024
2 93425 1 35024
2 93426 1 35028
2 93427 1 35028
2 93428 1 35028
2 93429 1 35050
2 93430 1 35050
2 93431 1 35051
2 93432 1 35051
2 93433 1 35051
2 93434 1 35051
2 93435 1 35061
2 93436 1 35061
2 93437 1 35062
2 93438 1 35062
2 93439 1 35063
2 93440 1 35063
2 93441 1 35065
2 93442 1 35065
2 93443 1 35065
2 93444 1 35070
2 93445 1 35070
2 93446 1 35075
2 93447 1 35075
2 93448 1 35121
2 93449 1 35121
2 93450 1 35131
2 93451 1 35131
2 93452 1 35133
2 93453 1 35133
2 93454 1 35162
2 93455 1 35162
2 93456 1 35172
2 93457 1 35172
2 93458 1 35179
2 93459 1 35179
2 93460 1 35181
2 93461 1 35181
2 93462 1 35182
2 93463 1 35182
2 93464 1 35182
2 93465 1 35184
2 93466 1 35184
2 93467 1 35186
2 93468 1 35186
2 93469 1 35190
2 93470 1 35190
2 93471 1 35229
2 93472 1 35229
2 93473 1 35265
2 93474 1 35265
2 93475 1 35274
2 93476 1 35274
2 93477 1 35278
2 93478 1 35278
2 93479 1 35303
2 93480 1 35303
2 93481 1 35323
2 93482 1 35323
2 93483 1 35331
2 93484 1 35331
2 93485 1 35342
2 93486 1 35342
2 93487 1 35349
2 93488 1 35349
2 93489 1 35349
2 93490 1 35349
2 93491 1 35349
2 93492 1 35351
2 93493 1 35351
2 93494 1 35351
2 93495 1 35353
2 93496 1 35353
2 93497 1 35355
2 93498 1 35355
2 93499 1 35355
2 93500 1 35368
2 93501 1 35368
2 93502 1 35373
2 93503 1 35373
2 93504 1 35423
2 93505 1 35423
2 93506 1 35424
2 93507 1 35424
2 93508 1 35433
2 93509 1 35433
2 93510 1 35433
2 93511 1 35451
2 93512 1 35451
2 93513 1 35452
2 93514 1 35452
2 93515 1 35472
2 93516 1 35472
2 93517 1 35485
2 93518 1 35485
2 93519 1 35485
2 93520 1 35504
2 93521 1 35504
2 93522 1 35531
2 93523 1 35531
2 93524 1 35531
2 93525 1 35538
2 93526 1 35538
2 93527 1 35561
2 93528 1 35561
2 93529 1 35565
2 93530 1 35565
2 93531 1 35566
2 93532 1 35566
2 93533 1 35568
2 93534 1 35568
2 93535 1 35572
2 93536 1 35572
2 93537 1 35572
2 93538 1 35576
2 93539 1 35576
2 93540 1 35581
2 93541 1 35581
2 93542 1 35582
2 93543 1 35582
2 93544 1 35590
2 93545 1 35590
2 93546 1 35591
2 93547 1 35591
2 93548 1 35591
2 93549 1 35617
2 93550 1 35617
2 93551 1 35632
2 93552 1 35632
2 93553 1 35633
2 93554 1 35633
2 93555 1 35633
2 93556 1 35662
2 93557 1 35662
2 93558 1 35672
2 93559 1 35672
2 93560 1 35673
2 93561 1 35673
2 93562 1 35681
2 93563 1 35681
2 93564 1 35703
2 93565 1 35703
2 93566 1 35719
2 93567 1 35719
2 93568 1 35720
2 93569 1 35720
2 93570 1 35720
2 93571 1 35720
2 93572 1 35722
2 93573 1 35722
2 93574 1 35739
2 93575 1 35739
2 93576 1 35739
2 93577 1 35739
2 93578 1 35739
2 93579 1 35741
2 93580 1 35741
2 93581 1 35747
2 93582 1 35747
2 93583 1 35760
2 93584 1 35760
2 93585 1 35772
2 93586 1 35772
2 93587 1 35774
2 93588 1 35774
2 93589 1 35788
2 93590 1 35788
2 93591 1 35795
2 93592 1 35795
2 93593 1 35816
2 93594 1 35816
2 93595 1 35828
2 93596 1 35828
2 93597 1 35860
2 93598 1 35860
2 93599 1 35861
2 93600 1 35861
2 93601 1 35861
2 93602 1 35861
2 93603 1 35861
2 93604 1 35861
2 93605 1 35863
2 93606 1 35863
2 93607 1 35883
2 93608 1 35883
2 93609 1 35894
2 93610 1 35894
2 93611 1 35894
2 93612 1 35895
2 93613 1 35895
2 93614 1 35905
2 93615 1 35905
2 93616 1 35928
2 93617 1 35928
2 93618 1 35931
2 93619 1 35931
2 93620 1 35988
2 93621 1 35988
2 93622 1 36006
2 93623 1 36006
2 93624 1 36006
2 93625 1 36070
2 93626 1 36070
2 93627 1 36071
2 93628 1 36071
2 93629 1 36073
2 93630 1 36073
2 93631 1 36105
2 93632 1 36105
2 93633 1 36129
2 93634 1 36129
2 93635 1 36135
2 93636 1 36135
2 93637 1 36140
2 93638 1 36140
2 93639 1 36144
2 93640 1 36144
2 93641 1 36163
2 93642 1 36163
2 93643 1 36180
2 93644 1 36180
2 93645 1 36180
2 93646 1 36181
2 93647 1 36181
2 93648 1 36204
2 93649 1 36204
2 93650 1 36218
2 93651 1 36218
2 93652 1 36225
2 93653 1 36225
2 93654 1 36228
2 93655 1 36228
2 93656 1 36236
2 93657 1 36236
2 93658 1 36236
2 93659 1 36237
2 93660 1 36237
2 93661 1 36237
2 93662 1 36307
2 93663 1 36307
2 93664 1 36335
2 93665 1 36335
2 93666 1 36335
2 93667 1 36335
2 93668 1 36370
2 93669 1 36370
2 93670 1 36370
2 93671 1 36375
2 93672 1 36375
2 93673 1 36377
2 93674 1 36377
2 93675 1 36381
2 93676 1 36381
2 93677 1 36381
2 93678 1 36395
2 93679 1 36395
2 93680 1 36409
2 93681 1 36409
2 93682 1 36417
2 93683 1 36417
2 93684 1 36462
2 93685 1 36462
2 93686 1 36472
2 93687 1 36472
2 93688 1 36503
2 93689 1 36503
2 93690 1 36522
2 93691 1 36522
2 93692 1 36625
2 93693 1 36625
2 93694 1 36628
2 93695 1 36628
2 93696 1 36629
2 93697 1 36629
2 93698 1 36632
2 93699 1 36632
2 93700 1 36671
2 93701 1 36671
2 93702 1 36676
2 93703 1 36676
2 93704 1 36677
2 93705 1 36677
2 93706 1 36705
2 93707 1 36705
2 93708 1 36705
2 93709 1 36706
2 93710 1 36706
2 93711 1 36727
2 93712 1 36727
2 93713 1 36729
2 93714 1 36729
2 93715 1 36730
2 93716 1 36730
2 93717 1 36731
2 93718 1 36731
2 93719 1 36732
2 93720 1 36732
2 93721 1 36732
2 93722 1 36732
2 93723 1 36732
2 93724 1 36732
2 93725 1 36747
2 93726 1 36747
2 93727 1 36747
2 93728 1 36747
2 93729 1 36759
2 93730 1 36759
2 93731 1 36763
2 93732 1 36763
2 93733 1 36777
2 93734 1 36777
2 93735 1 36778
2 93736 1 36778
2 93737 1 36778
2 93738 1 36812
2 93739 1 36812
2 93740 1 36825
2 93741 1 36825
2 93742 1 36842
2 93743 1 36842
2 93744 1 36843
2 93745 1 36843
2 93746 1 36845
2 93747 1 36845
2 93748 1 36845
2 93749 1 36855
2 93750 1 36855
2 93751 1 36876
2 93752 1 36876
2 93753 1 36899
2 93754 1 36899
2 93755 1 36899
2 93756 1 36906
2 93757 1 36906
2 93758 1 36943
2 93759 1 36943
2 93760 1 36943
2 93761 1 36943
2 93762 1 36954
2 93763 1 36954
2 93764 1 36962
2 93765 1 36962
2 93766 1 36975
2 93767 1 36975
2 93768 1 36975
2 93769 1 37009
2 93770 1 37009
2 93771 1 37012
2 93772 1 37012
2 93773 1 37013
2 93774 1 37013
2 93775 1 37014
2 93776 1 37014
2 93777 1 37014
2 93778 1 37035
2 93779 1 37035
2 93780 1 37037
2 93781 1 37037
2 93782 1 37054
2 93783 1 37054
2 93784 1 37064
2 93785 1 37064
2 93786 1 37064
2 93787 1 37073
2 93788 1 37073
2 93789 1 37084
2 93790 1 37084
2 93791 1 37097
2 93792 1 37097
2 93793 1 37142
2 93794 1 37142
2 93795 1 37142
2 93796 1 37185
2 93797 1 37185
2 93798 1 37213
2 93799 1 37213
2 93800 1 37231
2 93801 1 37231
2 93802 1 37252
2 93803 1 37252
2 93804 1 37283
2 93805 1 37283
2 93806 1 37283
2 93807 1 37292
2 93808 1 37292
2 93809 1 37295
2 93810 1 37295
2 93811 1 37295
2 93812 1 37296
2 93813 1 37296
2 93814 1 37328
2 93815 1 37328
2 93816 1 37338
2 93817 1 37338
2 93818 1 37352
2 93819 1 37352
2 93820 1 37354
2 93821 1 37354
2 93822 1 37380
2 93823 1 37380
2 93824 1 37381
2 93825 1 37381
2 93826 1 37382
2 93827 1 37382
2 93828 1 37401
2 93829 1 37401
2 93830 1 37401
2 93831 1 37401
2 93832 1 37409
2 93833 1 37409
2 93834 1 37457
2 93835 1 37457
2 93836 1 37457
2 93837 1 37488
2 93838 1 37488
2 93839 1 37516
2 93840 1 37516
2 93841 1 37516
2 93842 1 37517
2 93843 1 37517
2 93844 1 37541
2 93845 1 37541
2 93846 1 37544
2 93847 1 37544
2 93848 1 37583
2 93849 1 37583
2 93850 1 37583
2 93851 1 37583
2 93852 1 37583
2 93853 1 37623
2 93854 1 37623
2 93855 1 37636
2 93856 1 37636
2 93857 1 37657
2 93858 1 37657
2 93859 1 37657
2 93860 1 37657
2 93861 1 37677
2 93862 1 37677
2 93863 1 37678
2 93864 1 37678
2 93865 1 37755
2 93866 1 37755
2 93867 1 37759
2 93868 1 37759
2 93869 1 37772
2 93870 1 37772
2 93871 1 37796
2 93872 1 37796
2 93873 1 37798
2 93874 1 37798
2 93875 1 37798
2 93876 1 37802
2 93877 1 37802
2 93878 1 37803
2 93879 1 37803
2 93880 1 37806
2 93881 1 37806
2 93882 1 37811
2 93883 1 37811
2 93884 1 37814
2 93885 1 37814
2 93886 1 37814
2 93887 1 37814
2 93888 1 37838
2 93889 1 37838
2 93890 1 37838
2 93891 1 37838
2 93892 1 37842
2 93893 1 37842
2 93894 1 37847
2 93895 1 37847
2 93896 1 37847
2 93897 1 37881
2 93898 1 37881
2 93899 1 37886
2 93900 1 37886
2 93901 1 37892
2 93902 1 37892
2 93903 1 37908
2 93904 1 37908
2 93905 1 37912
2 93906 1 37912
2 93907 1 37922
2 93908 1 37922
2 93909 1 37936
2 93910 1 37936
2 93911 1 37943
2 93912 1 37943
2 93913 1 37943
2 93914 1 37943
2 93915 1 37943
2 93916 1 37943
2 93917 1 37943
2 93918 1 37970
2 93919 1 37970
2 93920 1 37987
2 93921 1 37987
2 93922 1 38025
2 93923 1 38025
2 93924 1 38025
2 93925 1 38025
2 93926 1 38026
2 93927 1 38026
2 93928 1 38026
2 93929 1 38026
2 93930 1 38046
2 93931 1 38046
2 93932 1 38067
2 93933 1 38067
2 93934 1 38069
2 93935 1 38069
2 93936 1 38081
2 93937 1 38081
2 93938 1 38081
2 93939 1 38082
2 93940 1 38082
2 93941 1 38082
2 93942 1 38083
2 93943 1 38083
2 93944 1 38083
2 93945 1 38091
2 93946 1 38091
2 93947 1 38091
2 93948 1 38094
2 93949 1 38094
2 93950 1 38096
2 93951 1 38096
2 93952 1 38096
2 93953 1 38097
2 93954 1 38097
2 93955 1 38097
2 93956 1 38099
2 93957 1 38099
2 93958 1 38111
2 93959 1 38111
2 93960 1 38115
2 93961 1 38115
2 93962 1 38180
2 93963 1 38180
2 93964 1 38205
2 93965 1 38205
2 93966 1 38205
2 93967 1 38205
2 93968 1 38205
2 93969 1 38205
2 93970 1 38217
2 93971 1 38217
2 93972 1 38217
2 93973 1 38229
2 93974 1 38229
2 93975 1 38229
2 93976 1 38229
2 93977 1 38229
2 93978 1 38229
2 93979 1 38260
2 93980 1 38260
2 93981 1 38261
2 93982 1 38261
2 93983 1 38273
2 93984 1 38273
2 93985 1 38274
2 93986 1 38274
2 93987 1 38274
2 93988 1 38274
2 93989 1 38283
2 93990 1 38283
2 93991 1 38286
2 93992 1 38286
2 93993 1 38290
2 93994 1 38290
2 93995 1 38291
2 93996 1 38291
2 93997 1 38304
2 93998 1 38304
2 93999 1 38341
2 94000 1 38341
2 94001 1 38346
2 94002 1 38346
2 94003 1 38359
2 94004 1 38359
2 94005 1 38359
2 94006 1 38375
2 94007 1 38375
2 94008 1 38397
2 94009 1 38397
2 94010 1 38400
2 94011 1 38400
2 94012 1 38401
2 94013 1 38401
2 94014 1 38405
2 94015 1 38405
2 94016 1 38405
2 94017 1 38406
2 94018 1 38406
2 94019 1 38408
2 94020 1 38408
2 94021 1 38408
2 94022 1 38409
2 94023 1 38409
2 94024 1 38423
2 94025 1 38423
2 94026 1 38423
2 94027 1 38424
2 94028 1 38424
2 94029 1 38424
2 94030 1 38432
2 94031 1 38432
2 94032 1 38433
2 94033 1 38433
2 94034 1 38502
2 94035 1 38502
2 94036 1 38515
2 94037 1 38515
2 94038 1 38515
2 94039 1 38515
2 94040 1 38516
2 94041 1 38516
2 94042 1 38517
2 94043 1 38517
2 94044 1 38535
2 94045 1 38535
2 94046 1 38551
2 94047 1 38551
2 94048 1 38551
2 94049 1 38551
2 94050 1 38552
2 94051 1 38552
2 94052 1 38577
2 94053 1 38577
2 94054 1 38578
2 94055 1 38578
2 94056 1 38578
2 94057 1 38578
2 94058 1 38589
2 94059 1 38589
2 94060 1 38590
2 94061 1 38590
2 94062 1 38590
2 94063 1 38606
2 94064 1 38606
2 94065 1 38607
2 94066 1 38607
2 94067 1 38607
2 94068 1 38615
2 94069 1 38615
2 94070 1 38620
2 94071 1 38620
2 94072 1 38621
2 94073 1 38621
2 94074 1 38657
2 94075 1 38657
2 94076 1 38664
2 94077 1 38664
2 94078 1 38682
2 94079 1 38682
2 94080 1 38685
2 94081 1 38685
2 94082 1 38685
2 94083 1 38687
2 94084 1 38687
2 94085 1 38695
2 94086 1 38695
2 94087 1 38699
2 94088 1 38699
2 94089 1 38699
2 94090 1 38700
2 94091 1 38700
2 94092 1 38721
2 94093 1 38721
2 94094 1 38724
2 94095 1 38724
2 94096 1 38730
2 94097 1 38730
2 94098 1 38732
2 94099 1 38732
2 94100 1 38741
2 94101 1 38741
2 94102 1 38745
2 94103 1 38745
2 94104 1 38745
2 94105 1 38747
2 94106 1 38747
2 94107 1 38751
2 94108 1 38751
2 94109 1 38751
2 94110 1 38754
2 94111 1 38754
2 94112 1 38756
2 94113 1 38756
2 94114 1 38756
2 94115 1 38756
2 94116 1 38772
2 94117 1 38772
2 94118 1 38772
2 94119 1 38775
2 94120 1 38775
2 94121 1 38782
2 94122 1 38782
2 94123 1 38819
2 94124 1 38819
2 94125 1 38853
2 94126 1 38853
2 94127 1 38854
2 94128 1 38854
2 94129 1 38863
2 94130 1 38863
2 94131 1 38863
2 94132 1 38885
2 94133 1 38885
2 94134 1 38886
2 94135 1 38886
2 94136 1 38909
2 94137 1 38909
2 94138 1 38939
2 94139 1 38939
2 94140 1 38972
2 94141 1 38972
2 94142 1 38972
2 94143 1 38972
2 94144 1 38972
2 94145 1 38972
2 94146 1 38972
2 94147 1 38979
2 94148 1 38979
2 94149 1 38984
2 94150 1 38984
2 94151 1 38984
2 94152 1 38984
2 94153 1 38985
2 94154 1 38985
2 94155 1 38985
2 94156 1 38985
2 94157 1 38985
2 94158 1 38985
2 94159 1 38985
2 94160 1 38987
2 94161 1 38987
2 94162 1 38990
2 94163 1 38990
2 94164 1 38990
2 94165 1 38991
2 94166 1 38991
2 94167 1 38999
2 94168 1 38999
2 94169 1 38999
2 94170 1 39000
2 94171 1 39000
2 94172 1 39026
2 94173 1 39026
2 94174 1 39029
2 94175 1 39029
2 94176 1 39045
2 94177 1 39045
2 94178 1 39045
2 94179 1 39045
2 94180 1 39061
2 94181 1 39061
2 94182 1 39061
2 94183 1 39064
2 94184 1 39064
2 94185 1 39074
2 94186 1 39074
2 94187 1 39075
2 94188 1 39075
2 94189 1 39075
2 94190 1 39088
2 94191 1 39088
2 94192 1 39088
2 94193 1 39139
2 94194 1 39139
2 94195 1 39141
2 94196 1 39141
2 94197 1 39141
2 94198 1 39149
2 94199 1 39149
2 94200 1 39149
2 94201 1 39151
2 94202 1 39151
2 94203 1 39151
2 94204 1 39158
2 94205 1 39158
2 94206 1 39161
2 94207 1 39161
2 94208 1 39161
2 94209 1 39161
2 94210 1 39165
2 94211 1 39165
2 94212 1 39165
2 94213 1 39171
2 94214 1 39171
2 94215 1 39171
2 94216 1 39171
2 94217 1 39174
2 94218 1 39174
2 94219 1 39174
2 94220 1 39175
2 94221 1 39175
2 94222 1 39175
2 94223 1 39183
2 94224 1 39183
2 94225 1 39183
2 94226 1 39192
2 94227 1 39192
2 94228 1 39206
2 94229 1 39206
2 94230 1 39206
2 94231 1 39206
2 94232 1 39206
2 94233 1 39206
2 94234 1 39207
2 94235 1 39207
2 94236 1 39226
2 94237 1 39226
2 94238 1 39226
2 94239 1 39226
2 94240 1 39226
2 94241 1 39226
2 94242 1 39227
2 94243 1 39227
2 94244 1 39244
2 94245 1 39244
2 94246 1 39244
2 94247 1 39245
2 94248 1 39245
2 94249 1 39259
2 94250 1 39259
2 94251 1 39274
2 94252 1 39274
2 94253 1 39274
2 94254 1 39275
2 94255 1 39275
2 94256 1 39283
2 94257 1 39283
2 94258 1 39284
2 94259 1 39284
2 94260 1 39287
2 94261 1 39287
2 94262 1 39331
2 94263 1 39331
2 94264 1 39354
2 94265 1 39354
2 94266 1 39359
2 94267 1 39359
2 94268 1 39371
2 94269 1 39371
2 94270 1 39379
2 94271 1 39379
2 94272 1 39409
2 94273 1 39409
2 94274 1 39413
2 94275 1 39413
2 94276 1 39417
2 94277 1 39417
2 94278 1 39417
2 94279 1 39431
2 94280 1 39431
2 94281 1 39454
2 94282 1 39454
2 94283 1 39468
2 94284 1 39468
2 94285 1 39468
2 94286 1 39468
2 94287 1 39468
2 94288 1 39491
2 94289 1 39491
2 94290 1 39511
2 94291 1 39511
2 94292 1 39511
2 94293 1 39529
2 94294 1 39529
2 94295 1 39530
2 94296 1 39530
2 94297 1 39530
2 94298 1 39530
2 94299 1 39531
2 94300 1 39531
2 94301 1 39531
2 94302 1 39532
2 94303 1 39532
2 94304 1 39568
2 94305 1 39568
2 94306 1 39568
2 94307 1 39577
2 94308 1 39577
2 94309 1 39578
2 94310 1 39578
2 94311 1 39581
2 94312 1 39581
2 94313 1 39596
2 94314 1 39596
2 94315 1 39596
2 94316 1 39620
2 94317 1 39620
2 94318 1 39624
2 94319 1 39624
2 94320 1 39624
2 94321 1 39642
2 94322 1 39642
2 94323 1 39650
2 94324 1 39650
2 94325 1 39658
2 94326 1 39658
2 94327 1 39680
2 94328 1 39680
2 94329 1 39692
2 94330 1 39692
2 94331 1 39716
2 94332 1 39716
2 94333 1 39755
2 94334 1 39755
2 94335 1 39756
2 94336 1 39756
2 94337 1 39758
2 94338 1 39758
2 94339 1 39758
2 94340 1 39771
2 94341 1 39771
2 94342 1 39771
2 94343 1 39779
2 94344 1 39779
2 94345 1 39801
2 94346 1 39801
2 94347 1 39801
2 94348 1 39801
2 94349 1 39802
2 94350 1 39802
2 94351 1 39860
2 94352 1 39860
2 94353 1 39868
2 94354 1 39868
2 94355 1 39897
2 94356 1 39897
2 94357 1 39898
2 94358 1 39898
2 94359 1 39917
2 94360 1 39917
2 94361 1 39925
2 94362 1 39925
2 94363 1 39926
2 94364 1 39926
2 94365 1 39965
2 94366 1 39965
2 94367 1 39992
2 94368 1 39992
2 94369 1 40063
2 94370 1 40063
2 94371 1 40066
2 94372 1 40066
2 94373 1 40094
2 94374 1 40094
2 94375 1 40094
2 94376 1 40115
2 94377 1 40115
2 94378 1 40129
2 94379 1 40129
2 94380 1 40129
2 94381 1 40130
2 94382 1 40130
2 94383 1 40130
2 94384 1 40130
2 94385 1 40130
2 94386 1 40131
2 94387 1 40131
2 94388 1 40167
2 94389 1 40167
2 94390 1 40173
2 94391 1 40173
2 94392 1 40196
2 94393 1 40196
2 94394 1 40203
2 94395 1 40203
2 94396 1 40218
2 94397 1 40218
2 94398 1 40220
2 94399 1 40220
2 94400 1 40242
2 94401 1 40242
2 94402 1 40242
2 94403 1 40243
2 94404 1 40243
2 94405 1 40249
2 94406 1 40249
2 94407 1 40249
2 94408 1 40249
2 94409 1 40250
2 94410 1 40250
2 94411 1 40318
2 94412 1 40318
2 94413 1 40327
2 94414 1 40327
2 94415 1 40357
2 94416 1 40357
2 94417 1 40372
2 94418 1 40372
2 94419 1 40373
2 94420 1 40373
2 94421 1 40394
2 94422 1 40394
2 94423 1 40394
2 94424 1 40394
2 94425 1 40394
2 94426 1 40400
2 94427 1 40400
2 94428 1 40412
2 94429 1 40412
2 94430 1 40412
2 94431 1 40417
2 94432 1 40417
2 94433 1 40450
2 94434 1 40450
2 94435 1 40450
2 94436 1 40454
2 94437 1 40454
2 94438 1 40464
2 94439 1 40464
2 94440 1 40501
2 94441 1 40501
2 94442 1 40501
2 94443 1 40515
2 94444 1 40515
2 94445 1 40522
2 94446 1 40522
2 94447 1 40534
2 94448 1 40534
2 94449 1 40552
2 94450 1 40552
2 94451 1 40560
2 94452 1 40560
2 94453 1 40563
2 94454 1 40563
2 94455 1 40564
2 94456 1 40564
2 94457 1 40576
2 94458 1 40576
2 94459 1 40579
2 94460 1 40579
2 94461 1 40582
2 94462 1 40582
2 94463 1 40620
2 94464 1 40620
2 94465 1 40629
2 94466 1 40629
2 94467 1 40629
2 94468 1 40639
2 94469 1 40639
2 94470 1 40653
2 94471 1 40653
2 94472 1 40653
2 94473 1 40657
2 94474 1 40657
2 94475 1 40663
2 94476 1 40663
2 94477 1 40663
2 94478 1 40674
2 94479 1 40674
2 94480 1 40723
2 94481 1 40723
2 94482 1 40725
2 94483 1 40725
2 94484 1 40735
2 94485 1 40735
2 94486 1 40735
2 94487 1 40735
2 94488 1 40743
2 94489 1 40743
2 94490 1 40794
2 94491 1 40794
2 94492 1 40830
2 94493 1 40830
2 94494 1 40838
2 94495 1 40838
2 94496 1 40838
2 94497 1 40849
2 94498 1 40849
2 94499 1 40878
2 94500 1 40878
2 94501 1 40878
2 94502 1 40878
2 94503 1 40878
2 94504 1 40896
2 94505 1 40896
2 94506 1 40896
2 94507 1 40924
2 94508 1 40924
2 94509 1 40928
2 94510 1 40928
2 94511 1 40928
2 94512 1 40935
2 94513 1 40935
2 94514 1 40935
2 94515 1 40935
2 94516 1 40942
2 94517 1 40942
2 94518 1 40942
2 94519 1 40942
2 94520 1 40942
2 94521 1 40942
2 94522 1 40943
2 94523 1 40943
2 94524 1 40943
2 94525 1 40943
2 94526 1 40944
2 94527 1 40944
2 94528 1 40944
2 94529 1 40971
2 94530 1 40971
2 94531 1 40972
2 94532 1 40972
2 94533 1 40975
2 94534 1 40975
2 94535 1 40982
2 94536 1 40982
2 94537 1 40982
2 94538 1 40982
2 94539 1 40982
2 94540 1 41008
2 94541 1 41008
2 94542 1 41008
2 94543 1 41008
2 94544 1 41020
2 94545 1 41020
2 94546 1 41021
2 94547 1 41021
2 94548 1 41021
2 94549 1 41022
2 94550 1 41022
2 94551 1 41032
2 94552 1 41032
2 94553 1 41032
2 94554 1 41045
2 94555 1 41045
2 94556 1 41068
2 94557 1 41068
2 94558 1 41119
2 94559 1 41119
2 94560 1 41126
2 94561 1 41126
2 94562 1 41155
2 94563 1 41155
2 94564 1 41166
2 94565 1 41166
2 94566 1 41169
2 94567 1 41169
2 94568 1 41201
2 94569 1 41201
2 94570 1 41201
2 94571 1 41308
2 94572 1 41308
2 94573 1 41347
2 94574 1 41347
2 94575 1 41356
2 94576 1 41356
2 94577 1 41383
2 94578 1 41383
2 94579 1 41384
2 94580 1 41384
2 94581 1 41477
2 94582 1 41477
2 94583 1 41481
2 94584 1 41481
2 94585 1 41492
2 94586 1 41492
2 94587 1 41499
2 94588 1 41499
2 94589 1 41558
2 94590 1 41558
2 94591 1 41573
2 94592 1 41573
2 94593 1 41580
2 94594 1 41580
2 94595 1 41581
2 94596 1 41581
2 94597 1 41581
2 94598 1 41582
2 94599 1 41582
2 94600 1 41586
2 94601 1 41586
2 94602 1 41598
2 94603 1 41598
2 94604 1 41611
2 94605 1 41611
2 94606 1 41611
2 94607 1 41613
2 94608 1 41613
2 94609 1 41699
2 94610 1 41699
2 94611 1 41700
2 94612 1 41700
2 94613 1 41700
2 94614 1 41723
2 94615 1 41723
2 94616 1 41734
2 94617 1 41734
2 94618 1 41738
2 94619 1 41738
2 94620 1 41762
2 94621 1 41762
2 94622 1 41773
2 94623 1 41773
2 94624 1 41795
2 94625 1 41795
2 94626 1 41797
2 94627 1 41797
2 94628 1 41806
2 94629 1 41806
2 94630 1 41827
2 94631 1 41827
2 94632 1 41827
2 94633 1 41827
2 94634 1 41827
2 94635 1 41827
2 94636 1 41828
2 94637 1 41828
2 94638 1 41828
2 94639 1 41828
2 94640 1 41866
2 94641 1 41866
2 94642 1 41866
2 94643 1 41876
2 94644 1 41876
2 94645 1 41876
2 94646 1 41877
2 94647 1 41877
2 94648 1 41896
2 94649 1 41896
2 94650 1 41919
2 94651 1 41919
2 94652 1 41919
2 94653 1 41919
2 94654 1 41919
2 94655 1 41919
2 94656 1 41919
2 94657 1 41919
2 94658 1 41919
2 94659 1 41928
2 94660 1 41928
2 94661 1 41930
2 94662 1 41930
2 94663 1 41930
2 94664 1 41934
2 94665 1 41934
2 94666 1 41940
2 94667 1 41940
2 94668 1 41940
2 94669 1 41941
2 94670 1 41941
2 94671 1 41946
2 94672 1 41946
2 94673 1 41946
2 94674 1 41960
2 94675 1 41960
2 94676 1 41962
2 94677 1 41962
2 94678 1 41980
2 94679 1 41980
2 94680 1 41986
2 94681 1 41986
2 94682 1 41996
2 94683 1 41996
2 94684 1 42034
2 94685 1 42034
2 94686 1 42035
2 94687 1 42035
2 94688 1 42035
2 94689 1 42035
2 94690 1 42036
2 94691 1 42036
2 94692 1 42071
2 94693 1 42071
2 94694 1 42087
2 94695 1 42087
2 94696 1 42087
2 94697 1 42099
2 94698 1 42099
2 94699 1 42099
2 94700 1 42099
2 94701 1 42100
2 94702 1 42100
2 94703 1 42106
2 94704 1 42106
2 94705 1 42124
2 94706 1 42124
2 94707 1 42124
2 94708 1 42141
2 94709 1 42141
2 94710 1 42145
2 94711 1 42145
2 94712 1 42164
2 94713 1 42164
2 94714 1 42164
2 94715 1 42164
2 94716 1 42165
2 94717 1 42165
2 94718 1 42195
2 94719 1 42195
2 94720 1 42211
2 94721 1 42211
2 94722 1 42231
2 94723 1 42231
2 94724 1 42244
2 94725 1 42244
2 94726 1 42263
2 94727 1 42263
2 94728 1 42293
2 94729 1 42293
2 94730 1 42293
2 94731 1 42295
2 94732 1 42295
2 94733 1 42295
2 94734 1 42299
2 94735 1 42299
2 94736 1 42318
2 94737 1 42318
2 94738 1 42319
2 94739 1 42319
2 94740 1 42320
2 94741 1 42320
2 94742 1 42341
2 94743 1 42341
2 94744 1 42345
2 94745 1 42345
2 94746 1 42345
2 94747 1 42345
2 94748 1 42345
2 94749 1 42345
2 94750 1 42375
2 94751 1 42375
2 94752 1 42379
2 94753 1 42379
2 94754 1 42446
2 94755 1 42446
2 94756 1 42468
2 94757 1 42468
2 94758 1 42476
2 94759 1 42476
2 94760 1 42481
2 94761 1 42481
2 94762 1 42514
2 94763 1 42514
2 94764 1 42525
2 94765 1 42525
2 94766 1 42568
2 94767 1 42568
2 94768 1 42568
2 94769 1 42592
2 94770 1 42592
2 94771 1 42641
2 94772 1 42641
2 94773 1 42666
2 94774 1 42666
2 94775 1 42669
2 94776 1 42669
2 94777 1 42675
2 94778 1 42675
2 94779 1 42714
2 94780 1 42714
2 94781 1 42720
2 94782 1 42720
2 94783 1 42723
2 94784 1 42723
2 94785 1 42796
2 94786 1 42796
2 94787 1 42850
2 94788 1 42850
2 94789 1 42910
2 94790 1 42910
2 94791 1 42915
2 94792 1 42915
2 94793 1 42918
2 94794 1 42918
2 94795 1 42927
2 94796 1 42927
2 94797 1 42929
2 94798 1 42929
2 94799 1 42943
2 94800 1 42943
2 94801 1 42943
2 94802 1 42943
2 94803 1 42944
2 94804 1 42944
2 94805 1 42944
2 94806 1 42966
2 94807 1 42966
2 94808 1 42975
2 94809 1 42975
2 94810 1 43002
2 94811 1 43002
2 94812 1 43006
2 94813 1 43006
2 94814 1 43016
2 94815 1 43016
2 94816 1 43030
2 94817 1 43030
2 94818 1 43034
2 94819 1 43034
2 94820 1 43039
2 94821 1 43039
2 94822 1 43059
2 94823 1 43059
2 94824 1 43085
2 94825 1 43085
2 94826 1 43106
2 94827 1 43106
2 94828 1 43106
2 94829 1 43106
2 94830 1 43112
2 94831 1 43112
2 94832 1 43152
2 94833 1 43152
2 94834 1 43169
2 94835 1 43169
2 94836 1 43183
2 94837 1 43183
2 94838 1 43184
2 94839 1 43184
2 94840 1 43213
2 94841 1 43213
2 94842 1 43213
2 94843 1 43221
2 94844 1 43221
2 94845 1 43222
2 94846 1 43222
2 94847 1 43224
2 94848 1 43224
2 94849 1 43225
2 94850 1 43225
2 94851 1 43225
2 94852 1 43225
2 94853 1 43225
2 94854 1 43225
2 94855 1 43225
2 94856 1 43225
2 94857 1 43225
2 94858 1 43228
2 94859 1 43228
2 94860 1 43236
2 94861 1 43236
2 94862 1 43255
2 94863 1 43255
2 94864 1 43258
2 94865 1 43258
2 94866 1 43264
2 94867 1 43264
2 94868 1 43264
2 94869 1 43265
2 94870 1 43265
2 94871 1 43265
2 94872 1 43271
2 94873 1 43271
2 94874 1 43298
2 94875 1 43298
2 94876 1 43344
2 94877 1 43344
2 94878 1 43350
2 94879 1 43350
2 94880 1 43350
2 94881 1 43350
2 94882 1 43370
2 94883 1 43370
2 94884 1 43389
2 94885 1 43389
2 94886 1 43389
2 94887 1 43417
2 94888 1 43417
2 94889 1 43441
2 94890 1 43441
2 94891 1 43521
2 94892 1 43521
2 94893 1 43541
2 94894 1 43541
2 94895 1 43601
2 94896 1 43601
2 94897 1 43616
2 94898 1 43616
2 94899 1 43620
2 94900 1 43620
2 94901 1 43632
2 94902 1 43632
2 94903 1 43637
2 94904 1 43637
2 94905 1 43639
2 94906 1 43639
2 94907 1 43656
2 94908 1 43656
2 94909 1 43675
2 94910 1 43675
2 94911 1 43678
2 94912 1 43678
2 94913 1 43688
2 94914 1 43688
2 94915 1 43748
2 94916 1 43748
2 94917 1 43748
2 94918 1 43749
2 94919 1 43749
2 94920 1 43766
2 94921 1 43766
2 94922 1 43819
2 94923 1 43819
2 94924 1 43836
2 94925 1 43836
2 94926 1 43837
2 94927 1 43837
2 94928 1 43837
2 94929 1 43846
2 94930 1 43846
2 94931 1 43846
2 94932 1 43846
2 94933 1 43846
2 94934 1 43846
2 94935 1 43846
2 94936 1 43847
2 94937 1 43847
2 94938 1 43848
2 94939 1 43848
2 94940 1 43876
2 94941 1 43876
2 94942 1 43876
2 94943 1 43896
2 94944 1 43896
2 94945 1 43898
2 94946 1 43898
2 94947 1 43908
2 94948 1 43908
2 94949 1 43938
2 94950 1 43938
2 94951 1 43979
2 94952 1 43979
2 94953 1 44006
2 94954 1 44006
2 94955 1 44006
2 94956 1 44016
2 94957 1 44016
2 94958 1 44016
2 94959 1 44029
2 94960 1 44029
2 94961 1 44032
2 94962 1 44032
2 94963 1 44048
2 94964 1 44048
2 94965 1 44048
2 94966 1 44056
2 94967 1 44056
2 94968 1 44056
2 94969 1 44056
2 94970 1 44062
2 94971 1 44062
2 94972 1 44062
2 94973 1 44116
2 94974 1 44116
2 94975 1 44118
2 94976 1 44118
2 94977 1 44137
2 94978 1 44137
2 94979 1 44167
2 94980 1 44167
2 94981 1 44167
2 94982 1 44167
2 94983 1 44167
2 94984 1 44170
2 94985 1 44170
2 94986 1 44179
2 94987 1 44179
2 94988 1 44182
2 94989 1 44182
2 94990 1 44205
2 94991 1 44205
2 94992 1 44218
2 94993 1 44218
2 94994 1 44218
2 94995 1 44230
2 94996 1 44230
2 94997 1 44257
2 94998 1 44257
2 94999 1 44260
2 95000 1 44260
2 95001 1 44260
2 95002 1 44276
2 95003 1 44276
2 95004 1 44281
2 95005 1 44281
2 95006 1 44316
2 95007 1 44316
2 95008 1 44342
2 95009 1 44342
2 95010 1 44359
2 95011 1 44359
2 95012 1 44359
2 95013 1 44366
2 95014 1 44366
2 95015 1 44374
2 95016 1 44374
2 95017 1 44374
2 95018 1 44376
2 95019 1 44376
2 95020 1 44378
2 95021 1 44378
2 95022 1 44378
2 95023 1 44406
2 95024 1 44406
2 95025 1 44407
2 95026 1 44407
2 95027 1 44407
2 95028 1 44407
2 95029 1 44443
2 95030 1 44443
2 95031 1 44511
2 95032 1 44511
2 95033 1 44562
2 95034 1 44562
2 95035 1 44676
2 95036 1 44676
2 95037 1 44677
2 95038 1 44677
2 95039 1 44677
2 95040 1 44681
2 95041 1 44681
2 95042 1 44690
2 95043 1 44690
2 95044 1 44690
2 95045 1 44692
2 95046 1 44692
2 95047 1 44696
2 95048 1 44696
2 95049 1 44700
2 95050 1 44700
2 95051 1 44717
2 95052 1 44717
2 95053 1 44724
2 95054 1 44724
2 95055 1 44736
2 95056 1 44736
2 95057 1 44776
2 95058 1 44776
2 95059 1 44788
2 95060 1 44788
2 95061 1 44927
2 95062 1 44927
2 95063 1 44937
2 95064 1 44937
2 95065 1 44952
2 95066 1 44952
2 95067 1 44952
2 95068 1 44953
2 95069 1 44953
2 95070 1 44961
2 95071 1 44961
2 95072 1 45024
2 95073 1 45024
2 95074 1 45044
2 95075 1 45044
2 95076 1 45053
2 95077 1 45053
2 95078 1 45121
2 95079 1 45121
2 95080 1 45159
2 95081 1 45159
2 95082 1 45189
2 95083 1 45189
2 95084 1 45192
2 95085 1 45192
2 95086 1 45227
2 95087 1 45227
2 95088 1 45244
2 95089 1 45244
2 95090 1 45267
2 95091 1 45267
2 95092 1 45373
2 95093 1 45373
2 95094 1 45382
2 95095 1 45382
2 95096 1 45387
2 95097 1 45387
2 95098 1 45390
2 95099 1 45390
2 95100 1 45390
2 95101 1 45390
2 95102 1 45391
2 95103 1 45391
2 95104 1 45391
2 95105 1 45450
2 95106 1 45450
2 95107 1 45451
2 95108 1 45451
2 95109 1 45464
2 95110 1 45464
2 95111 1 45464
2 95112 1 45524
2 95113 1 45524
2 95114 1 45569
2 95115 1 45569
2 95116 1 45570
2 95117 1 45570
2 95118 1 45613
2 95119 1 45613
2 95120 1 45619
2 95121 1 45619
2 95122 1 45619
2 95123 1 45685
2 95124 1 45685
2 95125 1 45686
2 95126 1 45686
2 95127 1 45687
2 95128 1 45687
2 95129 1 45720
2 95130 1 45720
2 95131 1 45747
2 95132 1 45747
2 95133 1 45840
2 95134 1 45840
2 95135 1 45862
2 95136 1 45862
2 95137 1 45864
2 95138 1 45864
2 95139 1 45868
2 95140 1 45868
2 95141 1 45868
2 95142 1 45868
2 95143 1 45871
2 95144 1 45871
2 95145 1 45873
2 95146 1 45873
2 95147 1 45887
2 95148 1 45887
2 95149 1 45887
2 95150 1 45887
2 95151 1 45887
2 95152 1 45902
2 95153 1 45902
2 95154 1 45905
2 95155 1 45905
2 95156 1 45913
2 95157 1 45913
2 95158 1 45926
2 95159 1 45926
2 95160 1 45927
2 95161 1 45927
2 95162 1 45942
2 95163 1 45942
2 95164 1 45979
2 95165 1 45979
2 95166 1 45979
2 95167 1 46000
2 95168 1 46000
2 95169 1 46008
2 95170 1 46008
2 95171 1 46019
2 95172 1 46019
2 95173 1 46182
2 95174 1 46182
2 95175 1 46182
2 95176 1 46194
2 95177 1 46194
2 95178 1 46202
2 95179 1 46202
2 95180 1 46328
2 95181 1 46328
2 95182 1 46379
2 95183 1 46379
2 95184 1 46408
2 95185 1 46408
2 95186 1 46408
2 95187 1 46420
2 95188 1 46420
2 95189 1 46445
2 95190 1 46445
2 95191 1 46470
2 95192 1 46470
2 95193 1 46480
2 95194 1 46480
2 95195 1 46480
2 95196 1 46516
2 95197 1 46516
2 95198 1 46516
2 95199 1 46629
2 95200 1 46629
2 95201 1 46630
2 95202 1 46630
2 95203 1 46633
2 95204 1 46633
2 95205 1 46669
2 95206 1 46669
2 95207 1 46669
2 95208 1 46670
2 95209 1 46670
2 95210 1 46671
2 95211 1 46671
2 95212 1 46682
2 95213 1 46682
2 95214 1 46727
2 95215 1 46727
2 95216 1 46727
2 95217 1 46764
2 95218 1 46764
2 95219 1 46764
2 95220 1 46776
2 95221 1 46776
2 95222 1 46784
2 95223 1 46784
2 95224 1 46789
2 95225 1 46789
2 95226 1 46802
2 95227 1 46802
2 95228 1 46802
2 95229 1 46802
2 95230 1 46802
2 95231 1 46808
2 95232 1 46808
2 95233 1 46816
2 95234 1 46816
2 95235 1 46816
2 95236 1 46942
2 95237 1 46942
2 95238 1 46982
2 95239 1 46982
2 95240 1 47005
2 95241 1 47005
2 95242 1 47023
2 95243 1 47023
2 95244 1 47057
2 95245 1 47057
2 95246 1 47057
2 95247 1 47057
2 95248 1 47057
2 95249 1 47057
2 95250 1 47085
2 95251 1 47085
2 95252 1 47145
2 95253 1 47145
2 95254 1 47154
2 95255 1 47154
2 95256 1 47154
2 95257 1 47164
2 95258 1 47164
2 95259 1 47168
2 95260 1 47168
2 95261 1 47188
2 95262 1 47188
2 95263 1 47188
2 95264 1 47188
2 95265 1 47188
2 95266 1 47188
2 95267 1 47188
2 95268 1 47189
2 95269 1 47189
2 95270 1 47201
2 95271 1 47201
2 95272 1 47202
2 95273 1 47202
2 95274 1 47214
2 95275 1 47214
2 95276 1 47214
2 95277 1 47239
2 95278 1 47239
2 95279 1 47239
2 95280 1 47263
2 95281 1 47263
2 95282 1 47276
2 95283 1 47276
2 95284 1 47298
2 95285 1 47298
2 95286 1 47305
2 95287 1 47305
2 95288 1 47305
2 95289 1 47312
2 95290 1 47312
2 95291 1 47312
2 95292 1 47317
2 95293 1 47317
2 95294 1 47324
2 95295 1 47324
2 95296 1 47324
2 95297 1 47350
2 95298 1 47350
2 95299 1 47352
2 95300 1 47352
2 95301 1 47354
2 95302 1 47354
2 95303 1 47384
2 95304 1 47384
2 95305 1 47385
2 95306 1 47385
2 95307 1 47388
2 95308 1 47388
2 95309 1 47388
2 95310 1 47390
2 95311 1 47390
2 95312 1 47396
2 95313 1 47396
2 95314 1 47396
2 95315 1 47396
2 95316 1 47397
2 95317 1 47397
2 95318 1 47463
2 95319 1 47463
2 95320 1 47468
2 95321 1 47468
2 95322 1 47518
2 95323 1 47518
2 95324 1 47518
2 95325 1 47551
2 95326 1 47551
2 95327 1 47613
2 95328 1 47613
2 95329 1 47626
2 95330 1 47626
2 95331 1 47651
2 95332 1 47651
2 95333 1 47651
2 95334 1 47651
2 95335 1 47651
2 95336 1 47675
2 95337 1 47675
2 95338 1 47681
2 95339 1 47681
2 95340 1 47698
2 95341 1 47698
2 95342 1 47715
2 95343 1 47715
2 95344 1 47716
2 95345 1 47716
2 95346 1 47742
2 95347 1 47742
2 95348 1 47743
2 95349 1 47743
2 95350 1 47744
2 95351 1 47744
2 95352 1 47752
2 95353 1 47752
2 95354 1 47765
2 95355 1 47765
2 95356 1 47765
2 95357 1 47765
2 95358 1 47765
2 95359 1 47765
2 95360 1 47774
2 95361 1 47774
2 95362 1 47774
2 95363 1 47802
2 95364 1 47802
2 95365 1 47820
2 95366 1 47820
2 95367 1 47856
2 95368 1 47856
2 95369 1 47856
2 95370 1 47856
2 95371 1 47860
2 95372 1 47860
2 95373 1 47954
2 95374 1 47954
2 95375 1 47980
2 95376 1 47980
2 95377 1 48007
2 95378 1 48007
2 95379 1 48019
2 95380 1 48019
2 95381 1 48028
2 95382 1 48028
2 95383 1 48038
2 95384 1 48038
2 95385 1 48039
2 95386 1 48039
2 95387 1 48039
2 95388 1 48110
2 95389 1 48110
2 95390 1 48111
2 95391 1 48111
2 95392 1 48125
2 95393 1 48125
2 95394 1 48126
2 95395 1 48126
2 95396 1 48135
2 95397 1 48135
2 95398 1 48188
2 95399 1 48188
2 95400 1 48192
2 95401 1 48192
2 95402 1 48199
2 95403 1 48199
2 95404 1 48213
2 95405 1 48213
2 95406 1 48213
2 95407 1 48229
2 95408 1 48229
2 95409 1 48317
2 95410 1 48317
2 95411 1 48359
2 95412 1 48359
2 95413 1 48360
2 95414 1 48360
2 95415 1 48368
2 95416 1 48368
2 95417 1 48368
2 95418 1 48368
2 95419 1 48368
2 95420 1 48402
2 95421 1 48402
2 95422 1 48410
2 95423 1 48410
2 95424 1 48413
2 95425 1 48413
2 95426 1 48457
2 95427 1 48457
2 95428 1 48457
2 95429 1 48470
2 95430 1 48470
2 95431 1 48509
2 95432 1 48509
2 95433 1 48521
2 95434 1 48521
2 95435 1 48548
2 95436 1 48548
2 95437 1 48550
2 95438 1 48550
2 95439 1 48569
2 95440 1 48569
2 95441 1 48597
2 95442 1 48597
2 95443 1 48601
2 95444 1 48601
2 95445 1 48601
2 95446 1 48611
2 95447 1 48611
2 95448 1 48615
2 95449 1 48615
2 95450 1 48639
2 95451 1 48639
2 95452 1 48639
2 95453 1 48675
2 95454 1 48675
2 95455 1 48689
2 95456 1 48689
2 95457 1 48689
2 95458 1 48689
2 95459 1 48692
2 95460 1 48692
2 95461 1 48693
2 95462 1 48693
2 95463 1 48706
2 95464 1 48706
2 95465 1 48707
2 95466 1 48707
2 95467 1 48732
2 95468 1 48732
2 95469 1 48732
2 95470 1 48733
2 95471 1 48733
2 95472 1 48760
2 95473 1 48760
2 95474 1 48768
2 95475 1 48768
2 95476 1 48788
2 95477 1 48788
2 95478 1 48788
2 95479 1 48799
2 95480 1 48799
2 95481 1 48800
2 95482 1 48800
2 95483 1 48802
2 95484 1 48802
2 95485 1 48802
2 95486 1 48822
2 95487 1 48822
2 95488 1 48824
2 95489 1 48824
2 95490 1 48824
2 95491 1 48850
2 95492 1 48850
2 95493 1 48850
2 95494 1 48862
2 95495 1 48862
2 95496 1 48862
2 95497 1 48862
2 95498 1 48862
2 95499 1 48874
2 95500 1 48874
2 95501 1 48874
2 95502 1 48875
2 95503 1 48875
2 95504 1 48878
2 95505 1 48878
2 95506 1 48929
2 95507 1 48929
2 95508 1 48961
2 95509 1 48961
2 95510 1 49009
2 95511 1 49009
2 95512 1 49068
2 95513 1 49068
2 95514 1 49114
2 95515 1 49114
2 95516 1 49114
2 95517 1 49147
2 95518 1 49147
2 95519 1 49197
2 95520 1 49197
2 95521 1 49221
2 95522 1 49221
2 95523 1 49236
2 95524 1 49236
2 95525 1 49237
2 95526 1 49237
2 95527 1 49237
2 95528 1 49254
2 95529 1 49254
2 95530 1 49257
2 95531 1 49257
2 95532 1 49271
2 95533 1 49271
2 95534 1 49286
2 95535 1 49286
2 95536 1 49286
2 95537 1 49286
2 95538 1 49289
2 95539 1 49289
2 95540 1 49289
2 95541 1 49337
2 95542 1 49337
2 95543 1 49361
2 95544 1 49361
2 95545 1 49383
2 95546 1 49383
2 95547 1 49391
2 95548 1 49391
2 95549 1 49399
2 95550 1 49399
2 95551 1 49399
2 95552 1 49409
2 95553 1 49409
2 95554 1 49440
2 95555 1 49440
2 95556 1 49440
2 95557 1 49456
2 95558 1 49456
2 95559 1 49478
2 95560 1 49478
2 95561 1 49518
2 95562 1 49518
2 95563 1 49539
2 95564 1 49539
2 95565 1 49594
2 95566 1 49594
2 95567 1 49605
2 95568 1 49605
2 95569 1 49655
2 95570 1 49655
2 95571 1 49668
2 95572 1 49668
2 95573 1 49670
2 95574 1 49670
2 95575 1 49685
2 95576 1 49685
2 95577 1 49780
2 95578 1 49780
2 95579 1 49793
2 95580 1 49793
2 95581 1 49915
2 95582 1 49915
2 95583 1 49955
2 95584 1 49955
2 95585 1 50021
2 95586 1 50021
2 95587 1 50055
2 95588 1 50055
2 95589 1 50058
2 95590 1 50058
2 95591 1 50094
2 95592 1 50094
2 95593 1 50102
2 95594 1 50102
2 95595 1 50115
2 95596 1 50115
2 95597 1 50115
2 95598 1 50126
2 95599 1 50126
2 95600 1 50138
2 95601 1 50138
2 95602 1 50154
2 95603 1 50154
2 95604 1 50231
2 95605 1 50231
2 95606 1 50262
2 95607 1 50262
2 95608 1 50262
2 95609 1 50263
2 95610 1 50263
2 95611 1 50263
2 95612 1 50388
2 95613 1 50388
2 95614 1 50466
2 95615 1 50466
2 95616 1 50480
2 95617 1 50480
2 95618 1 50480
2 95619 1 50484
2 95620 1 50484
2 95621 1 50485
2 95622 1 50485
2 95623 1 50505
2 95624 1 50505
2 95625 1 50630
2 95626 1 50630
2 95627 1 50631
2 95628 1 50631
2 95629 1 50656
2 95630 1 50656
2 95631 1 50761
2 95632 1 50761
2 95633 1 50873
2 95634 1 50873
2 95635 1 50926
2 95636 1 50926
2 95637 1 50933
2 95638 1 50933
2 95639 1 50962
2 95640 1 50962
2 95641 1 50965
2 95642 1 50965
2 95643 1 51040
2 95644 1 51040
2 95645 1 51123
2 95646 1 51123
2 95647 1 51184
2 95648 1 51184
2 95649 1 51196
2 95650 1 51196
2 95651 1 51215
2 95652 1 51215
2 95653 1 51290
2 95654 1 51290
2 95655 1 51290
2 95656 1 51306
2 95657 1 51306
2 95658 1 51313
2 95659 1 51313
2 95660 1 51313
2 95661 1 51314
2 95662 1 51314
2 95663 1 51316
2 95664 1 51316
2 95665 1 51328
2 95666 1 51328
2 95667 1 51338
2 95668 1 51338
2 95669 1 51355
2 95670 1 51355
2 95671 1 51356
2 95672 1 51356
2 95673 1 51356
2 95674 1 51376
2 95675 1 51376
2 95676 1 51382
2 95677 1 51382
2 95678 1 51471
2 95679 1 51471
2 95680 1 51479
2 95681 1 51479
2 95682 1 51487
2 95683 1 51487
2 95684 1 51487
2 95685 1 51493
2 95686 1 51493
2 95687 1 51541
2 95688 1 51541
2 95689 1 51546
2 95690 1 51546
2 95691 1 51549
2 95692 1 51549
2 95693 1 51554
2 95694 1 51554
2 95695 1 51555
2 95696 1 51555
2 95697 1 51555
2 95698 1 51561
2 95699 1 51561
2 95700 1 51566
2 95701 1 51566
2 95702 1 51576
2 95703 1 51576
2 95704 1 51581
2 95705 1 51581
2 95706 1 51585
2 95707 1 51585
2 95708 1 51591
2 95709 1 51591
2 95710 1 51592
2 95711 1 51592
2 95712 1 51597
2 95713 1 51597
2 95714 1 51606
2 95715 1 51606
2 95716 1 51612
2 95717 1 51612
2 95718 1 51613
2 95719 1 51613
2 95720 1 51615
2 95721 1 51615
2 95722 1 51621
2 95723 1 51621
2 95724 1 51629
2 95725 1 51629
2 95726 1 51635
2 95727 1 51635
2 95728 1 51664
2 95729 1 51664
2 95730 1 51719
2 95731 1 51719
2 95732 1 51719
2 95733 1 51731
2 95734 1 51731
2 95735 1 51731
2 95736 1 51735
2 95737 1 51735
2 95738 1 51743
2 95739 1 51743
2 95740 1 51801
2 95741 1 51801
2 95742 1 51815
2 95743 1 51815
2 95744 1 51815
2 95745 1 51815
2 95746 1 51822
2 95747 1 51822
2 95748 1 51852
2 95749 1 51852
2 95750 1 51859
2 95751 1 51859
2 95752 1 51887
2 95753 1 51887
2 95754 1 51919
2 95755 1 51919
2 95756 1 52024
2 95757 1 52024
2 95758 1 52031
2 95759 1 52031
2 95760 1 52034
2 95761 1 52034
2 95762 1 52035
2 95763 1 52035
2 95764 1 52035
2 95765 1 52035
2 95766 1 52037
2 95767 1 52037
2 95768 1 52055
2 95769 1 52055
2 95770 1 52059
2 95771 1 52059
2 95772 1 52072
2 95773 1 52072
2 95774 1 52080
2 95775 1 52080
2 95776 1 52091
2 95777 1 52091
2 95778 1 52112
2 95779 1 52112
2 95780 1 52125
2 95781 1 52125
2 95782 1 52126
2 95783 1 52126
2 95784 1 52147
2 95785 1 52147
2 95786 1 52196
2 95787 1 52196
2 95788 1 52199
2 95789 1 52199
2 95790 1 52215
2 95791 1 52215
2 95792 1 52215
2 95793 1 52243
2 95794 1 52243
2 95795 1 52260
2 95796 1 52260
2 95797 1 52265
2 95798 1 52265
2 95799 1 52286
2 95800 1 52286
2 95801 1 52286
2 95802 1 52320
2 95803 1 52320
2 95804 1 52321
2 95805 1 52321
2 95806 1 52330
2 95807 1 52330
2 95808 1 52330
2 95809 1 52361
2 95810 1 52361
2 95811 1 52423
2 95812 1 52423
2 95813 1 52439
2 95814 1 52439
2 95815 1 52469
2 95816 1 52469
2 95817 1 52476
2 95818 1 52476
2 95819 1 52476
2 95820 1 52478
2 95821 1 52478
2 95822 1 52479
2 95823 1 52479
2 95824 1 52479
2 95825 1 52533
2 95826 1 52533
2 95827 1 52533
2 95828 1 52541
2 95829 1 52541
2 95830 1 52542
2 95831 1 52542
2 95832 1 52569
2 95833 1 52569
2 95834 1 52663
2 95835 1 52663
2 95836 1 52675
2 95837 1 52675
2 95838 1 52711
2 95839 1 52711
2 95840 1 52728
2 95841 1 52728
2 95842 1 52730
2 95843 1 52730
2 95844 1 52760
2 95845 1 52760
2 95846 1 52760
2 95847 1 52833
2 95848 1 52833
2 95849 1 52853
2 95850 1 52853
2 95851 1 52856
2 95852 1 52856
2 95853 1 52856
2 95854 1 52856
2 95855 1 52939
2 95856 1 52939
2 95857 1 52940
2 95858 1 52940
2 95859 1 52959
2 95860 1 52959
2 95861 1 52970
2 95862 1 52970
2 95863 1 53016
2 95864 1 53016
2 95865 1 53016
2 95866 1 53017
2 95867 1 53017
2 95868 1 53017
2 95869 1 53017
2 95870 1 53028
2 95871 1 53028
2 95872 1 53049
2 95873 1 53049
2 95874 1 53096
2 95875 1 53096
2 95876 1 53105
2 95877 1 53105
2 95878 1 53112
2 95879 1 53112
2 95880 1 53144
2 95881 1 53144
2 95882 1 53204
2 95883 1 53204
2 95884 1 53204
2 95885 1 53206
2 95886 1 53206
2 95887 1 53220
2 95888 1 53220
2 95889 1 53220
2 95890 1 53220
2 95891 1 53221
2 95892 1 53221
2 95893 1 53228
2 95894 1 53228
2 95895 1 53228
2 95896 1 53228
2 95897 1 53245
2 95898 1 53245
2 95899 1 53309
2 95900 1 53309
2 95901 1 53354
2 95902 1 53354
2 95903 1 53357
2 95904 1 53357
2 95905 1 53364
2 95906 1 53364
2 95907 1 53380
2 95908 1 53380
2 95909 1 53380
2 95910 1 53385
2 95911 1 53385
2 95912 1 53385
2 95913 1 53385
2 95914 1 53385
2 95915 1 53397
2 95916 1 53397
2 95917 1 53399
2 95918 1 53399
2 95919 1 53405
2 95920 1 53405
2 95921 1 53472
2 95922 1 53472
2 95923 1 53480
2 95924 1 53480
2 95925 1 53511
2 95926 1 53511
2 95927 1 53539
2 95928 1 53539
2 95929 1 53576
2 95930 1 53576
2 95931 1 53576
2 95932 1 53576
2 95933 1 53576
2 95934 1 53583
2 95935 1 53583
2 95936 1 53585
2 95937 1 53585
2 95938 1 53648
2 95939 1 53648
2 95940 1 53729
2 95941 1 53729
2 95942 1 53756
2 95943 1 53756
2 95944 1 53759
2 95945 1 53759
2 95946 1 53837
2 95947 1 53837
2 95948 1 53837
2 95949 1 53837
2 95950 1 53840
2 95951 1 53840
2 95952 1 53849
2 95953 1 53849
2 95954 1 53954
2 95955 1 53954
2 95956 1 54021
2 95957 1 54021
2 95958 1 54028
2 95959 1 54028
2 95960 1 54051
2 95961 1 54051
2 95962 1 54051
2 95963 1 54052
2 95964 1 54052
2 95965 1 54052
2 95966 1 54052
2 95967 1 54052
2 95968 1 54052
2 95969 1 54141
2 95970 1 54141
2 95971 1 54157
2 95972 1 54157
2 95973 1 54162
2 95974 1 54162
2 95975 1 54196
2 95976 1 54196
2 95977 1 54267
2 95978 1 54267
2 95979 1 54383
2 95980 1 54383
2 95981 1 54432
2 95982 1 54432
2 95983 1 54433
2 95984 1 54433
2 95985 1 54457
2 95986 1 54457
2 95987 1 54458
2 95988 1 54458
2 95989 1 54465
2 95990 1 54465
2 95991 1 54466
2 95992 1 54466
2 95993 1 54578
2 95994 1 54578
2 95995 1 54578
2 95996 1 54594
2 95997 1 54594
2 95998 1 54594
2 95999 1 54667
2 96000 1 54667
2 96001 1 54774
2 96002 1 54774
2 96003 1 54774
2 96004 1 54789
2 96005 1 54789
2 96006 1 54789
2 96007 1 54803
2 96008 1 54803
2 96009 1 54838
2 96010 1 54838
2 96011 1 54838
2 96012 1 54838
2 96013 1 54906
2 96014 1 54906
2 96015 1 54946
2 96016 1 54946
2 96017 1 55063
2 96018 1 55063
2 96019 1 55098
2 96020 1 55098
2 96021 1 55156
2 96022 1 55156
2 96023 1 55372
2 96024 1 55372
2 96025 1 55431
2 96026 1 55431
2 96027 1 55467
2 96028 1 55467
2 96029 1 55486
2 96030 1 55486
2 96031 1 55627
2 96032 1 55627
2 96033 1 55680
2 96034 1 55680
2 96035 1 55806
2 96036 1 55806
2 96037 1 55825
2 96038 1 55825
2 96039 1 55825
2 96040 1 55861
2 96041 1 55861
2 96042 1 55909
2 96043 1 55909
2 96044 1 55916
2 96045 1 55916
2 96046 1 55939
2 96047 1 55939
2 96048 1 56069
2 96049 1 56069
2 96050 1 56161
2 96051 1 56161
2 96052 1 56183
2 96053 1 56183
2 96054 1 56184
2 96055 1 56184
2 96056 1 56184
2 96057 1 56184
2 96058 1 56199
2 96059 1 56199
2 96060 1 56200
2 96061 1 56200
2 96062 1 56460
2 96063 1 56460
2 96064 1 56644
2 96065 1 56644
2 96066 1 56645
2 96067 1 56645
2 96068 1 56645
2 96069 1 56741
2 96070 1 56741
2 96071 1 56793
2 96072 1 56793
2 96073 1 57024
2 96074 1 57024
2 96075 1 57122
2 96076 1 57122
0 27 5 140 1 25
0 28 5 259 1 57546
0 29 5 281 1 57823
0 30 5 301 1 58101
0 31 5 312 1 58376
0 32 5 125 1 58699
0 33 5 95 1 58821
0 34 5 77 1 58905
0 35 5 57 1 58918
0 36 5 134 1 59039
0 37 5 194 1 59179
0 38 5 314 1 59396
0 39 5 220 1 59709
0 40 5 107 1 59955
0 41 5 86 1 60083
0 42 5 60 1 60170
0 43 5 200 1 60202
0 44 5 257 1 60430
0 45 5 397 1 60705
0 46 5 350 1 61136
0 47 5 293 1 61503
0 48 5 132 1 61760
0 49 5 119 1 61874
0 50 5 84 1 62007
0 51 5 1 1 62142
0 52 7 60 2 63437 64653
0 53 5 8 1 66738
0 54 7 73 2 58700 59956
0 55 5 3 1 66806
0 56 7 70 2 66798 66879
0 57 5 2 1 66882
0 58 7 47 2 64760 66535
0 59 5 1 1 66954
0 60 7 15 2 57547 65106
0 61 5 11 1 67001
0 62 7 1 2 63925 67016
0 63 5 3 1 62
0 64 7 1 2 66955 67027
0 65 5 1 1 64
0 66 7 51 2 60084 61875
0 67 5 8 1 67030
0 68 7 1 2 26 67031
0 69 5 3 1 68
0 70 7 1 2 65 67089
0 71 5 1 1 70
0 72 7 1 2 57824 71
0 73 5 1 1 72
0 74 7 9 2 57548 59180
0 75 5 4 1 67092
0 76 7 6 2 65107 66536
0 77 7 5 2 64761 67105
0 78 7 1 2 67093 67111
0 79 5 1 1 78
0 80 7 7 2 57275 60085
0 81 7 3 2 61876 67116
0 82 5 1 1 67123
0 83 7 1 2 67028 67124
0 84 5 1 1 83
0 85 7 1 2 79 84
0 86 7 1 2 73 85
0 87 5 1 1 86
0 88 7 1 2 58822 87
0 89 5 1 1 88
0 90 7 110 2 62543 63926
0 91 5 181 1 67126
0 92 7 6 2 57549 67236
0 93 5 3 1 67417
0 94 7 4 2 63562 65108
0 95 7 8 2 60086 66537
0 96 7 1 2 67426 67430
0 97 7 1 2 67418 96
0 98 5 1 1 97
0 99 7 1 2 89 98
0 100 5 1 1 99
0 101 7 1 2 62008 100
0 102 5 1 1 101
0 103 7 9 2 57825 63563
0 104 7 2 2 59181 67438
0 105 7 43 2 66538 62009
0 106 7 3 2 60087 67449
0 107 5 4 1 67492
0 108 7 43 2 61877 66654
0 109 7 13 2 64762 67499
0 110 7 16 2 62284 60431
0 111 5 14 1 67555
0 112 7 1 2 57276 67571
0 113 7 1 2 67542 112
0 114 5 1 1 113
0 115 7 1 2 67495 114
0 116 5 1 1 115
0 117 7 1 2 67447 116
0 118 5 1 1 117
0 119 7 1 2 102 118
0 120 5 1 1 119
0 121 7 1 2 59040 120
0 122 5 1 1 121
0 123 7 2 2 62010 67237
0 124 7 16 2 57277 57550
0 125 5 7 1 67587
0 126 7 12 2 58823 67032
0 127 5 1 1 67610
0 128 7 1 2 67588 67611
0 129 7 1 2 67585 128
0 130 5 1 1 129
0 131 7 1 2 122 130
0 132 5 1 1 131
0 133 7 1 2 58919 132
0 134 5 1 1 133
0 135 7 84 2 57551 59041
0 136 5 103 1 67622
0 137 7 12 2 62544 67706
0 138 5 43 1 67809
0 139 7 2 2 63927 67707
0 140 5 7 1 67864
0 141 7 6 2 67821 67866
0 142 5 2 1 67873
0 143 7 19 2 67238 67874
0 144 5 2 1 67881
0 145 7 44 2 58824 60088
0 146 5 2 1 67902
0 147 7 14 2 61878 62011
0 148 7 5 2 67903 67948
0 149 7 1 2 67882 67962
0 150 5 1 1 149
0 151 7 1 2 134 150
0 152 5 1 1 151
0 153 7 1 2 64906 152
0 154 5 1 1 153
0 155 7 4 2 65109 62012
0 156 7 94 2 57826 59182
0 157 5 128 1 67971
0 158 7 2 2 67972 66956
0 159 5 1 1 68193
0 160 7 7 2 62144 63791
0 161 5 6 1 68195
0 162 7 1 2 67239 68202
0 163 7 1 2 67033 162
0 164 5 1 1 163
0 165 7 1 2 159 164
0 166 5 1 1 165
0 167 7 1 2 58825 166
0 168 5 1 1 167
0 169 7 1 2 67431 67448
0 170 5 1 1 169
0 171 7 1 2 168 170
0 172 5 1 1 171
0 173 7 1 2 57552 172
0 174 5 1 1 173
0 175 7 1 2 67973 67612
0 176 5 1 1 175
0 177 7 1 2 174 176
0 178 5 1 1 177
0 179 7 1 2 67967 178
0 180 5 1 1 179
0 181 7 1 2 154 180
0 182 5 2 1 181
0 183 7 1 2 63125 68208
0 184 5 1 1 183
0 185 7 81 2 62285 63792
0 186 5 134 1 68210
0 187 7 3 2 67974 68291
0 188 5 16 1 68425
0 189 7 103 2 62145 63734
0 190 5 103 1 68444
0 191 7 1 2 68547 67883
0 192 5 1 1 191
0 193 7 1 2 68428 192
0 194 5 7 1 193
0 195 7 11 2 58826 62013
0 196 7 23 2 60089 68657
0 197 5 11 1 68668
0 198 7 9 2 60432 61879
0 199 7 2 2 60203 68702
0 200 7 1 2 68669 68711
0 201 7 1 2 68650 200
0 202 5 2 1 201
0 203 7 1 2 184 68713
0 204 5 1 1 203
0 205 7 1 2 65363 204
0 206 5 1 1 205
0 207 7 99 2 57278 58920
0 208 5 83 1 68715
0 209 7 8 2 59042 68716
0 210 5 2 1 68897
0 211 7 5 2 58827 68898
0 212 7 12 2 59183 64907
0 213 5 2 1 68912
0 214 7 9 2 60706 61880
0 215 7 7 2 60090 68926
0 216 5 3 1 68935
0 217 7 1 2 68913 68936
0 218 7 2 2 68907 217
0 219 5 2 1 68945
0 220 7 17 2 59043 59184
0 221 5 2 1 68949
0 222 7 47 2 58921 64908
0 223 5 69 1 68968
0 224 7 3 2 59044 68969
0 225 5 4 1 69084
0 226 7 1 2 63928 69087
0 227 5 5 1 226
0 228 7 1 2 57279 69091
0 229 5 3 1 228
0 230 7 1 2 68966 69096
0 231 5 2 1 230
0 232 7 1 2 68937 69099
0 233 5 2 1 232
0 234 7 19 2 58922 59045
0 235 5 2 1 69103
0 236 7 8 2 64909 69104
0 237 7 3 2 66539 69124
0 238 7 7 2 59185 64763
0 239 7 1 2 63126 69135
0 240 7 1 2 69132 239
0 241 5 1 1 240
0 242 7 1 2 69101 241
0 243 5 1 1 242
0 244 7 1 2 58828 243
0 245 5 1 1 244
0 246 7 6 2 63564 58923
0 247 7 1 2 64910 69142
0 248 7 2 2 67432 247
0 249 5 1 1 69148
0 250 7 1 2 63127 68950
0 251 7 1 2 69149 250
0 252 5 1 1 251
0 253 7 1 2 245 252
0 254 5 1 1 253
0 255 7 1 2 57827 254
0 256 5 1 1 255
0 257 7 1 2 68947 256
0 258 5 1 1 257
0 259 7 1 2 57828 68946
0 260 5 1 1 259
0 261 7 1 2 67017 260
0 262 5 1 1 261
0 263 7 2 2 62014 262
0 264 7 1 2 258 69150
0 265 5 1 1 264
0 266 7 1 2 206 265
0 267 5 1 1 266
0 268 7 1 2 59397 267
0 269 5 1 1 268
0 270 7 6 2 65364 62015
0 271 7 10 2 65110 61881
0 272 7 5 2 69152 69158
0 273 7 26 2 57553 57829
0 274 5 3 1 69173
0 275 7 3 2 59186 69174
0 276 7 2 2 68908 69202
0 277 7 2 2 69168 69205
0 278 7 4 2 64119 60091
0 279 7 1 2 64911 69209
0 280 7 1 2 69207 279
0 281 5 1 1 280
0 282 7 1 2 269 281
0 283 5 1 1 282
0 284 7 1 2 58102 283
0 285 5 1 1 284
0 286 7 8 2 60092 60204
0 287 7 3 2 68658 69213
0 288 5 4 1 69221
0 289 7 23 2 64764 66655
0 290 7 52 2 63565 69228
0 291 7 13 2 59187 64120
0 292 7 1 2 68970 69303
0 293 7 1 2 69251 292
0 294 5 1 1 293
0 295 7 1 2 69224 294
0 296 5 1 1 295
0 297 7 1 2 57280 296
0 298 5 1 1 297
0 299 7 9 2 58924 60205
0 300 5 1 1 69316
0 301 7 1 2 69317 68670
0 302 5 1 1 301
0 303 7 1 2 298 302
0 304 5 1 1 303
0 305 7 1 2 59046 304
0 306 5 1 1 305
0 307 7 16 2 60093 62016
0 308 7 14 2 58829 69325
0 309 5 3 1 69341
0 310 7 6 2 59188 60206
0 311 5 2 1 69358
0 312 7 1 2 69342 69359
0 313 5 2 1 312
0 314 7 1 2 306 69366
0 315 5 1 1 314
0 316 7 1 2 60433 315
0 317 5 1 1 316
0 318 7 36 2 60207 60434
0 319 5 33 1 69368
0 320 7 1 2 59047 69404
0 321 5 2 1 320
0 322 7 6 2 60435 69015
0 323 5 30 1 69439
0 324 7 4 2 57281 69445
0 325 5 7 1 69475
0 326 7 1 2 69437 69479
0 327 5 1 1 326
0 328 7 4 2 58830 69210
0 329 7 1 2 62017 69486
0 330 7 1 2 327 329
0 331 5 1 1 330
0 332 7 1 2 65365 331
0 333 7 1 2 317 332
0 334 5 1 1 333
0 335 7 8 2 67904 67968
0 336 5 3 1 69490
0 337 7 1 2 69491 69100
0 338 5 1 1 337
0 339 7 8 2 64121 64912
0 340 5 2 1 69501
0 341 7 53 2 63566 64765
0 342 5 3 1 69511
0 343 7 20 2 66656 69512
0 344 5 1 1 69567
0 345 7 2 2 69502 69568
0 346 7 1 2 68899 69587
0 347 5 1 1 346
0 348 7 1 2 68691 347
0 349 5 1 1 348
0 350 7 1 2 58103 349
0 351 5 1 1 350
0 352 7 1 2 60707 351
0 353 7 1 2 338 352
0 354 5 1 1 353
0 355 7 1 2 57554 354
0 356 7 1 2 334 355
0 357 5 1 1 356
0 358 7 111 2 62018 67905
0 359 5 7 1 69589
0 360 7 11 2 58104 60708
0 361 5 7 1 69707
0 362 7 24 2 64122 65366
0 363 5 11 1 69725
0 364 7 2 2 59189 69726
0 365 5 3 1 69760
0 366 7 1 2 69718 69762
0 367 5 1 1 366
0 368 7 1 2 65111 367
0 369 5 1 1 368
0 370 7 1 2 59190 69369
0 371 5 4 1 370
0 372 7 9 2 58925 64123
0 373 7 2 2 59048 69769
0 374 7 1 2 64913 69778
0 375 5 1 1 374
0 376 7 1 2 69765 375
0 377 5 1 1 376
0 378 7 1 2 57282 377
0 379 5 1 1 378
0 380 7 12 2 63793 60208
0 381 5 5 1 69780
0 382 7 3 2 63735 69781
0 383 5 5 1 69797
0 384 7 2 2 59191 69800
0 385 5 3 1 69805
0 386 7 16 2 59398 64914
0 387 5 5 1 69810
0 388 7 23 2 60209 65112
0 389 5 4 1 69831
0 390 7 1 2 69826 69854
0 391 7 1 2 69806 390
0 392 5 1 1 391
0 393 7 3 2 58105 69370
0 394 5 2 1 69858
0 395 7 1 2 65367 69861
0 396 7 1 2 392 395
0 397 7 1 2 379 396
0 398 5 1 1 397
0 399 7 20 2 59049 64915
0 400 5 12 1 69863
0 401 7 5 2 58926 59192
0 402 7 2 2 69864 69895
0 403 5 2 1 69900
0 404 7 1 2 62824 69902
0 405 5 6 1 404
0 406 7 1 2 57283 69904
0 407 5 2 1 406
0 408 7 16 2 63794 63929
0 409 5 5 1 69912
0 410 7 1 2 58106 69928
0 411 5 2 1 410
0 412 7 1 2 60709 69933
0 413 7 1 2 69910 412
0 414 5 1 1 413
0 415 7 1 2 398 414
0 416 5 1 1 415
0 417 7 1 2 369 416
0 418 5 1 1 417
0 419 7 1 2 69590 418
0 420 5 1 1 419
0 421 7 6 2 62825 63567
0 422 7 6 2 69935 69229
0 423 7 1 2 64916 69941
0 424 7 28 2 59193 65113
0 425 5 6 1 69947
0 426 7 8 2 59050 64124
0 427 7 2 2 69948 69981
0 428 5 1 1 69989
0 429 7 9 2 58927 65368
0 430 5 4 1 69991
0 431 7 4 2 57284 69992
0 432 5 2 1 70004
0 433 7 1 2 69990 70005
0 434 7 1 2 423 433
0 435 5 1 1 434
0 436 7 1 2 420 435
0 437 7 1 2 357 436
0 438 5 1 1 437
0 439 7 1 2 57830 438
0 440 5 1 1 439
0 441 7 5 2 62286 63930
0 442 5 2 1 70010
0 443 7 8 2 63795 68445
0 444 5 4 1 70017
0 445 7 1 2 70011 70018
0 446 5 2 1 445
0 447 7 1 2 58107 70029
0 448 5 1 1 447
0 449 7 4 2 59051 68548
0 450 5 5 1 70031
0 451 7 3 2 67094 70032
0 452 5 1 1 70040
0 453 7 1 2 448 452
0 454 5 1 1 453
0 455 7 1 2 69371 454
0 456 5 1 1 455
0 457 7 3 2 60436 69883
0 458 5 5 1 70043
0 459 7 1 2 57555 69304
0 460 7 1 2 68203 459
0 461 7 1 2 70046 460
0 462 5 1 1 461
0 463 7 1 2 456 462
0 464 5 1 1 463
0 465 7 1 2 65369 464
0 466 5 1 1 465
0 467 7 12 2 58108 65114
0 468 5 7 1 70051
0 469 7 2 2 59194 70052
0 470 5 1 1 70070
0 471 7 1 2 58109 69092
0 472 5 2 1 471
0 473 7 1 2 67002 69905
0 474 5 1 1 473
0 475 7 1 2 70072 474
0 476 5 1 1 475
0 477 7 1 2 57285 476
0 478 5 1 1 477
0 479 7 1 2 470 478
0 480 5 1 1 479
0 481 7 1 2 60710 480
0 482 5 1 1 481
0 483 7 13 2 64917 68717
0 484 5 9 1 70074
0 485 7 1 2 69727 70075
0 486 5 1 1 485
0 487 7 1 2 69719 486
0 488 5 1 1 487
0 489 7 8 2 65115 67623
0 490 5 14 1 70096
0 491 7 5 2 59195 68292
0 492 5 4 1 70118
0 493 7 1 2 70104 70123
0 494 5 3 1 493
0 495 7 1 2 488 70127
0 496 5 1 1 495
0 497 7 1 2 482 496
0 498 7 1 2 466 497
0 499 5 1 1 498
0 500 7 1 2 69591 499
0 501 5 1 1 500
0 502 7 1 2 440 501
0 503 5 1 1 502
0 504 7 1 2 61882 503
0 505 5 1 1 504
0 506 7 48 2 59196 65370
0 507 5 58 1 70130
0 508 7 2 2 58110 70131
0 509 5 5 1 70236
0 510 7 5 2 62826 70178
0 511 5 17 1 70243
0 512 7 3 2 57831 70248
0 513 5 1 1 70265
0 514 7 1 2 67003 70266
0 515 5 1 1 514
0 516 7 1 2 70238 515
0 517 5 1 1 516
0 518 7 1 2 64125 517
0 519 5 1 1 518
0 520 7 43 2 60437 60711
0 521 5 26 1 70268
0 522 7 2 2 58111 70269
0 523 5 1 1 70337
0 524 7 17 2 57556 65371
0 525 5 4 1 70339
0 526 7 5 2 65116 70340
0 527 5 1 1 70360
0 528 7 1 2 64126 70361
0 529 5 1 1 528
0 530 7 1 2 523 529
0 531 5 1 1 530
0 532 7 1 2 67240 531
0 533 5 1 1 532
0 534 7 14 2 62827 68065
0 535 5 62 1 70365
0 536 7 3 2 64127 70379
0 537 7 2 2 60712 67018
0 538 5 2 1 70444
0 539 7 1 2 70441 70446
0 540 5 1 1 539
0 541 7 1 2 533 540
0 542 5 1 1 541
0 543 7 1 2 69125 542
0 544 5 1 1 543
0 545 7 1 2 519 544
0 546 5 1 1 545
0 547 7 12 2 58831 64766
0 548 5 1 1 70448
0 549 7 4 2 63568 60094
0 550 5 1 1 70460
0 551 7 2 2 548 550
0 552 5 79 1 70464
0 553 7 5 2 62019 70466
0 554 7 12 2 66540 70545
0 555 7 1 2 546 70550
0 556 5 1 1 555
0 557 7 21 2 66541 70467
0 558 7 9 2 57557 68549
0 559 5 60 1 70583
0 560 7 8 2 58112 63931
0 561 5 3 1 70652
0 562 7 15 2 60438 65372
0 563 5 4 1 70663
0 564 7 8 2 63796 59197
0 565 7 1 2 70664 70682
0 566 5 3 1 565
0 567 7 1 2 70660 70690
0 568 5 1 1 567
0 569 7 1 2 70592 568
0 570 5 1 1 569
0 571 7 10 2 57832 59052
0 572 5 7 1 70693
0 573 7 3 2 58113 70179
0 574 5 2 1 70710
0 575 7 1 2 70703 70711
0 576 5 1 1 575
0 577 7 8 2 57833 64918
0 578 5 3 1 70715
0 579 7 2 2 70716 69105
0 580 7 1 2 70270 70726
0 581 5 1 1 580
0 582 7 1 2 576 581
0 583 7 1 2 570 582
0 584 5 1 1 583
0 585 7 1 2 70562 584
0 586 5 1 1 585
0 587 7 1 2 62545 69405
0 588 5 3 1 587
0 589 7 10 2 62546 69913
0 590 5 1 1 70731
0 591 7 2 2 67556 68446
0 592 5 1 1 70741
0 593 7 1 2 70732 70742
0 594 5 4 1 593
0 595 7 55 2 59053 65117
0 596 5 55 1 70747
0 597 7 1 2 70748 70584
0 598 5 2 1 597
0 599 7 2 2 60210 70857
0 600 5 1 1 70859
0 601 7 1 2 70743 70860
0 602 5 1 1 601
0 603 7 2 2 65373 602
0 604 7 1 2 70728 70861
0 605 5 1 1 604
0 606 7 18 2 57286 64919
0 607 5 4 1 70863
0 608 7 1 2 60439 70881
0 609 5 3 1 608
0 610 7 3 2 58928 70885
0 611 5 2 1 70888
0 612 7 1 2 67127 67019
0 613 7 1 2 70891 612
0 614 5 1 1 613
0 615 7 1 2 59054 614
0 616 5 1 1 615
0 617 7 1 2 62547 67603
0 618 5 1 1 617
0 619 7 1 2 65118 618
0 620 5 1 1 619
0 621 7 3 2 62548 63736
0 622 5 2 1 70893
0 623 7 1 2 59198 70896
0 624 5 1 1 623
0 625 7 11 2 62828 60713
0 626 5 5 1 70898
0 627 7 17 2 62146 62287
0 628 5 10 1 70914
0 629 7 1 2 67241 70931
0 630 5 3 1 629
0 631 7 1 2 70899 70941
0 632 7 1 2 624 631
0 633 7 1 2 620 632
0 634 7 1 2 616 633
0 635 5 1 1 634
0 636 7 1 2 605 635
0 637 5 1 1 636
0 638 7 1 2 69862 637
0 639 5 1 1 638
0 640 7 1 2 67613 639
0 641 5 1 1 640
0 642 7 1 2 586 641
0 643 5 1 1 642
0 644 7 1 2 62020 643
0 645 5 1 1 644
0 646 7 10 2 63797 67557
0 647 5 21 1 70944
0 648 7 2 2 70954 68550
0 649 5 2 1 70975
0 650 7 2 2 59199 67572
0 651 5 5 1 70979
0 652 7 1 2 65374 70981
0 653 7 2 2 70977 652
0 654 7 1 2 62549 70986
0 655 5 2 1 654
0 656 7 1 2 62288 70683
0 657 5 2 1 656
0 658 7 3 2 63932 68293
0 659 7 1 2 68447 67708
0 660 5 4 1 659
0 661 7 1 2 70992 70995
0 662 5 2 1 661
0 663 7 9 2 60211 70593
0 664 5 2 1 71001
0 665 7 1 2 59200 71002
0 666 5 1 1 665
0 667 7 2 2 70999 666
0 668 5 1 1 71012
0 669 7 1 2 70990 71013
0 670 5 1 1 669
0 671 7 1 2 60440 670
0 672 5 2 1 671
0 673 7 2 2 62550 70749
0 674 5 2 1 71016
0 675 7 13 2 62289 68448
0 676 5 10 1 71020
0 677 7 2 2 65119 71033
0 678 5 1 1 71043
0 679 7 1 2 62551 678
0 680 5 3 1 679
0 681 7 1 2 63798 71045
0 682 5 1 1 681
0 683 7 1 2 71018 682
0 684 5 1 1 683
0 685 7 1 2 63933 684
0 686 5 2 1 685
0 687 7 1 2 71014 71048
0 688 5 1 1 687
0 689 7 1 2 60714 688
0 690 5 1 1 689
0 691 7 1 2 70988 690
0 692 5 1 1 691
0 693 7 13 2 58114 63569
0 694 7 5 2 64767 61883
0 695 7 19 2 66657 71063
0 696 7 2 2 71050 71068
0 697 7 1 2 692 71087
0 698 5 1 1 697
0 699 7 3 2 62552 70132
0 700 5 3 1 71089
0 701 7 1 2 69720 71092
0 702 5 2 1 701
0 703 7 1 2 70594 70551
0 704 5 1 1 703
0 705 7 3 2 64768 65120
0 706 7 5 2 67500 71097
0 707 7 2 2 64920 71100
0 708 7 6 2 62290 68196
0 709 5 4 1 71107
0 710 7 2 2 63570 63737
0 711 7 1 2 71108 71117
0 712 7 1 2 71105 711
0 713 5 1 1 712
0 714 7 1 2 704 713
0 715 5 1 1 714
0 716 7 1 2 71095 715
0 717 5 1 1 716
0 718 7 1 2 698 717
0 719 7 1 2 645 718
0 720 5 1 1 719
0 721 7 1 2 59399 720
0 722 5 1 1 721
0 723 7 1 2 556 722
0 724 7 1 2 505 723
0 725 5 1 1 724
0 726 7 1 2 58377 725
0 727 5 1 1 726
0 728 7 6 2 57834 63128
0 729 7 3 2 57558 68909
0 730 7 2 2 68914 69169
0 731 7 6 2 59400 60095
0 732 7 1 2 71128 71130
0 733 7 2 2 71125 732
0 734 7 1 2 71119 71136
0 735 5 1 1 734
0 736 7 1 2 727 735
0 737 7 1 2 285 736
0 738 5 1 1 737
0 739 7 1 2 59710 738
0 740 5 1 1 739
0 741 7 100 2 58115 59401
0 742 5 104 1 71138
0 743 7 1 2 64433 68209
0 744 5 1 1 743
0 745 7 1 2 68714 744
0 746 5 1 1 745
0 747 7 1 2 65375 746
0 748 5 1 1 747
0 749 7 4 2 58929 68951
0 750 5 1 1 71342
0 751 7 7 2 64434 64769
0 752 7 13 2 64921 66542
0 753 7 1 2 71346 71353
0 754 7 1 2 71343 753
0 755 5 1 1 754
0 756 7 1 2 69102 755
0 757 5 1 1 756
0 758 7 1 2 58832 757
0 759 5 1 1 758
0 760 7 3 2 68952 69143
0 761 7 9 2 64435 60096
0 762 7 2 2 71354 71369
0 763 7 1 2 71366 71378
0 764 5 1 1 763
0 765 7 1 2 759 764
0 766 5 1 1 765
0 767 7 1 2 57835 766
0 768 5 1 1 767
0 769 7 1 2 68948 768
0 770 5 1 1 769
0 771 7 1 2 69151 770
0 772 5 1 1 771
0 773 7 1 2 748 772
0 774 5 1 1 773
0 775 7 1 2 71139 774
0 776 5 1 1 775
0 777 7 77 2 62829 64128
0 778 5 115 1 71380
0 779 7 3 2 64922 71457
0 780 5 1 1 71572
0 781 7 1 2 71573 71370
0 782 7 1 2 69208 781
0 783 5 1 1 782
0 784 7 1 2 776 783
0 785 5 1 1 784
0 786 7 1 2 58378 785
0 787 5 1 1 786
0 788 7 1 2 740 787
0 789 5 1 1 788
0 790 7 1 2 65760 789
0 791 5 1 1 790
0 792 7 17 2 57836 58116
0 793 5 10 1 71575
0 794 7 1 2 71576 71137
0 795 5 1 1 794
0 796 7 6 2 59055 60715
0 797 5 1 1 71602
0 798 7 3 2 57559 71603
0 799 5 1 1 71608
0 800 7 6 2 60441 68814
0 801 5 13 1 71611
0 802 7 4 2 68551 71617
0 803 7 1 2 71609 71630
0 804 5 2 1 803
0 805 7 4 2 58930 68294
0 806 5 4 1 71636
0 807 7 6 2 57287 68295
0 808 5 2 1 71644
0 809 7 5 2 71640 71650
0 810 5 3 1 71652
0 811 7 7 2 67709 71653
0 812 5 2 1 71660
0 813 7 1 2 60212 71667
0 814 5 1 1 813
0 815 7 32 2 63738 60213
0 816 5 67 1 71669
0 817 7 5 2 71670 70915
0 818 5 5 1 71768
0 819 7 8 2 65121 67710
0 820 7 1 2 71773 71778
0 821 5 1 1 820
0 822 7 1 2 814 821
0 823 5 1 1 822
0 824 7 1 2 65376 823
0 825 5 1 1 824
0 826 7 1 2 71634 825
0 827 5 1 1 826
0 828 7 1 2 71069 827
0 829 5 1 1 828
0 830 7 53 2 63799 60442
0 831 5 98 1 71786
0 832 7 2 2 62147 71787
0 833 5 2 1 71937
0 834 7 1 2 57560 71939
0 835 5 2 1 834
0 836 7 1 2 60716 71941
0 837 5 1 1 836
0 838 7 13 2 66543 69326
0 839 7 1 2 837 71943
0 840 5 1 1 839
0 841 7 1 2 829 840
0 842 5 1 1 841
0 843 7 1 2 63571 842
0 844 5 1 1 843
0 845 7 6 2 64770 60717
0 846 7 1 2 71956 71942
0 847 5 1 1 846
0 848 7 1 2 67081 59
0 849 5 6 1 848
0 850 7 1 2 68659 71962
0 851 7 1 2 847 850
0 852 5 1 1 851
0 853 7 1 2 844 852
0 854 5 1 1 853
0 855 7 1 2 58117 854
0 856 5 1 1 855
0 857 7 3 2 70750 70341
0 858 5 4 1 71968
0 859 7 1 2 69993 69865
0 860 5 2 1 859
0 861 7 1 2 67020 71975
0 862 5 1 1 861
0 863 7 1 2 60718 69122
0 864 5 4 1 863
0 865 7 1 2 57288 71977
0 866 7 1 2 862 865
0 867 5 1 1 866
0 868 7 1 2 71971 867
0 869 5 1 1 868
0 870 7 1 2 67963 869
0 871 5 1 1 870
0 872 7 1 2 856 871
0 873 5 1 1 872
0 874 7 1 2 59201 873
0 875 5 1 1 874
0 876 7 1 2 69492 71978
0 877 5 1 1 876
0 878 7 22 2 60214 65377
0 879 5 1 1 71981
0 880 7 5 2 59202 70751
0 881 5 2 1 72003
0 882 7 1 2 71982 72004
0 883 5 1 1 882
0 884 7 28 2 64923 65378
0 885 5 13 1 72010
0 886 7 1 2 58118 72038
0 887 7 1 2 71979 886
0 888 5 1 1 887
0 889 7 1 2 883 888
0 890 5 1 1 889
0 891 7 1 2 69252 890
0 892 5 1 1 891
0 893 7 1 2 877 892
0 894 5 1 1 893
0 895 7 1 2 57561 894
0 896 5 1 1 895
0 897 7 12 2 65379 71839
0 898 5 39 1 72051
0 899 7 8 2 64771 60215
0 900 7 3 2 66658 72102
0 901 7 3 2 71051 72110
0 902 5 1 1 72113
0 903 7 1 2 72052 72114
0 904 5 1 1 903
0 905 7 6 2 67906 69153
0 906 5 6 1 72116
0 907 7 29 2 65122 60719
0 908 5 4 1 72128
0 909 7 11 2 69230 71052
0 910 5 1 1 72161
0 911 7 1 2 72129 72162
0 912 5 1 1 911
0 913 7 1 2 72122 912
0 914 5 1 1 913
0 915 7 1 2 69093 914
0 916 5 1 1 915
0 917 7 1 2 904 916
0 918 7 1 2 896 917
0 919 5 1 1 918
0 920 7 1 2 57289 919
0 921 5 1 1 920
0 922 7 5 2 58833 59203
0 923 7 3 2 69327 72172
0 924 5 6 1 72177
0 925 7 10 2 62291 63739
0 926 5 10 1 72186
0 927 7 1 2 72196 72115
0 928 5 1 1 927
0 929 7 1 2 72180 928
0 930 5 1 1 929
0 931 7 1 2 71840 930
0 932 5 1 1 931
0 933 7 1 2 59056 69949
0 934 5 2 1 933
0 935 7 1 2 62830 72206
0 936 5 6 1 935
0 937 7 2 2 57562 72208
0 938 5 3 1 72214
0 939 7 2 2 69318 69253
0 940 7 1 2 72215 72219
0 941 5 1 1 940
0 942 7 5 2 63934 70802
0 943 5 30 1 72221
0 944 7 5 2 57563 58834
0 945 7 1 2 69328 72256
0 946 5 5 1 945
0 947 7 1 2 72261 902
0 948 5 1 1 947
0 949 7 1 2 72226 948
0 950 5 1 1 949
0 951 7 1 2 941 950
0 952 7 1 2 932 951
0 953 5 1 1 952
0 954 7 1 2 65380 953
0 955 5 1 1 954
0 956 7 4 2 68815 68211
0 957 5 8 1 72266
0 958 7 11 2 59204 60720
0 959 5 6 1 72278
0 960 7 2 2 64924 70665
0 961 5 1 1 72295
0 962 7 1 2 72289 961
0 963 5 2 1 962
0 964 7 1 2 72163 72297
0 965 5 2 1 964
0 966 7 1 2 69950 68671
0 967 5 1 1 966
0 968 7 1 2 72299 967
0 969 5 1 1 968
0 970 7 1 2 72270 969
0 971 5 1 1 970
0 972 7 2 2 69951 69144
0 973 7 12 2 60721 66659
0 974 7 5 2 64772 72303
0 975 7 1 2 72301 72315
0 976 5 1 1 975
0 977 7 1 2 68692 976
0 978 5 1 1 977
0 979 7 1 2 58119 978
0 980 5 1 1 979
0 981 7 2 2 58835 69106
0 982 7 2 2 64925 62021
0 983 7 5 2 59205 60097
0 984 7 1 2 72322 72324
0 985 7 1 2 72320 984
0 986 5 1 1 985
0 987 7 1 2 980 986
0 988 7 1 2 971 987
0 989 7 1 2 955 988
0 990 7 1 2 921 989
0 991 5 1 1 990
0 992 7 1 2 61884 991
0 993 5 1 1 992
0 994 7 14 2 62148 60443
0 995 5 18 1 72329
0 996 7 3 2 57564 72343
0 997 5 2 1 72361
0 998 7 1 2 60722 72364
0 999 5 2 1 998
0 1000 7 1 2 69906 72366
0 1001 5 1 1 1000
0 1002 7 2 2 58120 67867
0 1003 5 2 1 72368
0 1004 7 9 2 64926 67624
0 1005 7 16 2 58931 65123
0 1006 5 10 1 72381
0 1007 7 8 2 65381 72382
0 1008 7 2 2 72372 72407
0 1009 5 1 1 72415
0 1010 7 1 2 72370 1009
0 1011 7 1 2 1001 1010
0 1012 5 1 1 1011
0 1013 7 1 2 70552 1012
0 1014 5 1 1 1013
0 1015 7 1 2 993 1014
0 1016 5 1 1 1015
0 1017 7 1 2 57837 1016
0 1018 5 1 1 1017
0 1019 7 1 2 875 1018
0 1020 5 1 1 1019
0 1021 7 1 2 59402 1020
0 1022 5 1 1 1021
0 1023 7 6 2 58121 62022
0 1024 7 1 2 65382 68204
0 1025 5 2 1 1024
0 1026 7 1 2 68905 72423
0 1027 5 1 1 1026
0 1028 7 1 2 67034 1027
0 1029 5 1 1 1028
0 1030 7 6 2 64773 65383
0 1031 7 1 2 69133 72425
0 1032 5 1 1 1031
0 1033 7 1 2 1029 1032
0 1034 5 1 1 1033
0 1035 7 1 2 58836 1034
0 1036 5 1 1 1035
0 1037 7 3 2 63572 69107
0 1038 7 11 2 60098 65384
0 1039 7 1 2 71355 72434
0 1040 7 1 2 72431 1039
0 1041 5 1 1 1040
0 1042 7 1 2 1036 1041
0 1043 5 1 1 1042
0 1044 7 1 2 67004 1043
0 1045 5 1 1 1044
0 1046 7 8 2 64927 61885
0 1047 7 2 2 72435 72445
0 1048 7 1 2 68910 72453
0 1049 5 1 1 1048
0 1050 7 1 2 1045 1049
0 1051 5 1 1 1050
0 1052 7 1 2 67242 1051
0 1053 5 1 1 1052
0 1054 7 33 2 65124 65385
0 1055 5 11 1 72455
0 1056 7 5 2 60099 72446
0 1057 5 3 1 72499
0 1058 7 1 2 72456 72500
0 1059 7 1 2 71126 1058
0 1060 5 1 1 1059
0 1061 7 1 2 1053 1060
0 1062 5 1 1 1061
0 1063 7 1 2 72417 1062
0 1064 5 1 1 1063
0 1065 7 9 2 64129 68066
0 1066 5 12 1 72507
0 1067 7 5 2 57290 60444
0 1068 7 2 2 68971 72528
0 1069 5 3 1 72533
0 1070 7 8 2 65125 68552
0 1071 5 13 1 72538
0 1072 7 1 2 60216 72539
0 1073 5 1 1 1072
0 1074 7 1 2 72535 1073
0 1075 5 1 1 1074
0 1076 7 8 2 63573 66660
0 1077 7 5 2 71064 72559
0 1078 7 2 2 65386 72567
0 1079 7 1 2 1075 72572
0 1080 5 1 1 1079
0 1081 7 1 2 68972 72344
0 1082 7 1 2 70553 1081
0 1083 5 1 1 1082
0 1084 7 1 2 1080 1083
0 1085 5 1 1 1084
0 1086 7 1 2 57565 1085
0 1087 5 1 1 1086
0 1088 7 12 2 65387 66544
0 1089 7 4 2 70468 72574
0 1090 5 2 1 72586
0 1091 7 1 2 127 72590
0 1092 5 1 1 1091
0 1093 7 1 2 68973 1092
0 1094 5 1 1 1093
0 1095 7 17 2 61886 67907
0 1096 7 1 2 70311 72592
0 1097 5 1 1 1096
0 1098 7 1 2 1094 1097
0 1099 5 1 1 1098
0 1100 7 1 2 62023 1099
0 1101 5 1 1 1100
0 1102 7 1 2 1087 1101
0 1103 5 1 1 1102
0 1104 7 1 2 59057 1103
0 1105 5 1 1 1104
0 1106 7 3 2 63574 65388
0 1107 7 2 2 67433 72609
0 1108 7 1 2 67005 72612
0 1109 5 1 1 1108
0 1110 7 2 2 60723 72397
0 1111 5 3 1 72614
0 1112 7 2 2 57291 72616
0 1113 5 3 1 72619
0 1114 7 1 2 65389 67573
0 1115 5 5 1 1114
0 1116 7 1 2 67021 72624
0 1117 7 1 2 72621 1116
0 1118 5 1 1 1117
0 1119 7 1 2 67035 1118
0 1120 5 1 1 1119
0 1121 7 4 2 64774 72575
0 1122 5 1 1 72629
0 1123 7 1 2 67006 72630
0 1124 5 1 1 1123
0 1125 7 1 2 1120 1124
0 1126 5 1 1 1125
0 1127 7 1 2 58837 1126
0 1128 5 1 1 1127
0 1129 7 1 2 1109 1128
0 1130 5 1 1 1129
0 1131 7 1 2 62024 1130
0 1132 5 1 1 1131
0 1133 7 1 2 1105 1132
0 1134 5 1 1 1133
0 1135 7 1 2 58122 1134
0 1136 5 1 1 1135
0 1137 7 3 2 57566 72011
0 1138 5 1 1 72633
0 1139 7 4 2 60100 65126
0 1140 7 2 2 67949 72636
0 1141 7 1 2 72634 72640
0 1142 7 1 2 68911 1141
0 1143 5 1 1 1142
0 1144 7 1 2 1136 1143
0 1145 5 1 1 1144
0 1146 7 1 2 72516 1145
0 1147 5 1 1 1146
0 1148 7 1 2 1064 1147
0 1149 7 1 2 1022 1148
0 1150 5 1 1 1149
0 1151 7 1 2 59711 1150
0 1152 5 1 1 1151
0 1153 7 1 2 795 1152
0 1154 5 1 1 1153
0 1155 7 1 2 58379 1154
0 1156 5 1 1 1155
0 1157 7 3 2 72457 71070
0 1158 7 17 2 58380 59403
0 1159 5 4 1 72645
0 1160 7 5 2 59206 59712
0 1161 7 2 2 72646 72666
0 1162 7 7 2 58123 64928
0 1163 5 2 1 72673
0 1164 7 1 2 63575 72674
0 1165 7 1 2 72671 1164
0 1166 7 1 2 72642 1165
0 1167 5 1 1 1166
0 1168 7 9 2 67450 67908
0 1169 7 1 2 70595 72682
0 1170 5 1 1 1169
0 1171 7 5 2 70469 67501
0 1172 7 1 2 71769 72691
0 1173 5 1 1 1172
0 1174 7 1 2 1170 1173
0 1175 5 1 1 1174
0 1176 7 1 2 72063 1175
0 1177 5 1 1 1176
0 1178 7 16 2 57567 64929
0 1179 5 19 1 72696
0 1180 7 20 2 61887 70470
0 1181 5 2 1 72731
0 1182 7 1 2 72712 72732
0 1183 5 1 1 1182
0 1184 7 4 2 63576 66957
0 1185 7 1 2 71021 72753
0 1186 5 1 1 1185
0 1187 7 1 2 1183 1186
0 1188 5 1 1 1187
0 1189 7 10 2 60724 71788
0 1190 5 3 1 72757
0 1191 7 1 2 66661 72758
0 1192 7 1 2 1188 1191
0 1193 5 1 1 1192
0 1194 7 1 2 1177 1193
0 1195 5 1 1 1194
0 1196 7 14 2 62831 63935
0 1197 5 4 1 72770
0 1198 7 15 2 63129 64130
0 1199 5 6 1 72788
0 1200 7 2 2 72771 72789
0 1201 7 1 2 64436 72809
0 1202 7 1 2 1195 1201
0 1203 5 1 1 1202
0 1204 7 1 2 1167 1203
0 1205 5 1 1 1204
0 1206 7 1 2 62553 1205
0 1207 5 1 1 1206
0 1208 7 14 2 57292 57838
0 1209 5 1 1 72811
0 1210 7 8 2 57568 58124
0 1211 5 1 1 72825
0 1212 7 3 2 72812 72826
0 1213 7 3 2 69108 72833
0 1214 7 2 2 72173 72836
0 1215 7 9 2 59713 64930
0 1216 7 1 2 72841 71131
0 1217 7 1 2 69170 1216
0 1218 7 1 2 72839 1217
0 1219 5 1 1 1218
0 1220 7 1 2 1207 1219
0 1221 7 1 2 1156 1220
0 1222 5 1 1 1221
0 1223 7 1 2 61137 1222
0 1224 5 1 1 1223
0 1225 7 36 2 64131 61138
0 1226 5 40 1 72850
0 1227 7 3 2 61139 70180
0 1228 5 9 1 72926
0 1229 7 6 2 64132 70181
0 1230 5 5 1 72938
0 1231 7 2 2 72929 72944
0 1232 7 3 2 72886 72949
0 1233 5 1 1 72951
0 1234 7 2 2 65761 70312
0 1235 5 8 1 72954
0 1236 7 1 2 59404 72955
0 1237 5 1 1 1236
0 1238 7 2 2 72952 1237
0 1239 7 1 2 70563 72964
0 1240 5 1 1 1239
0 1241 7 12 2 61140 61888
0 1242 7 15 2 59207 59405
0 1243 5 1 1 72978
0 1244 7 1 2 72979 67909
0 1245 7 1 2 72966 1244
0 1246 5 1 1 1245
0 1247 7 1 2 1240 1246
0 1248 5 1 1 1247
0 1249 7 1 2 68296 1248
0 1250 5 1 1 1249
0 1251 7 28 2 64133 65762
0 1252 5 8 1 72993
0 1253 7 1 2 70133 72994
0 1254 5 2 1 1253
0 1255 7 27 2 59406 61141
0 1256 5 16 1 73031
0 1257 7 3 2 73021 73058
0 1258 5 22 1 73074
0 1259 7 38 2 63936 60725
0 1260 5 47 1 73099
0 1261 7 2 2 67625 73137
0 1262 5 1 1 73184
0 1263 7 1 2 73077 73185
0 1264 5 1 1 1263
0 1265 7 1 2 73029 1264
0 1266 5 1 1 1265
0 1267 7 1 2 70471 67106
0 1268 7 1 2 1266 1267
0 1269 5 1 1 1268
0 1270 7 1 2 1250 1269
0 1271 5 1 1 1270
0 1272 7 1 2 57839 1271
0 1273 5 1 1 1272
0 1274 7 2 2 70752 70564
0 1275 5 1 1 73186
0 1276 7 4 2 65763 69305
0 1277 5 1 1 73188
0 1278 7 1 2 70342 73189
0 1279 7 1 2 73187 1278
0 1280 5 1 1 1279
0 1281 7 1 2 1273 1280
0 1282 5 1 1 1281
0 1283 7 1 2 57293 1282
0 1284 5 1 1 1283
0 1285 7 6 2 57840 61142
0 1286 7 2 2 72980 73192
0 1287 5 1 1 73198
0 1288 7 12 2 65127 68297
0 1289 5 10 1 73200
0 1290 7 1 2 73201 73078
0 1291 5 1 1 1290
0 1292 7 9 2 59058 59407
0 1293 5 1 1 73222
0 1294 7 4 2 57569 73223
0 1295 7 1 2 61143 73231
0 1296 5 1 1 1295
0 1297 7 1 2 1291 1296
0 1298 5 1 1 1297
0 1299 7 1 2 67243 1298
0 1300 5 1 1 1299
0 1301 7 1 2 1287 1300
0 1302 5 1 1 1301
0 1303 7 1 2 65390 1302
0 1304 5 1 1 1303
0 1305 7 38 2 60726 65764
0 1306 5 3 1 73235
0 1307 7 1 2 64134 72008
0 1308 5 3 1 1307
0 1309 7 1 2 57841 73276
0 1310 5 2 1 1309
0 1311 7 4 2 57570 71841
0 1312 5 12 1 73281
0 1313 7 1 2 73282 72517
0 1314 5 1 1 1313
0 1315 7 1 2 73279 1314
0 1316 5 1 1 1315
0 1317 7 1 2 73236 1316
0 1318 5 1 1 1317
0 1319 7 1 2 1304 1318
0 1320 5 1 1 1319
0 1321 7 1 2 72593 1320
0 1322 5 1 1 1321
0 1323 7 1 2 1284 1322
0 1324 5 1 1 1323
0 1325 7 1 2 62025 1324
0 1326 5 1 1 1325
0 1327 7 31 2 65391 65765
0 1328 5 8 1 73297
0 1329 7 3 2 64135 73298
0 1330 5 4 1 73336
0 1331 7 2 2 73337 71101
0 1332 7 5 2 57571 62832
0 1333 7 2 2 67439 73345
0 1334 7 1 2 68953 73350
0 1335 7 1 2 73343 1334
0 1336 5 1 1 1335
0 1337 7 1 2 1326 1336
0 1338 5 1 1 1337
0 1339 7 1 2 59714 1338
0 1340 5 1 1 1339
0 1341 7 7 2 63577 59059
0 1342 7 11 2 64437 61144
0 1343 5 2 1 73359
0 1344 7 19 2 59715 65392
0 1345 5 3 1 73372
0 1346 7 16 2 57842 65128
0 1347 5 5 1 73394
0 1348 7 1 2 73391 73395
0 1349 7 1 2 73370 1348
0 1350 7 3 2 65766 70182
0 1351 5 1 1 73415
0 1352 7 7 2 59408 64775
0 1353 7 2 2 67502 73418
0 1354 7 1 2 1351 73425
0 1355 7 2 2 1349 1354
0 1356 7 1 2 73352 73427
0 1357 5 1 1 1356
0 1358 7 5 2 59060 72458
0 1359 5 7 1 73429
0 1360 7 1 2 61145 73434
0 1361 5 7 1 1360
0 1362 7 2 2 72956 73441
0 1363 7 1 2 59208 73448
0 1364 5 1 1 1363
0 1365 7 7 2 60727 70803
0 1366 5 22 1 73450
0 1367 7 1 2 73457 73079
0 1368 5 1 1 1367
0 1369 7 1 2 1364 1368
0 1370 5 1 1 1369
0 1371 7 1 2 59716 1370
0 1372 5 1 1 1371
0 1373 7 5 2 72227 73458
0 1374 7 8 2 73138 73479
0 1375 5 1 1 73484
0 1376 7 12 2 59717 61146
0 1377 5 3 1 73492
0 1378 7 14 2 64438 65767
0 1379 5 3 1 73507
0 1380 7 1 2 59409 73508
0 1381 5 2 1 1380
0 1382 7 1 2 73504 73524
0 1383 5 2 1 1382
0 1384 7 1 2 73485 73526
0 1385 5 1 1 1384
0 1386 7 7 2 65768 70271
0 1387 7 1 2 59718 73528
0 1388 5 1 1 1387
0 1389 7 1 2 1385 1388
0 1390 5 1 1 1389
0 1391 7 1 2 57843 1390
0 1392 5 1 1 1391
0 1393 7 3 2 59061 72981
0 1394 7 18 2 64439 65393
0 1395 5 1 1 73538
0 1396 7 14 2 65129 65769
0 1397 5 5 1 73556
0 1398 7 2 2 73539 73557
0 1399 7 1 2 73535 73575
0 1400 5 1 1 1399
0 1401 7 1 2 1392 1400
0 1402 7 1 2 1372 1401
0 1403 5 1 1 1402
0 1404 7 1 2 57294 1403
0 1405 5 1 1 1404
0 1406 7 5 2 59410 67244
0 1407 5 18 1 73577
0 1408 7 1 2 73578 73493
0 1409 5 1 1 1408
0 1410 7 1 2 1405 1409
0 1411 5 1 1 1410
0 1412 7 1 2 70565 1411
0 1413 5 1 1 1412
0 1414 7 1 2 57295 73032
0 1415 5 3 1 1414
0 1416 7 33 2 65394 61147
0 1417 5 4 1 73603
0 1418 7 1 2 59209 73604
0 1419 5 2 1 1418
0 1420 7 1 2 73273 73640
0 1421 5 3 1 1420
0 1422 7 1 2 71842 73642
0 1423 5 1 1 1422
0 1424 7 1 2 73600 1423
0 1425 5 1 1 1424
0 1426 7 1 2 59719 1425
0 1427 5 1 1 1426
0 1428 7 40 2 59411 65770
0 1429 5 20 1 73645
0 1430 7 1 2 73646 72279
0 1431 5 1 1 1430
0 1432 7 1 2 61148 73373
0 1433 5 1 1 1432
0 1434 7 1 2 1431 1433
0 1435 5 2 1 1434
0 1436 7 1 2 71843 73705
0 1437 5 1 1 1436
0 1438 7 24 2 59412 64440
0 1439 5 2 1 73707
0 1440 7 5 2 65771 72459
0 1441 7 1 2 73708 73733
0 1442 5 2 1 1441
0 1443 7 6 2 57296 59210
0 1444 7 1 2 73494 73740
0 1445 5 1 1 1444
0 1446 7 1 2 73738 1445
0 1447 7 1 2 1437 1446
0 1448 5 1 1 1447
0 1449 7 1 2 57844 1448
0 1450 5 1 1 1449
0 1451 7 2 2 72982 73576
0 1452 5 1 1 73746
0 1453 7 1 2 1450 1452
0 1454 7 1 2 1427 1453
0 1455 5 1 1 1454
0 1456 7 1 2 72594 1455
0 1457 5 1 1 1456
0 1458 7 1 2 1413 1457
0 1459 5 1 1 1458
0 1460 7 1 2 62026 1459
0 1461 5 1 1 1460
0 1462 7 1 2 1357 1461
0 1463 5 1 1 1462
0 1464 7 1 2 57572 1463
0 1465 5 1 1 1464
0 1466 7 2 2 59413 72460
0 1467 5 1 1 73748
0 1468 7 18 2 59414 65130
0 1469 5 3 1 73750
0 1470 7 1 2 57845 72053
0 1471 5 1 1 1470
0 1472 7 1 2 73768 1471
0 1473 5 1 1 1472
0 1474 7 1 2 59211 1473
0 1475 5 1 1 1474
0 1476 7 1 2 1467 1475
0 1477 5 1 1 1476
0 1478 7 1 2 61149 1477
0 1479 5 1 1 1478
0 1480 7 14 2 60445 65772
0 1481 7 2 2 73771 71604
0 1482 5 2 1 73785
0 1483 7 1 2 67245 73786
0 1484 5 1 1 1483
0 1485 7 8 2 59062 65395
0 1486 5 5 1 73789
0 1487 7 1 2 73797 73410
0 1488 5 2 1 1487
0 1489 7 1 2 73080 73802
0 1490 5 1 1 1489
0 1491 7 1 2 1484 1490
0 1492 7 1 2 1479 1491
0 1493 5 1 1 1492
0 1494 7 1 2 59720 1493
0 1495 5 1 1 1494
0 1496 7 4 2 65773 67975
0 1497 5 2 1 73804
0 1498 7 2 2 59415 71844
0 1499 5 4 1 73810
0 1500 7 1 2 73540 73811
0 1501 7 1 2 73805 1500
0 1502 5 1 1 1501
0 1503 7 1 2 1495 1502
0 1504 5 1 1 1503
0 1505 7 1 2 57297 1504
0 1506 5 1 1 1505
0 1507 7 5 2 59063 67246
0 1508 5 4 1 73816
0 1509 7 21 2 59416 59721
0 1510 7 2 2 61150 73825
0 1511 7 1 2 73817 73846
0 1512 5 1 1 1511
0 1513 7 1 2 1506 1512
0 1514 5 1 1 1513
0 1515 7 1 2 70566 1514
0 1516 5 1 1 1515
0 1517 7 12 2 57298 59064
0 1518 5 3 1 73848
0 1519 7 1 2 60728 73860
0 1520 5 2 1 1519
0 1521 7 1 2 72518 73863
0 1522 5 1 1 1521
0 1523 7 17 2 65396 67247
0 1524 5 7 1 73865
0 1525 7 1 2 70753 73866
0 1526 5 1 1 1525
0 1527 7 1 2 1522 1526
0 1528 5 1 1 1527
0 1529 7 1 2 61151 1528
0 1530 5 1 1 1529
0 1531 7 3 2 62554 70804
0 1532 5 10 1 73889
0 1533 7 1 2 63937 73890
0 1534 5 13 1 1533
0 1535 7 1 2 73237 73902
0 1536 5 1 1 1535
0 1537 7 1 2 1530 1536
0 1538 5 1 1 1537
0 1539 7 1 2 59722 1538
0 1540 5 1 1 1539
0 1541 7 5 2 60729 68067
0 1542 5 7 1 73915
0 1543 7 21 2 67248 73920
0 1544 5 1 1 73927
0 1545 7 8 2 59065 65774
0 1546 5 3 1 73948
0 1547 7 1 2 73392 73949
0 1548 7 1 2 73751 1547
0 1549 7 1 2 73928 1548
0 1550 5 1 1 1549
0 1551 7 1 2 1540 1550
0 1552 5 1 1 1551
0 1553 7 1 2 72595 1552
0 1554 5 1 1 1553
0 1555 7 1 2 1516 1554
0 1556 5 1 1 1555
0 1557 7 1 2 62027 1556
0 1558 5 1 1 1557
0 1559 7 1 2 1465 1558
0 1560 5 1 1 1559
0 1561 7 1 2 58125 1560
0 1562 5 1 1 1561
0 1563 7 1 2 1340 1562
0 1564 5 1 1 1563
0 1565 7 1 2 58381 1564
0 1566 5 1 1 1565
0 1567 7 13 2 58126 59723
0 1568 5 1 1 73959
0 1569 7 2 2 73647 73960
0 1570 7 1 2 72257 68938
0 1571 5 1 1 1570
0 1572 7 10 2 57299 63130
0 1573 7 1 2 73974 72587
0 1574 5 1 1 1573
0 1575 7 1 2 1571 1574
0 1576 5 1 1 1575
0 1577 7 1 2 71845 1576
0 1578 5 1 1 1577
0 1579 7 2 2 70754 67910
0 1580 7 1 2 68927 73984
0 1581 5 1 1 1580
0 1582 7 5 2 57300 73459
0 1583 5 2 1 73986
0 1584 7 10 2 57573 63131
0 1585 7 1 2 73993 70567
0 1586 7 1 2 73987 1585
0 1587 5 1 1 1586
0 1588 7 1 2 1581 1587
0 1589 7 1 2 1578 1588
0 1590 5 1 1 1589
0 1591 7 1 2 67976 1590
0 1592 5 1 1 1591
0 1593 7 1 2 68298 67614
0 1594 5 1 1 1593
0 1595 7 7 2 59066 67589
0 1596 5 2 1 74003
0 1597 7 1 2 74004 70568
0 1598 5 1 1 1597
0 1599 7 1 2 1594 1598
0 1600 5 1 1 1599
0 1601 7 7 2 63132 65131
0 1602 7 1 2 74012 73867
0 1603 7 1 2 1600 1602
0 1604 5 1 1 1603
0 1605 7 1 2 1592 1604
0 1606 5 1 1 1605
0 1607 7 1 2 62028 1606
0 1608 5 1 1 1607
0 1609 7 2 2 63133 73353
0 1610 7 1 2 74019 69203
0 1611 7 1 2 72643 1610
0 1612 5 1 1 1611
0 1613 7 1 2 1608 1612
0 1614 5 1 1 1613
0 1615 7 1 2 73972 1614
0 1616 5 1 1 1615
0 1617 7 1 2 1566 1616
0 1618 5 1 1 1617
0 1619 7 1 2 71701 1618
0 1620 5 1 1 1619
0 1621 7 7 2 63800 69016
0 1622 5 15 1 74021
0 1623 7 3 2 63578 67590
0 1624 7 1 2 74043 73428
0 1625 5 1 1 1624
0 1626 7 1 2 67574 73706
0 1627 5 1 1 1626
0 1628 7 1 2 73739 1627
0 1629 5 1 1 1628
0 1630 7 1 2 57301 1629
0 1631 5 1 1 1630
0 1632 7 7 2 59212 61152
0 1633 5 1 1 74046
0 1634 7 4 2 57574 59724
0 1635 7 1 2 74047 74053
0 1636 5 1 1 1635
0 1637 7 1 2 1631 1636
0 1638 5 1 1 1637
0 1639 7 1 2 57846 1638
0 1640 5 1 1 1639
0 1641 7 2 2 57575 73033
0 1642 5 2 1 74057
0 1643 7 2 2 67575 73643
0 1644 7 1 2 57302 74061
0 1645 5 1 1 1644
0 1646 7 1 2 74059 1645
0 1647 5 1 1 1646
0 1648 7 1 2 59725 1647
0 1649 5 1 1 1648
0 1650 7 1 2 1640 1649
0 1651 5 1 1 1650
0 1652 7 1 2 72596 1651
0 1653 5 1 1 1652
0 1654 7 2 2 57303 58838
0 1655 7 3 2 67036 74063
0 1656 5 1 1 74065
0 1657 7 1 2 73747 74066
0 1658 5 1 1 1657
0 1659 7 1 2 59213 72345
0 1660 5 2 1 1659
0 1661 7 1 2 72625 74068
0 1662 5 1 1 1661
0 1663 7 1 2 73034 1662
0 1664 5 1 1 1663
0 1665 7 8 2 57576 65775
0 1666 5 3 1 74070
0 1667 7 1 2 59214 70272
0 1668 5 3 1 1667
0 1669 7 1 2 69749 74081
0 1670 5 1 1 1669
0 1671 7 1 2 74071 1670
0 1672 5 1 1 1671
0 1673 7 2 2 1664 1672
0 1674 5 1 1 74084
0 1675 7 1 2 73035 72346
0 1676 5 2 1 1675
0 1677 7 13 2 64136 65132
0 1678 5 4 1 74088
0 1679 7 1 2 57577 70273
0 1680 5 1 1 1679
0 1681 7 1 2 74101 1680
0 1682 5 2 1 1681
0 1683 7 1 2 65776 74105
0 1684 5 1 1 1683
0 1685 7 1 2 74086 1684
0 1686 5 1 1 1685
0 1687 7 1 2 57847 1686
0 1688 5 1 1 1687
0 1689 7 1 2 74085 1688
0 1690 5 1 1 1689
0 1691 7 1 2 59726 1690
0 1692 5 1 1 1691
0 1693 7 2 2 67576 70134
0 1694 5 1 1 74107
0 1695 7 1 2 57848 74108
0 1696 7 1 2 73527 1695
0 1697 5 1 1 1696
0 1698 7 1 2 1692 1697
0 1699 5 1 1 1698
0 1700 7 1 2 70569 1699
0 1701 5 1 1 1700
0 1702 7 1 2 1658 1701
0 1703 7 1 2 1653 1702
0 1704 5 1 1 1703
0 1705 7 1 2 62029 1704
0 1706 5 1 1 1705
0 1707 7 1 2 1625 1706
0 1708 5 1 1 1707
0 1709 7 1 2 58127 1708
0 1710 5 1 1 1709
0 1711 7 1 2 72461 73190
0 1712 5 3 1 1711
0 1713 7 1 2 57578 72965
0 1714 5 1 1 1713
0 1715 7 1 2 74109 1714
0 1716 5 1 1 1715
0 1717 7 1 2 70570 1716
0 1718 5 1 1 1717
0 1719 7 2 2 69728 73558
0 1720 5 3 1 74112
0 1721 7 23 2 59417 65397
0 1722 5 12 1 74117
0 1723 7 8 2 59215 65777
0 1724 5 1 1 74152
0 1725 7 1 2 74140 1724
0 1726 5 1 1 1725
0 1727 7 1 2 67577 73328
0 1728 7 1 2 1726 1727
0 1729 5 1 1 1728
0 1730 7 1 2 74114 1729
0 1731 5 1 1 1730
0 1732 7 1 2 57304 1731
0 1733 5 1 1 1732
0 1734 7 4 2 57579 59418
0 1735 7 1 2 74048 74160
0 1736 5 1 1 1735
0 1737 7 1 2 1733 1736
0 1738 5 1 1 1737
0 1739 7 1 2 72597 1738
0 1740 5 1 1 1739
0 1741 7 1 2 1718 1740
0 1742 5 1 1 1741
0 1743 7 1 2 57849 1742
0 1744 5 1 1 1743
0 1745 7 1 2 59419 74062
0 1746 5 1 1 1745
0 1747 7 1 2 74110 1746
0 1748 5 1 1 1747
0 1749 7 1 2 74067 1748
0 1750 5 1 1 1749
0 1751 7 1 2 1744 1750
0 1752 5 1 1 1751
0 1753 7 1 2 62030 1752
0 1754 5 1 1 1753
0 1755 7 5 2 63579 59216
0 1756 7 3 2 62833 74164
0 1757 7 5 2 57305 69175
0 1758 7 1 2 74169 74172
0 1759 7 1 2 73344 1758
0 1760 5 1 1 1759
0 1761 7 1 2 1754 1760
0 1762 5 1 1 1761
0 1763 7 1 2 59727 1762
0 1764 5 1 1 1763
0 1765 7 1 2 1710 1764
0 1766 5 1 1 1765
0 1767 7 1 2 58382 1766
0 1768 5 1 1 1767
0 1769 7 6 2 57306 60730
0 1770 7 1 2 74177 67615
0 1771 5 1 1 1770
0 1772 7 15 2 63134 65398
0 1773 5 6 1 74183
0 1774 7 1 2 74184 70571
0 1775 5 1 1 1774
0 1776 7 1 2 1771 1775
0 1777 5 1 1 1776
0 1778 7 1 2 62031 67578
0 1779 7 1 2 1777 1778
0 1780 5 1 1 1779
0 1781 7 5 2 63135 72462
0 1782 5 1 1 74204
0 1783 7 1 2 74205 74044
0 1784 7 1 2 71071 1783
0 1785 5 1 1 1784
0 1786 7 1 2 1780 1785
0 1787 5 1 1 1786
0 1788 7 1 2 59217 1787
0 1789 5 1 1 1788
0 1790 7 1 2 73975 67911
0 1791 7 1 2 69171 1790
0 1792 5 1 1 1791
0 1793 7 1 2 1789 1792
0 1794 5 1 1 1793
0 1795 7 1 2 57850 1794
0 1796 5 1 1 1795
0 1797 7 19 2 57307 65133
0 1798 5 4 1 74209
0 1799 7 4 2 63136 70135
0 1800 7 1 2 74210 74232
0 1801 7 1 2 67964 1800
0 1802 5 1 1 1801
0 1803 7 1 2 1796 1802
0 1804 5 1 1 1803
0 1805 7 1 2 73973 1804
0 1806 5 1 1 1805
0 1807 7 1 2 1768 1806
0 1808 5 1 1 1807
0 1809 7 1 2 74028 1808
0 1810 5 1 1 1809
0 1811 7 1 2 1620 1810
0 1812 7 1 2 1224 1811
0 1813 7 1 2 791 1812
0 1814 5 1 1 1813
0 1815 7 1 2 66883 1814
0 1816 5 1 1 1815
0 1817 7 3 2 59218 66739
0 1818 7 4 2 66662 68928
0 1819 7 1 2 74236 74239
0 1820 5 1 1 1819
0 1821 7 9 2 62032 66807
0 1822 7 32 2 66545 74243
0 1823 5 3 1 74252
0 1824 7 1 2 64931 74253
0 1825 5 1 1 1824
0 1826 7 1 2 1820 1825
0 1827 5 1 1 1826
0 1828 7 1 2 72347 1827
0 1829 5 1 1 1828
0 1830 7 17 2 65399 61889
0 1831 7 6 2 66663 66740
0 1832 7 3 2 74287 74304
0 1833 5 1 1 74310
0 1834 7 37 2 64932 65134
0 1835 5 36 1 74313
0 1836 7 1 2 74350 70886
0 1837 7 1 2 74311 1836
0 1838 5 1 1 1837
0 1839 7 1 2 1829 1838
0 1840 5 1 1 1839
0 1841 7 1 2 58932 1840
0 1842 5 1 1 1841
0 1843 7 1 2 59219 71983
0 1844 5 3 1 1843
0 1845 7 1 2 74228 74386
0 1846 5 1 1 1845
0 1847 7 1 2 72290 879
0 1848 5 8 1 1847
0 1849 7 17 2 66741 67503
0 1850 7 1 2 74389 74397
0 1851 7 1 2 1846 1850
0 1852 5 1 1 1851
0 1853 7 3 2 59220 59957
0 1854 7 6 2 58701 74414
0 1855 7 1 2 67451 74417
0 1856 5 1 1 1855
0 1857 7 1 2 1852 1856
0 1858 7 1 2 1842 1857
0 1859 5 1 1 1858
0 1860 7 1 2 59067 1859
0 1861 5 1 1 1860
0 1862 7 1 2 74284 1833
0 1863 5 2 1 1862
0 1864 7 1 2 64933 74285
0 1865 5 1 1 1864
0 1866 7 1 2 72348 1865
0 1867 7 1 2 74423 1866
0 1868 5 1 1 1867
0 1869 7 5 2 63438 58933
0 1870 7 4 2 64654 74425
0 1871 7 8 2 60217 61890
0 1872 7 2 2 65400 66664
0 1873 7 1 2 74434 74442
0 1874 7 1 2 74430 1873
0 1875 5 1 1 1874
0 1876 7 1 2 1868 1875
0 1877 5 1 1 1876
0 1878 7 1 2 59221 1877
0 1879 5 1 1 1878
0 1880 7 2 2 72463 74254
0 1881 5 2 1 74444
0 1882 7 1 2 1879 74446
0 1883 7 1 2 1861 1882
0 1884 5 1 1 1883
0 1885 7 1 2 61153 1884
0 1886 5 1 1 1885
0 1887 7 8 2 63801 65135
0 1888 5 6 1 74448
0 1889 7 1 2 60446 70025
0 1890 5 2 1 1889
0 1891 7 1 2 74456 74462
0 1892 5 1 1 1891
0 1893 7 8 2 64655 60731
0 1894 7 3 2 63439 74464
0 1895 7 10 2 63938 65778
0 1896 7 1 2 74475 67504
0 1897 7 1 2 74472 1896
0 1898 7 1 2 1892 1897
0 1899 5 1 1 1898
0 1900 7 1 2 1886 1899
0 1901 5 1 1 1900
0 1902 7 1 2 59420 1901
0 1903 5 1 1 1902
0 1904 7 4 2 66546 66808
0 1905 7 1 2 67969 74485
0 1906 5 1 1 1905
0 1907 7 4 2 58934 64656
0 1908 7 2 2 69866 74489
0 1909 7 5 2 60732 67505
0 1910 7 4 2 57308 63440
0 1911 7 1 2 74495 74500
0 1912 7 1 2 74493 1911
0 1913 5 1 1 1912
0 1914 7 1 2 1906 1913
0 1915 5 1 1 1914
0 1916 7 1 2 72995 1915
0 1917 5 1 1 1916
0 1918 7 17 2 64934 60447
0 1919 5 2 1 74504
0 1920 7 2 2 73849 69896
0 1921 5 1 1 74523
0 1922 7 1 2 64137 1921
0 1923 5 1 1 1922
0 1924 7 1 2 74505 1923
0 1925 5 1 1 1924
0 1926 7 1 2 68449 73812
0 1927 5 1 1 1926
0 1928 7 1 2 60218 73277
0 1929 7 1 2 1927 1928
0 1930 5 1 1 1929
0 1931 7 1 2 1925 1930
0 1932 5 1 1 1931
0 1933 7 1 2 65401 1932
0 1934 5 1 1 1933
0 1935 7 22 2 59421 60733
0 1936 5 7 1 74525
0 1937 7 4 2 57309 69109
0 1938 5 1 1 74554
0 1939 7 1 2 63939 1938
0 1940 5 1 1 1939
0 1941 7 1 2 74526 1940
0 1942 5 1 1 1941
0 1943 7 1 2 1934 1942
0 1944 5 1 1 1943
0 1945 7 1 2 74398 1944
0 1946 5 1 1 1945
0 1947 7 4 2 64935 73139
0 1948 5 1 1 74558
0 1949 7 1 2 69110 74559
0 1950 5 1 1 1949
0 1951 7 1 2 72939 1950
0 1952 5 1 1 1951
0 1953 7 1 2 65136 1952
0 1954 5 1 1 1953
0 1955 7 1 2 59422 68205
0 1956 5 1 1 1955
0 1957 7 1 2 1954 1956
0 1958 5 1 1 1957
0 1959 7 1 2 74255 1958
0 1960 5 1 1 1959
0 1961 7 1 2 1946 1960
0 1962 5 1 1 1961
0 1963 7 1 2 61154 1962
0 1964 5 1 1 1963
0 1965 7 1 2 1917 1964
0 1966 5 1 1 1965
0 1967 7 1 2 57851 1966
0 1968 5 1 1 1967
0 1969 7 3 2 74244 69134
0 1970 7 1 2 65137 73685
0 1971 7 1 2 72930 1970
0 1972 7 1 2 74562 1971
0 1973 5 1 1 1972
0 1974 7 1 2 1968 1973
0 1975 7 1 2 1903 1974
0 1976 5 1 1 1975
0 1977 7 1 2 57580 1976
0 1978 5 1 1 1977
0 1979 7 6 2 57852 68553
0 1980 5 1 1 74565
0 1981 7 2 2 67626 74566
0 1982 5 2 1 74571
0 1983 7 1 2 74573 73416
0 1984 5 1 1 1983
0 1985 7 1 2 73140 73193
0 1986 5 1 1 1985
0 1987 7 1 2 1984 1986
0 1988 5 1 1 1987
0 1989 7 1 2 74256 1988
0 1990 5 1 1 1989
0 1991 7 7 2 59068 60448
0 1992 5 1 1 74575
0 1993 7 2 2 1992 74457
0 1994 5 9 1 74582
0 1995 7 1 2 68554 74584
0 1996 5 1 1 1995
0 1997 7 2 2 57853 63802
0 1998 5 1 1 74593
0 1999 7 1 2 71019 1998
0 2000 7 1 2 1996 1999
0 2001 5 1 1 2000
0 2002 7 1 2 63940 2001
0 2003 5 1 1 2002
0 2004 7 5 2 63803 64936
0 2005 7 4 2 62292 74595
0 2006 5 2 1 74600
0 2007 7 1 2 65138 74601
0 2008 5 1 1 2007
0 2009 7 1 2 69766 2008
0 2010 5 1 1 2009
0 2011 7 1 2 68450 2010
0 2012 5 3 1 2011
0 2013 7 5 2 62293 59222
0 2014 7 1 2 70044 74609
0 2015 5 1 1 2014
0 2016 7 1 2 74606 2015
0 2017 7 1 2 2003 2016
0 2018 5 1 1 2017
0 2019 7 1 2 60734 2018
0 2020 5 1 1 2019
0 2021 7 1 2 65779 70989
0 2022 7 1 2 2020 2021
0 2023 5 1 1 2022
0 2024 7 1 2 72222 72546
0 2025 7 1 2 70035 2024
0 2026 5 1 1 2025
0 2027 7 1 2 71984 2026
0 2028 5 1 1 2027
0 2029 7 1 2 63804 68816
0 2030 5 4 1 2029
0 2031 7 1 2 74614 72298
0 2032 5 2 1 2031
0 2033 7 3 2 59223 72130
0 2034 5 1 1 74620
0 2035 7 1 2 58935 74621
0 2036 5 1 1 2035
0 2037 7 1 2 74618 2036
0 2038 7 1 2 2028 2037
0 2039 5 1 1 2038
0 2040 7 1 2 57854 2039
0 2041 5 1 1 2040
0 2042 7 2 2 60219 68555
0 2043 7 1 2 71846 74623
0 2044 5 1 1 2043
0 2045 7 7 2 57581 70694
0 2046 5 7 1 74625
0 2047 7 1 2 74314 74632
0 2048 5 2 1 2047
0 2049 7 1 2 2044 74639
0 2050 5 1 1 2049
0 2051 7 1 2 70136 2050
0 2052 5 1 1 2051
0 2053 7 1 2 61155 2052
0 2054 7 1 2 2041 2053
0 2055 5 1 1 2054
0 2056 7 1 2 2055 74399
0 2057 7 1 2 2023 2056
0 2058 5 1 1 2057
0 2059 7 1 2 1990 2058
0 2060 5 1 1 2059
0 2061 7 1 2 59423 2060
0 2062 5 1 1 2061
0 2063 7 4 2 72931 72957
0 2064 7 1 2 57855 74641
0 2065 5 1 1 2064
0 2066 7 1 2 59224 73529
0 2067 5 1 1 2066
0 2068 7 1 2 2065 2067
0 2069 5 2 1 2068
0 2070 7 1 2 74645 74563
0 2071 5 1 1 2070
0 2072 7 4 2 65402 73081
0 2073 7 1 2 74647 74257
0 2074 5 1 1 2073
0 2075 7 1 2 57856 74211
0 2076 7 9 2 64657 61156
0 2077 5 1 1 74651
0 2078 7 10 2 63441 59424
0 2079 7 1 2 74652 74660
0 2080 7 1 2 2075 2079
0 2081 7 1 2 74496 2080
0 2082 5 1 1 2081
0 2083 7 1 2 2074 2082
0 2084 5 1 1 2083
0 2085 7 1 2 69094 2084
0 2086 5 1 1 2085
0 2087 7 1 2 2071 2086
0 2088 7 1 2 2062 2087
0 2089 7 1 2 1978 2088
0 2090 5 1 1 2089
0 2091 7 1 2 58128 2090
0 2092 5 1 1 2091
0 2093 7 1 2 71458 74642
0 2094 5 1 1 2093
0 2095 7 1 2 2094 73030
0 2096 5 2 1 2095
0 2097 7 1 2 57310 74670
0 2098 5 1 1 2097
0 2099 7 5 2 58129 73036
0 2100 5 3 1 74672
0 2101 7 1 2 2098 74677
0 2102 5 2 1 2101
0 2103 7 1 2 59069 74680
0 2104 5 1 1 2103
0 2105 7 10 2 58130 61157
0 2106 5 6 1 74682
0 2107 7 1 2 73022 74692
0 2108 5 6 1 2107
0 2109 7 2 2 70137 74698
0 2110 5 1 1 74704
0 2111 7 2 2 58131 73082
0 2112 5 2 1 74706
0 2113 7 1 2 2110 74708
0 2114 5 1 1 2113
0 2115 7 2 2 65139 2114
0 2116 5 1 1 74710
0 2117 7 1 2 57311 74711
0 2118 5 1 1 2117
0 2119 7 1 2 2104 2118
0 2120 5 1 1 2119
0 2121 7 1 2 57857 2120
0 2122 5 1 1 2121
0 2123 7 2 2 73850 67095
0 2124 7 1 2 74113 74712
0 2125 5 1 1 2124
0 2126 7 1 2 57312 73530
0 2127 5 1 1 2126
0 2128 7 1 2 73059 2127
0 2129 5 1 1 2128
0 2130 7 1 2 59225 2129
0 2131 5 1 1 2130
0 2132 7 1 2 57313 74648
0 2133 5 1 1 2132
0 2134 7 1 2 2131 2133
0 2135 5 1 1 2134
0 2136 7 1 2 68299 2135
0 2137 5 1 1 2136
0 2138 7 2 2 67711 73100
0 2139 5 2 1 74714
0 2140 7 1 2 59425 74716
0 2141 5 1 1 2140
0 2142 7 1 2 67096 73790
0 2143 5 2 1 2142
0 2144 7 1 2 2141 74718
0 2145 5 1 1 2144
0 2146 7 1 2 61158 2145
0 2147 5 1 1 2146
0 2148 7 1 2 67627 72996
0 2149 5 2 1 2148
0 2150 7 1 2 2147 74720
0 2151 5 1 1 2150
0 2152 7 1 2 74212 2151
0 2153 5 1 1 2152
0 2154 7 1 2 2137 2153
0 2155 5 1 1 2154
0 2156 7 1 2 58132 2155
0 2157 5 1 1 2156
0 2158 7 1 2 2125 2157
0 2159 7 1 2 2122 2158
0 2160 5 1 1 2159
0 2161 7 1 2 74258 2160
0 2162 5 1 1 2161
0 2163 7 1 2 74259 74681
0 2164 5 1 1 2163
0 2165 7 8 2 65780 71381
0 2166 5 3 1 74722
0 2167 7 1 2 70138 74723
0 2168 5 1 1 2167
0 2169 7 1 2 60735 74673
0 2170 5 1 1 2169
0 2171 7 1 2 2168 2170
0 2172 5 1 1 2171
0 2173 7 2 2 74400 2172
0 2174 5 1 1 74733
0 2175 7 4 2 61159 71459
0 2176 5 3 1 74735
0 2177 7 1 2 73023 74739
0 2178 5 4 1 2177
0 2179 7 6 2 59958 67452
0 2180 7 2 2 58702 73141
0 2181 7 1 2 57314 74752
0 2182 7 1 2 74746 2181
0 2183 7 1 2 74742 2182
0 2184 5 1 1 2183
0 2185 7 1 2 2174 2184
0 2186 5 1 1 2185
0 2187 7 1 2 70755 2186
0 2188 5 1 1 2187
0 2189 7 1 2 2164 2188
0 2190 5 1 1 2189
0 2191 7 1 2 69176 2190
0 2192 5 1 1 2191
0 2193 7 1 2 2162 2192
0 2194 5 1 1 2193
0 2195 7 1 2 71702 2194
0 2196 5 1 1 2195
0 2197 7 1 2 74260 74671
0 2198 5 1 1 2197
0 2199 7 1 2 74213 74734
0 2200 5 1 1 2199
0 2201 7 1 2 2198 2200
0 2202 5 1 1 2201
0 2203 7 1 2 57582 2202
0 2204 5 1 1 2203
0 2205 7 3 2 61160 71140
0 2206 7 1 2 57315 74754
0 2207 5 1 1 2206
0 2208 7 1 2 2116 2207
0 2209 5 1 1 2208
0 2210 7 1 2 74261 2209
0 2211 5 1 1 2210
0 2212 7 1 2 2204 2211
0 2213 5 1 1 2212
0 2214 7 1 2 57858 2213
0 2215 5 1 1 2214
0 2216 7 8 2 58133 58703
0 2217 5 1 1 74757
0 2218 7 1 2 74758 74747
0 2219 7 1 2 1674 2218
0 2220 5 1 1 2219
0 2221 7 1 2 2215 2220
0 2222 5 1 1 2221
0 2223 7 1 2 74029 2222
0 2224 5 1 1 2223
0 2225 7 1 2 58936 69867
0 2226 5 2 1 2225
0 2227 7 1 2 67022 74765
0 2228 5 1 1 2227
0 2229 7 1 2 74262 2228
0 2230 5 1 1 2229
0 2231 7 2 2 64658 61891
0 2232 7 6 2 66665 74767
0 2233 7 2 2 63442 69111
0 2234 7 2 2 74769 74775
0 2235 7 5 2 62834 65140
0 2236 5 3 1 74779
0 2237 7 2 2 57583 60449
0 2238 5 1 1 74787
0 2239 7 1 2 74784 2238
0 2240 5 2 1 2239
0 2241 7 1 2 70864 74789
0 2242 7 1 2 74777 2241
0 2243 5 1 1 2242
0 2244 7 1 2 2230 2243
0 2245 5 1 1 2244
0 2246 7 1 2 57859 2245
0 2247 5 1 1 2246
0 2248 7 7 2 59959 62033
0 2249 7 3 2 66547 74791
0 2250 7 15 2 57584 58937
0 2251 5 5 1 74801
0 2252 7 7 2 58704 59070
0 2253 7 2 2 74802 74821
0 2254 7 1 2 74315 74828
0 2255 7 1 2 74798 2254
0 2256 5 1 1 2255
0 2257 7 1 2 64138 2256
0 2258 7 1 2 2247 2257
0 2259 5 1 1 2258
0 2260 7 12 2 63740 70916
0 2261 7 2 2 63443 74830
0 2262 7 7 2 64659 64937
0 2263 5 1 1 74844
0 2264 7 2 2 63805 74845
0 2265 7 3 2 66666 69159
0 2266 7 1 2 62555 74853
0 2267 7 1 2 74851 2266
0 2268 7 1 2 74842 2267
0 2269 5 1 1 2268
0 2270 7 7 2 57860 71847
0 2271 5 16 1 74856
0 2272 7 4 2 74863 70596
0 2273 5 2 1 74879
0 2274 7 1 2 74880 74263
0 2275 5 1 1 2274
0 2276 7 1 2 59426 2275
0 2277 7 1 2 2269 2276
0 2278 5 1 1 2277
0 2279 7 1 2 65781 2278
0 2280 7 1 2 2259 2279
0 2281 5 1 1 2280
0 2282 7 8 2 58705 62034
0 2283 7 6 2 58938 59960
0 2284 7 2 2 74885 74893
0 2285 7 1 2 71356 74899
0 2286 5 1 1 2285
0 2287 7 10 2 64660 60220
0 2288 5 1 1 74901
0 2289 7 7 2 63444 74902
0 2290 7 1 2 70585 74854
0 2291 7 1 2 74911 2290
0 2292 5 1 1 2291
0 2293 7 1 2 2286 2292
0 2294 5 1 1 2293
0 2295 7 1 2 73224 73194
0 2296 7 1 2 2294 2295
0 2297 5 1 1 2296
0 2298 7 1 2 2281 2297
0 2299 5 1 1 2298
0 2300 7 1 2 65403 2299
0 2301 5 1 1 2300
0 2302 7 1 2 64139 73559
0 2303 5 4 1 2302
0 2304 7 1 2 74918 74087
0 2305 5 1 1 2304
0 2306 7 1 2 69177 2305
0 2307 7 1 2 74564 2306
0 2308 5 1 1 2307
0 2309 7 1 2 2301 2308
0 2310 5 1 1 2309
0 2311 7 1 2 59226 2310
0 2312 5 1 1 2311
0 2313 7 1 2 74527 73772
0 2314 5 2 1 2313
0 2315 7 1 2 67007 74649
0 2316 5 1 1 2315
0 2317 7 1 2 74922 2316
0 2318 5 1 1 2317
0 2319 7 1 2 74264 70727
0 2320 7 1 2 2318 2319
0 2321 5 1 1 2320
0 2322 7 1 2 2312 2321
0 2323 7 1 2 2224 2322
0 2324 7 1 2 2196 2323
0 2325 7 1 2 2092 2324
0 2326 5 1 1 2325
0 2327 7 1 2 63137 2326
0 2328 5 1 1 2327
0 2329 7 6 2 63806 59427
0 2330 7 2 2 70274 74924
0 2331 5 3 1 74930
0 2332 7 11 2 62149 62556
0 2333 5 2 1 74935
0 2334 7 4 2 60221 72187
0 2335 5 1 1 74948
0 2336 7 2 2 74936 74949
0 2337 5 1 1 74952
0 2338 7 1 2 74931 74953
0 2339 5 1 1 2338
0 2340 7 3 2 62294 69884
0 2341 5 1 1 74954
0 2342 7 1 2 59227 74955
0 2343 5 1 1 2342
0 2344 7 1 2 71000 2343
0 2345 5 1 1 2344
0 2346 7 1 2 60450 2345
0 2347 5 2 1 2346
0 2348 7 1 2 69914 71046
0 2349 5 1 1 2348
0 2350 7 1 2 74957 2349
0 2351 5 1 1 2350
0 2352 7 1 2 60736 2351
0 2353 5 1 1 2352
0 2354 7 7 2 59228 60451
0 2355 5 2 1 74959
0 2356 7 31 2 60222 60737
0 2357 5 14 1 74968
0 2358 7 1 2 74960 74969
0 2359 5 2 1 2358
0 2360 7 11 2 63941 65404
0 2361 5 4 1 75015
0 2362 7 4 2 62557 75016
0 2363 5 7 1 75030
0 2364 7 1 2 75013 75034
0 2365 5 1 1 2364
0 2366 7 1 2 68451 2365
0 2367 5 1 1 2366
0 2368 7 4 2 59071 63942
0 2369 7 2 2 72131 75041
0 2370 5 4 1 75045
0 2371 7 2 2 68212 70666
0 2372 5 3 1 75051
0 2373 7 1 2 75047 75053
0 2374 5 1 1 2373
0 2375 7 1 2 62558 2374
0 2376 5 1 1 2375
0 2377 7 1 2 2367 2376
0 2378 7 1 2 2353 2377
0 2379 5 1 1 2378
0 2380 7 1 2 64140 2379
0 2381 5 1 1 2380
0 2382 7 1 2 2339 2381
0 2383 5 1 1 2382
0 2384 7 1 2 74401 2383
0 2385 5 1 1 2384
0 2386 7 4 2 64141 67128
0 2387 7 1 2 74265 75056
0 2388 5 1 1 2387
0 2389 7 6 2 72064 70597
0 2390 5 2 1 75060
0 2391 7 1 2 75061 74266
0 2392 5 2 1 2391
0 2393 7 7 2 65141 74596
0 2394 5 2 1 75070
0 2395 7 3 2 63445 63741
0 2396 7 1 2 75071 75079
0 2397 7 3 2 60738 70917
0 2398 5 1 1 75082
0 2399 7 1 2 74770 75083
0 2400 7 1 2 2396 2399
0 2401 5 1 1 2400
0 2402 7 1 2 75068 2401
0 2403 5 1 1 2402
0 2404 7 1 2 73582 2403
0 2405 5 1 1 2404
0 2406 7 1 2 2388 2405
0 2407 7 1 2 2385 2406
0 2408 5 1 1 2407
0 2409 7 1 2 62835 2408
0 2410 5 1 1 2409
0 2411 7 6 2 60452 70183
0 2412 5 1 1 75085
0 2413 7 1 2 75086 74267
0 2414 5 1 1 2413
0 2415 7 2 2 62295 74402
0 2416 7 3 2 59229 69406
0 2417 5 8 1 75093
0 2418 7 5 2 63943 74351
0 2419 5 6 1 75104
0 2420 7 2 2 60739 75109
0 2421 7 1 2 75096 75115
0 2422 7 1 2 75091 2421
0 2423 5 1 1 2422
0 2424 7 1 2 2414 2423
0 2425 5 1 1 2424
0 2426 7 1 2 68452 2425
0 2427 5 1 1 2426
0 2428 7 3 2 62035 70184
0 2429 7 1 2 67558 74486
0 2430 7 1 2 75117 2429
0 2431 5 1 1 2430
0 2432 7 1 2 2427 2431
0 2433 5 1 1 2432
0 2434 7 14 2 62559 63807
0 2435 5 1 1 75120
0 2436 7 1 2 64142 75121
0 2437 7 1 2 2433 2436
0 2438 5 1 1 2437
0 2439 7 1 2 2410 2438
0 2440 5 1 1 2439
0 2441 7 1 2 65782 2440
0 2442 5 1 1 2441
0 2443 7 16 2 62836 65405
0 2444 5 6 1 75134
0 2445 7 1 2 75150 75048
0 2446 5 1 1 2445
0 2447 7 1 2 68556 2446
0 2448 5 1 1 2447
0 2449 7 1 2 62837 72054
0 2450 5 1 1 2449
0 2451 7 1 2 2448 2450
0 2452 5 1 1 2451
0 2453 7 1 2 60223 2452
0 2454 5 1 1 2453
0 2455 7 2 2 65142 74615
0 2456 5 3 1 75156
0 2457 7 1 2 64938 75157
0 2458 5 1 1 2457
0 2459 7 1 2 63944 2458
0 2460 5 1 1 2459
0 2461 7 1 2 70900 2460
0 2462 5 1 1 2461
0 2463 7 1 2 62838 72012
0 2464 5 2 1 2463
0 2465 7 1 2 73101 68900
0 2466 5 1 1 2465
0 2467 7 1 2 75161 2466
0 2468 5 1 1 2467
0 2469 7 1 2 60453 2468
0 2470 5 1 1 2469
0 2471 7 1 2 2462 2470
0 2472 7 1 2 2454 2471
0 2473 5 1 1 2472
0 2474 7 1 2 69178 2473
0 2475 5 1 1 2474
0 2476 7 15 2 57316 68974
0 2477 5 17 1 75163
0 2478 7 2 2 60740 75178
0 2479 5 11 1 75195
0 2480 7 4 2 72039 75197
0 2481 7 1 2 70756 75208
0 2482 5 1 1 2481
0 2483 7 1 2 60224 72055
0 2484 5 1 1 2483
0 2485 7 1 2 2034 2484
0 2486 5 1 1 2485
0 2487 7 1 2 68557 2486
0 2488 5 1 1 2487
0 2489 7 1 2 74387 74619
0 2490 7 1 2 2488 2489
0 2491 7 1 2 2482 2490
0 2492 5 1 1 2491
0 2493 7 1 2 57861 2492
0 2494 5 1 1 2493
0 2495 7 8 2 65406 67628
0 2496 7 2 2 58939 69832
0 2497 5 1 1 75220
0 2498 7 2 2 58940 74506
0 2499 5 2 1 75222
0 2500 7 1 2 69855 75224
0 2501 5 2 1 2500
0 2502 7 1 2 57317 75226
0 2503 5 7 1 2502
0 2504 7 1 2 2497 75228
0 2505 5 8 1 2504
0 2506 7 1 2 75212 75235
0 2507 5 1 1 2506
0 2508 7 5 2 71789 70598
0 2509 5 1 1 75243
0 2510 7 1 2 60225 71034
0 2511 7 1 2 2509 2510
0 2512 5 2 1 2511
0 2513 7 1 2 74640 75248
0 2514 5 1 1 2513
0 2515 7 1 2 65407 2514
0 2516 5 1 1 2515
0 2517 7 1 2 71635 2516
0 2518 5 1 1 2517
0 2519 7 1 2 59230 2518
0 2520 5 1 1 2519
0 2521 7 1 2 2507 2520
0 2522 7 1 2 2494 2521
0 2523 5 1 1 2522
0 2524 7 1 2 62839 2523
0 2525 5 1 1 2524
0 2526 7 1 2 2475 2525
0 2527 5 1 1 2526
0 2528 7 1 2 74403 2527
0 2529 5 1 1 2528
0 2530 7 8 2 57318 71703
0 2531 5 9 1 75250
0 2532 7 12 2 69017 75258
0 2533 5 10 1 75267
0 2534 7 1 2 68213 75268
0 2535 5 4 1 2534
0 2536 7 1 2 65143 75289
0 2537 5 1 1 2536
0 2538 7 2 2 62560 2537
0 2539 5 1 1 75293
0 2540 7 1 2 62840 73142
0 2541 7 1 2 2539 2540
0 2542 5 1 1 2541
0 2543 7 6 2 60454 68300
0 2544 5 1 1 75295
0 2545 7 5 2 60741 67249
0 2546 5 3 1 75301
0 2547 7 1 2 57319 75017
0 2548 5 1 1 2547
0 2549 7 1 2 75306 2548
0 2550 5 1 1 2549
0 2551 7 1 2 75296 2550
0 2552 5 1 1 2551
0 2553 7 3 2 60742 67822
0 2554 5 1 1 75309
0 2555 7 2 2 63945 75310
0 2556 5 1 1 75312
0 2557 7 1 2 74214 75313
0 2558 5 1 1 2557
0 2559 7 1 2 2552 2558
0 2560 5 1 1 2559
0 2561 7 1 2 71704 2560
0 2562 5 1 1 2561
0 2563 7 1 2 63946 67810
0 2564 5 29 1 2563
0 2565 7 1 2 68975 69975
0 2566 7 1 2 72349 2565
0 2567 7 1 2 75314 2566
0 2568 5 2 1 2567
0 2569 7 1 2 60455 74626
0 2570 5 1 1 2569
0 2571 7 1 2 75343 2570
0 2572 5 1 1 2571
0 2573 7 1 2 60743 2572
0 2574 5 1 1 2573
0 2575 7 2 2 57320 75302
0 2576 5 1 1 75345
0 2577 7 2 2 68976 75018
0 2578 5 1 1 75347
0 2579 7 1 2 60456 2578
0 2580 7 1 2 2576 2579
0 2581 5 1 1 2580
0 2582 7 4 2 65144 73143
0 2583 5 2 1 75349
0 2584 7 6 2 62561 65145
0 2585 5 2 1 75355
0 2586 7 1 2 68301 75361
0 2587 7 1 2 75353 2586
0 2588 7 1 2 2581 2587
0 2589 5 1 1 2588
0 2590 7 1 2 2574 2589
0 2591 7 1 2 2562 2590
0 2592 7 2 2 2542 2591
0 2593 5 1 1 75363
0 2594 7 1 2 63808 70712
0 2595 5 1 1 2594
0 2596 7 1 2 75364 2595
0 2597 5 2 1 2596
0 2598 7 1 2 75365 74268
0 2599 5 1 1 2598
0 2600 7 1 2 64143 2599
0 2601 7 1 2 2529 2600
0 2602 5 1 1 2601
0 2603 7 4 2 63446 63809
0 2604 7 7 2 64661 60457
0 2605 5 1 1 75371
0 2606 7 1 2 72713 75372
0 2607 7 1 2 75367 2606
0 2608 7 2 2 74497 2607
0 2609 5 1 1 75378
0 2610 7 1 2 58134 75379
0 2611 5 1 1 2610
0 2612 7 1 2 75069 2611
0 2613 5 1 1 2612
0 2614 7 1 2 62562 2613
0 2615 5 1 1 2614
0 2616 7 1 2 70901 74269
0 2617 5 1 1 2616
0 2618 7 1 2 2615 2617
0 2619 5 1 1 2618
0 2620 7 1 2 63947 2619
0 2621 5 1 1 2620
0 2622 7 3 2 62841 58706
0 2623 7 1 2 70599 75380
0 2624 7 1 2 74799 2623
0 2625 5 1 1 2624
0 2626 7 2 2 68453 74240
0 2627 7 3 2 58135 66742
0 2628 7 17 2 63948 60226
0 2629 5 4 1 75388
0 2630 7 3 2 62296 75389
0 2631 5 2 1 75409
0 2632 7 1 2 75385 75410
0 2633 7 1 2 75383 2632
0 2634 5 1 1 2633
0 2635 7 1 2 2625 2634
0 2636 5 1 1 2635
0 2637 7 1 2 74864 2636
0 2638 5 1 1 2637
0 2639 7 1 2 59428 2638
0 2640 7 1 2 2621 2639
0 2641 5 1 1 2640
0 2642 7 1 2 61161 2641
0 2643 7 1 2 2602 2642
0 2644 5 1 1 2643
0 2645 7 1 2 2442 2644
0 2646 5 2 1 2645
0 2647 7 1 2 58383 75414
0 2648 5 1 1 2647
0 2649 7 5 2 64144 70275
0 2650 7 5 2 58707 64939
0 2651 7 1 2 74049 75421
0 2652 7 1 2 74748 2651
0 2653 7 1 2 75416 2652
0 2654 7 1 2 72837 2653
0 2655 5 1 1 2654
0 2656 7 1 2 64441 2655
0 2657 7 1 2 2648 2656
0 2658 7 1 2 2328 2657
0 2659 5 1 1 2658
0 2660 7 1 2 63138 75415
0 2661 5 1 1 2660
0 2662 7 25 2 58384 64145
0 2663 5 8 1 75426
0 2664 7 12 2 62842 61162
0 2665 5 1 1 75459
0 2666 7 3 2 67129 75460
0 2667 7 2 2 75427 75471
0 2668 5 1 1 75474
0 2669 7 14 2 62297 60227
0 2670 5 5 1 75476
0 2671 7 1 2 74404 75477
0 2672 5 1 1 2671
0 2673 7 1 2 74286 2672
0 2674 5 1 1 2673
0 2675 7 1 2 68454 2674
0 2676 5 1 1 2675
0 2677 7 1 2 62298 66809
0 2678 7 1 2 67453 2677
0 2679 5 1 1 2678
0 2680 7 1 2 2676 2679
0 2681 5 1 1 2680
0 2682 7 1 2 72065 2681
0 2683 5 1 1 2682
0 2684 7 1 2 2609 2683
0 2685 5 1 1 2684
0 2686 7 1 2 75475 2685
0 2687 5 1 1 2686
0 2688 7 1 2 59728 2687
0 2689 7 1 2 2661 2688
0 2690 5 1 1 2689
0 2691 7 1 2 70472 2690
0 2692 7 1 2 2659 2691
0 2693 5 1 1 2692
0 2694 7 71 2 63139 64442
0 2695 5 41 1 75495
0 2696 7 61 2 61892 66810
0 2697 5 5 1 75607
0 2698 7 2 2 70805 75179
0 2699 5 2 1 75673
0 2700 7 1 2 57585 75675
0 2701 5 1 1 2700
0 2702 7 1 2 69976 2701
0 2703 5 1 1 2702
0 2704 7 1 2 75608 2703
0 2705 5 1 1 2704
0 2706 7 12 2 58708 61893
0 2707 7 6 2 59961 64940
0 2708 7 4 2 75677 75689
0 2709 5 7 1 75695
0 2710 7 15 2 58941 67591
0 2711 5 3 1 75706
0 2712 7 19 2 64662 66548
0 2713 7 28 2 63447 75724
0 2714 7 1 2 75707 75743
0 2715 5 1 1 2714
0 2716 7 1 2 75699 2715
0 2717 5 1 1 2716
0 2718 7 1 2 72228 2717
0 2719 5 1 1 2718
0 2720 7 6 2 62299 68817
0 2721 5 17 1 75771
0 2722 7 3 2 71848 75777
0 2723 5 3 1 75794
0 2724 7 11 2 63448 59231
0 2725 7 2 2 75800 75725
0 2726 5 2 1 75811
0 2727 7 1 2 75700 75813
0 2728 5 3 1 2727
0 2729 7 1 2 75795 75815
0 2730 5 1 1 2729
0 2731 7 5 2 64663 67107
0 2732 7 4 2 63449 59072
0 2733 7 3 2 75818 75823
0 2734 5 1 1 75827
0 2735 7 1 2 59232 75828
0 2736 5 2 1 2735
0 2737 7 1 2 2730 75830
0 2738 7 1 2 2719 2737
0 2739 7 1 2 2705 2738
0 2740 5 1 1 2739
0 2741 7 1 2 57862 2740
0 2742 5 1 1 2741
0 2743 7 1 2 70757 67097
0 2744 5 2 1 2743
0 2745 7 10 2 60458 67712
0 2746 5 9 1 75834
0 2747 7 35 2 68302 75844
0 2748 5 1 1 75853
0 2749 7 4 2 59233 75854
0 2750 5 1 1 75888
0 2751 7 4 2 59234 71849
0 2752 5 20 1 75892
0 2753 7 4 2 57586 72229
0 2754 5 2 1 75916
0 2755 7 1 2 75896 75920
0 2756 5 7 1 2755
0 2757 7 1 2 68718 75922
0 2758 5 1 1 2757
0 2759 7 1 2 2750 2758
0 2760 5 2 1 2759
0 2761 7 1 2 64941 75929
0 2762 5 1 1 2761
0 2763 7 1 2 75832 2762
0 2764 5 1 1 2763
0 2765 7 1 2 75609 2764
0 2766 5 1 1 2765
0 2767 7 1 2 2742 2766
0 2768 5 1 1 2767
0 2769 7 1 2 65408 2768
0 2770 5 1 1 2769
0 2771 7 5 2 62563 60744
0 2772 5 12 1 75931
0 2773 7 1 2 75936 74426
0 2774 7 1 2 75819 2773
0 2775 7 1 2 74713 2774
0 2776 5 1 1 2775
0 2777 7 1 2 2770 2776
0 2778 5 1 1 2777
0 2779 7 1 2 69592 2778
0 2780 5 1 1 2779
0 2781 7 19 2 59962 61894
0 2782 7 22 2 58709 75948
0 2783 5 17 1 75967
0 2784 7 1 2 68303 75968
0 2785 5 2 1 2784
0 2786 7 1 2 72373 75744
0 2787 5 2 1 2786
0 2788 7 1 2 76006 76008
0 2789 5 1 1 2788
0 2790 7 1 2 67250 2789
0 2791 5 1 1 2790
0 2792 7 5 2 57863 75801
0 2793 7 4 2 64664 71357
0 2794 7 1 2 76010 76015
0 2795 5 2 1 2794
0 2796 7 1 2 2791 76019
0 2797 5 1 1 2796
0 2798 7 1 2 69593 2797
0 2799 5 1 1 2798
0 2800 7 18 2 59963 64776
0 2801 7 3 2 76021 67506
0 2802 7 2 2 63580 69179
0 2803 7 4 2 59073 60228
0 2804 5 1 1 76044
0 2805 7 6 2 58710 59235
0 2806 7 1 2 76045 76048
0 2807 7 1 2 76042 2806
0 2808 7 1 2 76039 2807
0 2809 5 1 1 2808
0 2810 7 1 2 2799 2809
0 2811 5 1 1 2810
0 2812 7 1 2 65146 2811
0 2813 5 1 1 2812
0 2814 7 12 2 64665 60101
0 2815 7 4 2 63450 76054
0 2816 5 1 1 76066
0 2817 7 1 2 67977 76067
0 2818 7 8 2 64942 68304
0 2819 5 5 1 76070
0 2820 7 3 2 58839 67454
0 2821 7 1 2 76071 76083
0 2822 7 1 2 2817 2821
0 2823 5 1 1 2822
0 2824 7 1 2 2813 2823
0 2825 5 1 1 2824
0 2826 7 1 2 65409 2825
0 2827 5 1 1 2826
0 2828 7 1 2 74846 72683
0 2829 7 7 2 65147 68954
0 2830 7 5 2 57864 63451
0 2831 7 4 2 57587 76093
0 2832 7 1 2 76086 76098
0 2833 7 1 2 2828 2832
0 2834 5 1 1 2833
0 2835 7 1 2 2827 2834
0 2836 5 1 1 2835
0 2837 7 1 2 68558 2836
0 2838 5 1 1 2837
0 2839 7 14 2 58711 63581
0 2840 7 1 2 60459 76102
0 2841 7 1 2 75690 2840
0 2842 7 4 2 67507 69136
0 2843 5 2 1 76116
0 2844 7 2 2 59074 69994
0 2845 7 1 2 74173 76122
0 2846 7 1 2 76117 2845
0 2847 7 1 2 2841 2846
0 2848 5 1 1 2847
0 2849 7 1 2 2838 2848
0 2850 7 1 2 2780 2849
0 2851 5 1 1 2850
0 2852 7 1 2 58136 2851
0 2853 5 1 1 2852
0 2854 7 12 2 69343 75745
0 2855 5 6 1 76124
0 2856 7 15 2 58137 67251
0 2857 5 80 1 76142
0 2858 7 1 2 68305 76143
0 2859 5 4 1 2858
0 2860 7 5 2 57588 73460
0 2861 5 7 1 76241
0 2862 7 1 2 73798 76246
0 2863 5 4 1 2862
0 2864 7 1 2 70380 76253
0 2865 5 1 1 2864
0 2866 7 5 2 58138 73144
0 2867 5 12 1 76257
0 2868 7 5 2 57589 73791
0 2869 5 7 1 76274
0 2870 7 1 2 62843 76279
0 2871 5 3 1 2870
0 2872 7 1 2 57865 76286
0 2873 5 1 1 2872
0 2874 7 1 2 76262 2873
0 2875 5 1 1 2874
0 2876 7 1 2 65148 2875
0 2877 5 1 1 2876
0 2878 7 1 2 2865 2877
0 2879 5 1 1 2878
0 2880 7 1 2 57321 2879
0 2881 5 1 1 2880
0 2882 7 1 2 76237 2881
0 2883 5 1 1 2882
0 2884 7 1 2 71705 2883
0 2885 5 1 1 2884
0 2886 7 1 2 57866 69907
0 2887 5 2 1 2886
0 2888 7 1 2 70073 76289
0 2889 5 1 1 2888
0 2890 7 1 2 72367 2889
0 2891 5 1 1 2890
0 2892 7 1 2 76144 67875
0 2893 5 2 1 2892
0 2894 7 14 2 65149 68977
0 2895 5 2 1 76293
0 2896 7 1 2 76294 74627
0 2897 5 2 1 2896
0 2898 7 1 2 62844 76309
0 2899 5 2 1 2898
0 2900 7 1 2 70362 76311
0 2901 5 1 1 2900
0 2902 7 1 2 76291 2901
0 2903 7 2 2 2891 2902
0 2904 5 1 1 76313
0 2905 7 3 2 57867 72350
0 2906 5 1 1 76315
0 2907 7 2 2 74069 2906
0 2908 5 1 1 76318
0 2909 7 1 2 72626 76319
0 2910 5 1 1 2909
0 2911 7 1 2 58139 2910
0 2912 5 1 1 2911
0 2913 7 15 2 57868 65410
0 2914 5 10 1 76320
0 2915 7 1 2 76321 67098
0 2916 5 2 1 2915
0 2917 7 1 2 2912 76345
0 2918 5 2 1 2917
0 2919 7 1 2 74030 76347
0 2920 5 1 1 2919
0 2921 7 1 2 76314 2920
0 2922 7 1 2 2885 2921
0 2923 5 1 1 2922
0 2924 7 1 2 76125 2923
0 2925 5 1 1 2924
0 2926 7 4 2 58942 74316
0 2927 5 6 1 76349
0 2928 7 4 2 60745 76353
0 2929 5 9 1 76359
0 2930 7 3 2 57322 76363
0 2931 5 2 1 76372
0 2932 7 1 2 76373 72040
0 2933 5 1 1 2932
0 2934 7 9 2 60460 71671
0 2935 5 2 1 76377
0 2936 7 4 2 65411 76386
0 2937 5 5 1 76388
0 2938 7 1 2 74352 76389
0 2939 5 1 1 2938
0 2940 7 2 2 2933 2939
0 2941 5 2 1 76397
0 2942 7 1 2 72291 76398
0 2943 5 1 1 2942
0 2944 7 1 2 72164 2943
0 2945 5 1 1 2944
0 2946 7 4 2 63949 72041
0 2947 5 2 1 76401
0 2948 7 1 2 70185 71612
0 2949 5 1 1 2948
0 2950 7 1 2 76405 2949
0 2951 5 1 1 2950
0 2952 7 1 2 68559 68915
0 2953 5 1 1 2952
0 2954 7 1 2 65412 72540
0 2955 5 2 1 2954
0 2956 7 1 2 2953 76407
0 2957 7 1 2 2951 2956
0 2958 5 1 1 2957
0 2959 7 1 2 69344 2958
0 2960 5 1 1 2959
0 2961 7 1 2 2945 2960
0 2962 5 1 1 2961
0 2963 7 1 2 57869 2962
0 2964 5 1 1 2963
0 2965 7 3 2 63582 69137
0 2966 7 2 2 60229 74443
0 2967 7 1 2 76409 76412
0 2968 5 2 1 2967
0 2969 7 2 2 67912 72323
0 2970 5 3 1 76416
0 2971 7 1 2 76414 76418
0 2972 5 1 1 2971
0 2973 7 1 2 58140 2972
0 2974 5 1 1 2973
0 2975 7 3 2 65150 70139
0 2976 5 1 1 76421
0 2977 7 1 2 76422 69345
0 2978 5 1 1 2977
0 2979 7 1 2 2974 2978
0 2980 5 1 1 2979
0 2981 7 1 2 68560 2980
0 2982 5 1 1 2981
0 2983 7 7 2 58141 65413
0 2984 5 4 1 76424
0 2985 7 1 2 76431 71613
0 2986 5 1 1 2985
0 2987 7 3 2 59236 72013
0 2988 5 1 1 76435
0 2989 7 1 2 62845 2988
0 2990 5 2 1 2989
0 2991 7 1 2 69346 76438
0 2992 7 1 2 2986 2991
0 2993 5 1 1 2992
0 2994 7 1 2 2982 2993
0 2995 7 1 2 2964 2994
0 2996 5 1 1 2995
0 2997 7 1 2 68306 2996
0 2998 5 1 1 2997
0 2999 7 4 2 57870 71706
0 3000 5 3 1 76440
0 3001 7 1 2 71605 76441
0 3002 5 1 1 3001
0 3003 7 1 2 74388 3002
0 3004 5 1 1 3003
0 3005 7 1 2 57590 3004
0 3006 5 1 1 3005
0 3007 7 8 2 62150 60230
0 3008 5 31 1 76447
0 3009 7 10 2 63742 76448
0 3010 5 22 1 76486
0 3011 7 3 2 65414 76496
0 3012 5 4 1 76518
0 3013 7 1 2 59237 69885
0 3014 7 1 2 76519 3013
0 3015 5 1 1 3014
0 3016 7 1 2 3006 3015
0 3017 5 1 1 3016
0 3018 7 1 2 65151 3017
0 3019 5 1 1 3018
0 3020 7 1 2 74628 71985
0 3021 5 1 1 3020
0 3022 7 1 2 3019 3021
0 3023 5 1 1 3022
0 3024 7 1 2 69254 3023
0 3025 5 1 1 3024
0 3026 7 1 2 72622 76402
0 3027 5 1 1 3026
0 3028 7 1 2 69594 3027
0 3029 5 1 1 3028
0 3030 7 1 2 3025 3029
0 3031 5 1 1 3030
0 3032 7 1 2 58142 3031
0 3033 5 1 1 3032
0 3034 7 10 2 59075 69180
0 3035 5 1 1 76525
0 3036 7 2 2 69952 69569
0 3037 5 1 1 76535
0 3038 7 1 2 60231 76536
0 3039 5 1 1 3038
0 3040 7 1 2 69700 3039
0 3041 5 1 1 3040
0 3042 7 1 2 57323 3041
0 3043 5 1 1 3042
0 3044 7 1 2 72111 72302
0 3045 5 1 1 3044
0 3046 7 1 2 76419 3045
0 3047 7 1 2 3043 3046
0 3048 5 1 1 3047
0 3049 7 1 2 65415 3048
0 3050 5 1 1 3049
0 3051 7 5 2 57324 72383
0 3052 5 9 1 76537
0 3053 7 1 2 63950 76542
0 3054 5 1 1 3053
0 3055 7 1 2 69595 3054
0 3056 5 1 1 3055
0 3057 7 1 2 3050 3056
0 3058 5 1 1 3057
0 3059 7 1 2 76526 3058
0 3060 5 1 1 3059
0 3061 7 1 2 69493 76406
0 3062 5 1 1 3061
0 3063 7 1 2 72300 3062
0 3064 5 1 1 3063
0 3065 7 1 2 68719 3064
0 3066 5 1 1 3065
0 3067 7 4 2 70053 69255
0 3068 5 1 1 76551
0 3069 7 1 2 74390 76552
0 3070 5 1 1 3069
0 3071 7 1 2 70140 69596
0 3072 5 1 1 3071
0 3073 7 1 2 3070 3072
0 3074 5 1 1 3073
0 3075 7 1 2 68561 3074
0 3076 5 1 1 3075
0 3077 7 1 2 75094 72117
0 3078 5 1 1 3077
0 3079 7 1 2 68693 76415
0 3080 5 1 1 3079
0 3081 7 1 2 58143 3080
0 3082 5 1 1 3081
0 3083 7 1 2 3078 3082
0 3084 7 1 2 3076 3083
0 3085 7 1 2 3066 3084
0 3086 5 1 1 3085
0 3087 7 1 2 67823 3086
0 3088 5 1 1 3087
0 3089 7 5 2 63743 60461
0 3090 5 11 1 76555
0 3091 7 1 2 76425 68672
0 3092 5 3 1 3091
0 3093 7 6 2 57325 58144
0 3094 5 1 1 76574
0 3095 7 2 2 69513 76575
0 3096 7 1 2 72304 76580
0 3097 5 1 1 3096
0 3098 7 1 2 72123 3097
0 3099 5 1 1 3098
0 3100 7 1 2 76527 3099
0 3101 5 1 1 3100
0 3102 7 1 2 76571 3101
0 3103 5 1 1 3102
0 3104 7 1 2 76560 3103
0 3105 5 1 1 3104
0 3106 7 4 2 60102 64943
0 3107 7 3 2 74064 76582
0 3108 7 3 2 65152 69154
0 3109 7 1 2 69897 76589
0 3110 7 1 2 76586 3109
0 3111 5 1 1 3110
0 3112 7 1 2 3105 3111
0 3113 7 1 2 3088 3112
0 3114 7 1 2 3060 3113
0 3115 7 1 2 3033 3114
0 3116 7 1 2 2998 3115
0 3117 5 1 1 3116
0 3118 7 1 2 3117 75610
0 3119 5 1 1 3118
0 3120 7 1 2 2925 3119
0 3121 5 1 1 3120
0 3122 7 1 2 59429 3121
0 3123 5 1 1 3122
0 3124 7 5 2 57871 67592
0 3125 7 2 2 72321 76592
0 3126 7 2 2 58712 76597
0 3127 7 12 2 59964 60103
0 3128 7 1 2 76601 71129
0 3129 7 1 2 76599 3128
0 3130 5 1 1 3129
0 3131 7 1 2 3123 3130
0 3132 7 1 2 2853 3131
0 3133 5 1 1 3132
0 3134 7 1 2 75496 3133
0 3135 5 1 1 3134
0 3136 7 52 2 58385 59729
0 3137 5 58 1 76613
0 3138 7 40 2 76665 75566
0 3139 5 2 1 76723
0 3140 7 1 2 76126 75366
0 3141 5 1 1 3140
0 3142 7 2 2 70704 67423
0 3143 5 1 1 76765
0 3144 7 1 2 68562 75315
0 3145 5 2 1 3144
0 3146 7 1 2 76766 76767
0 3147 5 1 1 3146
0 3148 7 1 2 60232 3147
0 3149 5 1 1 3148
0 3150 7 3 2 62564 64944
0 3151 7 1 2 59238 76769
0 3152 5 1 1 3151
0 3153 7 1 2 3149 3152
0 3154 5 1 1 3153
0 3155 7 1 2 65153 3154
0 3156 5 1 1 3155
0 3157 7 5 2 60233 67252
0 3158 5 1 1 76772
0 3159 7 1 2 68563 76773
0 3160 5 2 1 3159
0 3161 7 3 2 57872 74507
0 3162 5 1 1 76779
0 3163 7 1 2 76777 3162
0 3164 5 1 1 3163
0 3165 7 1 2 68307 3164
0 3166 5 1 1 3165
0 3167 7 1 2 69181 76046
0 3168 5 3 1 3167
0 3169 7 1 2 76782 69364
0 3170 7 1 2 72536 3169
0 3171 5 1 1 3170
0 3172 7 1 2 67824 3171
0 3173 5 1 1 3172
0 3174 7 1 2 3166 3173
0 3175 7 1 2 3156 3174
0 3176 5 1 1 3175
0 3177 7 1 2 69942 3176
0 3178 5 1 1 3177
0 3179 7 6 2 64777 64945
0 3180 5 1 1 76785
0 3181 7 2 2 66667 76786
0 3182 7 1 2 74170 76791
0 3183 5 1 1 3182
0 3184 7 1 2 69225 3183
0 3185 5 1 1 3184
0 3186 7 1 2 71779 3185
0 3187 5 1 1 3186
0 3188 7 2 2 58145 76497
0 3189 5 1 1 76793
0 3190 7 1 2 65154 3189
0 3191 5 1 1 3190
0 3192 7 9 2 68214 68455
0 3193 5 16 1 76795
0 3194 7 3 2 60462 76804
0 3195 5 2 1 76820
0 3196 7 1 2 60234 76821
0 3197 5 2 1 3196
0 3198 7 3 2 58146 71850
0 3199 5 2 1 76827
0 3200 7 1 2 64946 76830
0 3201 5 1 1 3200
0 3202 7 1 2 76825 3201
0 3203 7 1 2 3191 3202
0 3204 5 1 1 3203
0 3205 7 1 2 69347 3204
0 3206 5 1 1 3205
0 3207 7 1 2 3187 3206
0 3208 7 1 2 3178 3207
0 3209 5 1 1 3208
0 3210 7 1 2 65416 3209
0 3211 5 1 1 3210
0 3212 7 6 2 67253 69597
0 3213 7 1 2 69372 76832
0 3214 5 1 1 3213
0 3215 7 1 2 57873 74317
0 3216 7 1 2 69943 3215
0 3217 5 1 1 3216
0 3218 7 1 2 69355 3217
0 3219 5 1 1 3218
0 3220 7 1 2 68720 3219
0 3221 5 1 1 3220
0 3222 7 1 2 67978 69944
0 3223 5 1 1 3222
0 3224 7 1 2 69498 3223
0 3225 7 1 2 3221 3224
0 3226 5 1 1 3225
0 3227 7 1 2 68308 3226
0 3228 5 1 1 3227
0 3229 7 3 2 69231 67427
0 3230 7 7 2 62846 59239
0 3231 5 1 1 76841
0 3232 7 1 2 67825 76842
0 3233 5 1 1 3232
0 3234 7 1 2 76528 75390
0 3235 5 1 1 3234
0 3236 7 1 2 3233 3235
0 3237 5 1 1 3236
0 3238 7 1 2 76838 3237
0 3239 5 1 1 3238
0 3240 7 1 2 76072 68673
0 3241 5 1 1 3240
0 3242 7 1 2 3239 3241
0 3243 5 1 1 3242
0 3244 7 1 2 68564 3243
0 3245 5 1 1 3244
0 3246 7 3 2 68721 67913
0 3247 7 2 2 62036 76848
0 3248 5 1 1 76851
0 3249 7 2 2 64947 66668
0 3250 7 8 2 59076 64778
0 3251 5 1 1 76855
0 3252 7 1 2 76853 76856
0 3253 7 1 2 73351 3252
0 3254 5 1 1 3253
0 3255 7 1 2 3248 3254
0 3256 5 1 1 3255
0 3257 7 1 2 65155 3256
0 3258 5 1 1 3257
0 3259 7 4 2 57326 69898
0 3260 7 1 2 69945 76863
0 3261 5 1 1 3260
0 3262 7 1 2 69701 3261
0 3263 5 1 1 3262
0 3264 7 1 2 67826 3263
0 3265 5 1 1 3264
0 3266 7 4 2 60463 66669
0 3267 7 4 2 64779 76867
0 3268 7 1 2 75042 69145
0 3269 7 1 2 76871 3268
0 3270 7 1 2 74174 3269
0 3271 5 1 1 3270
0 3272 7 1 2 72181 3271
0 3273 7 1 2 3265 3272
0 3274 7 1 2 3258 3273
0 3275 7 1 2 3245 3274
0 3276 7 1 2 3228 3275
0 3277 5 1 1 3276
0 3278 7 1 2 60746 3277
0 3279 5 1 1 3278
0 3280 7 1 2 3214 3279
0 3281 7 1 2 3211 3280
0 3282 5 1 1 3281
0 3283 7 1 2 75611 3282
0 3284 5 1 1 3283
0 3285 7 1 2 3141 3284
0 3286 5 1 1 3285
0 3287 7 1 2 76724 3286
0 3288 5 1 1 3287
0 3289 7 14 2 62847 67130
0 3290 5 4 1 76875
0 3291 7 9 2 60464 68456
0 3292 5 9 1 76893
0 3293 7 2 2 69514 72305
0 3294 7 2 2 68215 76911
0 3295 5 1 1 76913
0 3296 7 1 2 76894 76914
0 3297 5 1 1 3296
0 3298 7 1 2 75062 69598
0 3299 5 1 1 3298
0 3300 7 1 2 3297 3299
0 3301 5 1 1 3300
0 3302 7 15 2 58386 63452
0 3303 7 2 2 76915 75726
0 3304 7 1 2 3301 76930
0 3305 5 1 1 3304
0 3306 7 5 2 60104 60465
0 3307 7 2 2 68660 76932
0 3308 5 2 1 76937
0 3309 7 1 2 71022 72066
0 3310 5 1 1 3309
0 3311 7 1 2 72767 3310
0 3312 5 2 1 3311
0 3313 7 1 2 69256 76941
0 3314 5 1 1 3313
0 3315 7 1 2 76939 3314
0 3316 5 1 1 3315
0 3317 7 1 2 58387 3316
0 3318 5 1 1 3317
0 3319 7 4 2 68565 67629
0 3320 5 23 1 76943
0 3321 7 4 2 65156 76947
0 3322 5 2 1 76970
0 3323 7 1 2 76971 72118
0 3324 5 1 1 3323
0 3325 7 1 2 3318 3324
0 3326 5 1 1 3325
0 3327 7 1 2 60235 3326
0 3328 5 1 1 3327
0 3329 7 5 2 58388 60747
0 3330 5 3 1 76976
0 3331 7 9 2 63810 65417
0 3332 7 3 2 74508 76984
0 3333 5 1 1 76993
0 3334 7 1 2 76981 3333
0 3335 5 2 1 3334
0 3336 7 1 2 76996 69599
0 3337 5 1 1 3336
0 3338 7 3 2 63583 63811
0 3339 7 9 2 58389 60466
0 3340 5 5 1 77001
0 3341 7 1 2 62300 77002
0 3342 7 1 2 76998 3341
0 3343 7 1 2 72316 3342
0 3344 5 1 1 3343
0 3345 7 1 2 3337 3344
0 3346 7 1 2 3328 3345
0 3347 5 1 1 3346
0 3348 7 1 2 75612 3347
0 3349 5 1 1 3348
0 3350 7 1 2 3305 3349
0 3351 5 1 1 3350
0 3352 7 1 2 76876 3351
0 3353 5 1 1 3352
0 3354 7 6 2 61895 76602
0 3355 7 5 2 58390 58840
0 3356 5 1 1 77021
0 3357 7 12 2 63812 60748
0 3358 5 4 1 77026
0 3359 7 1 2 58713 77027
0 3360 7 1 2 77022 3359
0 3361 7 1 2 77015 3360
0 3362 7 6 2 60467 76157
0 3363 5 1 1 77042
0 3364 7 3 2 62037 70600
0 3365 7 1 2 77043 77048
0 3366 7 1 2 3361 3365
0 3367 5 1 1 3366
0 3368 7 1 2 3353 3367
0 3369 5 1 1 3368
0 3370 7 1 2 59730 3369
0 3371 5 1 1 3370
0 3372 7 6 2 65418 69407
0 3373 5 22 1 77051
0 3374 7 1 2 77057 72620
0 3375 5 2 1 3374
0 3376 7 3 2 58943 69373
0 3377 5 1 1 77081
0 3378 7 1 2 65419 77082
0 3379 5 1 1 3378
0 3380 7 1 2 77079 3379
0 3381 5 2 1 3380
0 3382 7 2 2 67630 77084
0 3383 5 1 1 77086
0 3384 7 23 2 60236 68818
0 3385 5 8 1 77088
0 3386 7 47 2 68566 77111
0 3387 5 3 1 77119
0 3388 7 2 2 68309 77120
0 3389 5 3 1 77169
0 3390 7 6 2 67713 77171
0 3391 5 4 1 77174
0 3392 7 1 2 65157 72271
0 3393 5 1 1 3392
0 3394 7 1 2 77175 3393
0 3395 5 3 1 3394
0 3396 7 2 2 60749 77184
0 3397 5 2 1 77187
0 3398 7 6 2 60237 70667
0 3399 7 1 2 76805 77191
0 3400 5 1 1 3399
0 3401 7 1 2 77189 3400
0 3402 5 1 1 3401
0 3403 7 1 2 59240 3402
0 3404 5 1 1 3403
0 3405 7 1 2 3383 3404
0 3406 5 2 1 3405
0 3407 7 1 2 77197 75613
0 3408 5 1 1 3407
0 3409 7 2 2 68916 74555
0 3410 5 1 1 77199
0 3411 7 10 2 60468 66549
0 3412 7 3 2 77201 74465
0 3413 7 9 2 57591 63453
0 3414 7 1 2 77211 77214
0 3415 7 1 2 77200 3414
0 3416 5 1 1 3415
0 3417 7 1 2 3408 3416
0 3418 5 1 1 3417
0 3419 7 1 2 57874 3418
0 3420 5 1 1 3419
0 3421 7 2 2 59241 77087
0 3422 5 1 1 77223
0 3423 7 1 2 77224 75614
0 3424 5 1 1 3423
0 3425 7 1 2 3420 3424
0 3426 5 1 1 3425
0 3427 7 15 2 58147 64443
0 3428 7 1 2 77225 68674
0 3429 7 1 2 3426 3428
0 3430 5 1 1 3429
0 3431 7 1 2 3371 3430
0 3432 7 1 2 3288 3431
0 3433 5 1 1 3432
0 3434 7 1 2 64146 3433
0 3435 5 1 1 3434
0 3436 7 4 2 62565 58714
0 3437 7 2 2 75949 77240
0 3438 5 1 1 77244
0 3439 7 1 2 77058 77245
0 3440 5 1 1 3439
0 3441 7 32 2 66550 66743
0 3442 7 2 2 70902 77246
0 3443 5 1 1 77278
0 3444 7 1 2 3440 3443
0 3445 5 1 1 3444
0 3446 7 1 2 63951 3445
0 3447 5 1 1 3446
0 3448 7 4 2 64666 77202
0 3449 7 2 2 77280 75368
0 3450 5 2 1 77284
0 3451 7 1 2 76158 77285
0 3452 5 1 1 3451
0 3453 7 4 2 62566 66551
0 3454 7 4 2 66744 77288
0 3455 5 1 1 77292
0 3456 7 1 2 76263 77293
0 3457 5 1 1 3456
0 3458 7 3 2 63813 59965
0 3459 7 5 2 58715 77296
0 3460 7 1 2 60469 68929
0 3461 7 1 2 77299 3460
0 3462 5 1 1 3461
0 3463 7 1 2 3457 3462
0 3464 7 1 2 3452 3463
0 3465 5 1 1 3464
0 3466 7 1 2 70601 3465
0 3467 5 1 1 3466
0 3468 7 1 2 3447 3467
0 3469 5 1 1 3468
0 3470 7 1 2 59430 3469
0 3471 5 1 1 3470
0 3472 7 2 2 74521 69856
0 3473 5 9 1 77304
0 3474 7 4 2 63814 77306
0 3475 5 4 1 77315
0 3476 7 1 2 66811 74288
0 3477 7 1 2 77316 3476
0 3478 5 1 1 3477
0 3479 7 4 2 72464 75615
0 3480 5 1 1 77323
0 3481 7 2 2 60238 77324
0 3482 5 1 1 77327
0 3483 7 1 2 70602 77328
0 3484 5 1 1 3483
0 3485 7 1 2 3478 3484
0 3486 5 1 1 3485
0 3487 7 1 2 76159 3486
0 3488 5 1 1 3487
0 3489 7 1 2 3471 3488
0 3490 5 1 1 3489
0 3491 7 1 2 69600 3490
0 3492 5 1 1 3491
0 3493 7 2 2 66812 74435
0 3494 5 2 1 77329
0 3495 7 1 2 77286 77331
0 3496 5 1 1 3495
0 3497 7 1 2 62567 3496
0 3498 5 1 1 3497
0 3499 7 1 2 77300 68712
0 3500 5 1 1 3499
0 3501 7 1 2 3498 3500
0 3502 5 1 1 3501
0 3503 7 1 2 71023 3502
0 3504 5 1 1 3503
0 3505 7 2 2 58716 75122
0 3506 7 1 2 59966 72714
0 3507 7 1 2 68703 3506
0 3508 7 1 2 77333 3507
0 3509 5 1 1 3508
0 3510 7 1 2 3504 3509
0 3511 5 1 1 3510
0 3512 7 16 2 63952 59431
0 3513 7 2 2 71053 72317
0 3514 5 1 1 77351
0 3515 7 1 2 77335 77352
0 3516 7 1 2 3511 3515
0 3517 5 1 1 3516
0 3518 7 1 2 3492 3517
0 3519 5 1 1 3518
0 3520 7 1 2 76725 3519
0 3521 5 1 1 3520
0 3522 7 10 2 64444 64948
0 3523 5 3 1 77353
0 3524 7 1 2 77354 74233
0 3525 7 1 2 76553 3524
0 3526 5 2 1 3525
0 3527 7 8 2 59731 60105
0 3528 7 4 2 60750 62038
0 3529 7 1 2 60470 77376
0 3530 7 2 2 77368 3529
0 3531 7 5 2 58841 63953
0 3532 7 3 2 63815 77382
0 3533 7 11 2 62151 62848
0 3534 5 2 1 77390
0 3535 7 5 2 63744 77391
0 3536 5 1 1 77403
0 3537 7 1 2 77387 77404
0 3538 7 1 2 77380 3537
0 3539 5 1 1 3538
0 3540 7 1 2 77366 3539
0 3541 5 1 1 3540
0 3542 7 1 2 62568 3541
0 3543 5 1 1 3542
0 3544 7 24 2 62569 62849
0 3545 5 3 1 77408
0 3546 7 1 2 77409 77388
0 3547 7 1 2 77381 3546
0 3548 5 1 1 3547
0 3549 7 1 2 77367 3548
0 3550 5 1 1 3549
0 3551 7 1 2 62301 3550
0 3552 5 1 1 3551
0 3553 7 1 2 3543 3552
0 3554 5 1 1 3553
0 3555 7 1 2 59432 75969
0 3556 7 1 2 3554 3555
0 3557 5 1 1 3556
0 3558 7 1 2 61163 3557
0 3559 7 1 2 3521 3558
0 3560 7 1 2 3435 3559
0 3561 7 1 2 3135 3560
0 3562 5 1 1 3561
0 3563 7 4 2 57592 69982
0 3564 5 1 1 77435
0 3565 7 5 2 58944 72813
0 3566 7 2 2 77436 77439
0 3567 5 1 1 77444
0 3568 7 1 2 64949 77445
0 3569 5 1 1 3568
0 3570 7 1 2 74607 74958
0 3571 7 1 2 71049 3570
0 3572 5 1 1 3571
0 3573 7 1 2 59433 3572
0 3574 5 1 1 3573
0 3575 7 1 2 3569 3574
0 3576 5 1 1 3575
0 3577 7 1 2 60751 3576
0 3578 5 1 1 3577
0 3579 7 8 2 62570 59434
0 3580 5 1 1 77446
0 3581 7 1 2 77447 70987
0 3582 5 1 1 3581
0 3583 7 1 2 3578 3582
0 3584 5 1 1 3583
0 3585 7 1 2 75616 3584
0 3586 5 1 1 3585
0 3587 7 23 2 62302 62571
0 3588 5 1 1 77454
0 3589 7 8 2 62152 77455
0 3590 7 1 2 71986 77203
0 3591 7 2 2 77477 3590
0 3592 7 10 2 63745 63816
0 3593 5 2 1 77487
0 3594 7 2 2 59242 77488
0 3595 7 8 2 59435 64667
0 3596 5 1 1 77501
0 3597 7 5 2 63454 77502
0 3598 7 1 2 77499 77509
0 3599 7 1 2 77485 3598
0 3600 5 1 1 3599
0 3601 7 1 2 3586 3600
0 3602 5 1 1 3601
0 3603 7 1 2 58148 3602
0 3604 5 1 1 3603
0 3605 7 8 2 57875 64147
0 3606 5 1 1 77514
0 3607 7 2 2 63817 70087
0 3608 5 2 1 77522
0 3609 7 6 2 76498 77524
0 3610 5 3 1 77526
0 3611 7 1 2 77527 74780
0 3612 5 1 1 3611
0 3613 7 1 2 74509 68901
0 3614 5 1 1 3613
0 3615 7 1 2 3612 3614
0 3616 5 1 1 3615
0 3617 7 1 2 57593 3616
0 3618 5 1 1 3617
0 3619 7 3 2 59077 74318
0 3620 5 6 1 77535
0 3621 7 4 2 62850 58945
0 3622 7 2 2 57327 77544
0 3623 7 1 2 77536 77548
0 3624 5 1 1 3623
0 3625 7 1 2 3618 3624
0 3626 5 1 1 3625
0 3627 7 1 2 77515 3626
0 3628 5 1 1 3627
0 3629 7 7 2 74937 72188
0 3630 5 2 1 77550
0 3631 7 2 2 73752 74597
0 3632 5 1 1 77559
0 3633 7 1 2 77551 77560
0 3634 5 1 1 3633
0 3635 7 1 2 3628 3634
0 3636 5 1 1 3635
0 3637 7 3 2 70141 75970
0 3638 5 1 1 77561
0 3639 7 1 2 3636 77562
0 3640 5 1 1 3639
0 3641 7 1 2 3604 3640
0 3642 5 1 1 3641
0 3643 7 1 2 75497 3642
0 3644 5 1 1 3643
0 3645 7 3 2 64148 74319
0 3646 5 3 1 77564
0 3647 7 3 2 63954 74320
0 3648 5 1 1 77570
0 3649 7 4 2 59436 69374
0 3650 5 2 1 77573
0 3651 7 1 2 3648 77577
0 3652 5 1 1 3651
0 3653 7 1 2 62572 3652
0 3654 5 1 1 3653
0 3655 7 1 2 77567 3654
0 3656 5 1 1 3655
0 3657 7 1 2 68457 3656
0 3658 5 1 1 3657
0 3659 7 1 2 60471 69306
0 3660 5 1 1 3659
0 3661 7 1 2 3658 3660
0 3662 5 1 1 3661
0 3663 7 1 2 62303 3662
0 3664 5 1 1 3663
0 3665 7 17 2 63955 64149
0 3666 5 1 1 77579
0 3667 7 1 2 77580 71047
0 3668 5 1 1 3667
0 3669 7 1 2 3664 3668
0 3670 5 1 1 3669
0 3671 7 1 2 63818 3670
0 3672 5 1 1 3671
0 3673 7 1 2 60472 668
0 3674 5 1 1 3673
0 3675 7 4 2 65158 67131
0 3676 5 1 1 77596
0 3677 7 2 2 59078 77597
0 3678 5 1 1 77600
0 3679 7 1 2 3674 3678
0 3680 5 1 1 3679
0 3681 7 1 2 64150 3680
0 3682 5 1 1 3681
0 3683 7 1 2 60752 3682
0 3684 7 1 2 3672 3683
0 3685 5 1 1 3684
0 3686 7 9 2 62573 64151
0 3687 5 3 1 77602
0 3688 7 7 2 63746 63956
0 3689 5 2 1 77614
0 3690 7 1 2 62153 77615
0 3691 5 2 1 3690
0 3692 7 1 2 70955 77623
0 3693 5 1 1 3692
0 3694 7 1 2 77603 3693
0 3695 5 1 1 3694
0 3696 7 1 2 65420 3695
0 3697 5 1 1 3696
0 3698 7 1 2 62851 3697
0 3699 7 1 2 3685 3698
0 3700 5 1 1 3699
0 3701 7 2 2 68458 75097
0 3702 5 1 1 77625
0 3703 7 3 2 68216 77604
0 3704 7 1 2 77626 77627
0 3705 7 1 2 75116 3704
0 3706 5 1 1 3705
0 3707 7 1 2 3700 3706
0 3708 5 1 1 3707
0 3709 7 1 2 75617 3708
0 3710 5 1 1 3709
0 3711 7 6 2 64152 64668
0 3712 7 6 2 62852 63455
0 3713 7 2 2 77630 77636
0 3714 7 1 2 77500 77642
0 3715 7 1 2 77486 3714
0 3716 5 1 1 3715
0 3717 7 1 2 3710 3716
0 3718 5 1 1 3717
0 3719 7 1 2 76726 3718
0 3720 5 1 1 3719
0 3721 7 1 2 3644 3720
0 3722 5 1 1 3721
0 3723 7 1 2 69257 3722
0 3724 5 1 1 3723
0 3725 7 1 2 59437 74881
0 3726 5 2 1 3725
0 3727 7 8 2 57876 68310
0 3728 5 29 1 77646
0 3729 7 1 2 75845 77647
0 3730 5 4 1 3729
0 3731 7 2 2 62853 77683
0 3732 5 2 1 77687
0 3733 7 2 2 57594 73892
0 3734 5 2 1 77691
0 3735 7 4 2 74865 77693
0 3736 5 4 1 77695
0 3737 7 1 2 77121 77699
0 3738 5 1 1 3737
0 3739 7 1 2 77688 3738
0 3740 5 1 1 3739
0 3741 7 1 2 64153 3740
0 3742 5 1 1 3741
0 3743 7 1 2 77644 3742
0 3744 5 1 1 3743
0 3745 7 1 2 65421 3744
0 3746 5 1 1 3745
0 3747 7 8 2 58149 60473
0 3748 5 9 1 77703
0 3749 7 2 2 60753 77180
0 3750 5 1 1 77720
0 3751 7 1 2 77704 77721
0 3752 5 1 1 3751
0 3753 7 4 2 70586 77112
0 3754 5 14 1 77722
0 3755 7 1 2 69983 73396
0 3756 7 1 2 77723 3755
0 3757 5 1 1 3756
0 3758 7 1 2 3752 3757
0 3759 7 1 2 3746 3758
0 3760 5 1 1 3759
0 3761 7 1 2 59243 3760
0 3762 5 1 1 3761
0 3763 7 1 2 59079 69729
0 3764 5 2 1 3763
0 3765 7 2 2 60754 74576
0 3766 5 1 1 77742
0 3767 7 1 2 74102 3766
0 3768 5 3 1 3767
0 3769 7 1 2 57877 77744
0 3770 5 1 1 3769
0 3771 7 1 2 77740 3770
0 3772 5 1 1 3771
0 3773 7 1 2 58150 3772
0 3774 5 1 1 3773
0 3775 7 3 2 59438 70276
0 3776 5 2 1 77747
0 3777 7 1 2 70695 77748
0 3778 5 1 1 3777
0 3779 7 1 2 3774 3778
0 3780 5 1 1 3779
0 3781 7 1 2 57595 3780
0 3782 5 1 1 3781
0 3783 7 2 2 70696 70343
0 3784 5 1 1 77752
0 3785 7 1 2 58151 67827
0 3786 5 2 1 3785
0 3787 7 1 2 3784 77754
0 3788 5 1 1 3787
0 3789 7 1 2 74089 3788
0 3790 5 1 1 3789
0 3791 7 3 2 68311 71460
0 3792 5 2 1 77756
0 3793 7 11 2 57878 60755
0 3794 5 1 1 77761
0 3795 7 1 2 60474 77762
0 3796 5 1 1 3795
0 3797 7 1 2 69750 3796
0 3798 5 1 1 3797
0 3799 7 1 2 77757 3798
0 3800 5 1 1 3799
0 3801 7 1 2 3790 3800
0 3802 5 1 1 3801
0 3803 7 1 2 77122 3802
0 3804 5 1 1 3803
0 3805 7 2 2 70697 70054
0 3806 7 1 2 64154 77772
0 3807 5 1 1 3806
0 3808 7 1 2 3804 3807
0 3809 7 1 2 3782 3808
0 3810 7 1 2 3762 3809
0 3811 5 1 1 3810
0 3812 7 1 2 75498 3811
0 3813 5 1 1 3812
0 3814 7 12 2 58152 63140
0 3815 5 2 1 77774
0 3816 7 4 2 77775 73709
0 3817 5 2 1 77788
0 3818 7 14 2 63141 59732
0 3819 5 7 1 77794
0 3820 7 14 2 58391 64445
0 3821 5 8 1 77815
0 3822 7 7 2 77808 77829
0 3823 5 42 1 77837
0 3824 7 13 2 63819 64155
0 3825 5 1 1 77886
0 3826 7 4 2 60475 77887
0 3827 5 2 1 77899
0 3828 7 2 2 77844 77900
0 3829 5 1 1 77905
0 3830 7 1 2 62574 77906
0 3831 5 1 1 3830
0 3832 7 1 2 77792 3831
0 3833 5 1 1 3832
0 3834 7 1 2 70705 77789
0 3835 5 1 1 3834
0 3836 7 1 2 70587 3835
0 3837 5 1 1 3836
0 3838 7 1 2 70186 3837
0 3839 7 1 2 3833 3838
0 3840 5 1 1 3839
0 3841 7 5 2 62575 77581
0 3842 5 4 1 77907
0 3843 7 1 2 77912 75066
0 3844 5 1 1 3843
0 3845 7 5 2 62854 73583
0 3846 5 1 1 77916
0 3847 7 1 2 77845 77917
0 3848 7 1 2 3844 3847
0 3849 5 1 1 3848
0 3850 7 1 2 3840 3849
0 3851 7 1 2 3813 3850
0 3852 5 1 1 3851
0 3853 7 1 2 77247 3852
0 3854 5 1 1 3853
0 3855 7 1 2 62855 76948
0 3856 5 3 1 3855
0 3857 7 1 2 67254 77921
0 3858 5 2 1 3857
0 3859 7 2 2 70381 68312
0 3860 5 4 1 77926
0 3861 7 2 2 70382 68567
0 3862 5 1 1 77932
0 3863 7 1 2 77928 3862
0 3864 7 2 2 77924 3863
0 3865 5 2 1 77934
0 3866 7 1 2 60476 77936
0 3867 5 1 1 3866
0 3868 7 1 2 59439 70744
0 3869 7 1 2 70858 3868
0 3870 5 1 1 3869
0 3871 7 1 2 3867 3870
0 3872 5 1 1 3871
0 3873 7 1 2 65422 3872
0 3874 5 1 1 3873
0 3875 7 3 2 60477 71141
0 3876 5 1 1 77938
0 3877 7 1 2 64446 3876
0 3878 7 1 2 3874 3877
0 3879 5 1 1 3878
0 3880 7 11 2 63820 70277
0 3881 5 11 1 77941
0 3882 7 1 2 59440 77952
0 3883 5 8 1 3882
0 3884 7 1 2 62856 77963
0 3885 5 1 1 3884
0 3886 7 33 2 64156 60756
0 3887 5 12 1 77971
0 3888 7 7 2 71790 77972
0 3889 5 4 1 78016
0 3890 7 2 2 3885 78023
0 3891 5 5 1 78027
0 3892 7 1 2 71142 77953
0 3893 5 2 1 3892
0 3894 7 1 2 67132 78034
0 3895 5 1 1 3894
0 3896 7 1 2 78028 3895
0 3897 5 3 1 3896
0 3898 7 1 2 70603 78036
0 3899 5 1 1 3898
0 3900 7 12 2 60757 71238
0 3901 5 2 1 78039
0 3902 7 5 2 62576 60478
0 3903 5 5 1 78053
0 3904 7 1 2 70015 78058
0 3905 5 4 1 3904
0 3906 7 1 2 78040 78063
0 3907 5 1 1 3906
0 3908 7 1 2 59733 3907
0 3909 7 1 2 3899 3908
0 3910 5 1 1 3909
0 3911 7 1 2 63142 3910
0 3912 7 1 2 3879 3911
0 3913 5 1 1 3912
0 3914 7 24 2 64157 59734
0 3915 5 2 1 78067
0 3916 7 1 2 77942 78068
0 3917 5 2 1 3916
0 3918 7 8 2 64447 65159
0 3919 5 1 1 78095
0 3920 7 1 2 74118 78096
0 3921 5 1 1 3920
0 3922 7 1 2 78093 3921
0 3923 5 1 1 3922
0 3924 7 1 2 62857 3923
0 3925 5 1 1 3924
0 3926 7 2 2 58392 77964
0 3927 5 2 1 78103
0 3928 7 1 2 64448 78104
0 3929 5 1 1 3928
0 3930 7 1 2 3925 3929
0 3931 5 1 1 3930
0 3932 7 1 2 67133 3931
0 3933 5 1 1 3932
0 3934 7 1 2 77816 78029
0 3935 5 1 1 3934
0 3936 7 1 2 3933 3935
0 3937 5 1 1 3936
0 3938 7 1 2 70604 3937
0 3939 5 1 1 3938
0 3940 7 2 2 77973 77003
0 3941 5 1 1 78107
0 3942 7 1 2 73753 76985
0 3943 5 2 1 3942
0 3944 7 1 2 77010 78109
0 3945 5 3 1 3944
0 3946 7 1 2 72772 78111
0 3947 5 1 1 3946
0 3948 7 1 2 3941 3947
0 3949 5 1 1 3948
0 3950 7 1 2 62577 3949
0 3951 5 1 1 3950
0 3952 7 7 2 62304 58393
0 3953 7 3 2 60758 77582
0 3954 5 1 1 78121
0 3955 7 1 2 78114 78122
0 3956 5 1 1 3955
0 3957 7 1 2 3951 3956
0 3958 5 1 1 3957
0 3959 7 1 2 64449 3958
0 3960 5 1 1 3959
0 3961 7 1 2 3939 3960
0 3962 7 1 2 3913 3961
0 3963 5 1 1 3962
0 3964 7 1 2 60239 3963
0 3965 5 1 1 3964
0 3966 7 4 2 65423 71791
0 3967 7 1 2 69811 78124
0 3968 5 1 1 3967
0 3969 7 1 2 76982 3968
0 3970 5 2 1 3969
0 3971 7 1 2 62858 78128
0 3972 5 1 1 3971
0 3973 7 8 2 65424 68313
0 3974 5 12 1 78130
0 3975 7 1 2 75428 78138
0 3976 5 1 1 3975
0 3977 7 1 2 3972 3976
0 3978 5 1 1 3977
0 3979 7 1 2 63957 3978
0 3980 5 1 1 3979
0 3981 7 18 2 63143 59441
0 3982 5 11 1 78150
0 3983 7 1 2 78151 77052
0 3984 5 1 1 3983
0 3985 7 1 2 3980 3984
0 3986 5 1 1 3985
0 3987 7 1 2 64450 3986
0 3988 5 1 1 3987
0 3989 7 3 2 63958 71239
0 3990 5 2 1 78179
0 3991 7 1 2 77795 78180
0 3992 7 1 2 78139 3991
0 3993 5 1 1 3992
0 3994 7 1 2 3988 3993
0 3995 5 1 1 3994
0 3996 7 1 2 62578 3995
0 3997 5 1 1 3996
0 3998 7 1 2 71382 72009
0 3999 5 3 1 3998
0 4000 7 3 2 62305 71672
0 4001 5 5 1 78187
0 4002 7 2 2 57879 78190
0 4003 5 6 1 78195
0 4004 7 7 2 57596 68978
0 4005 5 8 1 78203
0 4006 7 1 2 62579 78210
0 4007 5 5 1 4006
0 4008 7 1 2 57328 78218
0 4009 5 3 1 4008
0 4010 7 4 2 78197 78223
0 4011 5 5 1 78226
0 4012 7 1 2 64158 69977
0 4013 5 1 1 4012
0 4014 7 1 2 58153 4013
0 4015 5 1 1 4014
0 4016 7 15 2 63959 60479
0 4017 5 7 1 78235
0 4018 7 1 2 57880 78250
0 4019 5 1 1 4018
0 4020 7 2 2 73821 4019
0 4021 7 1 2 4015 78257
0 4022 5 1 1 4021
0 4023 7 1 2 71461 4022
0 4024 5 1 1 4023
0 4025 7 1 2 78227 4024
0 4026 5 1 1 4025
0 4027 7 1 2 78184 4026
0 4028 5 1 1 4027
0 4029 7 2 2 64159 70366
0 4030 5 17 1 78259
0 4031 7 3 2 57597 71707
0 4032 5 20 1 78278
0 4033 7 5 2 62306 69018
0 4034 5 27 1 78301
0 4035 7 6 2 57329 78306
0 4036 5 4 1 78333
0 4037 7 12 2 78281 78339
0 4038 5 13 1 78343
0 4039 7 2 2 71851 78355
0 4040 5 2 1 78368
0 4041 7 1 2 78261 78369
0 4042 5 1 1 4041
0 4043 7 5 2 74803 72814
0 4044 5 1 1 78372
0 4045 7 1 2 62859 4044
0 4046 5 1 1 4045
0 4047 7 1 2 64950 4046
0 4048 5 1 1 4047
0 4049 7 1 2 71462 70932
0 4050 5 2 1 4049
0 4051 7 4 2 58946 71463
0 4052 5 3 1 78379
0 4053 7 1 2 78377 78383
0 4054 7 1 2 4048 4053
0 4055 5 1 1 4054
0 4056 7 1 2 72230 4055
0 4057 5 1 1 4056
0 4058 7 1 2 4042 4057
0 4059 7 1 2 4028 4058
0 4060 5 3 1 4059
0 4061 7 5 2 60759 75499
0 4062 7 1 2 78386 78389
0 4063 5 1 1 4062
0 4064 7 4 2 63144 73541
0 4065 5 2 1 78394
0 4066 7 2 2 75316 74215
0 4067 5 1 1 78400
0 4068 7 1 2 68979 78401
0 4069 5 2 1 4068
0 4070 7 1 2 67900 78402
0 4071 5 1 1 4070
0 4072 7 1 2 69408 4071
0 4073 5 1 1 4072
0 4074 7 3 2 60480 75180
0 4075 5 7 1 78404
0 4076 7 3 2 68314 76499
0 4077 5 4 1 78414
0 4078 7 2 2 78407 78415
0 4079 5 4 1 78421
0 4080 7 1 2 67255 78422
0 4081 5 2 1 4080
0 4082 7 1 2 4073 78427
0 4083 5 3 1 4082
0 4084 7 1 2 78395 78429
0 4085 5 1 1 4084
0 4086 7 4 2 62860 72067
0 4087 5 5 1 78432
0 4088 7 1 2 76727 78433
0 4089 5 1 1 4088
0 4090 7 1 2 4085 4089
0 4091 5 1 1 4090
0 4092 7 1 2 64160 4091
0 4093 5 1 1 4092
0 4094 7 1 2 4063 4093
0 4095 7 1 2 3997 4094
0 4096 7 1 2 3965 4095
0 4097 5 1 1 4096
0 4098 7 1 2 75618 4097
0 4099 5 1 1 4098
0 4100 7 1 2 3854 4099
0 4101 5 1 1 4100
0 4102 7 1 2 69601 4101
0 4103 5 1 1 4102
0 4104 7 1 2 65783 4103
0 4105 7 1 2 3724 4104
0 4106 5 1 1 4105
0 4107 7 1 2 3562 4106
0 4108 5 1 1 4107
0 4109 7 1 2 61504 4108
0 4110 7 1 2 2693 4109
0 4111 7 1 2 1816 4110
0 4112 5 1 1 4111
0 4113 7 12 2 62861 60481
0 4114 5 3 1 78441
0 4115 7 7 2 70019 77456
0 4116 5 3 1 78456
0 4117 7 1 2 78442 78463
0 4118 5 1 1 4117
0 4119 7 3 2 76160 76949
0 4120 5 2 1 78466
0 4121 7 1 2 65160 78467
0 4122 5 1 1 4121
0 4123 7 1 2 4118 4122
0 4124 5 1 1 4123
0 4125 7 1 2 65784 4124
0 4126 5 1 1 4125
0 4127 7 2 2 68722 73195
0 4128 5 1 1 78471
0 4129 7 1 2 75297 78472
0 4130 5 1 1 4129
0 4131 7 1 2 4126 4130
0 4132 5 1 1 4131
0 4133 7 1 2 64161 4132
0 4134 5 1 1 4133
0 4135 7 22 2 60482 61164
0 4136 5 1 1 78473
0 4137 7 11 2 62862 59442
0 4138 5 4 1 78495
0 4139 7 2 2 78474 78496
0 4140 5 1 1 78510
0 4141 7 3 2 63960 70605
0 4142 5 2 1 78512
0 4143 7 1 2 73037 78513
0 4144 5 1 1 4143
0 4145 7 16 2 59443 60483
0 4146 5 5 1 78517
0 4147 7 2 2 63821 78518
0 4148 5 2 1 78538
0 4149 7 2 2 63961 73560
0 4150 5 1 1 78542
0 4151 7 1 2 78540 4150
0 4152 5 1 1 4151
0 4153 7 1 2 70606 4152
0 4154 5 1 1 4153
0 4155 7 7 2 63962 65161
0 4156 5 1 1 78544
0 4157 7 4 2 63822 65785
0 4158 7 1 2 78545 78551
0 4159 5 1 1 4158
0 4160 7 1 2 71024 78519
0 4161 5 1 1 4160
0 4162 7 1 2 4159 4161
0 4163 7 1 2 4154 4162
0 4164 5 1 1 4163
0 4165 7 1 2 62863 4164
0 4166 5 1 1 4165
0 4167 7 1 2 4144 4166
0 4168 5 1 1 4167
0 4169 7 1 2 62580 4168
0 4170 5 1 1 4169
0 4171 7 1 2 4140 4170
0 4172 7 1 2 4134 4171
0 4173 5 1 1 4172
0 4174 7 1 2 60760 4173
0 4175 5 1 1 4174
0 4176 7 1 2 71240 74866
0 4177 7 2 2 72945 4176
0 4178 5 2 1 78555
0 4179 7 6 2 62581 71792
0 4180 5 3 1 78559
0 4181 7 2 2 77336 78560
0 4182 5 1 1 78568
0 4183 7 1 2 78557 4182
0 4184 5 1 1 4183
0 4185 7 1 2 70607 4184
0 4186 5 1 1 4185
0 4187 7 1 2 70653 77888
0 4188 5 1 1 4187
0 4189 7 1 2 4186 4188
0 4190 5 1 1 4189
0 4191 7 1 2 61165 4190
0 4192 5 1 1 4191
0 4193 7 5 2 60484 71383
0 4194 5 2 1 78570
0 4195 7 5 2 62307 64162
0 4196 5 1 1 78577
0 4197 7 1 2 78453 4196
0 4198 5 1 1 4197
0 4199 7 1 2 67134 4198
0 4200 5 1 1 4199
0 4201 7 1 2 78575 4200
0 4202 5 1 1 4201
0 4203 7 1 2 68459 4202
0 4204 5 1 1 4203
0 4205 7 1 2 67559 77918
0 4206 5 1 1 4205
0 4207 7 1 2 4204 4206
0 4208 5 1 1 4207
0 4209 7 1 2 65786 76986
0 4210 7 1 2 4208 4209
0 4211 5 1 1 4210
0 4212 7 1 2 4192 4211
0 4213 7 1 2 4175 4212
0 4214 5 1 1 4213
0 4215 7 1 2 60240 4214
0 4216 5 1 1 4215
0 4217 7 1 2 67811 76543
0 4218 5 2 1 4217
0 4219 7 1 2 73145 78582
0 4220 5 1 1 4219
0 4221 7 1 2 72541 68917
0 4222 5 1 1 4221
0 4223 7 1 2 4220 4222
0 4224 5 1 1 4223
0 4225 7 1 2 62864 4224
0 4226 5 1 1 4225
0 4227 7 2 2 76950 1980
0 4228 5 3 1 78584
0 4229 7 3 2 65162 77113
0 4230 5 8 1 78589
0 4231 7 2 2 78586 78590
0 4232 5 1 1 78600
0 4233 7 1 2 74633 4232
0 4234 5 1 1 4233
0 4235 7 1 2 73102 4234
0 4236 5 1 1 4235
0 4237 7 4 2 62582 73103
0 4238 5 15 1 78602
0 4239 7 3 2 68315 78606
0 4240 5 2 1 78621
0 4241 7 2 2 76264 78622
0 4242 7 15 2 64951 68568
0 4243 5 7 1 78628
0 4244 7 2 2 60485 78643
0 4245 5 4 1 78650
0 4246 7 1 2 78626 78652
0 4247 5 1 1 4246
0 4248 7 1 2 4236 4247
0 4249 7 1 2 4226 4248
0 4250 5 1 1 4249
0 4251 7 1 2 64163 4250
0 4252 5 1 1 4251
0 4253 7 2 2 71143 73146
0 4254 5 2 1 78656
0 4255 7 2 2 62583 78658
0 4256 5 1 1 78660
0 4257 7 1 2 71793 72946
0 4258 7 1 2 78661 4257
0 4259 5 1 1 4258
0 4260 7 1 2 73104 78497
0 4261 5 1 1 4260
0 4262 7 1 2 61166 4261
0 4263 7 1 2 4259 4262
0 4264 7 1 2 4252 4263
0 4265 5 1 1 4264
0 4266 7 5 2 67135 71241
0 4267 5 2 1 78662
0 4268 7 3 2 62865 69730
0 4269 5 2 1 78669
0 4270 7 17 2 64952 60761
0 4271 5 2 1 78674
0 4272 7 1 2 71794 78675
0 4273 5 2 1 4272
0 4274 7 1 2 78672 78693
0 4275 5 1 1 4274
0 4276 7 1 2 78663 4275
0 4277 5 1 1 4276
0 4278 7 7 2 62866 64953
0 4279 7 1 2 78017 78695
0 4280 5 1 1 4279
0 4281 7 1 2 65787 4280
0 4282 7 1 2 4277 4281
0 4283 5 1 1 4282
0 4284 7 1 2 4265 4283
0 4285 5 1 1 4284
0 4286 7 2 2 4216 4285
0 4287 5 1 1 78702
0 4288 7 1 2 59735 78703
0 4289 5 1 1 4288
0 4290 7 1 2 77648 70996
0 4291 5 2 1 4290
0 4292 7 1 2 65425 78704
0 4293 5 2 1 4292
0 4294 7 2 2 68217 77616
0 4295 7 1 2 74938 78708
0 4296 5 1 1 4295
0 4297 7 1 2 60762 4296
0 4298 5 1 1 4297
0 4299 7 1 2 78706 4298
0 4300 5 1 1 4299
0 4301 7 1 2 58154 4300
0 4302 5 1 1 4301
0 4303 7 4 2 60763 68569
0 4304 5 1 1 78710
0 4305 7 1 2 76529 78711
0 4306 5 1 1 4305
0 4307 7 1 2 4302 4306
0 4308 5 1 1 4307
0 4309 7 1 2 60486 4308
0 4310 5 1 1 4309
0 4311 7 6 2 62308 65426
0 4312 7 2 2 70020 78714
0 4313 5 1 1 78720
0 4314 7 1 2 69953 78721
0 4315 5 1 1 4314
0 4316 7 3 2 58155 70313
0 4317 5 3 1 78722
0 4318 7 2 2 70187 78723
0 4319 5 1 1 78728
0 4320 7 1 2 65163 71090
0 4321 5 1 1 4320
0 4322 7 1 2 4319 4321
0 4323 5 1 1 4322
0 4324 7 1 2 76951 4323
0 4325 5 1 1 4324
0 4326 7 1 2 4315 4325
0 4327 7 1 2 4310 4326
0 4328 5 1 1 4327
0 4329 7 1 2 60241 4328
0 4330 5 1 1 4329
0 4331 7 7 2 57598 73851
0 4332 5 4 1 78730
0 4333 7 5 2 78731 76295
0 4334 5 8 1 78741
0 4335 7 5 2 68980 74216
0 4336 5 12 1 78754
0 4337 7 2 2 78759 78423
0 4338 5 1 1 78771
0 4339 7 2 2 57599 69409
0 4340 5 3 1 78773
0 4341 7 2 2 59080 78774
0 4342 5 2 1 78778
0 4343 7 1 2 78772 78780
0 4344 5 1 1 4343
0 4345 7 1 2 57881 4344
0 4346 5 1 1 4345
0 4347 7 1 2 78746 4346
0 4348 5 1 1 4347
0 4349 7 1 2 73105 4348
0 4350 5 1 1 4349
0 4351 7 3 2 62584 72132
0 4352 5 2 1 78782
0 4353 7 1 2 78691 75026
0 4354 5 6 1 4353
0 4355 7 1 2 74867 78787
0 4356 5 3 1 4355
0 4357 7 1 2 78785 78793
0 4358 5 1 1 4357
0 4359 7 1 2 58156 4358
0 4360 5 1 1 4359
0 4361 7 8 2 62585 65427
0 4362 5 2 1 78796
0 4363 7 2 2 74510 78797
0 4364 5 1 1 78806
0 4365 7 2 2 70684 78807
0 4366 5 1 1 78808
0 4367 7 1 2 65788 4366
0 4368 7 1 2 4360 4367
0 4369 7 1 2 4350 4368
0 4370 7 1 2 4330 4369
0 4371 5 1 1 4370
0 4372 7 5 2 59081 67419
0 4373 5 5 1 78810
0 4374 7 9 2 65164 68723
0 4375 7 1 2 78811 78820
0 4376 5 1 1 4375
0 4377 7 2 2 76161 4376
0 4378 5 1 1 78829
0 4379 7 7 2 70806 73285
0 4380 7 4 2 62154 69019
0 4381 5 2 1 78838
0 4382 7 7 2 71708 78842
0 4383 5 37 1 78844
0 4384 7 1 2 70956 78845
0 4385 5 3 1 4384
0 4386 7 1 2 78831 78888
0 4387 5 2 1 4386
0 4388 7 1 2 58157 78891
0 4389 5 1 1 4388
0 4390 7 1 2 60764 4389
0 4391 5 1 1 4390
0 4392 7 1 2 4378 4391
0 4393 5 1 1 4392
0 4394 7 2 2 67714 76544
0 4395 5 2 1 78893
0 4396 7 2 2 73212 78894
0 4397 5 1 1 78897
0 4398 7 1 2 65428 4397
0 4399 5 1 1 4398
0 4400 7 1 2 76254 77123
0 4401 5 1 1 4400
0 4402 7 1 2 4399 4401
0 4403 5 3 1 4402
0 4404 7 1 2 70383 78899
0 4405 5 1 1 4404
0 4406 7 14 2 58158 67979
0 4407 5 8 1 78902
0 4408 7 1 2 61167 78916
0 4409 7 1 2 4405 4408
0 4410 7 1 2 4393 4409
0 4411 5 1 1 4410
0 4412 7 1 2 59444 4411
0 4413 7 1 2 4371 4412
0 4414 5 1 1 4413
0 4415 7 13 2 58159 64164
0 4416 5 3 1 78924
0 4417 7 3 2 65789 69410
0 4418 5 3 1 78940
0 4419 7 1 2 78925 78941
0 4420 5 1 1 4419
0 4421 7 9 2 57330 61168
0 4422 7 1 2 70055 78946
0 4423 5 2 1 4422
0 4424 7 1 2 73339 78955
0 4425 5 1 1 4424
0 4426 7 1 2 71709 4425
0 4427 5 1 1 4426
0 4428 7 2 2 57331 72997
0 4429 5 3 1 78957
0 4430 7 1 2 74693 78959
0 4431 5 2 1 4430
0 4432 7 1 2 76364 78962
0 4433 5 1 1 4432
0 4434 7 1 2 4433 74115
0 4435 7 1 2 4427 4434
0 4436 5 1 1 4435
0 4437 7 1 2 59244 4436
0 4438 5 1 1 4437
0 4439 7 1 2 4420 4438
0 4440 5 1 1 4439
0 4441 7 1 2 67631 4440
0 4442 5 1 1 4441
0 4443 7 11 2 57332 65429
0 4444 5 2 1 78964
0 4445 7 3 2 59245 78965
0 4446 7 1 2 61169 78977
0 4447 5 1 1 4446
0 4448 7 1 2 74919 4447
0 4449 5 1 1 4448
0 4450 7 1 2 58160 4449
0 4451 5 1 1 4450
0 4452 7 1 2 4451 74111
0 4453 5 1 1 4452
0 4454 7 1 2 71710 4453
0 4455 5 1 1 4454
0 4456 7 14 2 58161 65790
0 4457 5 9 1 78980
0 4458 7 1 2 69751 75014
0 4459 5 3 1 4458
0 4460 7 1 2 78981 79003
0 4461 5 1 1 4460
0 4462 7 1 2 70249 78958
0 4463 5 1 1 4462
0 4464 7 1 2 61170 70237
0 4465 5 1 1 4464
0 4466 7 1 2 4463 4465
0 4467 5 1 1 4466
0 4468 7 1 2 69446 4467
0 4469 5 1 1 4468
0 4470 7 1 2 4461 4469
0 4471 7 1 2 4455 4470
0 4472 5 1 1 4471
0 4473 7 1 2 68316 4472
0 4474 5 1 1 4473
0 4475 7 1 2 4442 4474
0 4476 5 1 1 4475
0 4477 7 1 2 57882 4476
0 4478 5 1 1 4477
0 4479 7 1 2 76375 70000
0 4480 5 3 1 4479
0 4481 7 1 2 67828 79006
0 4482 5 1 1 4481
0 4483 7 1 2 65430 75095
0 4484 5 2 1 4483
0 4485 7 1 2 4482 79009
0 4486 5 1 1 4485
0 4487 7 1 2 72998 4486
0 4488 5 1 1 4487
0 4489 7 4 2 73773 74970
0 4490 5 1 1 79011
0 4491 7 1 2 68570 79012
0 4492 5 1 1 4491
0 4493 7 1 2 78947 72408
0 4494 5 1 1 4493
0 4495 7 1 2 4492 4494
0 4496 5 1 1 4495
0 4497 7 1 2 67884 4496
0 4498 5 1 1 4497
0 4499 7 1 2 4488 4498
0 4500 5 1 1 4499
0 4501 7 1 2 58162 4500
0 4502 5 1 1 4501
0 4503 7 4 2 57333 69770
0 4504 7 2 2 64954 73734
0 4505 7 2 2 79015 79019
0 4506 5 1 1 79021
0 4507 7 1 2 67885 79022
0 4508 5 1 1 4507
0 4509 7 1 2 64451 4508
0 4510 7 1 2 4502 4509
0 4511 7 1 2 4478 4510
0 4512 7 1 2 4414 4511
0 4513 5 1 1 4512
0 4514 7 1 2 66884 4513
0 4515 7 1 2 4289 4514
0 4516 5 1 1 4515
0 4517 7 9 2 63456 59736
0 4518 5 2 1 79023
0 4519 7 10 2 64669 79024
0 4520 5 1 1 79034
0 4521 7 7 2 65791 71144
0 4522 7 8 2 60242 68460
0 4523 5 8 1 79051
0 4524 7 13 2 79059 78408
0 4525 5 10 1 79067
0 4526 7 1 2 70142 79068
0 4527 5 1 1 4526
0 4528 7 1 2 73147 76296
0 4529 5 2 1 4528
0 4530 7 1 2 70188 79090
0 4531 5 1 1 4530
0 4532 7 1 2 57334 4531
0 4533 5 3 1 4532
0 4534 7 1 2 59246 76390
0 4535 5 1 1 4534
0 4536 7 1 2 79092 4535
0 4537 5 3 1 4536
0 4538 7 1 2 59082 79095
0 4539 5 1 1 4538
0 4540 7 1 2 4527 4539
0 4541 5 1 1 4540
0 4542 7 1 2 57600 4541
0 4543 5 1 1 4542
0 4544 7 4 2 74031 69447
0 4545 7 5 2 57335 71852
0 4546 5 1 1 79102
0 4547 7 1 2 79098 79103
0 4548 5 2 1 4547
0 4549 7 4 2 59083 71711
0 4550 5 10 1 79109
0 4551 7 1 2 65165 79110
0 4552 5 3 1 4551
0 4553 7 2 2 79107 79123
0 4554 5 5 1 79126
0 4555 7 2 2 65431 79128
0 4556 5 1 1 79133
0 4557 7 1 2 59247 79134
0 4558 5 1 1 4557
0 4559 7 1 2 4543 4558
0 4560 5 1 1 4559
0 4561 7 1 2 57883 4560
0 4562 5 1 1 4561
0 4563 7 2 2 70143 78742
0 4564 5 1 1 79135
0 4565 7 1 2 4562 4564
0 4566 5 1 1 4565
0 4567 7 2 2 79044 4566
0 4568 7 1 2 79035 79137
0 4569 5 1 1 4568
0 4570 7 1 2 60243 75063
0 4571 5 1 1 4570
0 4572 7 1 2 72768 4571
0 4573 5 2 1 4572
0 4574 7 2 2 61171 79139
0 4575 7 5 2 58717 63963
0 4576 7 3 2 59967 79143
0 4577 7 20 2 64165 64452
0 4578 5 3 1 79151
0 4579 7 3 2 77410 79152
0 4580 7 1 2 79148 79174
0 4581 7 1 2 79141 4580
0 4582 5 1 1 4581
0 4583 7 1 2 4569 4582
0 4584 7 1 2 4516 4583
0 4585 5 1 1 4584
0 4586 7 1 2 70473 4585
0 4587 5 1 1 4586
0 4588 7 9 2 59737 64780
0 4589 7 5 2 63584 79177
0 4590 7 1 2 66813 79186
0 4591 7 1 2 79138 4590
0 4592 5 1 1 4591
0 4593 7 6 2 67136 71384
0 4594 7 7 2 58842 64453
0 4595 7 4 2 76068 79197
0 4596 7 1 2 79191 79204
0 4597 7 1 2 79142 4596
0 4598 5 1 1 4597
0 4599 7 1 2 4592 4598
0 4600 7 1 2 4587 4599
0 4601 5 1 1 4600
0 4602 7 1 2 62039 4601
0 4603 5 1 1 4602
0 4604 7 4 2 63747 69915
0 4605 7 1 2 77631 71347
0 4606 7 1 2 79208 4605
0 4607 7 11 2 62309 62867
0 4608 5 2 1 79212
0 4609 7 4 2 79213 74939
0 4610 7 9 2 63457 63585
0 4611 5 2 1 79229
0 4612 7 2 2 69375 79230
0 4613 7 5 2 61172 66670
0 4614 7 2 2 60765 79242
0 4615 7 1 2 79240 79247
0 4616 7 1 2 79225 4615
0 4617 7 1 2 4606 4616
0 4618 5 1 1 4617
0 4619 7 1 2 58394 4618
0 4620 7 1 2 4603 4619
0 4621 5 1 1 4620
0 4622 7 2 2 58947 70144
0 4623 5 1 1 79249
0 4624 7 1 2 79093 4623
0 4625 5 1 1 4624
0 4626 7 1 2 57601 4625
0 4627 5 1 1 4626
0 4628 7 1 2 78775 76432
0 4629 7 1 2 79080 4628
0 4630 5 1 1 4629
0 4631 7 1 2 70250 4630
0 4632 5 1 1 4631
0 4633 7 1 2 4627 4632
0 4634 5 1 1 4633
0 4635 7 20 2 59738 59968
0 4636 5 2 1 79251
0 4637 7 2 2 69329 79252
0 4638 7 1 2 4634 79273
0 4639 5 1 1 4638
0 4640 7 4 2 63748 64955
0 4641 5 1 1 79275
0 4642 7 2 2 300 4641
0 4643 5 4 1 79279
0 4644 7 1 2 62155 79280
0 4645 5 1 1 4644
0 4646 7 4 2 75259 4645
0 4647 7 4 2 64454 70278
0 4648 7 3 2 63964 79214
0 4649 7 10 2 64670 64781
0 4650 7 4 2 66671 79296
0 4651 7 1 2 79293 79306
0 4652 7 1 2 79289 4651
0 4653 7 1 2 79285 4652
0 4654 5 1 1 4653
0 4655 7 1 2 4639 4654
0 4656 5 1 1 4655
0 4657 7 1 2 64166 4656
0 4658 5 1 1 4657
0 4659 7 4 2 62040 76603
0 4660 7 1 2 57602 75350
0 4661 5 1 1 4660
0 4662 7 1 2 70189 4661
0 4663 5 2 1 4662
0 4664 7 1 2 68724 79314
0 4665 5 1 1 4664
0 4666 7 1 2 4665 1694
0 4667 5 1 1 4666
0 4668 7 1 2 64956 4667
0 4669 5 1 1 4668
0 4670 7 1 2 69954 70344
0 4671 5 2 1 4670
0 4672 7 1 2 4669 79316
0 4673 5 1 1 4672
0 4674 7 1 2 77226 4673
0 4675 5 1 1 4674
0 4676 7 1 2 70145 77227
0 4677 5 4 1 4676
0 4678 7 6 2 59739 60244
0 4679 7 2 2 70279 79322
0 4680 5 1 1 79328
0 4681 7 1 2 79318 4680
0 4682 5 1 1 4681
0 4683 7 1 2 57603 4682
0 4684 5 1 1 4683
0 4685 7 13 2 59740 60766
0 4686 5 3 1 79330
0 4687 7 3 2 63965 79331
0 4688 5 3 1 79346
0 4689 7 1 2 79319 79349
0 4690 5 1 1 4689
0 4691 7 1 2 65166 4690
0 4692 5 1 1 4691
0 4693 7 1 2 4684 4692
0 4694 5 1 1 4693
0 4695 7 1 2 68571 4694
0 4696 5 1 1 4695
0 4697 7 4 2 63966 72133
0 4698 7 1 2 79352 74054
0 4699 5 1 1 4698
0 4700 7 1 2 4696 4699
0 4701 7 1 2 4675 4700
0 4702 5 1 1 4701
0 4703 7 1 2 59445 4702
0 4704 5 1 1 4703
0 4705 7 11 2 60245 70280
0 4706 5 6 1 79356
0 4707 7 1 2 79357 73961
0 4708 7 1 2 78515 4707
0 4709 5 1 1 4708
0 4710 7 1 2 4704 4709
0 4711 5 1 1 4710
0 4712 7 1 2 79310 4711
0 4713 5 1 1 4712
0 4714 7 1 2 4658 4713
0 4715 5 1 1 4714
0 4716 7 1 2 63586 4715
0 4717 5 1 1 4716
0 4718 7 3 2 58163 69503
0 4719 5 1 1 79373
0 4720 7 7 2 60767 69376
0 4721 5 2 1 79376
0 4722 7 5 2 57336 71464
0 4723 5 2 1 79385
0 4724 7 2 2 78384 79390
0 4725 5 2 1 79392
0 4726 7 1 2 79377 79394
0 4727 5 1 1 4726
0 4728 7 1 2 4719 4727
0 4729 5 1 1 4728
0 4730 7 1 2 57604 4729
0 4731 5 1 1 4730
0 4732 7 1 2 78926 75198
0 4733 5 1 1 4732
0 4734 7 1 2 4731 4733
0 4735 5 1 1 4734
0 4736 7 1 2 59741 4735
0 4737 5 1 1 4736
0 4738 7 6 2 59248 64455
0 4739 7 3 2 74119 79396
0 4740 5 2 1 79402
0 4741 7 1 2 78091 79405
0 4742 5 1 1 4741
0 4743 7 1 2 58164 4742
0 4744 5 1 1 4743
0 4745 7 1 2 63967 74528
0 4746 5 5 1 4745
0 4747 7 1 2 69763 79407
0 4748 5 3 1 4747
0 4749 7 1 2 59742 79412
0 4750 5 1 1 4749
0 4751 7 1 2 4744 4750
0 4752 5 2 1 4751
0 4753 7 1 2 71035 79415
0 4754 5 1 1 4753
0 4755 7 1 2 73148 75708
0 4756 5 1 1 4755
0 4757 7 1 2 70190 1568
0 4758 7 1 2 4756 4757
0 4759 5 1 1 4758
0 4760 7 2 2 58165 73710
0 4761 5 5 1 79417
0 4762 7 1 2 78092 79419
0 4763 5 3 1 4762
0 4764 7 1 2 64957 79424
0 4765 7 1 2 4759 4764
0 4766 5 1 1 4765
0 4767 7 1 2 4754 4766
0 4768 5 1 1 4767
0 4769 7 1 2 65167 4768
0 4770 5 1 1 4769
0 4771 7 1 2 79332 69859
0 4772 5 1 1 4771
0 4773 7 1 2 65432 79425
0 4774 7 1 2 78356 4773
0 4775 5 1 1 4774
0 4776 7 1 2 4772 4775
0 4777 5 1 1 4776
0 4778 7 1 2 59249 4777
0 4779 5 1 1 4778
0 4780 7 1 2 4770 4779
0 4781 7 1 2 4737 4780
0 4782 5 2 1 4781
0 4783 7 1 2 70449 74792
0 4784 7 1 2 79427 4783
0 4785 5 1 1 4784
0 4786 7 1 2 4717 4785
0 4787 5 1 1 4786
0 4788 7 1 2 63458 4787
0 4789 5 1 1 4788
0 4790 7 9 2 58718 64671
0 4791 5 7 1 79429
0 4792 7 1 2 79430 70546
0 4793 7 1 2 79428 4792
0 4794 5 1 1 4793
0 4795 7 1 2 4789 4794
0 4796 5 1 1 4795
0 4797 7 1 2 59084 4796
0 4798 5 1 1 4797
0 4799 7 5 2 62868 64456
0 4800 7 14 2 58719 64167
0 4801 7 2 2 79445 79450
0 4802 7 2 2 59969 74971
0 4803 5 1 1 79466
0 4804 7 1 2 60487 79467
0 4805 7 1 2 79464 4804
0 4806 5 1 1 4805
0 4807 7 2 2 71618 75778
0 4808 5 1 1 79468
0 4809 7 1 2 64958 67579
0 4810 7 3 2 79469 4809
0 4811 5 1 1 79470
0 4812 7 1 2 70356 4811
0 4813 5 1 1 4812
0 4814 7 1 2 64168 4813
0 4815 5 1 1 4814
0 4816 7 1 2 64169 67101
0 4817 5 1 1 4816
0 4818 7 1 2 79378 4817
0 4819 5 1 1 4818
0 4820 7 1 2 4815 4819
0 4821 5 1 1 4820
0 4822 7 1 2 59743 4821
0 4823 5 1 1 4822
0 4824 7 1 2 79403 79471
0 4825 5 1 1 4824
0 4826 7 1 2 4823 4825
0 4827 5 1 1 4826
0 4828 7 1 2 58166 4827
0 4829 5 1 1 4828
0 4830 7 1 2 67008 79416
0 4831 5 1 1 4830
0 4832 7 1 2 73962 79004
0 4833 5 1 1 4832
0 4834 7 1 2 4831 4833
0 4835 5 1 1 4834
0 4836 7 1 2 68572 4835
0 4837 5 1 1 4836
0 4838 7 1 2 70146 78069
0 4839 7 1 2 79472 4838
0 4840 5 1 1 4839
0 4841 7 1 2 4837 4840
0 4842 7 1 2 4829 4841
0 4843 5 1 1 4842
0 4844 7 1 2 66885 4843
0 4845 5 1 1 4844
0 4846 7 1 2 4806 4845
0 4847 5 1 1 4846
0 4848 7 1 2 70474 4847
0 4849 5 1 1 4848
0 4850 7 2 2 60488 70903
0 4851 5 1 1 79473
0 4852 7 2 2 79474 69214
0 4853 7 4 2 66745 79153
0 4854 7 1 2 58843 79477
0 4855 7 1 2 79475 4854
0 4856 5 1 1 4855
0 4857 7 1 2 4849 4856
0 4858 5 1 1 4857
0 4859 7 1 2 62041 4858
0 4860 5 1 1 4859
0 4861 7 1 2 4798 4860
0 4862 5 1 1 4861
0 4863 7 1 2 57884 4862
0 4864 5 1 1 4863
0 4865 7 21 2 64170 60246
0 4866 5 4 1 79481
0 4867 7 3 2 67137 79482
0 4868 5 1 1 79506
0 4869 7 5 2 60768 67715
0 4870 5 9 1 79509
0 4871 7 3 2 65168 79510
0 4872 5 2 1 79523
0 4873 7 1 2 68461 70314
0 4874 7 1 2 78140 4873
0 4875 5 1 1 4874
0 4876 7 1 2 79526 4875
0 4877 5 1 1 4876
0 4878 7 1 2 79507 4877
0 4879 5 1 1 4878
0 4880 7 2 2 74972 76822
0 4881 5 1 1 79528
0 4882 7 1 2 75035 4881
0 4883 5 1 1 4882
0 4884 7 1 2 64171 4883
0 4885 5 1 1 4884
0 4886 7 2 2 63823 70668
0 4887 5 2 1 79530
0 4888 7 2 2 72157 79532
0 4889 5 7 1 79534
0 4890 7 3 2 60247 79536
0 4891 5 1 1 79543
0 4892 7 1 2 70588 77038
0 4893 5 1 1 4892
0 4894 7 1 2 79544 4893
0 4895 5 1 1 4894
0 4896 7 1 2 78694 4895
0 4897 7 1 2 4885 4896
0 4898 5 1 1 4897
0 4899 7 1 2 77919 4898
0 4900 5 1 1 4899
0 4901 7 1 2 4879 4900
0 4902 5 2 1 4901
0 4903 7 1 2 79205 79546
0 4904 5 1 1 4903
0 4905 7 14 2 58720 64457
0 4906 5 3 1 79548
0 4907 7 8 2 59970 79549
0 4908 5 1 1 79565
0 4909 7 1 2 79566 79547
0 4910 5 1 1 4909
0 4911 7 3 2 60769 68317
0 4912 5 1 1 79573
0 4913 7 1 2 78707 4912
0 4914 5 1 1 4913
0 4915 7 1 2 60489 4914
0 4916 5 1 1 4915
0 4917 7 1 2 76952 75019
0 4918 5 1 1 4917
0 4919 7 1 2 4916 4918
0 4920 5 1 1 4919
0 4921 7 1 2 60248 4920
0 4922 5 1 1 4921
0 4923 7 1 2 78794 4922
0 4924 5 1 1 4923
0 4925 7 1 2 59446 4924
0 4926 5 1 1 4925
0 4927 7 1 2 67632 79005
0 4928 5 1 1 4927
0 4929 7 1 2 78520 74973
0 4930 5 3 1 4929
0 4931 7 1 2 4928 79576
0 4932 5 1 1 4931
0 4933 7 1 2 68573 4932
0 4934 5 1 1 4933
0 4935 7 3 2 64172 72014
0 4936 5 4 1 79579
0 4937 7 1 2 79582 79577
0 4938 5 1 1 4937
0 4939 7 1 2 59250 4938
0 4940 5 1 1 4939
0 4941 7 1 2 4934 4940
0 4942 7 1 2 4926 4941
0 4943 5 1 1 4942
0 4944 7 1 2 58167 4943
0 4945 5 1 1 4944
0 4946 7 1 2 59447 78809
0 4947 5 1 1 4946
0 4948 7 4 2 77654 78585
0 4949 5 1 1 79586
0 4950 7 1 2 70147 79587
0 4951 5 1 1 4950
0 4952 7 1 2 69708 76953
0 4953 5 1 1 4952
0 4954 7 1 2 4951 4953
0 4955 5 1 1 4954
0 4956 7 1 2 60249 4955
0 4957 5 1 1 4956
0 4958 7 2 2 62586 69709
0 4959 5 1 1 79590
0 4960 7 1 2 59448 4959
0 4961 7 1 2 4957 4960
0 4962 5 1 1 4961
0 4963 7 2 2 64173 70239
0 4964 5 1 1 79592
0 4965 7 10 2 74804 73852
0 4966 5 9 1 79594
0 4967 7 2 2 64959 70251
0 4968 7 1 2 79595 79613
0 4969 5 1 1 4968
0 4970 7 1 2 79593 4969
0 4971 5 1 1 4970
0 4972 7 1 2 65169 4971
0 4973 7 1 2 4962 4972
0 4974 5 1 1 4973
0 4975 7 1 2 4947 4974
0 4976 7 1 2 4945 4975
0 4977 5 1 1 4976
0 4978 7 1 2 59744 4977
0 4979 5 1 1 4978
0 4980 7 5 2 70865 69995
0 4981 5 3 1 79615
0 4982 7 3 2 65170 79616
0 4983 5 3 1 79623
0 4984 7 4 2 59085 67099
0 4985 5 2 1 79629
0 4986 7 9 2 64458 71145
0 4987 5 2 1 79635
0 4988 7 1 2 79630 79636
0 4989 7 1 2 79624 4988
0 4990 5 1 1 4989
0 4991 7 1 2 4979 4990
0 4992 5 1 1 4991
0 4993 7 1 2 66886 4992
0 4994 5 1 1 4993
0 4995 7 1 2 4910 4994
0 4996 5 1 1 4995
0 4997 7 1 2 70475 4996
0 4998 5 1 1 4997
0 4999 7 1 2 4904 4998
0 5000 5 1 1 4999
0 5001 7 1 2 62042 5000
0 5002 5 1 1 5001
0 5003 7 1 2 65792 5002
0 5004 7 1 2 4864 5003
0 5005 5 1 1 5004
0 5006 7 5 2 64174 68725
0 5007 5 1 1 79646
0 5008 7 6 2 57885 64459
0 5009 7 1 2 62869 79651
0 5010 7 1 2 79647 5009
0 5011 7 1 2 75889 5010
0 5012 5 1 1 5011
0 5013 7 6 2 62870 78070
0 5014 5 2 1 79657
0 5015 7 1 2 79663 79420
0 5016 5 2 1 5015
0 5017 7 5 2 60490 68218
0 5018 5 4 1 79667
0 5019 7 4 2 67138 68462
0 5020 7 1 2 79668 79676
0 5021 7 1 2 79665 5020
0 5022 5 1 1 5021
0 5023 7 1 2 5012 5022
0 5024 5 1 1 5023
0 5025 7 1 2 60250 5024
0 5026 5 1 1 5025
0 5027 7 6 2 62310 70807
0 5028 5 5 1 79680
0 5029 7 1 2 57605 74583
0 5030 5 1 1 5029
0 5031 7 3 2 79686 5030
0 5032 7 3 2 69307 79652
0 5033 7 1 2 68574 78696
0 5034 7 1 2 79694 5033
0 5035 7 1 2 79691 5034
0 5036 5 1 1 5035
0 5037 7 1 2 5026 5036
0 5038 5 1 1 5037
0 5039 7 1 2 60770 5038
0 5040 5 1 1 5039
0 5041 7 3 2 57606 75043
0 5042 5 1 1 79697
0 5043 7 1 2 70991 5042
0 5044 5 2 1 5043
0 5045 7 1 2 68726 79700
0 5046 5 1 1 5045
0 5047 7 1 2 60251 76954
0 5048 7 1 2 70119 5047
0 5049 5 1 1 5048
0 5050 7 1 2 5046 5049
0 5051 5 1 1 5050
0 5052 7 1 2 60491 5051
0 5053 5 1 1 5052
0 5054 7 1 2 57337 63968
0 5055 7 1 2 74805 5054
0 5056 7 1 2 75072 5055
0 5057 5 1 1 5056
0 5058 7 1 2 5053 5057
0 5059 5 1 1 5058
0 5060 7 5 2 65433 71385
0 5061 7 1 2 79653 79702
0 5062 7 1 2 5059 5061
0 5063 5 1 1 5062
0 5064 7 1 2 5040 5063
0 5065 5 1 1 5064
0 5066 7 1 2 79307 5065
0 5067 5 1 1 5066
0 5068 7 4 2 57886 59449
0 5069 5 4 1 79707
0 5070 7 1 2 73461 78629
0 5071 5 2 1 5070
0 5072 7 1 2 73853 72384
0 5073 5 2 1 5072
0 5074 7 1 2 79715 79717
0 5075 5 1 1 5074
0 5076 7 1 2 57607 5075
0 5077 5 1 1 5076
0 5078 7 2 2 64960 73792
0 5079 5 1 1 79719
0 5080 7 1 2 68575 79720
0 5081 5 1 1 5080
0 5082 7 1 2 5077 5081
0 5083 5 1 1 5082
0 5084 7 1 2 59251 5083
0 5085 5 1 1 5084
0 5086 7 8 2 65434 70758
0 5087 5 1 1 79721
0 5088 7 1 2 75709 79722
0 5089 5 1 1 5088
0 5090 7 1 2 5085 5089
0 5091 5 1 1 5090
0 5092 7 1 2 79708 5091
0 5093 5 1 1 5092
0 5094 7 3 2 73286 73451
0 5095 5 4 1 79729
0 5096 7 1 2 78889 79730
0 5097 5 2 1 5096
0 5098 7 1 2 59450 79736
0 5099 5 1 1 5098
0 5100 7 2 2 67633 72385
0 5101 5 2 1 79738
0 5102 7 1 2 78966 79739
0 5103 5 1 1 5102
0 5104 7 1 2 5099 5103
0 5105 5 1 1 5104
0 5106 7 1 2 67256 5105
0 5107 5 1 1 5106
0 5108 7 4 2 57887 72983
0 5109 5 1 1 79742
0 5110 7 1 2 72519 78900
0 5111 5 1 1 5110
0 5112 7 1 2 5109 5111
0 5113 7 1 2 5107 5112
0 5114 5 1 1 5113
0 5115 7 1 2 58168 5114
0 5116 5 1 1 5115
0 5117 7 1 2 5093 5116
0 5118 5 3 1 5117
0 5119 7 1 2 79274 79746
0 5120 5 1 1 5119
0 5121 7 1 2 5067 5120
0 5122 5 1 1 5121
0 5123 7 1 2 63587 5122
0 5124 5 1 1 5123
0 5125 7 1 2 68318 78630
0 5126 5 2 1 5125
0 5127 7 2 2 67716 79749
0 5128 5 5 1 79751
0 5129 7 3 2 57888 79753
0 5130 5 1 1 79758
0 5131 7 2 2 67829 77124
0 5132 5 2 1 79761
0 5133 7 1 2 77655 79763
0 5134 5 2 1 5133
0 5135 7 1 2 65171 79765
0 5136 5 1 1 5135
0 5137 7 1 2 5130 5136
0 5138 5 1 1 5137
0 5139 7 1 2 60771 5138
0 5140 5 1 1 5139
0 5141 7 5 2 58169 63824
0 5142 7 2 2 60252 79767
0 5143 5 1 1 79772
0 5144 7 1 2 64175 5143
0 5145 7 1 2 5140 5144
0 5146 5 1 1 5145
0 5147 7 1 2 59451 70909
0 5148 5 5 1 5147
0 5149 7 1 2 64460 79774
0 5150 7 1 2 5146 5149
0 5151 5 1 1 5150
0 5152 7 1 2 73731 79664
0 5153 5 6 1 5152
0 5154 7 1 2 62587 79779
0 5155 7 1 2 79140 5154
0 5156 5 1 1 5155
0 5157 7 1 2 5151 5156
0 5158 5 1 1 5157
0 5159 7 1 2 63969 5158
0 5160 5 1 1 5159
0 5161 7 1 2 79752 75294
0 5162 5 1 1 5161
0 5163 7 1 2 62871 5162
0 5164 5 1 1 5163
0 5165 7 3 2 65435 74868
0 5166 7 1 2 71003 79785
0 5167 5 1 1 5166
0 5168 7 1 2 5164 5167
0 5169 5 1 1 5168
0 5170 7 1 2 59252 5169
0 5171 5 1 1 5170
0 5172 7 1 2 75135 78583
0 5173 5 1 1 5172
0 5174 7 9 2 57889 58948
0 5175 5 1 1 79788
0 5176 7 1 2 79358 79789
0 5177 5 1 1 5176
0 5178 7 1 2 75162 5177
0 5179 5 1 1 5178
0 5180 7 1 2 57338 5179
0 5181 5 1 1 5180
0 5182 7 7 2 65436 69448
0 5183 5 2 1 79797
0 5184 7 1 2 62872 79798
0 5185 5 1 1 5184
0 5186 7 1 2 5181 5185
0 5187 5 1 1 5186
0 5188 7 1 2 68319 5187
0 5189 5 1 1 5188
0 5190 7 1 2 5173 5189
0 5191 7 1 2 5171 5190
0 5192 5 1 1 5191
0 5193 7 1 2 64176 5192
0 5194 5 1 1 5193
0 5195 7 1 2 70315 74883
0 5196 5 1 1 5195
0 5197 7 1 2 60253 5196
0 5198 5 1 1 5197
0 5199 7 1 2 78565 5198
0 5200 5 1 1 5199
0 5201 7 1 2 78498 5200
0 5202 5 1 1 5201
0 5203 7 1 2 5194 5202
0 5204 5 1 1 5203
0 5205 7 1 2 64461 5204
0 5206 5 1 1 5205
0 5207 7 1 2 5160 5206
0 5208 5 2 1 5207
0 5209 7 1 2 76055 79806
0 5210 5 1 1 5209
0 5211 7 8 2 64782 79253
0 5212 5 1 1 79808
0 5213 7 1 2 79747 79809
0 5214 5 1 1 5213
0 5215 7 1 2 5210 5214
0 5216 5 1 1 5215
0 5217 7 1 2 68661 5216
0 5218 5 1 1 5217
0 5219 7 1 2 5124 5218
0 5220 5 1 1 5219
0 5221 7 1 2 63459 5220
0 5222 5 1 1 5221
0 5223 7 1 2 59971 79807
0 5224 5 1 1 5223
0 5225 7 17 2 59745 64672
0 5226 7 1 2 79816 79748
0 5227 5 1 1 5226
0 5228 7 1 2 5224 5227
0 5229 5 1 1 5228
0 5230 7 4 2 74886 70476
0 5231 7 1 2 5229 79833
0 5232 5 1 1 5231
0 5233 7 1 2 61173 5232
0 5234 7 1 2 5222 5233
0 5235 5 1 1 5234
0 5236 7 1 2 5005 5235
0 5237 5 1 1 5236
0 5238 7 7 2 63970 64961
0 5239 7 1 2 73238 79837
0 5240 5 2 1 5239
0 5241 7 1 2 73641 79844
0 5242 5 1 1 5241
0 5243 7 9 2 64177 59972
0 5244 7 6 2 64462 60492
0 5245 7 1 2 79846 79855
0 5246 7 1 2 77334 5245
0 5247 5 1 1 5246
0 5248 7 1 2 68727 77700
0 5249 5 1 1 5248
0 5250 7 1 2 77684 5249
0 5251 5 1 1 5250
0 5252 7 7 2 63460 59973
0 5253 5 1 1 79861
0 5254 7 4 2 79438 5253
0 5255 5 45 1 79868
0 5256 7 1 2 79872 73826
0 5257 7 1 2 5251 5256
0 5258 5 1 1 5257
0 5259 7 1 2 5247 5258
0 5260 5 1 1 5259
0 5261 7 1 2 70477 5260
0 5262 5 1 1 5261
0 5263 7 2 2 64463 76933
0 5264 7 2 2 62588 63461
0 5265 7 3 2 64673 79919
0 5266 7 2 2 58844 64178
0 5267 7 2 2 63825 79924
0 5268 7 1 2 79921 79926
0 5269 7 1 2 79917 5268
0 5270 5 1 1 5269
0 5271 7 1 2 5262 5270
0 5272 5 1 1 5271
0 5273 7 1 2 62043 5272
0 5274 5 1 1 5273
0 5275 7 6 2 63588 64464
0 5276 7 2 2 64783 79928
0 5277 7 2 2 77632 79934
0 5278 7 2 2 60493 77411
0 5279 5 1 1 79938
0 5280 7 6 2 63462 66672
0 5281 7 1 2 58949 79940
0 5282 7 1 2 79939 5281
0 5283 7 1 2 74005 5282
0 5284 7 1 2 79936 5283
0 5285 5 1 1 5284
0 5286 7 1 2 5274 5285
0 5287 5 1 1 5286
0 5288 7 1 2 5242 5287
0 5289 5 1 1 5288
0 5290 7 3 2 77448 71661
0 5291 5 1 1 79946
0 5292 7 7 2 66814 70478
0 5293 5 1 1 79949
0 5294 7 7 2 63463 58845
0 5295 7 6 2 76056 79956
0 5296 5 1 1 79963
0 5297 7 1 2 5293 5296
0 5298 5 10 1 5297
0 5299 7 11 2 64465 60772
0 5300 5 2 1 79979
0 5301 7 8 2 62873 60254
0 5302 5 3 1 79992
0 5303 7 6 2 60494 62044
0 5304 7 1 2 79993 80003
0 5305 7 1 2 79980 5304
0 5306 7 1 2 79969 5305
0 5307 7 1 2 79947 5306
0 5308 5 1 1 5307
0 5309 7 1 2 63145 5308
0 5310 7 1 2 5289 5309
0 5311 7 1 2 5237 5310
0 5312 5 1 1 5311
0 5313 7 1 2 4621 5312
0 5314 5 1 1 5313
0 5315 7 1 2 66552 5314
0 5316 5 1 1 5315
0 5317 7 3 2 72231 69602
0 5318 5 1 1 80009
0 5319 7 1 2 71853 69603
0 5320 5 4 1 5319
0 5321 7 2 2 62874 73354
0 5322 7 5 2 59253 69232
0 5323 7 2 2 65172 80018
0 5324 7 1 2 80016 80023
0 5325 5 1 1 5324
0 5326 7 1 2 80012 5325
0 5327 5 1 1 5326
0 5328 7 1 2 57608 5327
0 5329 5 1 1 5328
0 5330 7 1 2 5318 5329
0 5331 5 1 1 5330
0 5332 7 1 2 72999 5331
0 5333 5 1 1 5332
0 5334 7 2 2 68955 69258
0 5335 7 1 2 60495 80025
0 5336 5 1 1 5335
0 5337 7 1 2 69356 5336
0 5338 5 1 1 5337
0 5339 7 1 2 57609 5338
0 5340 5 1 1 5339
0 5341 7 1 2 80013 5340
0 5342 5 1 1 5341
0 5343 7 1 2 58170 5342
0 5344 5 1 1 5343
0 5345 7 2 2 57610 68675
0 5346 7 1 2 76087 80027
0 5347 5 1 1 5346
0 5348 7 1 2 5344 5347
0 5349 5 1 1 5348
0 5350 7 1 2 78948 5349
0 5351 5 1 1 5350
0 5352 7 1 2 5333 5351
0 5353 5 1 1 5352
0 5354 7 1 2 58950 5353
0 5355 5 1 1 5354
0 5356 7 4 2 61174 62045
0 5357 7 4 2 67914 80029
0 5358 7 1 2 72369 80033
0 5359 5 1 1 5358
0 5360 7 1 2 5355 5359
0 5361 5 1 1 5360
0 5362 7 1 2 64962 5361
0 5363 5 1 1 5362
0 5364 7 1 2 78956 1277
0 5365 5 1 1 5364
0 5366 7 1 2 68320 5365
0 5367 5 1 1 5366
0 5368 7 2 2 65173 67868
0 5369 5 1 1 80037
0 5370 7 1 2 78994 5369
0 5371 5 1 1 5370
0 5372 7 1 2 74699 5371
0 5373 5 1 1 5372
0 5374 7 1 2 5367 5373
0 5375 5 1 1 5374
0 5376 7 1 2 69604 5375
0 5377 5 1 1 5376
0 5378 7 1 2 5363 5377
0 5379 5 1 1 5378
0 5380 7 1 2 57890 5379
0 5381 5 1 1 5380
0 5382 7 2 2 72386 69868
0 5383 5 2 1 80039
0 5384 7 8 2 79099 71854
0 5385 5 3 1 80043
0 5386 7 1 2 57611 80044
0 5387 5 1 1 5386
0 5388 7 1 2 80041 5387
0 5389 5 7 1 5388
0 5390 7 1 2 80054 73191
0 5391 5 1 1 5390
0 5392 7 1 2 68981 75923
0 5393 5 1 1 5392
0 5394 7 1 2 59254 73202
0 5395 5 1 1 5394
0 5396 7 1 2 5393 5395
0 5397 5 1 1 5396
0 5398 7 1 2 57339 5397
0 5399 5 1 1 5398
0 5400 7 1 2 59255 78779
0 5401 5 1 1 5400
0 5402 7 1 2 61175 5401
0 5403 7 1 2 5399 5402
0 5404 5 1 1 5403
0 5405 7 1 2 69020 79669
0 5406 5 4 1 5405
0 5407 7 1 2 64179 80061
0 5408 5 2 1 5407
0 5409 7 1 2 65793 80065
0 5410 5 1 1 5409
0 5411 7 1 2 58171 5410
0 5412 7 1 2 5404 5411
0 5413 5 1 1 5412
0 5414 7 1 2 5391 5413
0 5415 5 1 1 5414
0 5416 7 1 2 69605 5415
0 5417 5 1 1 5416
0 5418 7 1 2 5381 5417
0 5419 5 1 1 5418
0 5420 7 1 2 65437 5419
0 5421 5 1 1 5420
0 5422 7 2 2 72158 70678
0 5423 5 6 1 80067
0 5424 7 3 2 60773 69021
0 5425 5 5 1 80075
0 5426 7 3 2 80069 80078
0 5427 7 1 2 72165 80083
0 5428 5 1 1 5427
0 5429 7 1 2 79799 69606
0 5430 5 1 1 5429
0 5431 7 1 2 5428 5430
0 5432 5 1 1 5431
0 5433 7 1 2 57340 5432
0 5434 5 1 1 5433
0 5435 7 5 2 58172 69607
0 5436 5 2 1 80086
0 5437 7 1 2 5434 80091
0 5438 5 1 1 5437
0 5439 7 1 2 68321 5438
0 5440 5 1 1 5439
0 5441 7 1 2 5440 76572
0 5442 5 1 1 5441
0 5443 7 1 2 67257 5442
0 5444 5 1 1 5443
0 5445 7 1 2 60774 69480
0 5446 5 4 1 5445
0 5447 7 2 2 68322 80093
0 5448 5 2 1 80097
0 5449 7 1 2 57891 80098
0 5450 5 1 1 5449
0 5451 7 1 2 79626 5450
0 5452 5 1 1 5451
0 5453 7 1 2 72178 5452
0 5454 5 1 1 5453
0 5455 7 2 2 62875 74634
0 5456 5 8 1 80101
0 5457 7 2 2 73149 68676
0 5458 7 1 2 72351 80111
0 5459 5 1 1 5458
0 5460 7 1 2 65438 76868
0 5461 7 1 2 76410 5460
0 5462 5 1 1 5461
0 5463 7 1 2 69499 5462
0 5464 5 2 1 5463
0 5465 7 1 2 70076 80113
0 5466 5 1 1 5465
0 5467 7 1 2 5459 5466
0 5468 5 1 1 5467
0 5469 7 1 2 80103 5468
0 5470 5 1 1 5469
0 5471 7 1 2 61176 5470
0 5472 7 1 2 5454 5471
0 5473 7 1 2 5444 5472
0 5474 7 4 2 57612 63589
0 5475 7 4 2 69233 80115
0 5476 7 1 2 77705 80119
0 5477 5 1 1 5476
0 5478 7 1 2 73203 69608
0 5479 5 1 1 5478
0 5480 7 1 2 5477 5479
0 5481 5 1 1 5480
0 5482 7 1 2 67258 5481
0 5483 5 1 1 5482
0 5484 7 2 2 76872 71054
0 5485 5 1 1 80123
0 5486 7 1 2 72262 5485
0 5487 5 1 1 5486
0 5488 7 1 2 70698 5487
0 5489 5 1 1 5488
0 5490 7 1 2 80092 5489
0 5491 7 1 2 5483 5490
0 5492 5 1 1 5491
0 5493 7 1 2 65439 5492
0 5494 5 1 1 5493
0 5495 7 1 2 72223 67023
0 5496 5 1 1 5495
0 5497 7 1 2 69348 5496
0 5498 5 1 1 5497
0 5499 7 3 2 60775 72232
0 5500 7 2 2 69182 69259
0 5501 7 1 2 80125 80128
0 5502 5 1 1 5501
0 5503 7 2 2 71606 67440
0 5504 7 1 2 80019 80130
0 5505 5 1 1 5504
0 5506 7 1 2 5502 5505
0 5507 7 1 2 5498 5506
0 5508 5 1 1 5507
0 5509 7 1 2 58173 5508
0 5510 5 1 1 5509
0 5511 7 1 2 70252 69609
0 5512 5 1 1 5511
0 5513 7 5 2 70191 73150
0 5514 5 1 1 80132
0 5515 7 4 2 62156 63971
0 5516 5 2 1 80137
0 5517 7 1 2 80133 80141
0 5518 7 1 2 76554 5517
0 5519 5 1 1 5518
0 5520 7 1 2 5512 5519
0 5521 5 1 1 5520
0 5522 7 1 2 67830 5521
0 5523 5 1 1 5522
0 5524 7 2 2 75846 68426
0 5525 5 4 1 80143
0 5526 7 1 2 80144 69610
0 5527 5 1 1 5526
0 5528 7 1 2 5523 5527
0 5529 7 1 2 5510 5528
0 5530 7 1 2 5494 5529
0 5531 5 1 1 5530
0 5532 7 1 2 71712 5531
0 5533 5 1 1 5532
0 5534 7 2 2 69234 73355
0 5535 7 1 2 57613 70669
0 5536 5 3 1 5535
0 5537 7 1 2 60776 70933
0 5538 7 1 2 80142 5537
0 5539 7 1 2 67029 5538
0 5540 5 1 1 5539
0 5541 7 1 2 80151 5540
0 5542 5 1 1 5541
0 5543 7 1 2 57892 5542
0 5544 5 1 1 5543
0 5545 7 8 2 62157 79276
0 5546 5 4 1 80154
0 5547 7 1 2 70148 80155
0 5548 5 1 1 5547
0 5549 7 2 2 60496 70149
0 5550 5 1 1 80166
0 5551 7 1 2 78676 76593
0 5552 5 1 1 5551
0 5553 7 1 2 5550 5552
0 5554 5 1 1 5553
0 5555 7 1 2 58951 5554
0 5556 5 1 1 5555
0 5557 7 1 2 5548 5556
0 5558 7 1 2 5544 5557
0 5559 5 1 1 5558
0 5560 7 1 2 80149 5559
0 5561 5 1 1 5560
0 5562 7 1 2 68068 80099
0 5563 5 1 1 5562
0 5564 7 1 2 69611 5563
0 5565 5 1 1 5564
0 5566 7 4 2 66673 71957
0 5567 7 1 2 67980 80168
0 5568 7 1 2 74045 5567
0 5569 5 1 1 5568
0 5570 7 1 2 5565 5569
0 5571 7 1 2 5561 5570
0 5572 5 1 1 5571
0 5573 7 1 2 58174 5572
0 5574 5 1 1 5573
0 5575 7 2 2 70679 72292
0 5576 5 6 1 80172
0 5577 7 2 2 66674 80174
0 5578 7 1 2 69449 69515
0 5579 7 1 2 80180 5578
0 5580 5 1 1 5579
0 5581 7 1 2 69702 5580
0 5582 5 1 1 5581
0 5583 7 1 2 57341 5582
0 5584 5 1 1 5583
0 5585 7 1 2 75348 76839
0 5586 5 1 1 5585
0 5587 7 1 2 5584 5586
0 5588 5 1 1 5587
0 5589 7 1 2 58175 5588
0 5590 5 1 1 5589
0 5591 7 4 2 59256 72465
0 5592 5 1 1 80182
0 5593 7 1 2 70063 5592
0 5594 7 1 2 79094 5593
0 5595 5 1 1 5594
0 5596 7 1 2 69349 5595
0 5597 5 1 1 5596
0 5598 7 1 2 5590 5597
0 5599 5 1 1 5598
0 5600 7 1 2 67831 5599
0 5601 5 1 1 5600
0 5602 7 1 2 5574 5601
0 5603 7 1 2 5533 5602
0 5604 7 1 2 5473 5603
0 5605 5 1 1 5604
0 5606 7 1 2 70993 80124
0 5607 5 1 1 5606
0 5608 7 2 2 62589 73213
0 5609 7 2 2 67717 80186
0 5610 5 7 1 80188
0 5611 7 1 2 80190 69612
0 5612 5 1 1 5611
0 5613 7 1 2 5607 5612
0 5614 5 1 1 5613
0 5615 7 1 2 77125 5614
0 5616 5 1 1 5615
0 5617 7 3 2 62876 74869
0 5618 5 1 1 80197
0 5619 7 1 2 69978 77694
0 5620 7 1 2 80198 5619
0 5621 5 1 1 5620
0 5622 7 1 2 69613 5621
0 5623 5 1 1 5622
0 5624 7 1 2 60777 5623
0 5625 7 1 2 5616 5624
0 5626 5 1 1 5625
0 5627 7 6 2 63826 78236
0 5628 5 4 1 80200
0 5629 7 1 2 80201 72166
0 5630 5 1 1 5629
0 5631 7 1 2 72182 5630
0 5632 5 1 1 5631
0 5633 7 1 2 62590 5632
0 5634 5 1 1 5633
0 5635 7 2 2 70685 69614
0 5636 5 1 1 80210
0 5637 7 1 2 60497 80211
0 5638 5 1 1 5637
0 5639 7 1 2 65440 5638
0 5640 7 1 2 5634 5639
0 5641 5 1 1 5640
0 5642 7 1 2 5626 5641
0 5643 5 1 1 5642
0 5644 7 3 2 63972 71987
0 5645 5 1 1 80212
0 5646 7 1 2 72293 5645
0 5647 5 1 1 5646
0 5648 7 1 2 62591 5647
0 5649 5 1 1 5648
0 5650 7 1 2 75049 5649
0 5651 5 2 1 5650
0 5652 7 1 2 80215 72167
0 5653 5 1 1 5652
0 5654 7 1 2 74966 74458
0 5655 5 2 1 5654
0 5656 7 1 2 80217 72119
0 5657 5 1 1 5656
0 5658 7 1 2 78715 69494
0 5659 5 1 1 5658
0 5660 7 4 2 64784 60498
0 5661 7 2 2 72306 80219
0 5662 7 1 2 70686 71055
0 5663 7 1 2 80223 5662
0 5664 5 1 1 5663
0 5665 7 1 2 5659 5664
0 5666 5 1 1 5665
0 5667 7 1 2 68463 5666
0 5668 5 1 1 5667
0 5669 7 1 2 5657 5668
0 5670 7 1 2 5653 5669
0 5671 5 1 1 5670
0 5672 7 1 2 70608 5671
0 5673 5 1 1 5672
0 5674 7 1 2 63973 80087
0 5675 5 1 1 5674
0 5676 7 1 2 65794 5675
0 5677 7 1 2 5673 5676
0 5678 7 1 2 5643 5677
0 5679 5 1 1 5678
0 5680 7 1 2 59452 5679
0 5681 7 1 2 5605 5680
0 5682 5 1 1 5681
0 5683 7 1 2 73204 78963
0 5684 5 1 1 5683
0 5685 7 4 2 57342 67634
0 5686 7 1 2 73000 80225
0 5687 5 1 1 5686
0 5688 7 1 2 5684 5687
0 5689 5 1 1 5688
0 5690 7 1 2 65441 5689
0 5691 5 1 1 5690
0 5692 7 2 2 65795 69710
0 5693 5 1 1 80229
0 5694 7 1 2 57343 80230
0 5695 5 1 1 5694
0 5696 7 1 2 5691 5695
0 5697 5 1 1 5696
0 5698 7 1 2 67259 5697
0 5699 5 1 1 5698
0 5700 7 3 2 60778 75855
0 5701 5 1 1 80231
0 5702 7 1 2 69752 5701
0 5703 5 1 1 5702
0 5704 7 2 2 65796 70384
0 5705 7 1 2 57344 80234
0 5706 7 1 2 5703 5705
0 5707 5 1 1 5706
0 5708 7 1 2 5699 5707
0 5709 5 1 1 5708
0 5710 7 1 2 71713 5709
0 5711 5 1 1 5710
0 5712 7 3 2 58176 72233
0 5713 5 1 1 80236
0 5714 7 1 2 57893 72209
0 5715 5 1 1 5714
0 5716 7 1 2 5713 5715
0 5717 5 4 1 5716
0 5718 7 1 2 80239 78307
0 5719 5 1 1 5718
0 5720 7 4 2 64963 70385
0 5721 5 1 1 80243
0 5722 7 1 2 74806 80244
0 5723 5 1 1 5722
0 5724 7 1 2 76162 5723
0 5725 5 2 1 5724
0 5726 7 1 2 71855 80247
0 5727 5 1 1 5726
0 5728 7 1 2 78917 5727
0 5729 7 1 2 5719 5728
0 5730 5 1 1 5729
0 5731 7 1 2 73239 5730
0 5732 5 1 1 5731
0 5733 7 1 2 5711 5732
0 5734 5 1 1 5733
0 5735 7 1 2 69615 5734
0 5736 5 1 1 5735
0 5737 7 1 2 66675 73735
0 5738 7 2 2 74175 5737
0 5739 7 2 2 59257 71714
0 5740 5 1 1 80251
0 5741 7 3 2 64180 64785
0 5742 7 1 2 80017 80253
0 5743 7 1 2 80252 5742
0 5744 7 1 2 80249 5743
0 5745 5 1 1 5744
0 5746 7 1 2 5736 5745
0 5747 7 1 2 5682 5746
0 5748 7 1 2 5421 5747
0 5749 5 1 1 5748
0 5750 7 1 2 76728 5749
0 5751 5 1 1 5750
0 5752 7 1 2 71036 72056
0 5753 5 2 1 5752
0 5754 7 1 2 67139 80256
0 5755 5 1 1 5754
0 5756 7 4 2 63827 70918
0 5757 7 2 2 70281 80258
0 5758 5 1 1 80262
0 5759 7 1 2 63749 80263
0 5760 5 1 1 5759
0 5761 7 1 2 5755 5760
0 5762 5 1 1 5761
0 5763 7 1 2 69616 5762
0 5764 5 2 1 5763
0 5765 7 13 2 68819 78644
0 5766 5 7 1 80266
0 5767 7 2 2 63974 80279
0 5768 5 1 1 80286
0 5769 7 1 2 79574 80287
0 5770 5 1 1 5769
0 5771 7 1 2 63828 76335
0 5772 7 1 2 4304 5771
0 5773 7 1 2 80134 5772
0 5774 5 1 1 5773
0 5775 7 1 2 5770 5774
0 5776 5 1 1 5775
0 5777 7 2 2 60499 5776
0 5778 5 1 1 80288
0 5779 7 1 2 70609 80216
0 5780 5 1 1 5779
0 5781 7 1 2 5778 5780
0 5782 5 1 1 5781
0 5783 7 1 2 69260 5782
0 5784 5 1 1 5783
0 5785 7 1 2 69617 80257
0 5786 5 1 1 5785
0 5787 7 1 2 5784 5786
0 5788 5 2 1 5787
0 5789 7 1 2 62877 80290
0 5790 5 1 1 5789
0 5791 7 1 2 80264 5790
0 5792 5 1 1 5791
0 5793 7 1 2 64181 5792
0 5794 5 1 1 5793
0 5795 7 1 2 73106 77412
0 5796 5 3 1 5795
0 5797 7 8 2 62592 72773
0 5798 5 1 1 80295
0 5799 7 6 2 60779 76163
0 5800 5 1 1 80303
0 5801 7 1 2 68219 80304
0 5802 5 1 1 5801
0 5803 7 1 2 5798 5802
0 5804 5 1 1 5803
0 5805 7 2 2 60500 5804
0 5806 7 1 2 68464 80309
0 5807 5 1 1 5806
0 5808 7 1 2 80292 5807
0 5809 5 1 1 5808
0 5810 7 1 2 69618 5809
0 5811 5 1 1 5810
0 5812 7 1 2 65797 5811
0 5813 7 1 2 5794 5812
0 5814 5 1 1 5813
0 5815 7 2 2 59086 78237
0 5816 5 1 1 80311
0 5817 7 1 2 74785 5816
0 5818 5 1 1 5817
0 5819 7 2 2 75164 5818
0 5820 5 1 1 80313
0 5821 7 1 2 59087 76843
0 5822 5 1 1 5821
0 5823 7 1 2 5820 5822
0 5824 5 1 1 5823
0 5825 7 1 2 80120 5824
0 5826 5 1 1 5825
0 5827 7 2 2 68220 78238
0 5828 5 1 1 80315
0 5829 7 1 2 68677 5828
0 5830 5 1 1 5829
0 5831 7 1 2 5826 5830
0 5832 5 1 1 5831
0 5833 7 1 2 57894 5832
0 5834 5 1 1 5833
0 5835 7 2 2 62593 72207
0 5836 5 3 1 80317
0 5837 7 10 2 72234 80319
0 5838 5 1 1 80322
0 5839 7 1 2 80323 69946
0 5840 5 1 1 5839
0 5841 7 1 2 5840 80014
0 5842 5 1 1 5841
0 5843 7 1 2 78357 5842
0 5844 5 1 1 5843
0 5845 7 1 2 78224 76444
0 5846 5 1 1 5845
0 5847 7 1 2 71856 69235
0 5848 7 1 2 74171 5847
0 5849 5 1 1 5848
0 5850 7 1 2 69703 5849
0 5851 5 1 1 5850
0 5852 7 1 2 5846 5851
0 5853 5 1 1 5852
0 5854 7 1 2 71025 68967
0 5855 5 1 1 5854
0 5856 7 1 2 80010 5855
0 5857 5 1 1 5856
0 5858 7 1 2 64182 5857
0 5859 7 1 2 5853 5858
0 5860 7 1 2 5844 5859
0 5861 7 1 2 5834 5860
0 5862 5 1 1 5861
0 5863 7 4 2 60106 69377
0 5864 7 2 2 68662 80332
0 5865 5 1 1 80336
0 5866 7 5 2 74321 69236
0 5867 7 3 2 63590 63975
0 5868 7 1 2 77457 80343
0 5869 7 1 2 80338 5868
0 5870 5 1 1 5869
0 5871 7 1 2 5865 5870
0 5872 5 1 1 5871
0 5873 7 1 2 68465 5872
0 5874 5 1 1 5873
0 5875 7 1 2 67140 72168
0 5876 5 1 1 5875
0 5877 7 1 2 69226 5876
0 5878 5 1 1 5877
0 5879 7 1 2 67560 5878
0 5880 5 1 1 5879
0 5881 7 1 2 5874 5880
0 5882 5 1 1 5881
0 5883 7 1 2 63829 5882
0 5884 5 1 1 5883
0 5885 7 2 2 67141 69619
0 5886 5 1 1 80346
0 5887 7 1 2 59453 5886
0 5888 7 1 2 5884 5887
0 5889 5 1 1 5888
0 5890 7 1 2 5862 5889
0 5891 5 1 1 5890
0 5892 7 1 2 60780 5891
0 5893 5 1 1 5892
0 5894 7 1 2 60501 3143
0 5895 5 1 1 5894
0 5896 7 3 2 57345 67832
0 5897 7 1 2 78546 80348
0 5898 5 1 1 5897
0 5899 7 1 2 5895 5898
0 5900 5 1 1 5899
0 5901 7 1 2 71715 5900
0 5902 5 1 1 5901
0 5903 7 2 2 67260 71645
0 5904 5 1 1 80351
0 5905 7 1 2 3035 750
0 5906 7 1 2 5904 5905
0 5907 5 1 1 5906
0 5908 7 1 2 60502 5907
0 5909 5 1 1 5908
0 5910 7 7 2 64964 68466
0 5911 5 2 1 80353
0 5912 7 1 2 68956 80354
0 5913 5 1 1 5912
0 5914 7 1 2 75344 5913
0 5915 7 1 2 5909 5914
0 5916 7 1 2 5902 5915
0 5917 5 2 1 5916
0 5918 7 2 2 80362 69237
0 5919 7 1 2 64183 69936
0 5920 7 1 2 80364 5919
0 5921 5 1 1 5920
0 5922 7 1 2 63830 74511
0 5923 5 1 1 5922
0 5924 7 1 2 68467 69833
0 5925 5 3 1 5924
0 5926 7 1 2 5923 80366
0 5927 5 2 1 5926
0 5928 7 1 2 76164 80369
0 5929 5 1 1 5928
0 5930 7 7 2 60255 72547
0 5931 5 2 1 80371
0 5932 7 1 2 70745 80372
0 5933 5 1 1 5932
0 5934 7 2 2 62878 69411
0 5935 5 5 1 80380
0 5936 7 1 2 80382 70729
0 5937 7 1 2 5933 5936
0 5938 5 2 1 5937
0 5939 7 1 2 64184 80387
0 5940 5 1 1 5939
0 5941 7 1 2 5929 5940
0 5942 5 1 1 5941
0 5943 7 1 2 69620 5942
0 5944 5 1 1 5943
0 5945 7 1 2 65442 5944
0 5946 7 1 2 5921 5945
0 5947 5 1 1 5946
0 5948 7 1 2 5893 5947
0 5949 5 1 1 5948
0 5950 7 2 2 60256 77337
0 5951 5 1 1 80389
0 5952 7 1 2 78054 68678
0 5953 7 1 2 80390 5952
0 5954 5 1 1 5953
0 5955 7 1 2 61177 5954
0 5956 7 1 2 5949 5955
0 5957 5 1 1 5956
0 5958 7 1 2 58395 5957
0 5959 7 1 2 5814 5958
0 5960 5 1 1 5959
0 5961 7 2 2 69330 77023
0 5962 7 11 2 65174 61178
0 5963 5 1 1 80393
0 5964 7 1 2 80394 71988
0 5965 5 2 1 5964
0 5966 7 1 2 65798 78443
0 5967 5 1 1 5966
0 5968 7 1 2 80404 5967
0 5969 5 1 1 5968
0 5970 7 1 2 80391 5969
0 5971 5 1 1 5970
0 5972 7 2 2 59454 68468
0 5973 7 3 2 73299 68679
0 5974 5 1 1 80408
0 5975 7 1 2 74781 80409
0 5976 5 1 1 5975
0 5977 7 34 2 60781 61179
0 5978 5 7 1 80411
0 5979 7 3 2 58177 80412
0 5980 7 9 2 58396 63591
0 5981 7 2 2 80455 76873
0 5982 7 1 2 80452 80464
0 5983 5 1 1 5982
0 5984 7 1 2 5976 5983
0 5985 5 1 1 5984
0 5986 7 1 2 80406 5985
0 5987 5 1 1 5986
0 5988 7 1 2 5971 5987
0 5989 5 1 1 5988
0 5990 7 1 2 67142 5989
0 5991 5 1 1 5990
0 5992 7 4 2 65443 69834
0 5993 5 1 1 80466
0 5994 7 2 2 69621 80467
0 5995 7 2 2 58397 71242
0 5996 5 1 1 80472
0 5997 7 1 2 61180 80473
0 5998 7 1 2 80470 5997
0 5999 5 1 1 5998
0 6000 7 1 2 5991 5999
0 6001 5 1 1 6000
0 6002 7 1 2 67718 6001
0 6003 5 1 1 6002
0 6004 7 5 2 58178 72851
0 6005 5 4 1 80474
0 6006 7 3 2 76449 76556
0 6007 5 15 1 80483
0 6008 7 1 2 80486 71610
0 6009 5 1 1 6008
0 6010 7 8 2 65175 71716
0 6011 5 18 1 80501
0 6012 7 4 2 60782 80509
0 6013 5 1 1 80527
0 6014 7 2 2 69481 80528
0 6015 5 3 1 80531
0 6016 7 1 2 68323 77059
0 6017 7 1 2 80533 6016
0 6018 5 1 1 6017
0 6019 7 1 2 6009 6018
0 6020 5 1 1 6019
0 6021 7 1 2 67981 6020
0 6022 5 1 1 6021
0 6023 7 2 2 77060 79007
0 6024 7 1 2 67886 80536
0 6025 5 1 1 6024
0 6026 7 1 2 6022 6025
0 6027 5 2 1 6026
0 6028 7 1 2 80475 80538
0 6029 5 1 1 6028
0 6030 7 3 2 79215 75123
0 6031 7 6 2 65176 73300
0 6032 7 1 2 77338 80543
0 6033 7 1 2 80540 6032
0 6034 5 1 1 6033
0 6035 7 1 2 6029 6034
0 6036 5 1 1 6035
0 6037 7 1 2 69622 6036
0 6038 5 1 1 6037
0 6039 7 1 2 6003 6038
0 6040 7 1 2 5960 6039
0 6041 5 1 1 6040
0 6042 7 1 2 59746 6041
0 6043 5 1 1 6042
0 6044 7 18 2 58398 61181
0 6045 5 5 1 80549
0 6046 7 2 2 57895 69955
0 6047 5 4 1 80572
0 6048 7 1 2 67261 79008
0 6049 5 1 1 6048
0 6050 7 1 2 80574 6049
0 6051 5 1 1 6050
0 6052 7 1 2 59088 6051
0 6053 5 1 1 6052
0 6054 7 1 2 67982 75199
0 6055 5 1 1 6054
0 6056 7 1 2 6053 6055
0 6057 5 1 1 6056
0 6058 7 1 2 57614 6057
0 6059 5 1 1 6058
0 6060 7 1 2 57346 70759
0 6061 5 4 1 6060
0 6062 7 1 2 65444 70026
0 6063 5 2 1 6062
0 6064 7 1 2 80578 80582
0 6065 5 1 1 6064
0 6066 7 1 2 67983 6065
0 6067 5 1 1 6066
0 6068 7 1 2 6059 6067
0 6069 5 1 1 6068
0 6070 7 1 2 80550 6069
0 6071 5 1 1 6070
0 6072 7 6 2 58399 65445
0 6073 5 6 1 80584
0 6074 7 2 2 80590 73648
0 6075 7 2 2 60783 78211
0 6076 5 3 1 80598
0 6077 7 1 2 80596 80600
0 6078 5 1 1 6077
0 6079 7 1 2 78334 80551
0 6080 5 1 1 6079
0 6081 7 1 2 6078 6080
0 6082 5 1 1 6081
0 6083 7 1 2 59258 6082
0 6084 5 1 1 6083
0 6085 7 5 2 58952 65799
0 6086 5 2 1 80603
0 6087 7 1 2 78152 80604
0 6088 7 1 2 72635 6087
0 6089 5 1 1 6088
0 6090 7 1 2 6084 6089
0 6091 5 1 1 6090
0 6092 7 1 2 57896 6091
0 6093 5 1 1 6092
0 6094 7 3 2 68982 70345
0 6095 5 1 1 80610
0 6096 7 1 2 78153 74153
0 6097 7 1 2 80611 6096
0 6098 5 1 1 6097
0 6099 7 1 2 6093 6098
0 6100 5 1 1 6099
0 6101 7 1 2 71857 6100
0 6102 5 1 1 6101
0 6103 7 2 2 69956 73605
0 6104 5 1 1 80613
0 6105 7 2 2 57347 79790
0 6106 5 1 1 80615
0 6107 7 1 2 80616 72374
0 6108 7 1 2 80614 6107
0 6109 5 2 1 6108
0 6110 7 3 2 57897 73151
0 6111 5 7 1 80619
0 6112 7 2 2 73480 80620
0 6113 5 1 1 80629
0 6114 7 1 2 80591 80630
0 6115 5 1 1 6114
0 6116 7 3 2 63146 59259
0 6117 7 1 2 80631 79723
0 6118 5 1 1 6117
0 6119 7 1 2 6115 6118
0 6120 5 1 1 6119
0 6121 7 1 2 65800 78308
0 6122 7 1 2 6120 6121
0 6123 5 1 1 6122
0 6124 7 1 2 80617 6123
0 6125 5 1 1 6124
0 6126 7 1 2 59455 6125
0 6127 5 1 1 6126
0 6128 7 1 2 6102 6127
0 6129 7 1 2 6071 6128
0 6130 5 1 1 6129
0 6131 7 1 2 69623 6130
0 6132 5 1 1 6131
0 6133 7 5 2 58400 59260
0 6134 7 2 2 73196 80634
0 6135 5 1 1 80639
0 6136 7 1 2 57348 80597
0 6137 7 1 2 73929 6136
0 6138 5 1 1 6137
0 6139 7 1 2 6135 6138
0 6140 5 1 1 6139
0 6141 7 1 2 75856 6140
0 6142 5 1 1 6141
0 6143 7 3 2 57349 71120
0 6144 7 1 2 70150 73649
0 6145 7 1 2 80641 6144
0 6146 5 1 1 6145
0 6147 7 1 2 6142 6146
0 6148 5 1 1 6147
0 6149 7 1 2 69624 6148
0 6150 5 1 1 6149
0 6151 7 2 2 59261 73419
0 6152 7 1 2 74020 80644
0 6153 7 1 2 80250 6152
0 6154 5 1 1 6153
0 6155 7 1 2 6150 6154
0 6156 5 1 1 6155
0 6157 7 1 2 71717 6156
0 6158 5 1 1 6157
0 6159 7 3 2 59456 73301
0 6160 7 1 2 80646 80339
0 6161 7 3 2 57615 71121
0 6162 7 1 2 80649 71367
0 6163 7 1 2 6160 6162
0 6164 5 1 1 6163
0 6165 7 1 2 6158 6164
0 6166 7 1 2 6132 6165
0 6167 5 1 1 6166
0 6168 7 1 2 77228 6167
0 6169 5 1 1 6168
0 6170 7 1 2 6043 6169
0 6171 7 1 2 5751 6170
0 6172 5 1 1 6171
0 6173 7 1 2 66887 6172
0 6174 5 1 1 6173
0 6175 7 2 2 71989 73509
0 6176 5 1 1 80652
0 6177 7 1 2 72759 73495
0 6178 5 1 1 6177
0 6179 7 1 2 6176 6178
0 6180 5 1 1 6179
0 6181 7 1 2 63147 6180
0 6182 5 1 1 6181
0 6183 7 3 2 70282 80552
0 6184 5 1 1 80654
0 6185 7 6 2 63831 64466
0 6186 7 1 2 80655 80657
0 6187 5 1 1 6186
0 6188 7 1 2 6182 6187
0 6189 5 1 1 6188
0 6190 7 1 2 63976 6189
0 6191 5 1 1 6190
0 6192 7 5 2 63148 73240
0 6193 5 1 1 80663
0 6194 7 1 2 79397 80664
0 6195 5 1 1 6194
0 6196 7 1 2 6191 6195
0 6197 5 1 1 6196
0 6198 7 1 2 71386 6197
0 6199 5 1 1 6198
0 6200 7 7 2 63977 61182
0 6201 7 2 2 77943 80668
0 6202 7 1 2 77790 80675
0 6203 5 1 1 6202
0 6204 7 1 2 6199 6203
0 6205 5 1 1 6204
0 6206 7 1 2 62594 6205
0 6207 5 1 1 6206
0 6208 7 7 2 71387 75500
0 6209 7 1 2 73950 80677
0 6210 7 1 2 79353 6209
0 6211 5 1 1 6210
0 6212 7 1 2 6207 6211
0 6213 5 1 1 6212
0 6214 7 1 2 70610 6213
0 6215 5 1 1 6214
0 6216 7 1 2 77711 75077
0 6217 5 1 1 6216
0 6218 7 1 2 77458 80407
0 6219 7 1 2 6217 6218
0 6220 5 1 1 6219
0 6221 7 3 2 68983 73854
0 6222 5 3 1 80684
0 6223 7 1 2 77516 74788
0 6224 7 1 2 80685 6223
0 6225 5 1 1 6224
0 6226 7 1 2 6220 6225
0 6227 5 1 1 6226
0 6228 7 1 2 63978 6227
0 6229 5 1 1 6228
0 6230 7 2 2 62595 69088
0 6231 5 1 1 80690
0 6232 7 1 2 57350 6231
0 6233 5 2 1 6232
0 6234 7 1 2 76445 80692
0 6235 5 2 1 6234
0 6236 7 1 2 67580 80694
0 6237 5 1 1 6236
0 6238 7 4 2 57898 76500
0 6239 5 5 1 80696
0 6240 7 1 2 77525 80697
0 6241 5 2 1 6240
0 6242 7 1 2 74635 80705
0 6243 7 1 2 6237 6242
0 6244 5 1 1 6243
0 6245 7 1 2 59262 6244
0 6246 5 1 1 6245
0 6247 7 2 2 57616 77528
0 6248 5 1 1 80707
0 6249 7 8 2 65177 67262
0 6250 5 2 1 80709
0 6251 7 1 2 80708 80710
0 6252 5 1 1 6251
0 6253 7 2 2 76297 72815
0 6254 5 1 1 80719
0 6255 7 2 2 59089 80720
0 6256 5 1 1 80721
0 6257 7 1 2 6252 6256
0 6258 7 1 2 6246 6257
0 6259 5 1 1 6258
0 6260 7 1 2 71388 6259
0 6261 5 1 1 6260
0 6262 7 1 2 6229 6261
0 6263 5 1 1 6262
0 6264 7 1 2 60784 6263
0 6265 5 1 1 6264
0 6266 7 1 2 78670 80363
0 6267 5 1 1 6266
0 6268 7 1 2 6265 6267
0 6269 5 1 1 6268
0 6270 7 1 2 61183 6269
0 6271 5 1 1 6270
0 6272 7 1 2 74724 80289
0 6273 5 1 1 6272
0 6274 7 1 2 6271 6273
0 6275 5 1 1 6274
0 6276 7 1 2 75501 6275
0 6277 5 1 1 6276
0 6278 7 1 2 6215 6277
0 6279 5 1 1 6278
0 6280 7 1 2 74305 6279
0 6281 5 1 1 6280
0 6282 7 1 2 75847 77170
0 6283 5 1 1 6282
0 6284 7 1 2 70105 6283
0 6285 5 7 1 6284
0 6286 7 3 2 73302 80723
0 6287 7 1 2 67263 80730
0 6288 5 1 1 6287
0 6289 7 4 2 58953 70760
0 6290 5 1 1 80733
0 6291 7 1 2 70866 80734
0 6292 5 4 1 6291
0 6293 7 1 2 61184 80737
0 6294 5 2 1 6293
0 6295 7 1 2 65446 80741
0 6296 5 1 1 6295
0 6297 7 2 2 65801 71858
0 6298 5 2 1 80743
0 6299 7 1 2 70808 75269
0 6300 5 2 1 6299
0 6301 7 1 2 80744 80747
0 6302 5 1 1 6301
0 6303 7 1 2 6296 6302
0 6304 5 1 1 6303
0 6305 7 1 2 57617 6304
0 6306 5 1 1 6305
0 6307 7 3 2 65802 73462
0 6308 7 1 2 72068 75270
0 6309 5 1 1 6308
0 6310 7 1 2 80749 6309
0 6311 5 1 1 6310
0 6312 7 1 2 6306 6311
0 6313 5 1 1 6312
0 6314 7 1 2 67984 6313
0 6315 5 1 1 6314
0 6316 7 1 2 6288 6315
0 6317 5 2 1 6316
0 6318 7 2 2 72647 74759
0 6319 7 2 2 74793 80754
0 6320 7 1 2 59747 80756
0 6321 7 1 2 80752 6320
0 6322 5 1 1 6321
0 6323 7 1 2 6281 6322
0 6324 5 1 1 6323
0 6325 7 1 2 70479 6324
0 6326 5 1 1 6325
0 6327 7 7 2 62879 72790
0 6328 5 1 1 80758
0 6329 7 1 2 79929 80759
0 6330 7 1 2 80365 6329
0 6331 5 1 1 6330
0 6332 7 8 2 58179 75567
0 6333 5 4 1 80765
0 6334 7 3 2 59457 75568
0 6335 5 1 1 80777
0 6336 7 4 2 80773 6335
0 6337 5 1 1 80780
0 6338 7 9 2 76666 80781
0 6339 7 1 2 67143 80784
0 6340 5 2 1 6339
0 6341 7 28 2 62880 63149
0 6342 5 8 1 80795
0 6343 7 4 2 64467 80796
0 6344 5 1 1 80831
0 6345 7 1 2 80793 6344
0 6346 5 1 1 6345
0 6347 7 1 2 80370 6346
0 6348 5 1 1 6347
0 6349 7 6 2 64468 72791
0 6350 7 1 2 80835 80388
0 6351 5 1 1 6350
0 6352 7 1 2 6348 6351
0 6353 5 1 1 6352
0 6354 7 1 2 69625 6353
0 6355 5 1 1 6354
0 6356 7 1 2 65447 6355
0 6357 7 1 2 6331 6356
0 6358 5 1 1 6357
0 6359 7 2 2 76667 76877
0 6360 5 1 1 80841
0 6361 7 1 2 75569 6360
0 6362 5 4 1 6361
0 6363 7 1 2 79171 80843
0 6364 5 1 1 6363
0 6365 7 5 2 64185 77846
0 6366 5 2 1 80847
0 6367 7 1 2 76165 80848
0 6368 5 2 1 6367
0 6369 7 1 2 6364 80854
0 6370 5 2 1 6369
0 6371 7 1 2 80856 69222
0 6372 5 1 1 6371
0 6373 7 21 2 63979 77413
0 6374 5 3 1 80858
0 6375 7 1 2 80859 69570
0 6376 7 1 2 80849 6375
0 6377 5 1 1 6376
0 6378 7 1 2 6372 6377
0 6379 5 1 1 6378
0 6380 7 1 2 70611 6379
0 6381 5 1 1 6380
0 6382 7 5 2 75502 69571
0 6383 5 1 1 80882
0 6384 7 4 2 62596 58180
0 6385 7 3 2 62311 77339
0 6386 7 1 2 80887 80891
0 6387 7 1 2 80883 6386
0 6388 5 1 1 6387
0 6389 7 1 2 6381 6388
0 6390 5 1 1 6389
0 6391 7 1 2 60503 6390
0 6392 5 1 1 6391
0 6393 7 7 2 63150 73711
0 6394 5 1 1 80894
0 6395 7 1 2 63980 71118
0 6396 7 2 2 80895 6395
0 6397 7 1 2 77478 80340
0 6398 7 1 2 80901 6397
0 6399 5 1 1 6398
0 6400 7 1 2 6392 6399
0 6401 5 1 1 6400
0 6402 7 1 2 63832 6401
0 6403 5 1 1 6402
0 6404 7 1 2 57618 79129
0 6405 5 1 1 6404
0 6406 7 5 2 6405 80738
0 6407 5 11 1 80903
0 6408 7 1 2 80908 76844
0 6409 5 1 1 6408
0 6410 7 1 2 57619 80314
0 6411 5 1 1 6410
0 6412 7 1 2 62312 75897
0 6413 5 4 1 6412
0 6414 7 1 2 79060 80919
0 6415 5 1 1 6414
0 6416 7 1 2 70088 79633
0 6417 7 1 2 6415 6416
0 6418 5 1 1 6417
0 6419 7 1 2 62881 72235
0 6420 7 1 2 6418 6419
0 6421 5 1 1 6420
0 6422 7 1 2 6411 6421
0 6423 5 1 1 6422
0 6424 7 1 2 57899 6423
0 6425 5 1 1 6424
0 6426 7 1 2 6409 6425
0 6427 5 1 1 6426
0 6428 7 1 2 6427 80884
0 6429 5 1 1 6428
0 6430 7 1 2 70761 72197
0 6431 5 1 1 6430
0 6432 7 1 2 59263 78464
0 6433 5 1 1 6432
0 6434 7 1 2 6431 6433
0 6435 7 1 2 70809 78212
0 6436 5 1 1 6435
0 6437 7 1 2 57351 6436
0 6438 5 2 1 6437
0 6439 7 14 2 62158 71673
0 6440 7 6 2 62313 71795
0 6441 5 1 1 80939
0 6442 7 1 2 80925 80940
0 6443 5 5 1 6442
0 6444 7 2 2 57900 80945
0 6445 5 1 1 80950
0 6446 7 1 2 80923 6445
0 6447 7 1 2 6434 6446
0 6448 7 2 2 78370 6447
0 6449 5 1 1 80952
0 6450 7 1 2 75503 6449
0 6451 5 1 1 6450
0 6452 7 1 2 77847 80296
0 6453 5 1 1 6452
0 6454 7 1 2 6451 6453
0 6455 5 1 1 6454
0 6456 7 1 2 69626 6455
0 6457 5 1 1 6456
0 6458 7 1 2 6429 6457
0 6459 5 1 1 6458
0 6460 7 1 2 64186 6459
0 6461 5 1 1 6460
0 6462 7 2 2 67144 73712
0 6463 5 1 1 80954
0 6464 7 5 2 63151 58846
0 6465 7 3 2 69331 80956
0 6466 7 1 2 80955 80961
0 6467 5 1 1 6466
0 6468 7 1 2 60785 6467
0 6469 7 1 2 6461 6468
0 6470 7 1 2 6403 6469
0 6471 5 1 1 6470
0 6472 7 1 2 6358 6471
0 6473 5 1 1 6472
0 6474 7 3 2 62882 80850
0 6475 5 2 1 80964
0 6476 7 1 2 6394 80967
0 6477 5 7 1 6476
0 6478 7 2 2 69378 80969
0 6479 5 1 1 80976
0 6480 7 1 2 80977 80347
0 6481 5 1 1 6480
0 6482 7 2 2 71243 75504
0 6483 5 8 1 80978
0 6484 7 1 2 80794 80980
0 6485 5 5 1 6484
0 6486 7 1 2 80988 80471
0 6487 5 1 1 6486
0 6488 7 2 2 62159 80888
0 6489 7 1 2 80993 80224
0 6490 7 1 2 80902 6489
0 6491 5 1 1 6490
0 6492 7 1 2 6487 6491
0 6493 5 1 1 6492
0 6494 7 1 2 67719 6493
0 6495 5 1 1 6494
0 6496 7 1 2 6481 6495
0 6497 7 1 2 6473 6496
0 6498 5 1 1 6497
0 6499 7 1 2 61185 6498
0 6500 5 1 1 6499
0 6501 7 1 2 64187 80291
0 6502 5 1 1 6501
0 6503 7 1 2 6502 80265
0 6504 5 1 1 6503
0 6505 7 1 2 62883 6504
0 6506 5 1 1 6505
0 6507 7 4 2 64188 72069
0 6508 5 1 1 80995
0 6509 7 2 2 77965 74831
0 6510 5 1 1 80999
0 6511 7 1 2 6508 6510
0 6512 5 3 1 6511
0 6513 7 1 2 67145 81001
0 6514 5 1 1 6513
0 6515 7 1 2 71026 78018
0 6516 5 2 1 6515
0 6517 7 1 2 6514 81004
0 6518 5 1 1 6517
0 6519 7 1 2 69627 6518
0 6520 5 1 1 6519
0 6521 7 1 2 6506 6520
0 6522 5 1 1 6521
0 6523 7 1 2 75505 6522
0 6524 5 1 1 6523
0 6525 7 9 2 62884 63750
0 6526 5 1 1 81006
0 6527 7 1 2 77889 81007
0 6528 7 1 2 77383 6527
0 6529 7 8 2 62597 70919
0 6530 7 7 2 60107 60786
0 6531 7 2 2 81023 80004
0 6532 7 1 2 81015 81030
0 6533 7 1 2 6528 6532
0 6534 5 1 1 6533
0 6535 7 1 2 6524 6534
0 6536 5 1 1 6535
0 6537 7 1 2 65803 76668
0 6538 7 1 2 6536 6537
0 6539 5 1 1 6538
0 6540 7 1 2 6500 6539
0 6541 5 1 1 6540
0 6542 7 1 2 66815 6541
0 6543 5 1 1 6542
0 6544 7 16 2 58181 58401
0 6545 5 1 1 81032
0 6546 7 4 2 63464 73827
0 6547 7 4 2 81033 81048
0 6548 7 3 2 64674 81052
0 6549 5 1 1 81056
0 6550 7 2 2 70762 67985
0 6551 5 2 1 81059
0 6552 7 2 2 70346 69261
0 6553 5 1 1 81063
0 6554 7 1 2 81060 81064
0 6555 5 1 1 6554
0 6556 7 8 2 65448 67986
0 6557 5 11 1 81065
0 6558 7 2 2 71859 79687
0 6559 5 5 1 81084
0 6560 7 1 2 73930 81085
0 6561 5 1 1 6560
0 6562 7 1 2 81073 6561
0 6563 5 2 1 6562
0 6564 7 1 2 81091 69628
0 6565 5 1 1 6564
0 6566 7 1 2 6555 6565
0 6567 5 1 1 6566
0 6568 7 1 2 77126 6567
0 6569 5 1 1 6568
0 6570 7 2 2 69957 75213
0 6571 5 1 1 81093
0 6572 7 1 2 57620 73486
0 6573 5 1 1 6572
0 6574 7 2 2 65449 75893
0 6575 5 5 1 81095
0 6576 7 3 2 6573 81097
0 6577 5 2 1 81102
0 6578 7 1 2 57901 81105
0 6579 5 1 1 6578
0 6580 7 1 2 6571 6579
0 6581 5 1 1 6580
0 6582 7 1 2 69629 6581
0 6583 5 1 1 6582
0 6584 7 1 2 6569 6583
0 6585 5 1 1 6584
0 6586 7 1 2 65804 6585
0 6587 5 1 1 6586
0 6588 7 1 2 60108 68918
0 6589 7 1 2 76590 6588
0 6590 7 1 2 76598 6589
0 6591 5 1 1 6590
0 6592 7 1 2 6587 6591
0 6593 5 1 1 6592
0 6594 7 1 2 81057 6593
0 6595 5 1 1 6594
0 6596 7 1 2 61896 6595
0 6597 7 1 2 6543 6596
0 6598 7 1 2 6326 6597
0 6599 7 1 2 6174 6598
0 6600 5 1 1 6599
0 6601 7 1 2 5316 6600
0 6602 5 1 1 6601
0 6603 7 1 2 66110 6602
0 6604 5 1 1 6603
0 6605 7 1 2 66403 6604
0 6606 7 1 2 4112 6605
0 6607 5 1 1 6606
0 6608 7 1 2 71774 69929
0 6609 5 2 1 6608
0 6610 7 14 2 61505 61897
0 6611 7 5 2 66676 81109
0 6612 7 1 2 70283 81123
0 6613 7 2 2 81107 6612
0 6614 7 1 2 80797 77605
0 6615 7 1 2 81128 6614
0 6616 5 1 1 6615
0 6617 7 1 2 71465 79096
0 6618 5 1 1 6617
0 6619 7 1 2 71146 80487
0 6620 5 1 1 6619
0 6621 7 1 2 6618 6620
0 6622 5 1 1 6621
0 6623 7 1 2 57902 6622
0 6624 5 1 1 6623
0 6625 7 1 2 72947 78755
0 6626 5 1 1 6625
0 6627 7 3 2 59458 73152
0 6628 5 15 1 81130
0 6629 7 1 2 80488 81131
0 6630 5 1 1 6629
0 6631 7 1 2 6626 6630
0 6632 5 1 1 6631
0 6633 7 1 2 58182 6632
0 6634 5 1 1 6633
0 6635 7 1 2 6624 6634
0 6636 5 1 1 6635
0 6637 7 1 2 68324 6636
0 6638 5 2 1 6637
0 6639 7 1 2 79069 72948
0 6640 5 1 1 6639
0 6641 7 1 2 81133 6640
0 6642 5 1 1 6641
0 6643 7 1 2 67833 6642
0 6644 5 1 1 6643
0 6645 7 1 2 59459 74629
0 6646 5 1 1 6645
0 6647 7 1 2 6644 6646
0 6648 5 1 1 6647
0 6649 7 1 2 58183 6648
0 6650 5 1 1 6649
0 6651 7 1 2 57903 71466
0 6652 5 3 1 6651
0 6653 7 1 2 71244 81150
0 6654 5 2 1 6653
0 6655 7 1 2 63833 71245
0 6656 5 2 1 6655
0 6657 7 4 2 62314 71246
0 6658 5 4 1 81157
0 6659 7 2 2 81155 81161
0 6660 5 3 1 81165
0 6661 7 2 2 81153 81166
0 6662 7 2 2 73153 79070
0 6663 5 1 1 81172
0 6664 7 1 2 70192 6663
0 6665 5 2 1 6664
0 6666 7 1 2 81170 81174
0 6667 5 1 1 6666
0 6668 7 1 2 72398 69482
0 6669 5 3 1 6668
0 6670 7 1 2 70151 67834
0 6671 7 2 2 81176 6670
0 6672 5 2 1 81179
0 6673 7 1 2 59460 81180
0 6674 5 1 1 6673
0 6675 7 1 2 6667 6674
0 6676 7 1 2 6650 6675
0 6677 7 1 2 81148 6676
0 6678 5 1 1 6677
0 6679 7 6 2 58402 66111
0 6680 5 4 1 81183
0 6681 7 1 2 67455 81184
0 6682 7 1 2 6678 6681
0 6683 5 1 1 6682
0 6684 7 1 2 6616 6683
0 6685 5 1 1 6684
0 6686 7 1 2 64469 6685
0 6687 5 1 1 6686
0 6688 7 2 2 68820 70106
0 6689 5 1 1 81193
0 6690 7 5 2 75857 6689
0 6691 5 3 1 81195
0 6692 7 1 2 74234 81196
0 6693 5 2 1 6692
0 6694 7 1 2 63152 81106
0 6695 5 2 1 6694
0 6696 7 1 2 63153 73487
0 6697 5 2 1 6696
0 6698 7 1 2 63154 75351
0 6699 5 2 1 6698
0 6700 7 1 2 59264 75417
0 6701 5 1 1 6700
0 6702 7 1 2 74198 6701
0 6703 5 1 1 6702
0 6704 7 1 2 59090 6703
0 6705 5 1 1 6704
0 6706 7 1 2 81209 6705
0 6707 5 1 1 6706
0 6708 7 1 2 57621 6707
0 6709 5 1 1 6708
0 6710 7 1 2 81207 6709
0 6711 5 1 1 6710
0 6712 7 1 2 68728 6711
0 6713 5 1 1 6712
0 6714 7 1 2 81205 6713
0 6715 5 1 1 6714
0 6716 7 1 2 57904 6715
0 6717 5 1 1 6716
0 6718 7 1 2 81203 6717
0 6719 5 1 1 6718
0 6720 7 1 2 64965 6719
0 6721 5 1 1 6720
0 6722 7 1 2 75924 74185
0 6723 5 2 1 6722
0 6724 7 6 2 60257 67635
0 6725 5 2 1 81213
0 6726 7 1 2 74622 81214
0 6727 5 1 1 6726
0 6728 7 1 2 81211 6727
0 6729 5 1 1 6728
0 6730 7 1 2 57905 6729
0 6731 5 1 1 6730
0 6732 7 4 2 59091 73994
0 6733 5 1 1 81221
0 6734 7 1 2 81222 76423
0 6735 5 3 1 6734
0 6736 7 1 2 6731 81225
0 6737 5 1 1 6736
0 6738 7 1 2 68576 6737
0 6739 5 1 1 6738
0 6740 7 2 2 57906 80632
0 6741 5 1 1 81228
0 6742 7 3 2 72057 79688
0 6743 5 6 1 81230
0 6744 7 1 2 81229 81231
0 6745 5 2 1 6744
0 6746 7 2 2 6739 81239
0 6747 5 1 1 81241
0 6748 7 1 2 59461 81226
0 6749 7 1 2 81240 6748
0 6750 7 1 2 81212 6749
0 6751 5 1 1 6750
0 6752 7 1 2 6747 6751
0 6753 5 1 1 6752
0 6754 7 1 2 6721 6753
0 6755 5 1 1 6754
0 6756 7 1 2 58184 66112
0 6757 7 1 2 6755 6756
0 6758 5 1 1 6757
0 6759 7 23 2 58403 61506
0 6760 5 8 1 81243
0 6761 7 1 2 62885 80622
0 6762 5 1 1 6761
0 6763 7 1 2 75858 6762
0 6764 5 1 1 6763
0 6765 7 5 2 76265 513
0 6766 5 1 1 81274
0 6767 7 1 2 81275 74719
0 6768 7 1 2 6764 6767
0 6769 5 1 1 6768
0 6770 7 1 2 75279 6769
0 6771 5 1 1 6770
0 6772 7 2 2 62886 70107
0 6773 5 2 1 81279
0 6774 7 1 2 57907 81281
0 6775 5 2 1 6774
0 6776 7 1 2 70064 81283
0 6777 5 1 1 6776
0 6778 7 1 2 73154 6777
0 6779 5 1 1 6778
0 6780 7 3 2 65178 67835
0 6781 5 1 1 81285
0 6782 7 1 2 58185 81286
0 6783 5 1 1 6782
0 6784 7 1 2 74217 79250
0 6785 5 2 1 6784
0 6786 7 1 2 81276 81288
0 6787 5 1 1 6786
0 6788 7 1 2 68325 6787
0 6789 5 1 1 6788
0 6790 7 1 2 6783 6789
0 6791 7 1 2 6779 6790
0 6792 7 1 2 6771 6791
0 6793 5 1 1 6792
0 6794 7 1 2 81244 6793
0 6795 5 1 1 6794
0 6796 7 1 2 57352 80062
0 6797 5 1 1 6796
0 6798 7 1 2 71718 70957
0 6799 5 2 1 6798
0 6800 7 2 2 6797 81290
0 6801 7 4 2 78832 81292
0 6802 5 3 1 81294
0 6803 7 1 2 81298 78607
0 6804 5 1 1 6803
0 6805 7 8 2 70193 80623
0 6806 7 1 2 80904 81301
0 6807 7 1 2 6804 6806
0 6808 5 1 1 6807
0 6809 7 1 2 58186 6808
0 6810 5 1 1 6809
0 6811 7 1 2 68326 79097
0 6812 5 1 1 6811
0 6813 7 1 2 67636 81175
0 6814 5 1 1 6813
0 6815 7 1 2 6812 6814
0 6816 5 1 1 6815
0 6817 7 1 2 57908 6816
0 6818 5 1 1 6817
0 6819 7 1 2 63155 81181
0 6820 7 1 2 6818 6819
0 6821 7 1 2 6810 6820
0 6822 5 1 1 6821
0 6823 7 2 2 67146 72070
0 6824 5 1 1 81309
0 6825 7 2 2 5618 6824
0 6826 5 1 1 81311
0 6827 7 2 2 58187 77954
0 6828 5 2 1 81313
0 6829 7 3 2 68469 81315
0 6830 5 1 1 81317
0 6831 7 1 2 70316 77624
0 6832 5 1 1 6831
0 6833 7 1 2 62598 6832
0 6834 5 1 1 6833
0 6835 7 1 2 6830 6834
0 6836 5 1 1 6835
0 6837 7 1 2 62315 6836
0 6838 5 1 1 6837
0 6839 7 1 2 81312 6838
0 6840 5 1 1 6839
0 6841 7 1 2 60258 6840
0 6842 5 1 1 6841
0 6843 7 2 2 62599 72488
0 6844 5 1 1 81320
0 6845 7 1 2 62316 72071
0 6846 5 1 1 6845
0 6847 7 1 2 6844 6846
0 6848 5 1 1 6847
0 6849 7 1 2 62887 6848
0 6850 5 1 1 6849
0 6851 7 1 2 73107 77459
0 6852 5 1 1 6851
0 6853 7 1 2 58404 6852
0 6854 7 1 2 6850 6853
0 6855 7 1 2 6842 6854
0 6856 5 1 1 6855
0 6857 7 1 2 66113 6856
0 6858 7 1 2 6822 6857
0 6859 5 1 1 6858
0 6860 7 1 2 6795 6859
0 6861 5 1 1 6860
0 6862 7 1 2 59462 6861
0 6863 5 1 1 6862
0 6864 7 21 2 64189 66114
0 6865 7 1 2 2556 3231
0 6866 5 1 1 6865
0 6867 7 1 2 81322 6866
0 6868 5 1 1 6867
0 6869 7 1 2 64190 67812
0 6870 5 1 1 6869
0 6871 7 1 2 3846 6870
0 6872 5 1 1 6871
0 6873 7 2 2 66115 6872
0 6874 5 1 1 81343
0 6875 7 5 2 61507 68327
0 6876 7 1 2 68577 76145
0 6877 7 1 2 81345 6876
0 6878 5 1 1 6877
0 6879 7 1 2 6874 6878
0 6880 5 1 1 6879
0 6881 7 1 2 65450 6880
0 6882 5 1 1 6881
0 6883 7 1 2 6868 6882
0 6884 5 1 1 6883
0 6885 7 1 2 64966 6884
0 6886 5 1 1 6885
0 6887 7 8 2 59265 61508
0 6888 7 5 2 58188 81350
0 6889 7 1 2 74567 81358
0 6890 5 1 1 6889
0 6891 7 6 2 66116 77974
0 6892 5 1 1 81363
0 6893 7 2 2 63981 68729
0 6894 7 1 2 81364 81369
0 6895 5 1 1 6894
0 6896 7 1 2 6890 6895
0 6897 5 1 1 6896
0 6898 7 1 2 64967 6897
0 6899 5 1 1 6898
0 6900 7 4 2 58954 76576
0 6901 7 4 2 61509 67264
0 6902 7 1 2 73921 81375
0 6903 7 1 2 81371 6902
0 6904 5 1 1 6903
0 6905 7 33 2 60787 66117
0 6906 7 4 2 79483 81379
0 6907 5 1 1 81412
0 6908 7 1 2 57909 81413
0 6909 5 1 1 6908
0 6910 7 1 2 6904 6909
0 6911 7 1 2 6899 6910
0 6912 5 1 1 6911
0 6913 7 1 2 68328 6912
0 6914 5 1 1 6913
0 6915 7 3 2 70699 72827
0 6916 5 1 1 81416
0 6917 7 3 2 61510 73155
0 6918 7 1 2 81417 81419
0 6919 5 1 1 6918
0 6920 7 13 2 58189 61511
0 6921 7 1 2 70152 81422
0 6922 5 2 1 6921
0 6923 7 1 2 68578 81414
0 6924 5 1 1 6923
0 6925 7 1 2 81435 6924
0 6926 5 1 1 6925
0 6927 7 1 2 67836 6926
0 6928 5 1 1 6927
0 6929 7 1 2 6919 6928
0 6930 7 1 2 6914 6929
0 6931 7 1 2 6886 6930
0 6932 5 1 1 6931
0 6933 7 1 2 65179 6932
0 6934 5 1 1 6933
0 6935 7 1 2 68329 81415
0 6936 5 1 1 6935
0 6937 7 1 2 70194 1262
0 6938 5 2 1 6937
0 6939 7 10 2 64968 61512
0 6940 5 1 1 81439
0 6941 7 1 2 58190 81440
0 6942 7 1 2 81437 6941
0 6943 5 1 1 6942
0 6944 7 1 2 6936 6943
0 6945 5 1 1 6944
0 6946 7 1 2 68579 6945
0 6947 5 1 1 6946
0 6948 7 1 2 81420 81372
0 6949 5 1 1 6948
0 6950 7 1 2 6907 6949
0 6951 5 1 1 6950
0 6952 7 1 2 67637 6951
0 6953 5 1 1 6952
0 6954 7 1 2 74512 81365
0 6955 5 1 1 6954
0 6956 7 1 2 81436 6955
0 6957 5 1 1 6956
0 6958 7 1 2 72272 6957
0 6959 5 1 1 6958
0 6960 7 1 2 6953 6959
0 6961 7 1 2 6947 6960
0 6962 5 1 1 6961
0 6963 7 1 2 57910 6962
0 6964 5 1 1 6963
0 6965 7 3 2 67638 75165
0 6966 5 7 1 81449
0 6967 7 1 2 62888 81452
0 6968 5 2 1 6967
0 6969 7 16 2 60504 66118
0 6970 7 1 2 77975 81461
0 6971 7 1 2 81459 6970
0 6972 5 1 1 6971
0 6973 7 1 2 76275 81359
0 6974 7 1 2 80280 6973
0 6975 5 1 1 6974
0 6976 7 1 2 6972 6975
0 6977 7 1 2 6964 6976
0 6978 7 1 2 6934 6977
0 6979 5 1 1 6978
0 6980 7 1 2 58405 6979
0 6981 5 1 1 6980
0 6982 7 1 2 6863 6981
0 6983 7 1 2 6758 6982
0 6984 5 1 1 6983
0 6985 7 2 2 59748 66553
0 6986 7 1 2 62046 81477
0 6987 7 1 2 6984 6986
0 6988 5 1 1 6987
0 6989 7 1 2 6687 6988
0 6990 5 1 1 6989
0 6991 7 1 2 66816 6990
0 6992 5 1 1 6991
0 6993 7 1 2 62889 69899
0 6994 5 1 1 6993
0 6995 7 6 2 57911 63982
0 6996 5 1 1 81479
0 6997 7 1 2 71719 81480
0 6998 5 1 1 6997
0 6999 7 1 2 6994 6998
0 7000 5 1 1 6999
0 7001 7 1 2 60788 7000
0 7002 5 1 1 7001
0 7003 7 3 2 62890 71990
0 7004 5 1 1 81485
0 7005 7 1 2 58955 81486
0 7006 5 1 1 7005
0 7007 7 1 2 7002 7006
0 7008 5 2 1 7007
0 7009 7 1 2 81323 81488
0 7010 5 1 1 7009
0 7011 7 24 2 65451 61513
0 7012 7 4 2 59266 81490
0 7013 7 1 2 71577 81514
0 7014 5 1 1 7013
0 7015 7 1 2 7010 7014
0 7016 5 1 1 7015
0 7017 7 1 2 57353 7016
0 7018 5 1 1 7017
0 7019 7 2 2 69771 79838
0 7020 7 1 2 81380 81518
0 7021 5 1 1 7020
0 7022 7 4 2 58191 71720
0 7023 5 2 1 81520
0 7024 7 1 2 81521 81515
0 7025 5 1 1 7024
0 7026 7 1 2 7021 7025
0 7027 5 1 1 7026
0 7028 7 1 2 57912 7027
0 7029 5 1 1 7028
0 7030 7 1 2 7018 7029
0 7031 5 1 1 7030
0 7032 7 1 2 57622 7031
0 7033 5 1 1 7032
0 7034 7 6 2 58192 59267
0 7035 5 3 1 81526
0 7036 7 2 2 76322 81527
0 7037 5 1 1 81535
0 7038 7 2 2 61514 75166
0 7039 7 1 2 81536 81537
0 7040 5 1 1 7039
0 7041 7 1 2 7033 7040
0 7042 5 1 1 7041
0 7043 7 1 2 71860 7042
0 7044 5 1 1 7043
0 7045 7 1 2 73488 78204
0 7046 5 2 1 7045
0 7047 7 2 2 69958 73793
0 7048 5 2 1 81541
0 7049 7 1 2 81539 81543
0 7050 5 1 1 7049
0 7051 7 1 2 81423 7050
0 7052 5 1 1 7051
0 7053 7 1 2 74353 75136
0 7054 5 1 1 7053
0 7055 7 1 2 80126 81532
0 7056 5 1 1 7055
0 7057 7 1 2 7054 7056
0 7058 5 1 1 7057
0 7059 7 3 2 66119 71721
0 7060 7 1 2 64191 81545
0 7061 7 1 2 7058 7060
0 7062 5 1 1 7061
0 7063 7 1 2 7052 7062
0 7064 5 1 1 7063
0 7065 7 1 2 57913 7064
0 7066 5 1 1 7065
0 7067 7 14 2 66120 71389
0 7068 7 1 2 72697 80175
0 7069 5 1 1 7068
0 7070 7 1 2 72387 74391
0 7071 5 1 1 7070
0 7072 7 1 2 7069 7071
0 7073 5 1 1 7072
0 7074 7 1 2 81548 7073
0 7075 5 1 1 7074
0 7076 7 2 2 74322 81491
0 7077 7 1 2 74807 81528
0 7078 7 1 2 81562 7077
0 7079 5 1 1 7078
0 7080 7 1 2 7075 7079
0 7081 5 1 1 7080
0 7082 7 1 2 59092 7081
0 7083 5 1 1 7082
0 7084 7 1 2 7066 7083
0 7085 5 1 1 7084
0 7086 7 1 2 57354 7085
0 7087 5 1 1 7086
0 7088 7 7 2 64969 66121
0 7089 7 2 2 81564 80176
0 7090 7 2 2 73346 69779
0 7091 7 1 2 81571 81573
0 7092 5 1 1 7091
0 7093 7 1 2 78309 75046
0 7094 5 1 1 7093
0 7095 7 2 2 62891 72489
0 7096 5 1 1 81575
0 7097 7 2 2 69022 68221
0 7098 5 7 1 81577
0 7099 7 1 2 73156 81579
0 7100 7 1 2 81576 7099
0 7101 5 1 1 7100
0 7102 7 1 2 7094 7101
0 7103 5 1 1 7102
0 7104 7 1 2 81324 7103
0 7105 5 1 1 7104
0 7106 7 2 2 65452 78191
0 7107 5 2 1 81586
0 7108 7 2 2 70763 81587
0 7109 5 1 1 81590
0 7110 7 1 2 81360 81591
0 7111 5 1 1 7110
0 7112 7 1 2 7105 7111
0 7113 5 1 1 7112
0 7114 7 1 2 57914 7113
0 7115 5 1 1 7114
0 7116 7 1 2 7092 7115
0 7117 7 1 2 7087 7116
0 7118 7 2 2 7044 7117
0 7119 7 2 2 63834 69440
0 7120 5 11 1 81594
0 7121 7 1 2 57355 81596
0 7122 5 2 1 7121
0 7123 7 3 2 60259 76557
0 7124 5 6 1 81609
0 7125 7 5 2 63835 80510
0 7126 5 2 1 81618
0 7127 7 1 2 81612 81623
0 7128 5 4 1 7127
0 7129 7 1 2 81607 81625
0 7130 5 1 1 7129
0 7131 7 1 2 57623 7130
0 7132 5 1 1 7131
0 7133 7 3 2 79127 7132
0 7134 5 9 1 81629
0 7135 7 1 2 67265 81632
0 7136 5 2 1 7135
0 7137 7 1 2 65453 81633
0 7138 5 2 1 7137
0 7139 7 1 2 73157 80951
0 7140 5 1 1 7139
0 7141 7 1 2 78747 79010
0 7142 7 1 2 7140 7141
0 7143 7 1 2 81643 7142
0 7144 7 1 2 81641 7143
0 7145 5 2 1 7144
0 7146 7 1 2 58193 81645
0 7147 5 1 1 7146
0 7148 7 2 2 77440 72375
0 7149 5 1 1 81647
0 7150 7 1 2 75352 81648
0 7151 5 1 1 7150
0 7152 7 1 2 7147 7151
0 7153 5 1 1 7152
0 7154 7 1 2 61515 7153
0 7155 5 2 1 7154
0 7156 7 9 2 62892 63836
0 7157 5 2 1 81651
0 7158 7 2 2 62600 81652
0 7159 7 1 2 71991 81662
0 7160 5 1 1 7159
0 7161 7 1 2 58194 71796
0 7162 5 1 1 7161
0 7163 7 1 2 75362 7162
0 7164 5 1 1 7163
0 7165 7 8 2 63751 60789
0 7166 5 2 1 81664
0 7167 7 1 2 81665 80138
0 7168 7 1 2 7164 7167
0 7169 5 1 1 7168
0 7170 7 1 2 7160 7169
0 7171 5 1 1 7170
0 7172 7 1 2 62317 7171
0 7173 5 1 1 7172
0 7174 7 3 2 62601 79768
0 7175 7 2 2 63983 70284
0 7176 7 1 2 81674 81677
0 7177 5 1 1 7176
0 7178 7 1 2 7173 7177
0 7179 5 1 1 7178
0 7180 7 1 2 66122 7179
0 7181 5 1 1 7180
0 7182 7 1 2 81649 7181
0 7183 5 1 1 7182
0 7184 7 1 2 59463 7183
0 7185 5 1 1 7184
0 7186 7 1 2 81592 7185
0 7187 5 1 1 7186
0 7188 7 1 2 59749 7187
0 7189 5 1 1 7188
0 7190 7 1 2 67837 78631
0 7191 5 2 1 7190
0 7192 7 1 2 77656 81679
0 7193 5 1 1 7192
0 7194 7 1 2 80177 7193
0 7195 5 2 1 7194
0 7196 7 1 2 67639 72134
0 7197 5 2 1 7196
0 7198 7 2 2 58956 74392
0 7199 7 1 2 57356 81685
0 7200 5 1 1 7199
0 7201 7 1 2 81683 7200
0 7202 5 1 1 7201
0 7203 7 1 2 57915 7202
0 7204 5 1 1 7203
0 7205 7 1 2 81681 7204
0 7206 5 1 1 7205
0 7207 7 1 2 59464 7206
0 7208 5 1 1 7207
0 7209 7 1 2 74529 80281
0 7210 5 1 1 7209
0 7211 7 6 2 57357 69319
0 7212 5 1 1 81687
0 7213 7 1 2 70153 81688
0 7214 5 1 1 7213
0 7215 7 1 2 7210 7214
0 7216 5 1 1 7215
0 7217 7 1 2 57916 7216
0 7218 5 1 1 7217
0 7219 7 10 2 58957 59465
0 7220 5 6 1 81693
0 7221 7 3 2 57358 81694
0 7222 5 2 1 81709
0 7223 7 1 2 74393 81710
0 7224 5 1 1 7223
0 7225 7 1 2 7218 7224
0 7226 5 1 1 7225
0 7227 7 1 2 75859 7226
0 7228 5 1 1 7227
0 7229 7 1 2 74568 72376
0 7230 7 1 2 80167 7229
0 7231 5 1 1 7230
0 7232 7 1 2 7228 7231
0 7233 7 1 2 7208 7232
0 7234 5 2 1 7233
0 7235 7 2 2 66123 81714
0 7236 7 1 2 77229 81716
0 7237 5 1 1 7236
0 7238 7 1 2 7189 7237
0 7239 5 1 1 7238
0 7240 7 1 2 58406 7239
0 7241 5 1 1 7240
0 7242 7 1 2 59750 77776
0 7243 7 1 2 81717 7242
0 7244 5 1 1 7243
0 7245 7 1 2 7241 7244
0 7246 5 1 1 7245
0 7247 7 1 2 74405 7246
0 7248 5 1 1 7247
0 7249 7 1 2 6992 7248
0 7250 5 1 1 7249
0 7251 7 1 2 70480 7250
0 7252 5 1 1 7251
0 7253 7 5 2 57359 61898
0 7254 7 3 2 66817 81718
0 7255 5 2 1 81723
0 7256 7 2 2 76016 74427
0 7257 5 1 1 81728
0 7258 7 1 2 75989 7257
0 7259 5 3 1 7258
0 7260 7 1 2 57624 81730
0 7261 5 1 1 7260
0 7262 7 2 2 81726 7261
0 7263 7 1 2 67593 75746
0 7264 5 1 1 7263
0 7265 7 1 2 75668 7264
0 7266 5 2 1 7265
0 7267 7 1 2 71722 81735
0 7268 5 1 1 7267
0 7269 7 1 2 81733 7268
0 7270 5 1 1 7269
0 7271 7 1 2 57917 7270
0 7272 5 1 1 7271
0 7273 7 6 2 57625 58721
0 7274 7 3 2 75950 81737
0 7275 5 3 1 81743
0 7276 7 1 2 75167 81744
0 7277 5 1 1 7276
0 7278 7 1 2 7272 7277
0 7279 5 1 1 7278
0 7280 7 1 2 71861 7279
0 7281 5 1 1 7280
0 7282 7 1 2 57918 75829
0 7283 5 1 1 7282
0 7284 7 1 2 73893 81724
0 7285 5 1 1 7284
0 7286 7 1 2 7283 7285
0 7287 5 1 1 7286
0 7288 7 1 2 78310 7287
0 7289 5 1 1 7288
0 7290 7 3 2 74218 75747
0 7291 5 1 1 81749
0 7292 7 1 2 70700 81750
0 7293 5 1 1 7292
0 7294 7 1 2 77692 75971
0 7295 5 1 1 7294
0 7296 7 1 2 7293 7295
0 7297 5 1 1 7296
0 7298 7 1 2 71723 7297
0 7299 5 1 1 7298
0 7300 7 7 2 59974 65180
0 7301 7 2 2 61899 81752
0 7302 7 1 2 57919 74822
0 7303 7 1 2 81759 7302
0 7304 5 1 1 7303
0 7305 7 1 2 7299 7304
0 7306 7 1 2 7289 7305
0 7307 7 1 2 7281 7306
0 7308 5 1 1 7307
0 7309 7 1 2 69630 7308
0 7310 5 1 1 7309
0 7311 7 10 2 69262 75972
0 7312 7 2 2 57920 78743
0 7313 5 2 1 81771
0 7314 7 1 2 81761 81772
0 7315 5 1 1 7314
0 7316 7 1 2 7310 7315
0 7317 5 1 1 7316
0 7318 7 1 2 73158 7317
0 7319 5 2 1 7318
0 7320 7 4 2 66818 69160
0 7321 5 3 1 81777
0 7322 7 2 2 67838 75748
0 7323 7 1 2 57360 81784
0 7324 5 1 1 7323
0 7325 7 1 2 81781 7324
0 7326 5 1 1 7325
0 7327 7 1 2 71724 7326
0 7328 5 1 1 7327
0 7329 7 1 2 68984 81785
0 7330 5 1 1 7329
0 7331 7 1 2 67813 69483
0 7332 5 1 1 7331
0 7333 7 1 2 75619 7332
0 7334 5 1 1 7333
0 7335 7 1 2 7330 7334
0 7336 7 1 2 7328 7335
0 7337 5 1 1 7336
0 7338 7 1 2 70154 7337
0 7339 5 1 1 7338
0 7340 7 3 2 74237 72576
0 7341 5 1 1 81786
0 7342 7 2 2 75691 69161
0 7343 7 4 2 58722 58958
0 7344 7 1 2 57361 81791
0 7345 7 1 2 81789 7344
0 7346 5 1 1 7345
0 7347 7 1 2 7341 7346
0 7348 5 1 1 7347
0 7349 7 1 2 57921 7348
0 7350 5 1 1 7349
0 7351 7 1 2 80489 75973
0 7352 5 1 1 7351
0 7353 7 1 2 76538 75749
0 7354 5 1 1 7353
0 7355 7 1 2 7352 7354
0 7356 5 1 1 7355
0 7357 7 1 2 70155 7356
0 7358 5 1 1 7357
0 7359 7 1 2 7350 7358
0 7360 5 1 1 7359
0 7361 7 1 2 68330 7360
0 7362 5 1 1 7361
0 7363 7 3 2 59093 69450
0 7364 5 7 1 81795
0 7365 7 1 2 76594 75974
0 7366 7 1 2 81796 7365
0 7367 5 1 1 7366
0 7368 7 3 2 59094 59975
0 7369 7 4 2 81805 81738
0 7370 7 1 2 76442 69162
0 7371 7 1 2 81808 7370
0 7372 5 1 1 7371
0 7373 7 1 2 7367 7372
0 7374 7 1 2 7362 7373
0 7375 7 1 2 7339 7374
0 7376 5 1 1 7375
0 7377 7 1 2 69631 7376
0 7378 5 1 1 7377
0 7379 7 1 2 81775 7378
0 7380 5 1 1 7379
0 7381 7 1 2 59466 7380
0 7382 5 1 1 7381
0 7383 7 1 2 61516 7382
0 7384 5 1 1 7383
0 7385 7 1 2 77204 74912
0 7386 5 1 1 7385
0 7387 7 1 2 75669 7386
0 7388 5 2 1 7387
0 7389 7 1 2 68470 81812
0 7390 5 2 1 7389
0 7391 7 3 2 58723 60505
0 7392 5 2 1 81816
0 7393 7 2 2 75951 81817
0 7394 5 1 1 81821
0 7395 7 2 2 81814 7394
0 7396 5 1 1 81823
0 7397 7 1 2 60790 7396
0 7398 5 1 1 7397
0 7399 7 1 2 77281 77637
0 7400 5 1 1 7399
0 7401 7 1 2 7398 7400
0 7402 5 1 1 7401
0 7403 7 1 2 63837 7402
0 7404 5 1 1 7403
0 7405 7 3 2 64675 77638
0 7406 7 2 2 66554 76521
0 7407 7 1 2 81825 81828
0 7408 5 1 1 7407
0 7409 7 1 2 7404 7408
0 7410 5 1 1 7409
0 7411 7 1 2 62318 7410
0 7412 5 1 1 7411
0 7413 7 2 2 58195 75405
0 7414 5 1 1 81830
0 7415 7 1 2 77294 7414
0 7416 5 1 1 7415
0 7417 7 9 2 63838 69379
0 7418 5 7 1 81832
0 7419 7 1 2 67266 81841
0 7420 5 1 1 7419
0 7421 7 1 2 75620 7420
0 7422 5 1 1 7421
0 7423 7 1 2 7416 7422
0 7424 5 1 1 7423
0 7425 7 1 2 60791 7424
0 7426 5 1 1 7425
0 7427 7 4 2 62893 71797
0 7428 5 1 1 81848
0 7429 7 3 2 58196 80206
0 7430 5 6 1 81852
0 7431 7 1 2 62602 81855
0 7432 5 2 1 7431
0 7433 7 1 2 7428 81861
0 7434 5 2 1 7433
0 7435 7 1 2 60260 81863
0 7436 5 2 1 7435
0 7437 7 1 2 81865 5279
0 7438 5 1 1 7437
0 7439 7 1 2 77248 7438
0 7440 5 1 1 7439
0 7441 7 1 2 7426 7440
0 7442 7 1 2 7412 7441
0 7443 5 1 1 7442
0 7444 7 1 2 69632 7443
0 7445 5 1 1 7444
0 7446 7 11 2 59467 66124
0 7447 5 1 1 81867
0 7448 7 7 2 58847 64676
0 7449 7 7 2 63465 81878
0 7450 5 1 1 81885
0 7451 7 7 2 60792 66555
0 7452 7 4 2 69332 81892
0 7453 5 1 1 81899
0 7454 7 1 2 81886 81900
0 7455 5 2 1 7454
0 7456 7 2 2 72135 81762
0 7457 5 1 1 81905
0 7458 7 4 2 69333 79957
0 7459 5 1 1 81907
0 7460 7 8 2 60261 66556
0 7461 7 5 2 64677 81911
0 7462 7 1 2 81908 81919
0 7463 5 3 1 7462
0 7464 7 1 2 7457 81924
0 7465 5 1 1 7464
0 7466 7 1 2 68471 7465
0 7467 5 1 1 7466
0 7468 7 1 2 81903 7467
0 7469 5 1 1 7468
0 7470 7 1 2 63984 7469
0 7471 5 1 1 7470
0 7472 7 2 2 80005 81893
0 7473 7 1 2 79964 81927
0 7474 5 1 1 7473
0 7475 7 3 2 69516 77301
0 7476 7 1 2 75137 67508
0 7477 7 1 2 81929 7476
0 7478 5 1 1 7477
0 7479 7 1 2 7474 7478
0 7480 5 1 1 7479
0 7481 7 1 2 60262 7480
0 7482 5 1 1 7481
0 7483 7 1 2 7471 7482
0 7484 5 1 1 7483
0 7485 7 1 2 77460 7484
0 7486 5 1 1 7485
0 7487 7 1 2 81868 7486
0 7488 7 1 2 7445 7487
0 7489 5 1 1 7488
0 7490 7 5 2 57922 60263
0 7491 5 4 1 81932
0 7492 7 2 2 68985 78547
0 7493 5 1 1 81941
0 7494 7 1 2 81937 7493
0 7495 5 1 1 7494
0 7496 7 1 2 57362 7495
0 7497 5 1 1 7496
0 7498 7 2 2 74354 81613
0 7499 7 1 2 57923 81943
0 7500 5 1 1 7499
0 7501 7 1 2 7497 7500
0 7502 5 3 1 7501
0 7503 7 1 2 81945 77249
0 7504 5 1 1 7503
0 7505 7 7 2 69441 75260
0 7506 5 11 1 81948
0 7507 7 1 2 81955 75621
0 7508 5 1 1 7507
0 7509 7 1 2 7504 7508
0 7510 5 1 1 7509
0 7511 7 1 2 68331 7510
0 7512 5 1 1 7511
0 7513 7 1 2 80502 68924
0 7514 5 1 1 7513
0 7515 7 1 2 75229 7514
0 7516 5 2 1 7515
0 7517 7 1 2 81966 77250
0 7518 5 1 1 7517
0 7519 7 1 2 75990 7518
0 7520 5 1 1 7519
0 7521 7 1 2 67839 7520
0 7522 5 1 1 7521
0 7523 7 1 2 77127 81778
0 7524 5 1 1 7523
0 7525 7 4 2 59095 64678
0 7526 5 1 1 81968
0 7527 7 1 2 81912 81969
0 7528 7 1 2 76099 7527
0 7529 5 1 1 7528
0 7530 7 1 2 7524 7529
0 7531 7 1 2 7522 7530
0 7532 7 1 2 7512 7531
0 7533 5 1 1 7532
0 7534 7 1 2 60793 7533
0 7535 5 1 1 7534
0 7536 7 3 2 64679 65181
0 7537 5 1 1 81972
0 7538 7 3 2 71358 81973
0 7539 7 3 2 62894 75802
0 7540 5 1 1 81978
0 7541 7 6 2 63466 65454
0 7542 5 1 1 81981
0 7543 7 1 2 67814 81982
0 7544 5 1 1 7543
0 7545 7 1 2 7540 7544
0 7546 5 1 1 7545
0 7547 7 1 2 81975 7546
0 7548 5 1 1 7547
0 7549 7 1 2 70706 75622
0 7550 5 2 1 7549
0 7551 7 3 2 74323 75750
0 7552 5 1 1 81989
0 7553 7 1 2 75991 7552
0 7554 5 1 1 7553
0 7555 7 1 2 62895 7554
0 7556 5 1 1 7555
0 7557 7 1 2 81987 7556
0 7558 5 1 1 7557
0 7559 7 1 2 65455 7558
0 7560 5 1 1 7559
0 7561 7 1 2 7548 7560
0 7562 7 1 2 7535 7561
0 7563 5 1 1 7562
0 7564 7 1 2 69633 7563
0 7565 5 1 1 7564
0 7566 7 1 2 57363 81489
0 7567 5 1 1 7566
0 7568 7 2 2 63985 78677
0 7569 5 2 1 81992
0 7570 7 1 2 79791 81993
0 7571 5 1 1 7570
0 7572 7 1 2 7567 7571
0 7573 5 1 1 7572
0 7574 7 1 2 75860 7573
0 7575 5 1 1 7574
0 7576 7 1 2 72816 81686
0 7577 5 1 1 7576
0 7578 7 1 2 81682 7577
0 7579 5 1 1 7578
0 7580 7 1 2 62896 7579
0 7581 5 1 1 7580
0 7582 7 1 2 76530 79354
0 7583 5 1 1 7582
0 7584 7 1 2 7581 7583
0 7585 7 1 2 7575 7584
0 7586 5 1 1 7585
0 7587 7 1 2 75623 7586
0 7588 5 1 1 7587
0 7589 7 1 2 57626 77279
0 7590 7 1 2 80722 7589
0 7591 5 1 1 7590
0 7592 7 1 2 7588 7591
0 7593 5 1 1 7592
0 7594 7 1 2 69263 7593
0 7595 5 1 1 7594
0 7596 7 1 2 64192 7595
0 7597 7 1 2 7565 7596
0 7598 5 1 1 7597
0 7599 7 1 2 7489 7598
0 7600 5 1 1 7599
0 7601 7 10 2 64970 72466
0 7602 5 4 1 81996
0 7603 7 19 2 62047 67434
0 7604 5 1 1 82010
0 7605 7 3 2 81997 82011
0 7606 7 2 2 67147 81879
0 7607 7 1 2 77639 82032
0 7608 7 1 2 82029 7607
0 7609 5 1 1 7608
0 7610 7 1 2 7600 7609
0 7611 5 1 1 7610
0 7612 7 1 2 7384 7611
0 7613 5 1 1 7612
0 7614 7 5 2 58848 67950
0 7615 7 2 2 57924 58724
0 7616 7 2 2 76604 82039
0 7617 7 1 2 82034 82041
0 7618 7 2 2 80909 7617
0 7619 5 1 1 82043
0 7620 7 1 2 81516 82044
0 7621 5 1 1 7620
0 7622 7 2 2 75727 76094
0 7623 5 2 1 82045
0 7624 7 1 2 82047 81734
0 7625 5 1 1 7624
0 7626 7 1 2 69634 7625
0 7627 5 1 1 7626
0 7628 7 3 2 74245 67616
0 7629 5 2 1 82049
0 7630 7 3 2 75728 74501
0 7631 7 1 2 69350 82054
0 7632 5 1 1 7631
0 7633 7 3 2 75952 82040
0 7634 5 1 1 82057
0 7635 7 1 2 69264 82058
0 7636 5 1 1 7635
0 7637 7 1 2 7632 7636
0 7638 5 1 1 7637
0 7639 7 1 2 57627 7638
0 7640 5 1 1 7639
0 7641 7 1 2 82052 7640
0 7642 5 1 1 7641
0 7643 7 1 2 71725 7642
0 7644 5 1 1 7643
0 7645 7 2 2 78311 67509
0 7646 7 9 2 76022 76103
0 7647 5 1 1 82062
0 7648 7 1 2 82063 72817
0 7649 7 1 2 82060 7648
0 7650 5 1 1 7649
0 7651 7 1 2 7644 7650
0 7652 7 1 2 7627 7651
0 7653 5 1 1 7652
0 7654 7 1 2 71862 7653
0 7655 5 1 1 7654
0 7656 7 3 2 68730 76104
0 7657 7 1 2 76040 82071
0 7658 5 1 1 7657
0 7659 7 1 2 76136 7658
0 7660 5 1 1 7659
0 7661 7 2 2 57628 7660
0 7662 5 1 1 82074
0 7663 7 1 2 60264 76137
0 7664 5 1 1 7663
0 7665 7 1 2 82075 7664
0 7666 5 1 1 7665
0 7667 7 1 2 75280 77251
0 7668 5 1 1 7667
0 7669 7 1 2 75992 7668
0 7670 5 1 1 7669
0 7671 7 1 2 69635 7670
0 7672 5 1 1 7671
0 7673 7 1 2 7666 7672
0 7674 5 1 1 7673
0 7675 7 1 2 73894 7674
0 7676 5 1 1 7675
0 7677 7 1 2 78358 68680
0 7678 5 1 1 7677
0 7679 7 1 2 71775 73397
0 7680 7 1 2 80150 7679
0 7681 5 1 1 7680
0 7682 7 1 2 7678 7681
0 7683 5 1 1 7682
0 7684 7 1 2 75624 7683
0 7685 5 1 1 7684
0 7686 7 1 2 7676 7685
0 7687 7 1 2 7655 7686
0 7688 5 1 1 7687
0 7689 7 1 2 70156 7688
0 7690 5 1 1 7689
0 7691 7 1 2 7619 7690
0 7692 7 1 2 81776 7691
0 7693 5 1 1 7692
0 7694 7 1 2 61517 7693
0 7695 5 1 1 7694
0 7696 7 3 2 69916 81462
0 7697 7 1 2 75993 3455
0 7698 5 1 1 7697
0 7699 7 1 2 74832 7698
0 7700 5 1 1 7699
0 7701 7 1 2 3438 7700
0 7702 5 1 1 7701
0 7703 7 1 2 82076 7702
0 7704 5 1 1 7703
0 7705 7 1 2 70764 72698
0 7706 5 3 1 7705
0 7707 7 1 2 58959 70128
0 7708 5 1 1 7707
0 7709 7 1 2 82079 7708
0 7710 5 2 1 7709
0 7711 7 1 2 67009 69085
0 7712 5 4 1 7711
0 7713 7 1 2 62160 82084
0 7714 5 1 1 7713
0 7715 7 2 2 82082 7714
0 7716 7 25 2 61518 66557
0 7717 7 6 2 64680 82090
0 7718 7 1 2 76095 82115
0 7719 7 1 2 82088 7718
0 7720 5 1 1 7719
0 7721 7 1 2 7704 7720
0 7722 5 1 1 7721
0 7723 7 1 2 60794 7722
0 7724 5 1 1 7723
0 7725 7 4 2 60795 67148
0 7726 5 6 1 82121
0 7727 7 1 2 2748 80624
0 7728 5 1 1 7727
0 7729 7 2 2 82125 7728
0 7730 5 1 1 82131
0 7731 7 1 2 75625 82132
0 7732 5 1 1 7731
0 7733 7 3 2 63467 74847
0 7734 7 2 2 62319 82133
0 7735 7 3 2 63839 69959
0 7736 5 1 1 82138
0 7737 7 1 2 72577 82139
0 7738 7 1 2 82136 7737
0 7739 5 1 1 7738
0 7740 7 1 2 7732 7739
0 7741 5 1 1 7740
0 7742 7 1 2 68580 7741
0 7743 5 1 1 7742
0 7744 7 2 2 67640 78608
0 7745 5 2 1 82141
0 7746 7 2 2 82143 81302
0 7747 5 1 1 82145
0 7748 7 2 2 67149 79511
0 7749 5 2 1 82147
0 7750 7 1 2 70077 82149
0 7751 5 1 1 7750
0 7752 7 1 2 82146 7751
0 7753 5 1 1 7752
0 7754 7 1 2 75626 7753
0 7755 5 1 1 7754
0 7756 7 10 2 60265 68731
0 7757 5 2 1 82151
0 7758 7 2 2 63840 82152
0 7759 5 1 1 82163
0 7760 7 1 2 81787 82164
0 7761 5 1 1 7760
0 7762 7 1 2 7755 7761
0 7763 5 1 1 7762
0 7764 7 1 2 65182 7763
0 7765 5 1 1 7764
0 7766 7 1 2 75696 7747
0 7767 5 1 1 7766
0 7768 7 2 2 76323 75751
0 7769 5 1 1 82165
0 7770 7 1 2 60506 82153
0 7771 7 1 2 82166 7770
0 7772 5 1 1 7771
0 7773 7 3 2 64971 71619
0 7774 5 3 1 82167
0 7775 7 1 2 80625 82170
0 7776 5 1 1 7775
0 7777 7 1 2 78609 75975
0 7778 7 1 2 7776 7777
0 7779 5 1 1 7778
0 7780 7 1 2 7772 7779
0 7781 5 1 1 7780
0 7782 7 1 2 68332 7781
0 7783 5 1 1 7782
0 7784 7 1 2 7767 7783
0 7785 7 1 2 7765 7784
0 7786 7 1 2 7743 7785
0 7787 5 1 1 7786
0 7788 7 1 2 61519 7787
0 7789 5 1 1 7788
0 7790 7 1 2 7724 7789
0 7791 5 1 1 7790
0 7792 7 1 2 69265 7791
0 7793 5 1 1 7792
0 7794 7 1 2 71863 81736
0 7795 5 1 1 7794
0 7796 7 2 2 67150 73452
0 7797 5 2 1 82173
0 7798 7 1 2 82175 82055
0 7799 5 1 1 7798
0 7800 7 1 2 7799 81746
0 7801 7 1 2 7795 7800
0 7802 5 1 1 7801
0 7803 7 1 2 71726 7802
0 7804 5 1 1 7803
0 7805 7 1 2 82126 75752
0 7806 5 1 1 7805
0 7807 7 1 2 81727 7806
0 7808 5 1 1 7807
0 7809 7 1 2 80063 7808
0 7810 5 1 1 7809
0 7811 7 1 2 75861 81731
0 7812 5 1 1 7811
0 7813 7 1 2 75994 82048
0 7814 5 1 1 7813
0 7815 7 1 2 73159 7814
0 7816 5 1 1 7815
0 7817 7 3 2 57629 75824
0 7818 7 1 2 75820 82177
0 7819 5 1 1 7818
0 7820 7 1 2 7634 7819
0 7821 7 1 2 7816 7820
0 7822 7 1 2 7812 7821
0 7823 7 1 2 7810 7822
0 7824 7 1 2 7804 7823
0 7825 5 1 1 7824
0 7826 7 7 2 61520 62048
0 7827 7 1 2 67915 82180
0 7828 7 1 2 7825 7827
0 7829 5 1 1 7828
0 7830 7 1 2 7793 7829
0 7831 5 1 1 7830
0 7832 7 1 2 59468 7831
0 7833 5 1 1 7832
0 7834 7 4 2 66125 66746
0 7835 7 1 2 82187 72684
0 7836 7 1 2 75418 7835
0 7837 5 1 1 7836
0 7838 7 1 2 7833 7837
0 7839 7 1 2 7695 7838
0 7840 5 1 1 7839
0 7841 7 1 2 58197 7840
0 7842 5 1 1 7841
0 7843 7 1 2 7621 7842
0 7844 7 1 2 7613 7843
0 7845 5 1 1 7844
0 7846 7 1 2 59751 7845
0 7847 5 1 1 7846
0 7848 7 29 2 64470 66126
0 7849 5 5 1 82191
0 7850 7 2 2 77128 75627
0 7851 5 2 1 82225
0 7852 7 1 2 62161 75670
0 7853 5 1 1 7852
0 7854 7 3 2 81732 7853
0 7855 7 1 2 57630 82229
0 7856 5 1 1 7855
0 7857 7 1 2 82227 7856
0 7858 5 1 1 7857
0 7859 7 1 2 73160 7858
0 7860 5 1 1 7859
0 7861 7 1 2 71037 81788
0 7862 5 1 1 7861
0 7863 7 1 2 7860 7862
0 7864 5 1 1 7863
0 7865 7 1 2 57925 7864
0 7866 5 1 1 7865
0 7867 7 2 2 78302 75261
0 7868 5 9 1 82232
0 7869 7 1 2 82234 77563
0 7870 5 1 1 7869
0 7871 7 1 2 7866 7870
0 7872 5 1 1 7871
0 7873 7 2 2 58849 59469
0 7874 7 6 2 69334 82243
0 7875 5 1 1 82245
0 7876 7 1 2 7872 82246
0 7877 5 1 1 7876
0 7878 7 1 2 76017 81909
0 7879 5 3 1 7878
0 7880 7 1 2 71992 81763
0 7881 5 1 1 7880
0 7882 7 1 2 82251 7881
0 7883 5 1 1 7882
0 7884 7 1 2 57631 7883
0 7885 5 1 1 7884
0 7886 7 1 2 82053 7885
0 7887 5 1 1 7886
0 7888 7 1 2 58960 7887
0 7889 5 1 1 7888
0 7890 7 2 2 75729 81983
0 7891 5 2 1 82254
0 7892 7 1 2 75701 82256
0 7893 5 1 1 7892
0 7894 7 1 2 69636 7893
0 7895 5 1 1 7894
0 7896 7 1 2 7889 7895
0 7897 5 1 1 7896
0 7898 7 1 2 57364 7897
0 7899 5 1 1 7898
0 7900 7 1 2 75995 82257
0 7901 5 1 1 7900
0 7902 7 1 2 57632 7901
0 7903 5 1 1 7902
0 7904 7 4 2 65456 71727
0 7905 5 1 1 82258
0 7906 7 1 2 82259 75753
0 7907 5 1 1 7906
0 7908 7 2 2 58725 74894
0 7909 7 1 2 72447 82262
0 7910 5 1 1 7909
0 7911 7 1 2 7907 7910
0 7912 7 1 2 7903 7911
0 7913 5 1 1 7912
0 7914 7 1 2 69637 7913
0 7915 5 1 1 7914
0 7916 7 1 2 7899 7915
0 7917 5 1 1 7916
0 7918 7 1 2 72520 7917
0 7919 5 1 1 7918
0 7920 7 1 2 72699 77252
0 7921 5 1 1 7920
0 7922 7 1 2 75996 7921
0 7923 5 2 1 7922
0 7924 7 1 2 68732 82264
0 7925 5 1 1 7924
0 7926 7 1 2 81747 7925
0 7927 5 1 1 7926
0 7928 7 1 2 65457 7927
0 7929 5 1 1 7928
0 7930 7 2 2 75730 74661
0 7931 5 1 1 82266
0 7932 7 1 2 75490 82267
0 7933 5 1 1 7932
0 7934 7 1 2 7929 7933
0 7935 5 1 1 7934
0 7936 7 1 2 69638 7935
0 7937 5 1 1 7936
0 7938 7 1 2 76105 75710
0 7939 7 8 2 59470 59976
0 7940 7 3 2 64786 82268
0 7941 7 1 2 74498 82276
0 7942 7 1 2 7938 7941
0 7943 5 1 1 7942
0 7944 7 1 2 7937 7943
0 7945 5 1 1 7944
0 7946 7 1 2 67267 7945
0 7947 5 1 1 7946
0 7948 7 3 2 72015 66819
0 7949 7 1 2 61900 82279
0 7950 5 1 1 7949
0 7951 7 1 2 7931 7950
0 7952 5 1 1 7951
0 7953 7 1 2 76833 7952
0 7954 5 1 1 7953
0 7955 7 1 2 69812 76023
0 7956 7 1 2 72307 75678
0 7957 7 1 2 7955 7956
0 7958 7 1 2 76043 7957
0 7959 5 1 1 7958
0 7960 7 1 2 7954 7959
0 7961 5 1 1 7960
0 7962 7 1 2 68581 7961
0 7963 5 1 1 7962
0 7964 7 1 2 7947 7963
0 7965 7 1 2 7919 7964
0 7966 5 1 1 7965
0 7967 7 1 2 58198 7966
0 7968 5 1 1 7967
0 7969 7 1 2 7877 7968
0 7970 5 1 1 7969
0 7971 7 1 2 82192 7970
0 7972 5 1 1 7971
0 7973 7 1 2 81492 67951
0 7974 7 1 2 72834 7973
0 7975 7 2 2 75692 71132
0 7976 7 2 2 72174 81792
0 7977 7 1 2 82282 82284
0 7978 7 1 2 7974 7977
0 7979 5 1 1 7978
0 7980 7 1 2 7972 7979
0 7981 5 1 1 7980
0 7982 7 1 2 71864 7981
0 7983 5 1 1 7982
0 7984 7 1 2 57926 80114
0 7985 5 1 1 7984
0 7986 7 1 2 72467 69639
0 7987 5 1 1 7986
0 7988 7 4 2 63592 59471
0 7989 7 1 2 69238 82286
0 7990 7 1 2 80178 7989
0 7991 5 1 1 7990
0 7992 7 1 2 7987 7991
0 7993 7 1 2 7985 7992
0 7994 5 1 1 7993
0 7995 7 1 2 59096 7994
0 7996 5 1 1 7995
0 7997 7 1 2 73931 68681
0 7998 5 1 1 7997
0 7999 7 1 2 7996 7998
0 8000 5 1 1 7999
0 8001 7 1 2 58199 8000
0 8002 5 1 1 8001
0 8003 7 1 2 60796 80318
0 8004 5 1 1 8003
0 8005 7 1 2 72236 82247
0 8006 7 1 2 8004 8005
0 8007 5 1 1 8006
0 8008 7 1 2 8002 8007
0 8009 5 1 1 8008
0 8010 7 1 2 75697 8009
0 8011 5 1 1 8010
0 8012 7 4 2 65458 71467
0 8013 5 2 1 82290
0 8014 7 1 2 57927 82291
0 8015 5 1 1 8014
0 8016 7 2 2 71247 8015
0 8017 5 2 1 82296
0 8018 7 1 2 72237 82298
0 8019 5 1 1 8018
0 8020 7 2 2 59472 68957
0 8021 7 1 2 65183 75937
0 8022 7 1 2 82300 8021
0 8023 5 1 1 8022
0 8024 7 1 2 8019 8023
0 8025 5 1 1 8024
0 8026 7 1 2 76127 8025
0 8027 5 1 1 8026
0 8028 7 1 2 8011 8027
0 8029 5 1 1 8028
0 8030 7 1 2 57633 8029
0 8031 5 1 1 8030
0 8032 7 3 2 59097 72136
0 8033 5 2 1 82302
0 8034 7 1 2 80173 82305
0 8035 5 1 1 8034
0 8036 7 4 2 67510 76787
0 8037 7 3 2 58200 82269
0 8038 7 1 2 58726 67441
0 8039 7 1 2 82311 8038
0 8040 7 1 2 82307 8039
0 8041 7 1 2 8035 8040
0 8042 5 1 1 8041
0 8043 7 1 2 8031 8042
0 8044 5 1 1 8043
0 8045 7 1 2 68582 8044
0 8046 5 1 1 8045
0 8047 7 3 2 72016 77253
0 8048 5 1 1 82314
0 8049 7 1 2 8048 81748
0 8050 5 1 1 8049
0 8051 7 1 2 68733 8050
0 8052 5 1 1 8051
0 8053 7 1 2 65459 82265
0 8054 5 1 1 8053
0 8055 7 1 2 8052 8054
0 8056 5 1 1 8055
0 8057 7 1 2 57928 8056
0 8058 5 1 1 8057
0 8059 7 1 2 70006 81745
0 8060 5 1 1 8059
0 8061 7 1 2 8058 8060
0 8062 5 1 1 8061
0 8063 7 1 2 72238 8062
0 8064 5 1 1 8063
0 8065 7 1 2 70347 79792
0 8066 7 1 2 81725 8065
0 8067 5 1 1 8066
0 8068 7 1 2 8064 8067
0 8069 5 1 1 8068
0 8070 7 1 2 80088 8069
0 8071 5 1 1 8070
0 8072 7 4 2 68734 75976
0 8073 5 2 1 82317
0 8074 7 1 2 72263 3514
0 8075 5 1 1 8074
0 8076 7 1 2 82318 8075
0 8077 5 1 1 8076
0 8078 7 1 2 58201 76128
0 8079 5 1 1 8078
0 8080 7 1 2 8077 8079
0 8081 5 1 1 8080
0 8082 7 1 2 72239 8081
0 8083 5 1 1 8082
0 8084 7 2 2 70097 71056
0 8085 7 1 2 72318 82323
0 8086 5 1 1 8085
0 8087 7 1 2 73481 80112
0 8088 5 1 1 8087
0 8089 7 1 2 8086 8088
0 8090 5 1 1 8089
0 8091 7 1 2 82230 8090
0 8092 5 1 1 8091
0 8093 7 3 2 67456 76583
0 8094 5 1 1 82325
0 8095 7 2 2 79958 82326
0 8096 7 5 2 64681 65460
0 8097 5 1 1 82330
0 8098 7 3 2 59268 82331
0 8099 5 2 1 82335
0 8100 7 1 2 82328 82336
0 8101 5 1 1 8100
0 8102 7 4 2 58202 69517
0 8103 7 1 2 75628 82340
0 8104 7 1 2 80181 8103
0 8105 5 1 1 8104
0 8106 7 1 2 8101 8105
0 8107 5 1 1 8106
0 8108 7 1 2 68333 8107
0 8109 5 1 1 8108
0 8110 7 1 2 57634 74560
0 8111 5 1 1 8110
0 8112 7 1 2 70195 8111
0 8113 5 1 1 8112
0 8114 7 1 2 79959 81970
0 8115 7 2 2 82012 8114
0 8116 5 1 1 82344
0 8117 7 1 2 65184 82345
0 8118 7 1 2 8113 8117
0 8119 5 1 1 8118
0 8120 7 1 2 8109 8119
0 8121 7 1 2 8092 8120
0 8122 7 1 2 8083 8121
0 8123 5 1 1 8122
0 8124 7 1 2 57929 8123
0 8125 5 1 1 8124
0 8126 7 2 2 64972 75779
0 8127 5 2 1 82346
0 8128 7 1 2 60797 82348
0 8129 5 1 1 8128
0 8130 7 1 2 77254 8129
0 8131 5 1 1 8130
0 8132 7 1 2 75997 75831
0 8133 7 1 2 8131 8132
0 8134 5 1 1 8133
0 8135 7 1 2 80011 8134
0 8136 5 1 1 8135
0 8137 7 1 2 66677 74394
0 8138 7 4 2 58727 64787
0 8139 7 3 2 63593 82350
0 8140 7 1 2 68902 81760
0 8141 7 1 2 82354 8140
0 8142 7 1 2 8137 8141
0 8143 5 1 1 8142
0 8144 7 1 2 8136 8143
0 8145 5 1 1 8144
0 8146 7 1 2 58203 8145
0 8147 5 1 1 8146
0 8148 7 1 2 68958 82315
0 8149 5 1 1 8148
0 8150 7 1 2 73489 75629
0 8151 5 1 1 8150
0 8152 7 1 2 8149 8151
0 8153 5 1 1 8152
0 8154 7 1 2 75711 8153
0 8155 5 1 1 8154
0 8156 7 1 2 70765 70157
0 8157 7 1 2 75630 8156
0 8158 5 1 1 8157
0 8159 7 1 2 8155 8158
0 8160 5 1 1 8159
0 8161 7 1 2 69640 8160
0 8162 5 1 1 8161
0 8163 7 1 2 8147 8162
0 8164 7 1 2 8125 8163
0 8165 5 1 1 8164
0 8166 7 1 2 59473 8165
0 8167 5 1 1 8166
0 8168 7 1 2 65461 69183
0 8169 7 1 2 82226 8168
0 8170 5 1 1 8169
0 8171 7 1 2 75938 82231
0 8172 5 1 1 8171
0 8173 7 1 2 76501 75939
0 8174 7 1 2 75754 8173
0 8175 5 1 1 8174
0 8176 7 1 2 82228 8175
0 8177 5 1 1 8176
0 8178 7 1 2 57635 8177
0 8179 5 1 1 8178
0 8180 7 1 2 7769 8179
0 8181 7 1 2 8172 8180
0 8182 5 1 1 8181
0 8183 7 1 2 58204 8182
0 8184 5 1 1 8183
0 8185 7 1 2 8170 8184
0 8186 5 1 1 8185
0 8187 7 1 2 69641 8186
0 8188 5 1 1 8187
0 8189 7 2 2 71578 82072
0 8190 7 2 2 67511 72103
0 8191 7 8 2 59977 65462
0 8192 7 1 2 82359 82361
0 8193 7 1 2 82357 8192
0 8194 5 1 1 8193
0 8195 7 1 2 8188 8194
0 8196 7 1 2 8167 8195
0 8197 5 1 1 8196
0 8198 7 1 2 73278 8197
0 8199 5 1 1 8198
0 8200 7 1 2 8071 8199
0 8201 7 1 2 8046 8200
0 8202 5 1 1 8201
0 8203 7 1 2 82193 8202
0 8204 5 1 1 8203
0 8205 7 1 2 61901 79311
0 8206 7 2 2 57930 72468
0 8207 7 2 2 72175 74823
0 8208 7 17 2 59474 61521
0 8209 5 4 1 82373
0 8210 7 4 2 58205 82374
0 8211 5 3 1 82394
0 8212 7 1 2 82371 82395
0 8213 7 1 2 82369 8212
0 8214 7 1 2 8205 8213
0 8215 7 1 2 78359 8214
0 8216 5 1 1 8215
0 8217 7 1 2 8204 8216
0 8218 7 1 2 7983 8217
0 8219 7 1 2 7847 8218
0 8220 5 1 1 8219
0 8221 7 1 2 58407 8220
0 8222 5 1 1 8221
0 8223 7 1 2 79175 81129
0 8224 5 1 1 8223
0 8225 7 31 2 59752 66127
0 8226 5 2 1 82401
0 8227 7 5 2 67457 82402
0 8228 7 10 2 59269 74630
0 8229 5 4 1 82439
0 8230 7 1 2 79071 67887
0 8231 5 1 1 8230
0 8232 7 1 2 82449 8231
0 8233 5 1 1 8232
0 8234 7 1 2 65463 8233
0 8235 5 1 1 8234
0 8236 7 2 2 72377 80573
0 8237 5 1 1 82453
0 8238 7 1 2 8235 8237
0 8239 5 1 1 8238
0 8240 7 1 2 58206 8239
0 8241 5 1 1 8240
0 8242 7 1 2 73108 77755
0 8243 5 1 1 8242
0 8244 7 2 2 80104 8243
0 8245 7 1 2 79072 82455
0 8246 5 1 1 8245
0 8247 7 1 2 67641 70267
0 8248 5 1 1 8247
0 8249 7 1 2 67840 76258
0 8250 5 1 1 8249
0 8251 7 1 2 70240 8250
0 8252 7 1 2 8248 8251
0 8253 7 1 2 81182 8252
0 8254 7 1 2 8246 8253
0 8255 5 1 1 8254
0 8256 7 1 2 59475 8255
0 8257 5 1 1 8256
0 8258 7 1 2 8241 8257
0 8259 7 1 2 81149 8258
0 8260 5 1 1 8259
0 8261 7 1 2 82434 8260
0 8262 5 1 1 8261
0 8263 7 1 2 8224 8262
0 8264 5 1 1 8263
0 8265 7 1 2 66747 8264
0 8266 5 1 1 8265
0 8267 7 1 2 62897 81002
0 8268 5 1 1 8267
0 8269 7 1 2 81005 8268
0 8270 5 1 1 8269
0 8271 7 1 2 67151 8270
0 8272 5 1 1 8271
0 8273 7 3 2 72189 77392
0 8274 7 1 2 82457 78019
0 8275 5 1 1 8274
0 8276 7 1 2 8272 8275
0 8277 5 1 1 8276
0 8278 7 1 2 64471 82091
0 8279 7 1 2 8277 8278
0 8280 5 1 1 8279
0 8281 7 2 2 61902 82403
0 8282 7 2 2 65464 70958
0 8283 5 2 1 82462
0 8284 7 4 2 70108 82464
0 8285 5 7 1 82466
0 8286 7 1 2 59476 82470
0 8287 5 1 1 8286
0 8288 7 1 2 58207 72469
0 8289 5 1 1 8288
0 8290 7 1 2 8287 8289
0 8291 5 1 1 8290
0 8292 7 1 2 67268 8291
0 8293 5 1 1 8292
0 8294 7 1 2 64193 73435
0 8295 5 2 1 8294
0 8296 7 1 2 57636 82477
0 8297 5 1 1 8296
0 8298 7 1 2 73813 8297
0 8299 5 1 1 8298
0 8300 7 1 2 70386 8299
0 8301 5 1 1 8300
0 8302 7 1 2 73754 76276
0 8303 5 2 1 8302
0 8304 7 1 2 8301 82479
0 8305 7 1 2 8293 8304
0 8306 5 1 1 8305
0 8307 7 1 2 77129 8306
0 8308 5 1 1 8307
0 8309 7 2 2 70244 80626
0 8310 5 3 1 82481
0 8311 7 1 2 75862 82483
0 8312 5 1 1 8311
0 8313 7 2 2 81277 8312
0 8314 5 1 1 82486
0 8315 7 1 2 59477 8314
0 8316 5 1 1 8315
0 8317 7 4 2 68069 73214
0 8318 5 1 1 82488
0 8319 7 1 2 58208 73868
0 8320 7 1 2 8318 8319
0 8321 5 1 1 8320
0 8322 7 1 2 8316 8321
0 8323 7 1 2 8308 8322
0 8324 5 1 1 8323
0 8325 7 1 2 82460 8324
0 8326 5 1 1 8325
0 8327 7 1 2 8280 8326
0 8328 5 1 1 8327
0 8329 7 1 2 74246 8328
0 8330 5 1 1 8329
0 8331 7 1 2 8266 8330
0 8332 5 1 1 8331
0 8333 7 1 2 63156 8332
0 8334 5 1 1 8333
0 8335 7 3 2 66128 69308
0 8336 7 1 2 57637 72137
0 8337 5 1 1 8336
0 8338 7 1 2 70680 8337
0 8339 5 2 1 8338
0 8340 7 1 2 63841 80152
0 8341 5 1 1 8340
0 8342 7 4 2 82495 8341
0 8343 7 1 2 68735 82497
0 8344 5 1 1 8343
0 8345 7 1 2 60507 76277
0 8346 5 1 1 8345
0 8347 7 1 2 8344 8346
0 8348 5 1 1 8347
0 8349 7 1 2 82492 8348
0 8350 5 1 1 8349
0 8351 7 2 2 74090 81381
0 8352 5 3 1 82501
0 8353 7 4 2 64194 81382
0 8354 5 1 1 82506
0 8355 7 1 2 81998 82375
0 8356 5 1 1 8355
0 8357 7 1 2 8354 8356
0 8358 5 2 1 8357
0 8359 7 1 2 68736 82510
0 8360 5 1 1 8359
0 8361 7 1 2 82503 8360
0 8362 5 1 1 8361
0 8363 7 1 2 59270 8362
0 8364 5 1 1 8363
0 8365 7 1 2 65465 81463
0 8366 7 1 2 79016 8365
0 8367 5 1 1 8366
0 8368 7 1 2 8364 8367
0 8369 5 1 1 8368
0 8370 7 1 2 68334 8369
0 8371 5 1 1 8370
0 8372 7 1 2 82502 76864
0 8373 5 1 1 8372
0 8374 7 3 2 64973 81493
0 8375 5 1 1 82512
0 8376 7 1 2 72984 82513
0 8377 5 1 1 8376
0 8378 7 1 2 82504 8377
0 8379 5 1 1 8378
0 8380 7 1 2 68737 8379
0 8381 5 1 1 8380
0 8382 7 4 2 64195 81464
0 8383 5 1 1 82515
0 8384 7 1 2 65466 82516
0 8385 5 1 1 8384
0 8386 7 1 2 59271 82511
0 8387 5 1 1 8386
0 8388 7 1 2 8385 8387
0 8389 7 1 2 8381 8388
0 8390 5 1 1 8389
0 8391 7 1 2 67642 8390
0 8392 5 1 1 8391
0 8393 7 1 2 8373 8392
0 8394 7 1 2 8371 8393
0 8395 5 1 1 8394
0 8396 7 1 2 57931 8395
0 8397 5 1 1 8396
0 8398 7 1 2 8350 8397
0 8399 5 1 1 8398
0 8400 7 1 2 59753 8399
0 8401 5 1 1 8400
0 8402 7 4 2 80226 79793
0 8403 5 1 1 82519
0 8404 7 14 2 65467 66129
0 8405 7 4 2 65185 82523
0 8406 7 4 2 59272 73713
0 8407 7 1 2 82537 82541
0 8408 7 1 2 82520 8407
0 8409 5 1 1 8408
0 8410 7 1 2 8401 8409
0 8411 5 1 1 8410
0 8412 7 1 2 75631 8411
0 8413 5 1 1 8412
0 8414 7 2 2 65468 72985
0 8415 7 42 2 59754 61522
0 8416 5 12 1 82547
0 8417 7 2 2 64472 81565
0 8418 5 2 1 82601
0 8419 7 1 2 82589 82603
0 8420 5 5 1 8419
0 8421 7 1 2 82545 82605
0 8422 5 1 1 8421
0 8423 7 3 2 59755 81566
0 8424 7 1 2 77976 82610
0 8425 5 2 1 8424
0 8426 7 1 2 8422 82613
0 8427 5 1 1 8426
0 8428 7 1 2 70766 8427
0 8429 5 1 1 8428
0 8430 7 1 2 78071 81572
0 8431 5 1 1 8430
0 8432 7 1 2 8429 8431
0 8433 5 1 1 8432
0 8434 7 1 2 57638 8433
0 8435 5 1 1 8434
0 8436 7 1 2 71865 69504
0 8437 7 1 2 82404 8436
0 8438 7 1 2 80179 8437
0 8439 5 1 1 8438
0 8440 7 1 2 8435 8439
0 8441 5 1 1 8440
0 8442 7 1 2 57932 8441
0 8443 5 1 1 8442
0 8444 7 1 2 72842 82493
0 8445 7 1 2 82498 8444
0 8446 5 1 1 8445
0 8447 7 1 2 8443 8446
0 8448 5 1 1 8447
0 8449 7 1 2 75632 8448
0 8450 5 1 1 8449
0 8451 7 7 2 63468 66558
0 8452 7 1 2 69184 82615
0 8453 7 1 2 82303 8452
0 8454 7 4 2 60266 79817
0 8455 7 1 2 82494 82622
0 8456 7 1 2 8453 8455
0 8457 5 1 1 8456
0 8458 7 1 2 8450 8457
0 8459 5 1 1 8458
0 8460 7 1 2 68583 8459
0 8461 5 1 1 8460
0 8462 7 2 2 78205 72818
0 8463 5 1 1 82626
0 8464 7 8 2 59273 64682
0 8465 7 1 2 82628 79333
0 8466 7 1 2 81325 77205
0 8467 7 1 2 75825 8466
0 8468 7 1 2 8465 8467
0 8469 7 1 2 82627 8468
0 8470 5 1 1 8469
0 8471 7 1 2 8461 8470
0 8472 7 1 2 8413 8471
0 8473 5 1 1 8472
0 8474 7 1 2 72418 8473
0 8475 5 1 1 8474
0 8476 7 1 2 8334 8475
0 8477 5 1 1 8476
0 8478 7 1 2 67916 8477
0 8479 5 1 1 8478
0 8480 7 1 2 76614 76106
0 8481 7 1 2 82277 8480
0 8482 5 1 1 8481
0 8483 7 12 2 58408 64683
0 8484 7 1 2 70481 82636
0 8485 7 1 2 81049 8484
0 8486 5 1 1 8485
0 8487 7 1 2 8482 8486
0 8488 5 1 1 8487
0 8489 7 19 2 66130 61903
0 8490 7 1 2 77712 74459
0 8491 5 2 1 8490
0 8492 7 1 2 82648 82667
0 8493 7 1 2 8488 8492
0 8494 5 1 1 8493
0 8495 7 1 2 75998 77287
0 8496 5 2 1 8495
0 8497 7 1 2 70482 82669
0 8498 5 1 1 8497
0 8499 7 1 2 77206 81930
0 8500 5 1 1 8499
0 8501 7 2 2 61904 79965
0 8502 5 1 1 82671
0 8503 7 1 2 8500 8502
0 8504 7 1 2 8498 8503
0 8505 5 1 1 8504
0 8506 7 18 2 60267 61523
0 8507 7 1 2 82673 80678
0 8508 7 1 2 8505 8507
0 8509 5 1 1 8508
0 8510 7 1 2 8494 8509
0 8511 5 1 1 8510
0 8512 7 1 2 72308 8511
0 8513 5 1 1 8512
0 8514 7 3 2 66131 79254
0 8515 7 2 2 69155 82691
0 8516 7 2 2 67037 77024
0 8517 7 1 2 58728 82696
0 8518 7 1 2 82694 8517
0 8519 5 1 1 8518
0 8520 7 1 2 8513 8519
0 8521 5 1 1 8520
0 8522 7 1 2 67152 8521
0 8523 5 1 1 8522
0 8524 7 2 2 65469 71248
0 8525 5 1 1 82698
0 8526 7 1 2 79578 8525
0 8527 5 1 1 8526
0 8528 7 1 2 80392 75679
0 8529 7 1 2 82692 8528
0 8530 7 1 2 8527 8529
0 8531 5 1 1 8530
0 8532 7 1 2 8523 8531
0 8533 5 1 1 8532
0 8534 7 1 2 70612 8533
0 8535 5 1 1 8534
0 8536 7 1 2 75633 81715
0 8537 5 1 1 8536
0 8538 7 1 2 66559 72138
0 8539 7 2 2 74776 8538
0 8540 7 2 2 69185 74848
0 8541 7 3 2 57365 59478
0 8542 5 2 1 82704
0 8543 7 1 2 82702 82705
0 8544 7 1 2 82700 8543
0 8545 5 1 1 8544
0 8546 7 1 2 8537 8545
0 8547 5 1 1 8546
0 8548 7 8 2 64788 66132
0 8549 7 5 2 63594 59756
0 8550 7 2 2 82709 82717
0 8551 7 1 2 66678 77777
0 8552 7 1 2 82722 8551
0 8553 7 1 2 8547 8552
0 8554 5 1 1 8553
0 8555 7 1 2 8535 8554
0 8556 7 1 2 8479 8555
0 8557 7 1 2 8222 8556
0 8558 7 1 2 7252 8557
0 8559 5 1 1 8558
0 8560 7 1 2 61186 8559
0 8561 5 1 1 8560
0 8562 7 1 2 77649 79648
0 8563 5 1 1 8562
0 8564 7 1 2 5291 8563
0 8565 5 1 1 8564
0 8566 7 1 2 65186 8565
0 8567 5 1 1 8566
0 8568 7 1 2 3567 8567
0 8569 5 1 1 8568
0 8570 7 1 2 59274 8569
0 8571 5 1 1 8570
0 8572 7 1 2 69930 78059
0 8573 5 1 1 8572
0 8574 7 1 2 70613 8573
0 8575 5 1 1 8574
0 8576 7 1 2 57933 71038
0 8577 5 2 1 8576
0 8578 7 1 2 75898 82724
0 8579 5 1 1 8578
0 8580 7 1 2 8575 8579
0 8581 5 2 1 8580
0 8582 7 1 2 71147 82726
0 8583 5 1 1 8582
0 8584 7 1 2 8571 8583
0 8585 5 1 1 8584
0 8586 7 1 2 60268 8585
0 8587 5 1 1 8586
0 8588 7 1 2 69931 80920
0 8589 5 2 1 8588
0 8590 7 2 2 62603 82728
0 8591 5 1 1 82730
0 8592 7 1 2 71148 82731
0 8593 5 1 1 8592
0 8594 7 1 2 8587 8593
0 8595 5 1 1 8594
0 8596 7 1 2 69266 8595
0 8597 5 1 1 8596
0 8598 7 2 2 59479 74574
0 8599 5 1 1 82732
0 8600 7 2 2 69984 67010
0 8601 5 1 1 82734
0 8602 7 2 2 67269 73769
0 8603 7 1 2 70959 82736
0 8604 5 1 1 8603
0 8605 7 1 2 8601 8604
0 8606 5 2 1 8605
0 8607 7 1 2 58961 82738
0 8608 5 1 1 8607
0 8609 7 4 2 60508 67270
0 8610 5 3 1 82740
0 8611 7 1 2 72700 82741
0 8612 5 1 1 8611
0 8613 7 1 2 8608 8612
0 8614 5 1 1 8613
0 8615 7 1 2 57366 8614
0 8616 5 1 1 8615
0 8617 7 1 2 8599 8616
0 8618 5 1 1 8617
0 8619 7 1 2 69642 8618
0 8620 5 1 1 8619
0 8621 7 1 2 8597 8620
0 8622 5 1 1 8621
0 8623 7 1 2 75634 8622
0 8624 5 1 1 8623
0 8625 7 3 2 64974 67271
0 8626 5 1 1 82747
0 8627 7 1 2 71620 82748
0 8628 5 1 1 8627
0 8629 7 1 2 70367 8628
0 8630 5 1 1 8629
0 8631 7 1 2 57639 8630
0 8632 5 1 1 8631
0 8633 7 3 2 57934 69412
0 8634 5 2 1 82750
0 8635 7 1 2 59275 82751
0 8636 5 1 1 8635
0 8637 7 1 2 81524 8636
0 8638 7 1 2 8632 8637
0 8639 5 1 1 8638
0 8640 7 1 2 59098 8639
0 8641 5 1 1 8640
0 8642 7 2 2 62320 74355
0 8643 5 1 1 82755
0 8644 7 1 2 8643 82752
0 8645 5 1 1 8644
0 8646 7 1 2 62898 8645
0 8647 5 1 1 8646
0 8648 7 1 2 59276 8647
0 8649 5 1 1 8648
0 8650 7 1 2 67581 72675
0 8651 5 1 1 8650
0 8652 7 1 2 64196 8651
0 8653 7 1 2 8649 8652
0 8654 7 1 2 8641 8653
0 8655 5 1 1 8654
0 8656 7 1 2 60509 79698
0 8657 5 1 1 8656
0 8658 7 2 2 74608 8657
0 8659 7 1 2 57935 70047
0 8660 5 1 1 8659
0 8661 7 1 2 74610 8660
0 8662 5 1 1 8661
0 8663 7 1 2 59480 8662
0 8664 7 1 2 82757 8663
0 8665 5 1 1 8664
0 8666 7 1 2 69643 8665
0 8667 7 1 2 8655 8666
0 8668 5 1 1 8667
0 8669 7 1 2 79277 80220
0 8670 7 1 2 82287 8669
0 8671 7 1 2 66679 70920
0 8672 7 1 2 81675 8671
0 8673 7 1 2 8670 8672
0 8674 5 1 1 8673
0 8675 7 1 2 8668 8674
0 8676 5 1 1 8675
0 8677 7 1 2 77255 8676
0 8678 5 1 1 8677
0 8679 7 1 2 8624 8678
0 8680 5 1 1 8679
0 8681 7 1 2 58409 8680
0 8682 5 1 1 8681
0 8683 7 1 2 7662 82252
0 8684 5 1 1 8683
0 8685 7 1 2 71866 8684
0 8686 5 1 1 8685
0 8687 7 1 2 60269 70810
0 8688 5 2 1 8687
0 8689 7 2 2 79689 82759
0 8690 7 1 2 76129 82761
0 8691 5 1 1 8690
0 8692 7 2 2 57367 59978
0 8693 7 2 2 82351 82763
0 8694 7 2 2 67512 67428
0 8695 7 1 2 69112 82767
0 8696 7 1 2 82765 8695
0 8697 5 1 1 8696
0 8698 7 1 2 8691 8697
0 8699 7 1 2 8686 8698
0 8700 5 1 1 8699
0 8701 7 1 2 59277 8700
0 8702 5 1 1 8701
0 8703 7 3 2 67643 75755
0 8704 5 1 1 82769
0 8705 7 1 2 82168 82770
0 8706 5 1 1 8705
0 8707 7 1 2 65187 82319
0 8708 5 1 1 8707
0 8709 7 1 2 8706 8708
0 8710 5 1 1 8709
0 8711 7 1 2 69644 8710
0 8712 5 1 1 8711
0 8713 7 1 2 8702 8712
0 8714 5 1 1 8713
0 8715 7 1 2 57936 8714
0 8716 5 1 1 8715
0 8717 7 1 2 69960 75977
0 8718 5 2 1 8717
0 8719 7 1 2 75803 76018
0 8720 5 1 1 8719
0 8721 7 1 2 81782 8720
0 8722 5 2 1 8721
0 8723 7 1 2 67644 82774
0 8724 5 1 1 8723
0 8725 7 1 2 82772 8724
0 8726 5 1 1 8725
0 8727 7 1 2 68738 8726
0 8728 5 1 1 8727
0 8729 7 2 2 68959 77215
0 8730 7 1 2 81976 82776
0 8731 5 1 1 8730
0 8732 7 1 2 8728 8731
0 8733 5 1 1 8732
0 8734 7 1 2 69645 8733
0 8735 5 1 1 8734
0 8736 7 1 2 8716 8735
0 8737 5 1 1 8736
0 8738 7 1 2 63157 8737
0 8739 5 1 1 8738
0 8740 7 1 2 78282 69123
0 8741 5 1 1 8740
0 8742 7 3 2 59979 67272
0 8743 7 9 2 57368 58729
0 8744 5 2 1 82781
0 8745 7 1 2 60510 82782
0 8746 7 1 2 67965 8745
0 8747 7 1 2 82778 8746
0 8748 7 1 2 8741 8747
0 8749 5 1 1 8748
0 8750 7 1 2 8739 8749
0 8751 5 1 1 8750
0 8752 7 1 2 59481 8751
0 8753 5 1 1 8752
0 8754 7 3 2 59278 67038
0 8755 5 1 1 82792
0 8756 7 1 2 74091 74794
0 8757 7 1 2 82793 8756
0 8758 7 1 2 76600 8757
0 8759 5 1 1 8758
0 8760 7 1 2 8753 8759
0 8761 5 1 1 8760
0 8762 7 1 2 58209 8761
0 8763 5 1 1 8762
0 8764 7 17 2 63158 58730
0 8765 7 2 2 82795 82270
0 8766 7 1 2 72641 82812
0 8767 7 1 2 69206 8766
0 8768 5 1 1 8767
0 8769 7 1 2 8763 8768
0 8770 7 1 2 8682 8769
0 8771 5 1 1 8770
0 8772 7 1 2 66133 8771
0 8773 5 1 1 8772
0 8774 7 1 2 67987 75756
0 8775 5 2 1 8774
0 8776 7 1 2 69869 81779
0 8777 5 1 1 8776
0 8778 7 1 2 82814 8777
0 8779 5 1 1 8778
0 8780 7 1 2 57640 8779
0 8781 5 1 1 8780
0 8782 7 1 2 76011 75821
0 8783 5 1 1 8782
0 8784 7 1 2 8781 8783
0 8785 5 1 1 8784
0 8786 7 1 2 63159 8785
0 8787 5 1 1 8786
0 8788 7 2 2 69870 66820
0 8789 7 2 2 67273 68704
0 8790 7 1 2 82816 82818
0 8791 5 1 1 8790
0 8792 7 1 2 8787 8791
0 8793 5 1 1 8792
0 8794 7 1 2 59482 8793
0 8795 5 1 1 8794
0 8796 7 2 2 59099 79847
0 8797 7 2 2 59279 75422
0 8798 7 1 2 69186 69163
0 8799 7 1 2 82822 8798
0 8800 7 2 2 82820 8799
0 8801 5 1 1 82824
0 8802 7 1 2 8795 8801
0 8803 5 1 1 8802
0 8804 7 1 2 58210 8803
0 8805 5 1 1 8804
0 8806 7 3 2 57641 70387
0 8807 5 1 1 82826
0 8808 7 1 2 80575 8807
0 8809 5 1 1 8808
0 8810 7 1 2 64197 8809
0 8811 5 1 1 8810
0 8812 7 1 2 78521 70994
0 8813 5 1 1 8812
0 8814 7 1 2 8811 8813
0 8815 5 1 1 8814
0 8816 7 1 2 77256 8815
0 8817 5 1 1 8816
0 8818 7 2 2 64198 67011
0 8819 5 1 1 82829
0 8820 7 1 2 8819 82744
0 8821 5 1 1 8820
0 8822 7 1 2 69871 75978
0 8823 7 1 2 8821 8822
0 8824 5 1 1 8823
0 8825 7 1 2 8817 8824
0 8826 5 1 1 8825
0 8827 7 1 2 58410 8826
0 8828 5 1 1 8827
0 8829 7 2 2 70767 75680
0 8830 7 1 2 59280 70717
0 8831 7 1 2 73995 82271
0 8832 7 1 2 8830 8831
0 8833 7 1 2 82831 8832
0 8834 5 1 1 8833
0 8835 7 1 2 8828 8834
0 8836 7 1 2 8805 8835
0 8837 5 1 1 8836
0 8838 7 1 2 66134 8837
0 8839 5 1 1 8838
0 8840 7 4 2 66560 75386
0 8841 7 1 2 79743 82833
0 8842 5 1 1 8841
0 8843 7 2 2 62604 71249
0 8844 5 3 1 82837
0 8845 7 7 2 82839 78182
0 8846 5 5 1 82842
0 8847 7 6 2 71468 82843
0 8848 5 2 1 82854
0 8849 7 1 2 72378 75979
0 8850 7 1 2 82855 8849
0 8851 5 1 1 8850
0 8852 7 1 2 8842 8851
0 8853 5 1 1 8852
0 8854 7 1 2 65188 81245
0 8855 7 1 2 8853 8854
0 8856 5 1 1 8855
0 8857 7 1 2 8839 8856
0 8858 5 1 1 8857
0 8859 7 1 2 69646 8858
0 8860 5 1 1 8859
0 8861 7 3 2 66135 75429
0 8862 7 1 2 74790 82862
0 8863 5 1 1 8862
0 8864 7 22 2 63160 66136
0 8865 5 3 1 82865
0 8866 7 2 2 81266 82887
0 8867 5 4 1 82890
0 8868 7 2 2 71149 82892
0 8869 5 2 1 82896
0 8870 7 1 2 67582 82897
0 8871 5 1 1 8870
0 8872 7 1 2 8863 8871
0 8873 5 1 1 8872
0 8874 7 2 2 57937 73356
0 8875 7 1 2 74418 82308
0 8876 7 1 2 82900 8875
0 8877 7 1 2 8873 8876
0 8878 5 1 1 8877
0 8879 7 1 2 8860 8878
0 8880 5 1 1 8879
0 8881 7 1 2 68584 8880
0 8882 5 1 1 8881
0 8883 7 3 2 58211 78154
0 8884 5 7 1 82902
0 8885 7 1 2 75451 82905
0 8886 5 5 1 8885
0 8887 7 1 2 82912 81751
0 8888 5 1 1 8887
0 8889 7 17 2 63161 71250
0 8890 5 54 1 82917
0 8891 7 2 2 60511 82934
0 8892 5 1 1 82988
0 8893 7 1 2 75980 82989
0 8894 5 1 1 8893
0 8895 7 1 2 8888 8894
0 8896 5 1 1 8895
0 8897 7 1 2 66137 8896
0 8898 5 1 1 8897
0 8899 7 4 2 58411 76577
0 8900 7 2 2 65189 82092
0 8901 7 8 2 64684 74662
0 8902 7 1 2 82994 82996
0 8903 7 1 2 82990 8902
0 8904 5 1 1 8903
0 8905 7 1 2 8898 8904
0 8906 5 1 1 8905
0 8907 7 1 2 76834 8906
0 8908 5 1 1 8907
0 8909 7 1 2 58412 81549
0 8910 5 1 1 8909
0 8911 7 1 2 82898 8910
0 8912 5 1 1 8911
0 8913 7 5 2 57938 76049
0 8914 7 2 2 76024 83004
0 8915 5 1 1 83009
0 8916 7 1 2 82768 83010
0 8917 7 1 2 8912 8916
0 8918 5 1 1 8917
0 8919 7 1 2 8908 8918
0 8920 5 1 1 8919
0 8921 7 1 2 57642 8920
0 8922 5 1 1 8921
0 8923 7 1 2 75757 73741
0 8924 5 1 1 8923
0 8925 7 1 2 81783 8924
0 8926 5 1 1 8925
0 8927 7 1 2 57939 8926
0 8928 5 1 1 8927
0 8929 7 1 2 8928 82773
0 8930 5 1 1 8929
0 8931 7 1 2 82913 8930
0 8932 5 1 1 8931
0 8933 7 5 2 63469 77633
0 8934 7 1 2 66561 82991
0 8935 7 1 2 83011 8934
0 8936 5 1 1 8935
0 8937 7 1 2 8932 8936
0 8938 5 1 1 8937
0 8939 7 12 2 66138 62049
0 8940 7 4 2 83016 67917
0 8941 7 1 2 8938 83028
0 8942 5 1 1 8941
0 8943 7 1 2 8922 8942
0 8944 5 1 1 8943
0 8945 7 1 2 74032 8944
0 8946 5 1 1 8945
0 8947 7 1 2 75863 81764
0 8948 5 1 1 8947
0 8949 7 1 2 76138 8948
0 8950 5 1 1 8949
0 8951 7 1 2 68739 8950
0 8952 5 1 1 8951
0 8953 7 1 2 63842 82756
0 8954 5 2 1 8953
0 8955 7 1 2 77257 83032
0 8956 5 1 1 8955
0 8957 7 1 2 75999 8956
0 8958 5 1 1 8957
0 8959 7 1 2 69647 8958
0 8960 5 1 1 8959
0 8961 7 1 2 8952 8960
0 8962 5 1 1 8961
0 8963 7 1 2 67988 8962
0 8964 5 1 1 8963
0 8965 7 1 2 76000 2734
0 8966 5 1 1 8965
0 8967 7 1 2 57643 8966
0 8968 5 1 1 8967
0 8969 7 1 2 63843 72399
0 8970 5 1 1 8969
0 8971 7 1 2 75635 8970
0 8972 5 1 1 8971
0 8973 7 1 2 8968 8972
0 8974 5 1 1 8973
0 8975 7 1 2 64975 8974
0 8976 5 1 1 8975
0 8977 7 1 2 66748 72352
0 8978 7 5 2 57644 66562
0 8979 7 1 2 69113 83034
0 8980 7 1 2 8977 8979
0 8981 5 1 1 8980
0 8982 7 1 2 8976 8981
0 8983 5 1 1 8982
0 8984 7 1 2 76835 8983
0 8985 5 1 1 8984
0 8986 7 1 2 8964 8985
0 8987 5 1 1 8986
0 8988 7 2 2 71150 81246
0 8989 5 3 1 83039
0 8990 7 1 2 8987 83040
0 8991 5 1 1 8990
0 8992 7 1 2 69114 75758
0 8993 5 1 1 8992
0 8994 7 1 2 75671 8993
0 8995 5 1 1 8994
0 8996 7 1 2 67100 69572
0 8997 5 1 1 8996
0 8998 7 1 2 69704 8997
0 8999 5 1 1 8998
0 9000 7 1 2 57940 8999
0 9001 5 1 1 9000
0 9002 7 1 2 72183 9001
0 9003 5 1 1 9002
0 9004 7 1 2 58212 68694
0 9005 5 1 1 9004
0 9006 7 1 2 82863 9005
0 9007 5 1 1 9006
0 9008 7 1 2 82899 9007
0 9009 5 1 1 9008
0 9010 7 1 2 70867 9009
0 9011 7 1 2 9003 9010
0 9012 5 1 1 9011
0 9013 7 2 2 67274 82914
0 9014 5 1 1 83044
0 9015 7 6 2 57645 66139
0 9016 7 1 2 69648 83046
0 9017 7 1 2 83045 9016
0 9018 5 1 1 9017
0 9019 7 1 2 9012 9018
0 9020 5 1 1 9019
0 9021 7 1 2 65190 9020
0 9022 5 1 1 9021
0 9023 7 2 2 67989 69649
0 9024 7 1 2 66140 82915
0 9025 7 1 2 83052 9024
0 9026 5 1 1 9025
0 9027 7 1 2 9022 9026
0 9028 5 1 1 9027
0 9029 7 1 2 8995 9028
0 9030 5 1 1 9029
0 9031 7 1 2 8991 9030
0 9032 7 1 2 8946 9031
0 9033 7 1 2 8882 9032
0 9034 7 1 2 8773 9033
0 9035 5 1 1 9034
0 9036 7 1 2 65470 9035
0 9037 5 1 1 9036
0 9038 7 3 2 58213 68335
0 9039 5 1 1 83054
0 9040 7 1 2 68740 80105
0 9041 5 1 1 9040
0 9042 7 1 2 9039 9041
0 9043 5 1 1 9042
0 9044 7 1 2 59281 9043
0 9045 5 1 1 9044
0 9046 7 1 2 71579 75780
0 9047 5 1 1 9046
0 9048 7 1 2 9045 9047
0 9049 5 1 1 9048
0 9050 7 1 2 64976 9049
0 9051 5 1 1 9050
0 9052 7 1 2 78918 9051
0 9053 5 1 1 9052
0 9054 7 1 2 60512 9053
0 9055 5 1 1 9054
0 9056 7 1 2 76047 70071
0 9057 5 1 1 9056
0 9058 7 1 2 9055 9057
0 9059 5 1 1 9058
0 9060 7 1 2 77258 9059
0 9061 5 1 1 9060
0 9062 7 8 2 58214 63470
0 9063 7 1 2 83057 81920
0 9064 5 3 1 9063
0 9065 7 1 2 75712 75636
0 9066 5 1 1 9065
0 9067 7 1 2 83065 9066
0 9068 5 1 1 9067
0 9069 7 1 2 57941 9068
0 9070 5 1 1 9069
0 9071 7 2 2 75953 74760
0 9072 5 1 1 83068
0 9073 7 1 2 9070 9072
0 9074 5 1 1 9073
0 9075 7 1 2 72240 9074
0 9076 5 1 1 9075
0 9077 7 1 2 72210 75637
0 9078 5 1 1 9077
0 9079 7 2 2 64977 82834
0 9080 7 1 2 74577 83070
0 9081 5 1 1 9080
0 9082 7 1 2 9078 9081
0 9083 5 1 1 9082
0 9084 7 6 2 57646 68741
0 9085 5 9 1 83072
0 9086 7 2 2 62605 83078
0 9087 5 2 1 83087
0 9088 7 1 2 9083 83089
0 9089 5 1 1 9088
0 9090 7 1 2 9076 9089
0 9091 7 1 2 9061 9090
0 9092 5 1 1 9091
0 9093 7 1 2 69650 9092
0 9094 5 1 1 9093
0 9095 7 2 2 76831 72216
0 9096 5 1 1 83091
0 9097 7 2 2 81933 75759
0 9098 5 1 1 83093
0 9099 7 1 2 75702 9098
0 9100 5 1 1 9099
0 9101 7 1 2 9096 9100
0 9102 5 1 1 9101
0 9103 7 1 2 70718 75981
0 9104 5 1 1 9103
0 9105 7 1 2 83066 9104
0 9106 5 1 1 9105
0 9107 7 1 2 75925 9106
0 9108 5 1 1 9107
0 9109 7 1 2 9102 9108
0 9110 5 1 1 9109
0 9111 7 1 2 69651 9110
0 9112 5 1 1 9111
0 9113 7 3 2 79848 67543
0 9114 7 1 2 64978 72828
0 9115 7 1 2 67442 74824
0 9116 7 1 2 9114 9115
0 9117 7 1 2 83095 9116
0 9118 5 1 1 9117
0 9119 7 1 2 9112 9118
0 9120 5 1 1 9119
0 9121 7 1 2 68585 9120
0 9122 5 1 1 9121
0 9123 7 3 2 57369 71580
0 9124 7 2 2 74808 83098
0 9125 7 2 2 76107 83096
0 9126 7 1 2 83101 83103
0 9127 5 1 1 9126
0 9128 7 1 2 76146 83035
0 9129 7 1 2 74913 9128
0 9130 5 1 1 9129
0 9131 7 2 2 58731 70388
0 9132 7 2 2 59980 75781
0 9133 7 1 2 61905 83107
0 9134 7 1 2 83105 9133
0 9135 5 1 1 9134
0 9136 7 1 2 9130 9135
0 9137 5 1 1 9136
0 9138 7 1 2 69652 9137
0 9139 5 1 1 9138
0 9140 7 1 2 9127 9139
0 9141 5 1 1 9140
0 9142 7 1 2 71867 9141
0 9143 5 1 1 9142
0 9144 7 1 2 71102 82821
0 9145 7 1 2 82358 9144
0 9146 5 1 1 9145
0 9147 7 1 2 9143 9146
0 9148 7 1 2 9122 9147
0 9149 7 1 2 9094 9148
0 9150 5 1 1 9149
0 9151 7 1 2 60798 9150
0 9152 5 1 1 9151
0 9153 7 1 2 74903 82616
0 9154 7 1 2 75317 9153
0 9155 5 1 1 9154
0 9156 7 1 2 75703 9155
0 9157 5 1 1 9156
0 9158 7 1 2 68586 9157
0 9159 5 1 1 9158
0 9160 7 1 2 68336 83094
0 9161 5 1 1 9160
0 9162 7 2 2 75804 81921
0 9163 5 1 1 83109
0 9164 7 1 2 57647 83110
0 9165 5 1 1 9164
0 9166 7 1 2 76007 82321
0 9167 7 1 2 9165 9166
0 9168 7 1 2 9161 9167
0 9169 7 1 2 9159 9168
0 9170 5 1 1 9169
0 9171 7 1 2 68682 9170
0 9172 5 1 1 9171
0 9173 7 2 2 82629 82329
0 9174 5 1 1 83111
0 9175 7 1 2 66821 71057
0 9176 7 1 2 82360 9175
0 9177 5 1 1 9176
0 9178 7 1 2 9174 9177
0 9179 5 1 1 9178
0 9180 7 1 2 62606 9179
0 9181 5 1 1 9180
0 9182 7 2 2 77302 82341
0 9183 7 1 2 67513 75478
0 9184 7 1 2 83113 9183
0 9185 5 1 1 9184
0 9186 7 1 2 9181 9185
0 9187 7 1 2 9172 9186
0 9188 5 1 1 9187
0 9189 7 1 2 65191 9188
0 9190 5 1 1 9189
0 9191 7 1 2 77414 77176
0 9192 5 1 1 9191
0 9193 7 1 2 75638 9192
0 9194 5 1 1 9193
0 9195 7 1 2 76774 71668
0 9196 5 1 1 9195
0 9197 7 1 2 75223 80349
0 9198 5 1 1 9197
0 9199 7 1 2 70389 74356
0 9200 5 2 1 9199
0 9201 7 1 2 75298 76443
0 9202 5 1 1 9201
0 9203 7 1 2 83115 9202
0 9204 7 1 2 9198 9203
0 9205 7 1 2 9196 9204
0 9206 5 1 1 9205
0 9207 7 1 2 77259 9206
0 9208 5 1 1 9207
0 9209 7 1 2 9194 9208
0 9210 5 1 1 9209
0 9211 7 1 2 69653 9210
0 9212 5 1 1 9211
0 9213 7 1 2 9190 9212
0 9214 5 1 1 9213
0 9215 7 1 2 60799 9214
0 9216 5 1 1 9215
0 9217 7 1 2 80700 81906
0 9218 5 1 1 9217
0 9219 7 2 2 63471 77384
0 9220 7 2 2 76057 67458
0 9221 7 1 2 83117 83119
0 9222 5 1 1 9221
0 9223 7 1 2 9218 9222
0 9224 5 1 1 9223
0 9225 7 1 2 58215 9224
0 9226 5 1 1 9225
0 9227 7 5 2 59282 74324
0 9228 5 1 1 83121
0 9229 7 3 2 66749 81894
0 9230 5 1 1 83126
0 9231 7 2 2 69654 83127
0 9232 7 1 2 83122 83129
0 9233 5 1 1 9232
0 9234 7 1 2 9226 9233
0 9235 5 1 1 9234
0 9236 7 1 2 67720 9235
0 9237 5 1 1 9236
0 9238 7 1 2 83058 71944
0 9239 7 1 2 82033 9238
0 9240 5 1 1 9239
0 9241 7 1 2 9237 9240
0 9242 7 1 2 9216 9241
0 9243 5 1 1 9242
0 9244 7 1 2 59483 9243
0 9245 5 1 1 9244
0 9246 7 2 2 75782 74616
0 9247 5 1 1 83131
0 9248 7 6 2 68337 83132
0 9249 5 6 1 83133
0 9250 7 1 2 71592 83139
0 9251 5 1 1 9250
0 9252 7 3 2 62050 67108
0 9253 7 1 2 76584 81887
0 9254 7 1 2 83145 9253
0 9255 7 1 2 70442 9254
0 9256 7 1 2 9251 9255
0 9257 5 1 1 9256
0 9258 7 1 2 9245 9257
0 9259 7 1 2 9152 9258
0 9260 5 1 1 9259
0 9261 7 1 2 58413 9260
0 9262 5 1 1 9261
0 9263 7 1 2 75713 72005
0 9264 5 2 1 9263
0 9265 7 1 2 57942 75930
0 9266 5 1 1 9265
0 9267 7 1 2 83148 9266
0 9268 5 1 1 9267
0 9269 7 1 2 75639 9268
0 9270 5 1 1 9269
0 9271 7 1 2 75926 75698
0 9272 5 1 1 9271
0 9273 7 1 2 69835 75731
0 9274 7 1 2 82777 9273
0 9275 5 1 1 9274
0 9276 7 1 2 9272 9275
0 9277 5 1 1 9276
0 9278 7 1 2 57943 9277
0 9279 5 1 1 9278
0 9280 7 1 2 58732 79631
0 9281 7 1 2 81790 9280
0 9282 5 1 1 9281
0 9283 7 1 2 9279 9282
0 9284 5 1 1 9283
0 9285 7 1 2 68587 9284
0 9286 5 1 1 9285
0 9287 7 1 2 74513 75812
0 9288 7 1 2 82521 9287
0 9289 5 1 1 9288
0 9290 7 1 2 9286 9289
0 9291 7 1 2 9270 9290
0 9292 5 1 1 9291
0 9293 7 1 2 60800 9292
0 9294 5 1 1 9293
0 9295 7 1 2 75805 71122
0 9296 7 1 2 81977 9295
0 9297 7 1 2 83134 9296
0 9298 5 1 1 9297
0 9299 7 1 2 9294 9298
0 9300 5 1 1 9299
0 9301 7 1 2 71151 68683
0 9302 7 1 2 9300 9301
0 9303 5 1 1 9302
0 9304 7 1 2 9262 9303
0 9305 5 1 1 9304
0 9306 7 1 2 66141 9305
0 9307 5 1 1 9306
0 9308 7 4 2 69239 75982
0 9309 7 1 2 72432 83150
0 9310 5 1 1 9309
0 9311 7 1 2 76139 9310
0 9312 5 1 1 9311
0 9313 7 1 2 57648 9312
0 9314 5 1 1 9313
0 9315 7 1 2 9314 8116
0 9316 5 1 1 9315
0 9317 7 1 2 57370 9316
0 9318 5 1 1 9317
0 9319 7 1 2 66750 71637
0 9320 7 1 2 72685 9319
0 9321 5 1 1 9320
0 9322 7 1 2 9318 9321
0 9323 5 1 1 9322
0 9324 7 1 2 64979 9323
0 9325 5 1 1 9324
0 9326 7 2 2 72258 75826
0 9327 7 1 2 83120 83154
0 9328 5 1 1 9327
0 9329 7 1 2 9325 9328
0 9330 5 1 1 9329
0 9331 7 20 2 67990 81034
0 9332 5 2 1 83156
0 9333 7 3 2 61524 73755
0 9334 7 1 2 83157 83178
0 9335 7 1 2 9330 9334
0 9336 5 1 1 9335
0 9337 7 1 2 64473 9336
0 9338 7 1 2 9307 9337
0 9339 7 1 2 9037 9338
0 9340 5 1 1 9339
0 9341 7 5 2 62607 59283
0 9342 5 3 1 83181
0 9343 7 1 2 75067 592
0 9344 5 1 1 9343
0 9345 7 2 2 60270 9344
0 9346 5 1 1 83189
0 9347 7 1 2 83182 83190
0 9348 5 2 1 9347
0 9349 7 1 2 62608 70001
0 9350 5 1 1 9349
0 9351 7 1 2 69380 9350
0 9352 5 1 1 9351
0 9353 7 1 2 77080 9352
0 9354 5 1 1 9353
0 9355 7 1 2 62321 9354
0 9356 5 1 1 9355
0 9357 7 2 2 65471 68588
0 9358 5 2 1 83193
0 9359 7 3 2 80070 83195
0 9360 5 1 1 83197
0 9361 7 1 2 57649 83198
0 9362 5 1 1 9361
0 9363 7 3 2 65472 75356
0 9364 5 1 1 83200
0 9365 7 1 2 9362 9364
0 9366 5 1 1 9365
0 9367 7 1 2 60271 9366
0 9368 5 1 1 9367
0 9369 7 2 2 4364 9368
0 9370 7 1 2 9356 83203
0 9371 5 1 1 9370
0 9372 7 1 2 63844 9371
0 9373 5 1 1 9372
0 9374 7 1 2 78804 797
0 9375 5 2 1 9374
0 9376 7 2 2 65192 70614
0 9377 5 2 1 83207
0 9378 7 1 2 83205 83208
0 9379 5 1 1 9378
0 9380 7 2 2 68472 78716
0 9381 7 1 2 74578 83211
0 9382 5 1 1 9381
0 9383 7 1 2 9379 9382
0 9384 5 1 1 9383
0 9385 7 1 2 60272 9384
0 9386 5 1 1 9385
0 9387 7 2 2 62609 59100
0 9388 5 1 1 83213
0 9389 7 1 2 72139 83214
0 9390 5 2 1 9389
0 9391 7 1 2 9386 83215
0 9392 7 1 2 9373 9391
0 9393 5 1 1 9392
0 9394 7 1 2 63986 9393
0 9395 5 1 1 9394
0 9396 7 1 2 83191 9395
0 9397 5 1 1 9396
0 9398 7 1 2 72169 9397
0 9399 5 1 1 9398
0 9400 7 6 2 74357 80282
0 9401 5 1 1 83217
0 9402 7 2 2 65193 74636
0 9403 5 2 1 83223
0 9404 7 2 2 9401 83225
0 9405 5 1 1 83227
0 9406 7 1 2 60801 83228
0 9407 5 1 1 9406
0 9408 7 2 2 62610 74358
0 9409 5 4 1 83229
0 9410 7 1 2 71868 71039
0 9411 5 3 1 9410
0 9412 7 1 2 60273 83235
0 9413 5 3 1 9412
0 9414 7 2 2 83231 83238
0 9415 5 1 1 83241
0 9416 7 1 2 65473 83242
0 9417 5 1 1 9416
0 9418 7 1 2 59284 9417
0 9419 7 1 2 9407 9418
0 9420 5 1 1 9419
0 9421 7 4 2 60802 74359
0 9422 5 14 1 83243
0 9423 7 1 2 83244 79762
0 9424 5 1 1 9423
0 9425 7 3 2 58216 74360
0 9426 5 1 1 83261
0 9427 7 3 2 57371 76561
0 9428 5 5 1 83264
0 9429 7 1 2 74361 83265
0 9430 5 3 1 9429
0 9431 7 2 2 62611 71674
0 9432 5 2 1 83275
0 9433 7 1 2 70723 78060
0 9434 7 1 2 83277 9433
0 9435 5 1 1 9434
0 9436 7 1 2 83272 9435
0 9437 5 1 1 9436
0 9438 7 1 2 65474 9437
0 9439 5 1 1 9438
0 9440 7 1 2 9426 9439
0 9441 5 1 1 9440
0 9442 7 1 2 63987 9441
0 9443 5 1 1 9442
0 9444 7 1 2 9424 9443
0 9445 7 1 2 9420 9444
0 9446 5 1 1 9445
0 9447 7 1 2 69655 9446
0 9448 5 1 1 9447
0 9449 7 1 2 9399 9448
0 9450 5 1 1 9449
0 9451 7 1 2 59484 9450
0 9452 5 1 1 9451
0 9453 7 4 2 57372 64199
0 9454 7 2 2 70348 69115
0 9455 5 1 1 83283
0 9456 7 1 2 83279 83284
0 9457 5 1 1 9456
0 9458 7 3 2 60803 83262
0 9459 5 1 1 83285
0 9460 7 1 2 80283 83286
0 9461 5 1 1 9460
0 9462 7 1 2 9457 9461
0 9463 5 1 1 9462
0 9464 7 1 2 67275 9463
0 9465 5 1 1 9464
0 9466 7 4 2 65475 68742
0 9467 5 2 1 83288
0 9468 7 2 2 83292 70109
0 9469 5 2 1 83294
0 9470 7 1 2 64200 83296
0 9471 5 1 1 9470
0 9472 7 2 2 77114 76944
0 9473 5 6 1 83298
0 9474 7 1 2 83245 83299
0 9475 5 1 1 9474
0 9476 7 1 2 9471 9475
0 9477 5 1 1 9476
0 9478 7 1 2 70390 9477
0 9479 5 1 1 9478
0 9480 7 1 2 62612 76408
0 9481 5 1 1 9480
0 9482 7 1 2 64201 78724
0 9483 7 1 2 9481 9482
0 9484 5 1 1 9483
0 9485 7 1 2 9479 9484
0 9486 7 1 2 9465 9485
0 9487 5 1 1 9486
0 9488 7 1 2 69656 9487
0 9489 5 1 1 9488
0 9490 7 1 2 9452 9489
0 9491 5 1 1 9490
0 9492 7 1 2 77260 9491
0 9493 5 1 1 9492
0 9494 7 2 2 70368 78815
0 9495 5 5 1 83306
0 9496 7 1 2 64202 83307
0 9497 5 1 1 9496
0 9498 7 1 2 60804 79073
0 9499 7 1 2 9497 9498
0 9500 5 1 1 9499
0 9501 7 1 2 73869 81215
0 9502 5 1 1 9501
0 9503 7 3 2 65476 77307
0 9504 7 2 2 75318 83313
0 9505 5 2 1 83316
0 9506 7 1 2 68743 83317
0 9507 5 1 1 9506
0 9508 7 1 2 9502 9507
0 9509 7 1 2 9500 9508
0 9510 5 1 1 9509
0 9511 7 1 2 69657 9510
0 9512 5 1 1 9511
0 9513 7 1 2 76531 81956
0 9514 5 1 1 9513
0 9515 7 1 2 70065 9514
0 9516 5 1 1 9515
0 9517 7 1 2 64203 9516
0 9518 5 1 1 9517
0 9519 7 1 2 65194 79948
0 9520 5 1 1 9519
0 9521 7 1 2 9518 9520
0 9522 5 1 1 9521
0 9523 7 1 2 59285 9522
0 9524 5 1 1 9523
0 9525 7 1 2 70036 78064
0 9526 5 2 1 9525
0 9527 7 2 2 57944 70027
0 9528 5 1 1 83322
0 9529 7 2 2 60513 9528
0 9530 5 1 1 83324
0 9531 7 1 2 62322 83325
0 9532 5 1 1 9531
0 9533 7 1 2 83320 9532
0 9534 5 1 1 9533
0 9535 7 1 2 71152 9534
0 9536 5 1 1 9535
0 9537 7 1 2 9524 9536
0 9538 5 1 1 9537
0 9539 7 1 2 65477 9538
0 9540 5 1 1 9539
0 9541 7 4 2 62323 59485
0 9542 7 2 2 60805 83326
0 9543 7 1 2 74460 80162
0 9544 5 2 1 9543
0 9545 7 1 2 83330 83332
0 9546 5 2 1 9545
0 9547 7 3 2 62613 76354
0 9548 5 1 1 83336
0 9549 7 1 2 57373 9548
0 9550 5 2 1 9549
0 9551 7 2 2 57945 81614
0 9552 5 3 1 83341
0 9553 7 1 2 83339 83343
0 9554 5 1 1 9553
0 9555 7 1 2 67645 9554
0 9556 5 1 1 9555
0 9557 7 2 2 6254 9556
0 9558 5 1 1 83346
0 9559 7 1 2 64204 9558
0 9560 5 1 1 9559
0 9561 7 1 2 83334 9560
0 9562 5 1 1 9561
0 9563 7 1 2 58217 9562
0 9564 5 1 1 9563
0 9565 7 5 2 59286 70701
0 9566 7 5 2 75714 83348
0 9567 5 2 1 83353
0 9568 7 1 2 77565 83354
0 9569 5 2 1 9568
0 9570 7 1 2 9564 83360
0 9571 7 1 2 9540 9570
0 9572 5 1 1 9571
0 9573 7 1 2 69573 9572
0 9574 5 1 1 9573
0 9575 7 1 2 9512 9574
0 9576 5 1 1 9575
0 9577 7 1 2 75640 9576
0 9578 5 1 1 9577
0 9579 7 1 2 9493 9578
0 9580 5 1 1 9579
0 9581 7 1 2 58414 9580
0 9582 5 1 1 9581
0 9583 7 1 2 77212 76012
0 9584 5 1 1 9583
0 9585 7 6 2 59981 74289
0 9586 7 3 2 82796 83362
0 9587 5 1 1 83368
0 9588 7 1 2 65195 83369
0 9589 5 1 1 9588
0 9590 7 1 2 9584 9589
0 9591 5 1 1 9590
0 9592 7 1 2 64980 9591
0 9593 5 1 1 9592
0 9594 7 2 2 66822 68930
0 9595 5 5 1 83371
0 9596 7 1 2 74186 77261
0 9597 5 1 1 9596
0 9598 7 1 2 83373 9597
0 9599 5 2 1 9598
0 9600 7 1 2 80711 83378
0 9601 5 1 1 9600
0 9602 7 1 2 9593 9601
0 9603 5 1 1 9602
0 9604 7 1 2 67646 9603
0 9605 5 1 1 9604
0 9606 7 4 2 59982 68931
0 9607 7 2 2 83005 83380
0 9608 5 1 1 83384
0 9609 7 1 2 57946 75816
0 9610 5 1 1 9609
0 9611 7 1 2 68919 75983
0 9612 5 3 1 9611
0 9613 7 1 2 9610 83386
0 9614 5 1 1 9613
0 9615 7 1 2 74187 9614
0 9616 5 1 1 9615
0 9617 7 1 2 9608 9616
0 9618 5 1 1 9617
0 9619 7 1 2 65196 9618
0 9620 5 1 1 9619
0 9621 7 1 2 9605 9620
0 9622 5 1 1 9621
0 9623 7 1 2 59486 9622
0 9624 5 1 1 9623
0 9625 7 1 2 65478 82825
0 9626 5 1 1 9625
0 9627 7 1 2 9624 9626
0 9628 5 1 1 9627
0 9629 7 1 2 69658 9628
0 9630 5 1 1 9629
0 9631 7 2 2 73996 70702
0 9632 7 5 2 59487 66680
0 9633 7 1 2 76025 83391
0 9634 7 1 2 83389 9633
0 9635 7 3 2 64981 74290
0 9636 7 2 2 58733 74165
0 9637 7 1 2 83396 83399
0 9638 7 1 2 9634 9637
0 9639 5 1 1 9638
0 9640 7 1 2 9630 9639
0 9641 5 1 1 9640
0 9642 7 1 2 58218 9641
0 9643 5 1 1 9642
0 9644 7 1 2 80650 69172
0 9645 7 1 2 82283 82372
0 9646 7 1 2 9644 9645
0 9647 5 1 1 9646
0 9648 7 1 2 9643 9647
0 9649 5 1 1 9648
0 9650 7 1 2 68589 9649
0 9651 5 1 1 9650
0 9652 7 1 2 67888 78678
0 9653 5 1 1 9652
0 9654 7 1 2 83318 9653
0 9655 5 1 1 9654
0 9656 7 1 2 68744 9655
0 9657 5 1 1 9656
0 9658 7 7 2 59287 67647
0 9659 7 2 2 77763 83401
0 9660 5 1 1 83408
0 9661 7 1 2 67991 80592
0 9662 5 1 1 9661
0 9663 7 1 2 78812 72042
0 9664 5 1 1 9663
0 9665 7 1 2 9662 9664
0 9666 5 1 1 9665
0 9667 7 1 2 83247 9666
0 9668 5 1 1 9667
0 9669 7 1 2 9660 9668
0 9670 7 1 2 9657 9669
0 9671 5 1 1 9670
0 9672 7 1 2 75641 9671
0 9673 5 1 1 9672
0 9674 7 1 2 83402 73398
0 9675 5 2 1 9674
0 9676 7 2 2 65479 67889
0 9677 7 1 2 77115 71621
0 9678 7 1 2 83412 9677
0 9679 5 1 1 9678
0 9680 7 1 2 83410 9679
0 9681 5 1 1 9680
0 9682 7 1 2 63162 9681
0 9683 5 1 1 9682
0 9684 7 1 2 74974 83355
0 9685 5 1 1 9684
0 9686 7 1 2 9683 9685
0 9687 5 1 1 9686
0 9688 7 1 2 77262 9687
0 9689 5 1 1 9688
0 9690 7 1 2 9673 9689
0 9691 5 1 1 9690
0 9692 7 1 2 69659 9691
0 9693 5 1 1 9692
0 9694 7 1 2 83248 75642
0 9695 5 1 1 9694
0 9696 7 7 2 63472 64982
0 9697 5 1 1 83414
0 9698 7 1 2 65480 83415
0 9699 7 1 2 75822 9698
0 9700 5 1 1 9699
0 9701 7 1 2 9695 9700
0 9702 5 1 1 9701
0 9703 7 1 2 68745 9702
0 9704 5 1 1 9703
0 9705 7 1 2 3480 9704
0 9706 5 1 1 9705
0 9707 7 5 2 63163 63595
0 9708 7 3 2 83421 69240
0 9709 7 1 2 82440 83426
0 9710 7 1 2 9706 9709
0 9711 5 1 1 9710
0 9712 7 1 2 9693 9711
0 9713 5 1 1 9712
0 9714 7 1 2 71153 9713
0 9715 5 1 1 9714
0 9716 7 2 2 67918 74795
0 9717 7 3 2 59288 71469
0 9718 7 1 2 74291 83431
0 9719 7 1 2 83429 9718
0 9720 7 3 2 57947 77308
0 9721 5 2 1 83434
0 9722 7 8 2 57650 69116
0 9723 5 2 1 83439
0 9724 7 2 2 83440 82783
0 9725 7 1 2 83435 83449
0 9726 7 1 2 9719 9725
0 9727 5 1 1 9726
0 9728 7 1 2 61525 9727
0 9729 7 1 2 9715 9728
0 9730 7 1 2 9651 9729
0 9731 7 1 2 9582 9730
0 9732 5 1 1 9731
0 9733 7 1 2 72159 75027
0 9734 5 7 1 9733
0 9735 7 1 2 80701 83451
0 9736 5 1 1 9735
0 9737 7 1 2 62614 77192
0 9738 5 1 1 9737
0 9739 7 1 2 9736 9738
0 9740 5 1 1 9739
0 9741 7 1 2 58219 9740
0 9742 5 1 1 9741
0 9743 7 6 2 63752 74940
0 9744 7 1 2 69961 71993
0 9745 7 1 2 83458 9744
0 9746 5 1 1 9745
0 9747 7 1 2 9742 9746
0 9748 5 1 1 9747
0 9749 7 1 2 67721 9748
0 9750 5 1 1 9749
0 9751 7 4 2 62324 75124
0 9752 5 7 1 83464
0 9753 7 2 2 69836 83465
0 9754 5 1 1 83475
0 9755 7 1 2 70158 83476
0 9756 5 1 1 9755
0 9757 7 2 2 65481 77461
0 9758 5 1 1 83477
0 9759 7 1 2 71798 83478
0 9760 5 1 1 9759
0 9761 7 1 2 75028 9360
0 9762 5 1 1 9761
0 9763 7 1 2 60274 77657
0 9764 7 1 2 9762 9763
0 9765 5 1 1 9764
0 9766 7 1 2 9760 9765
0 9767 5 1 1 9766
0 9768 7 1 2 58220 9767
0 9769 5 1 1 9768
0 9770 7 1 2 9756 9769
0 9771 7 1 2 9750 9770
0 9772 5 1 1 9771
0 9773 7 1 2 75643 9772
0 9774 5 1 1 9773
0 9775 7 5 2 58221 63753
0 9776 7 1 2 76994 83479
0 9777 7 1 2 81016 77263
0 9778 7 1 2 9776 9777
0 9779 5 1 1 9778
0 9780 7 1 2 9774 9779
0 9781 5 1 1 9780
0 9782 7 1 2 69267 9781
0 9783 5 1 1 9782
0 9784 7 2 2 78591 78712
0 9785 5 1 1 83484
0 9786 7 3 2 63754 65482
0 9787 5 1 1 83486
0 9788 7 3 2 62162 83487
0 9789 5 2 1 83489
0 9790 7 1 2 9785 83492
0 9791 5 1 1 9790
0 9792 7 1 2 75644 9791
0 9793 5 1 1 9792
0 9794 7 1 2 69962 78679
0 9795 5 1 1 9794
0 9796 7 1 2 70661 9795
0 9797 5 1 1 9796
0 9798 7 1 2 74637 9797
0 9799 5 2 1 9798
0 9800 7 1 2 74611 82753
0 9801 5 1 1 9800
0 9802 7 1 2 65483 9801
0 9803 7 1 2 82758 9802
0 9804 5 1 1 9803
0 9805 7 1 2 59289 71044
0 9806 5 2 1 9805
0 9807 7 1 2 80102 83496
0 9808 5 1 1 9807
0 9809 7 1 2 60275 9808
0 9810 5 1 1 9809
0 9811 7 1 2 63988 72400
0 9812 5 1 1 9811
0 9813 7 1 2 60276 9812
0 9814 5 1 1 9813
0 9815 7 1 2 75230 9814
0 9816 5 1 1 9815
0 9817 7 1 2 67841 9816
0 9818 5 1 1 9817
0 9819 7 1 2 57948 74961
0 9820 5 4 1 9819
0 9821 7 1 2 60806 83498
0 9822 7 1 2 9818 9821
0 9823 7 1 2 9810 9822
0 9824 5 1 1 9823
0 9825 7 1 2 9804 9824
0 9826 5 1 1 9825
0 9827 7 1 2 83494 9826
0 9828 5 1 1 9827
0 9829 7 1 2 75760 9828
0 9830 5 1 1 9829
0 9831 7 1 2 9793 9830
0 9832 5 1 1 9831
0 9833 7 1 2 69660 9832
0 9834 5 1 1 9833
0 9835 7 1 2 9783 9834
0 9836 5 1 1 9835
0 9837 7 1 2 59488 9836
0 9838 5 1 1 9837
0 9839 7 1 2 69837 76130
0 9840 5 1 1 9839
0 9841 7 1 2 69588 82059
0 9842 5 1 1 9841
0 9843 7 1 2 9840 9842
0 9844 5 1 1 9843
0 9845 7 1 2 58222 9844
0 9846 5 1 1 9845
0 9847 7 1 2 75704 9163
0 9848 5 2 1 9847
0 9849 7 1 2 57949 83502
0 9850 5 1 1 9849
0 9851 7 1 2 83387 9850
0 9852 5 1 1 9851
0 9853 7 1 2 69495 9852
0 9854 5 1 1 9853
0 9855 7 1 2 9846 9854
0 9856 5 1 1 9855
0 9857 7 1 2 60807 9856
0 9858 5 1 1 9857
0 9859 7 2 2 65484 83104
0 9860 5 1 1 83504
0 9861 7 5 2 57950 60514
0 9862 5 2 1 83506
0 9863 7 1 2 68920 83507
0 9864 7 1 2 83505 9863
0 9865 5 1 1 9864
0 9866 7 1 2 9858 9865
0 9867 5 1 1 9866
0 9868 7 1 2 68590 9867
0 9869 5 1 1 9868
0 9870 7 1 2 69360 81765
0 9871 5 1 1 9870
0 9872 7 1 2 82253 9871
0 9873 5 1 1 9872
0 9874 7 1 2 68746 9873
0 9875 5 2 1 9874
0 9876 7 6 2 63596 66823
0 9877 5 1 1 83515
0 9878 7 1 2 74782 67544
0 9879 7 1 2 83516 9878
0 9880 5 1 1 9879
0 9881 7 1 2 76140 9880
0 9882 5 1 1 9881
0 9883 7 1 2 59290 9882
0 9884 5 1 1 9883
0 9885 7 1 2 83513 9884
0 9886 5 1 1 9885
0 9887 7 1 2 65485 9886
0 9888 5 1 1 9887
0 9889 7 1 2 65197 83112
0 9890 5 1 1 9889
0 9891 7 1 2 9888 9890
0 9892 5 1 1 9891
0 9893 7 1 2 64205 9892
0 9894 5 1 1 9893
0 9895 7 1 2 70670 82050
0 9896 5 1 1 9895
0 9897 7 1 2 82073 83097
0 9898 5 1 1 9897
0 9899 7 1 2 81925 9898
0 9900 5 1 1 9899
0 9901 7 1 2 58223 9900
0 9902 5 2 1 9901
0 9903 7 1 2 65198 76001
0 9904 5 1 1 9903
0 9905 7 1 2 76852 9904
0 9906 7 1 2 82775 9905
0 9907 5 1 1 9906
0 9908 7 1 2 83521 9907
0 9909 5 1 1 9908
0 9910 7 1 2 60808 9909
0 9911 5 1 1 9910
0 9912 7 1 2 9896 9911
0 9913 7 1 2 9894 9912
0 9914 5 1 1 9913
0 9915 7 1 2 57951 9914
0 9916 5 1 1 9915
0 9917 7 1 2 9869 9916
0 9918 5 1 1 9917
0 9919 7 1 2 67648 9918
0 9920 5 1 1 9919
0 9921 7 1 2 64206 77325
0 9922 5 1 1 9921
0 9923 7 2 2 83059 77282
0 9924 5 1 1 83523
0 9925 7 1 2 78680 83524
0 9926 5 1 1 9925
0 9927 7 1 2 9922 9926
0 9928 5 1 1 9927
0 9929 7 1 2 67276 9928
0 9930 5 1 1 9929
0 9931 7 1 2 79580 75761
0 9932 5 2 1 9931
0 9933 7 1 2 72140 75984
0 9934 5 1 1 9933
0 9935 7 1 2 83525 9934
0 9936 5 1 1 9935
0 9937 7 1 2 70391 9936
0 9938 5 1 1 9937
0 9939 7 1 2 9930 9938
0 9940 5 1 1 9939
0 9941 7 1 2 68747 9940
0 9942 5 1 1 9941
0 9943 7 1 2 69309 82316
0 9944 5 1 1 9943
0 9945 7 2 2 73161 74141
0 9946 7 1 2 83527 81780
0 9947 5 1 1 9946
0 9948 7 1 2 9944 9947
0 9949 5 1 1 9948
0 9950 7 1 2 68748 9949
0 9951 5 1 1 9950
0 9952 7 1 2 68749 72676
0 9953 7 1 2 83128 9952
0 9954 5 1 1 9953
0 9955 7 1 2 3638 9954
0 9956 5 1 1 9955
0 9957 7 1 2 60515 9956
0 9958 5 1 1 9957
0 9959 7 1 2 9951 9958
0 9960 5 1 1 9959
0 9961 7 1 2 67649 9960
0 9962 5 1 1 9961
0 9963 7 1 2 59291 74975
0 9964 5 4 1 9963
0 9965 7 1 2 77568 83529
0 9966 5 1 1 9965
0 9967 7 1 2 67842 9966
0 9968 5 1 1 9967
0 9969 7 1 2 67722 75105
0 9970 5 1 1 9969
0 9971 7 1 2 69731 9970
0 9972 5 1 1 9971
0 9973 7 1 2 9968 9972
0 9974 5 1 1 9973
0 9975 7 1 2 82835 9974
0 9976 5 1 1 9975
0 9977 7 1 2 9962 9976
0 9978 7 1 2 9942 9977
0 9979 5 1 1 9978
0 9980 7 1 2 69661 9979
0 9981 5 1 1 9980
0 9982 7 1 2 83067 83388
0 9983 5 1 1 9982
0 9984 7 1 2 57952 9983
0 9985 5 1 1 9984
0 9986 7 1 2 58224 83503
0 9987 5 1 1 9986
0 9988 7 1 2 9985 9987
0 9989 5 1 1 9988
0 9990 7 6 2 67919 77377
0 9991 5 1 1 83533
0 9992 7 1 2 72542 83534
0 9993 7 1 2 9989 9992
0 9994 5 1 1 9993
0 9995 7 1 2 63164 9994
0 9996 7 1 2 9981 9995
0 9997 7 1 2 9920 9996
0 9998 7 1 2 9838 9997
0 9999 5 1 1 9998
0 10000 7 2 2 75354 1948
0 10001 7 1 2 70196 76131
0 10002 7 1 2 83539 10001
0 10003 5 2 1 10002
0 10004 7 1 2 78548 72104
0 10005 7 1 2 83517 10004
0 10006 7 1 2 75384 10005
0 10007 5 1 1 10006
0 10008 7 1 2 83541 10007
0 10009 5 1 1 10008
0 10010 7 1 2 67723 10009
0 10011 5 1 1 10010
0 10012 7 1 2 69932 74999
0 10013 5 1 1 10012
0 10014 7 1 2 68473 10013
0 10015 5 2 1 10014
0 10016 7 1 2 77955 83543
0 10017 5 1 1 10016
0 10018 7 1 2 77264 10017
0 10019 5 1 1 10018
0 10020 7 1 2 63989 75985
0 10021 5 1 1 10020
0 10022 7 1 2 10019 10021
0 10023 5 1 1 10022
0 10024 7 1 2 62325 10023
0 10025 5 1 1 10024
0 10026 7 1 2 83374 81815
0 10027 5 1 1 10026
0 10028 7 1 2 63990 10027
0 10029 5 1 1 10028
0 10030 7 1 2 10025 10029
0 10031 5 1 1 10030
0 10032 7 1 2 69662 10031
0 10033 5 1 1 10032
0 10034 7 1 2 10011 10033
0 10035 5 1 1 10034
0 10036 7 1 2 64207 10035
0 10037 5 1 1 10036
0 10038 7 1 2 74843 81922
0 10039 5 1 1 10038
0 10040 7 1 2 70615 75986
0 10041 5 1 1 10040
0 10042 7 1 2 10039 10041
0 10043 5 1 1 10042
0 10044 7 2 2 81031 10043
0 10045 7 1 2 77389 83545
0 10046 5 1 1 10045
0 10047 7 1 2 10037 10046
0 10048 5 1 1 10047
0 10049 7 1 2 62615 10048
0 10050 5 1 1 10049
0 10051 7 1 2 79927 83546
0 10052 5 1 1 10051
0 10053 7 1 2 58415 10052
0 10054 7 1 2 10050 10053
0 10055 5 1 1 10054
0 10056 7 1 2 9999 10055
0 10057 5 1 1 10056
0 10058 7 1 2 78004 70197
0 10059 7 1 2 77330 10058
0 10060 5 1 1 10059
0 10061 7 1 2 83526 10060
0 10062 5 1 1 10061
0 10063 7 1 2 80465 10062
0 10064 5 1 1 10063
0 10065 7 1 2 77385 77510
0 10066 7 1 2 82030 10065
0 10067 5 1 1 10066
0 10068 7 1 2 10064 10067
0 10069 5 1 1 10068
0 10070 7 1 2 68474 10069
0 10071 5 1 1 10070
0 10072 7 1 2 60516 69732
0 10073 5 1 1 10072
0 10074 7 1 2 72141 75391
0 10075 5 2 1 10074
0 10076 7 1 2 10073 83547
0 10077 5 1 1 10076
0 10078 7 1 2 80456 83151
0 10079 7 1 2 10077 10078
0 10080 5 1 1 10079
0 10081 7 1 2 10071 10080
0 10082 5 1 1 10081
0 10083 7 1 2 68222 10082
0 10084 5 1 1 10083
0 10085 7 8 2 58734 58850
0 10086 5 1 1 83549
0 10087 7 6 2 76605 83550
0 10088 7 2 2 77340 83557
0 10089 7 1 2 74292 77049
0 10090 7 1 2 83563 10089
0 10091 5 1 1 10090
0 10092 7 1 2 10084 10091
0 10093 5 1 1 10092
0 10094 7 1 2 62616 10093
0 10095 5 1 1 10094
0 10096 7 1 2 77283 81910
0 10097 5 1 1 10096
0 10098 7 1 2 72142 67514
0 10099 7 1 2 81931 10098
0 10100 5 1 1 10099
0 10101 7 1 2 10097 10100
0 10102 5 1 1 10101
0 10103 7 1 2 68475 10102
0 10104 5 1 1 10103
0 10105 7 1 2 72072 76132
0 10106 5 2 1 10105
0 10107 7 1 2 9860 83565
0 10108 7 1 2 10104 10107
0 10109 5 1 1 10108
0 10110 7 1 2 60277 10109
0 10111 5 1 1 10110
0 10112 7 1 2 64208 76133
0 10113 5 1 1 10112
0 10114 7 2 2 69241 72610
0 10115 7 1 2 77890 83567
0 10116 5 1 1 10115
0 10117 7 1 2 9991 10116
0 10118 5 1 1 10117
0 10119 7 1 2 75645 10118
0 10120 5 1 1 10119
0 10121 7 1 2 10113 10120
0 10122 7 1 2 10111 10121
0 10123 5 1 1 10122
0 10124 7 1 2 63991 10123
0 10125 5 1 1 10124
0 10126 7 1 2 79527 4891
0 10127 5 1 1 10126
0 10128 7 1 2 81766 10127
0 10129 5 1 1 10128
0 10130 7 1 2 81904 10129
0 10131 5 1 1 10130
0 10132 7 1 2 64209 10131
0 10133 5 1 1 10132
0 10134 7 3 2 62163 81666
0 10135 5 4 1 83569
0 10136 7 1 2 69838 83570
0 10137 5 1 1 10136
0 10138 7 1 2 69753 10137
0 10139 5 1 1 10138
0 10140 7 1 2 80344 83152
0 10141 7 1 2 10139 10140
0 10142 5 1 1 10141
0 10143 7 1 2 83542 10142
0 10144 5 1 1 10143
0 10145 7 1 2 62326 10144
0 10146 5 1 1 10145
0 10147 7 1 2 10133 10146
0 10148 7 1 2 10125 10147
0 10149 5 1 1 10148
0 10150 7 1 2 62617 10149
0 10151 5 1 1 10150
0 10152 7 1 2 63845 76134
0 10153 5 1 1 10152
0 10154 7 1 2 79545 81767
0 10155 5 1 1 10154
0 10156 7 1 2 10153 10155
0 10157 5 1 1 10156
0 10158 7 1 2 68476 10157
0 10159 5 1 1 10158
0 10160 7 1 2 83566 10159
0 10161 5 1 1 10160
0 10162 7 1 2 62327 10161
0 10163 5 1 1 10162
0 10164 7 2 2 63846 75098
0 10165 5 2 1 83576
0 10166 7 1 2 75762 83577
0 10167 5 1 1 10166
0 10168 7 1 2 83375 10167
0 10169 5 1 1 10168
0 10170 7 1 2 69663 10169
0 10171 5 1 1 10170
0 10172 7 1 2 10163 10171
0 10173 5 1 1 10172
0 10174 7 1 2 64210 10173
0 10175 5 1 1 10174
0 10176 7 1 2 77966 69664
0 10177 5 1 1 10176
0 10178 7 2 2 66681 83452
0 10179 7 1 2 64211 69782
0 10180 7 1 2 69518 10179
0 10181 7 1 2 83580 10180
0 10182 5 1 1 10181
0 10183 7 1 2 10177 10182
0 10184 5 1 1 10183
0 10185 7 1 2 75646 10184
0 10186 5 1 1 10185
0 10187 7 6 2 64212 69381
0 10188 7 1 2 67459 83582
0 10189 7 1 2 79966 10188
0 10190 5 1 1 10189
0 10191 7 1 2 10186 10190
0 10192 5 1 1 10191
0 10193 7 1 2 70616 10192
0 10194 5 1 1 10193
0 10195 7 1 2 76796 69215
0 10196 7 1 2 81888 81928
0 10197 7 1 2 10195 10196
0 10198 5 1 1 10197
0 10199 7 1 2 10194 10198
0 10200 7 1 2 10175 10199
0 10201 7 1 2 10151 10200
0 10202 5 1 1 10201
0 10203 7 1 2 58416 10202
0 10204 5 1 1 10203
0 10205 7 1 2 10095 10204
0 10206 5 1 1 10205
0 10207 7 1 2 62899 10206
0 10208 5 1 1 10207
0 10209 7 1 2 66142 10208
0 10210 7 1 2 10057 10209
0 10211 5 1 1 10210
0 10212 7 1 2 9732 10211
0 10213 5 1 1 10212
0 10214 7 1 2 70078 80712
0 10215 5 1 1 10214
0 10216 7 1 2 70369 10215
0 10217 5 1 1 10216
0 10218 7 1 2 64213 10217
0 10219 5 1 1 10218
0 10220 7 1 2 5951 10219
0 10221 5 1 1 10220
0 10222 7 1 2 69665 10221
0 10223 5 1 1 10222
0 10224 7 3 2 63992 69382
0 10225 5 2 1 83588
0 10226 7 1 2 77449 83589
0 10227 7 1 2 72170 10226
0 10228 5 1 1 10227
0 10229 7 1 2 10223 10228
0 10230 5 1 1 10229
0 10231 7 1 2 65486 10230
0 10232 5 1 1 10231
0 10233 7 1 2 72819 75221
0 10234 5 1 1 10233
0 10235 7 1 2 77713 10234
0 10236 5 1 1 10235
0 10237 7 1 2 59292 10236
0 10238 5 1 1 10237
0 10239 7 1 2 68750 69839
0 10240 5 2 1 10239
0 10241 7 1 2 83511 83593
0 10242 5 1 1 10241
0 10243 7 1 2 71470 10242
0 10244 5 1 1 10243
0 10245 7 1 2 10238 10244
0 10246 5 1 1 10245
0 10247 7 1 2 10246 83535
0 10248 5 1 1 10247
0 10249 7 1 2 10232 10248
0 10250 5 1 1 10249
0 10251 7 1 2 77265 10250
0 10252 5 1 1 10251
0 10253 7 1 2 60809 76545
0 10254 5 3 1 10253
0 10255 7 2 2 64983 83595
0 10256 5 1 1 83598
0 10257 7 1 2 74142 83599
0 10258 5 1 1 10257
0 10259 7 1 2 5993 10258
0 10260 5 1 1 10259
0 10261 7 1 2 67277 10260
0 10262 5 1 1 10261
0 10263 7 4 2 60810 69413
0 10264 5 1 1 83600
0 10265 7 1 2 78262 83601
0 10266 5 1 1 10265
0 10267 7 1 2 10262 10266
0 10268 5 1 1 10267
0 10269 7 1 2 69666 10268
0 10270 5 1 1 10269
0 10271 7 1 2 71622 72677
0 10272 5 1 1 10271
0 10273 7 1 2 81289 10272
0 10274 5 1 1 10273
0 10275 7 1 2 77517 69574
0 10276 7 1 2 10274 10275
0 10277 5 1 1 10276
0 10278 7 1 2 10270 10277
0 10279 5 1 1 10278
0 10280 7 1 2 75647 10279
0 10281 5 1 1 10280
0 10282 7 1 2 10252 10281
0 10283 5 1 1 10282
0 10284 7 1 2 58417 10283
0 10285 5 1 1 10284
0 10286 7 1 2 64984 83372
0 10287 5 3 1 10286
0 10288 7 2 2 64985 74188
0 10289 5 1 1 83607
0 10290 7 1 2 83530 10289
0 10291 5 1 1 10290
0 10292 7 1 2 77266 10291
0 10293 5 1 1 10292
0 10294 7 1 2 83604 10293
0 10295 5 1 1 10294
0 10296 7 1 2 68751 10295
0 10297 5 1 1 10296
0 10298 7 1 2 74395 75648
0 10299 5 1 1 10298
0 10300 7 1 2 10297 10299
0 10301 5 1 1 10300
0 10302 7 1 2 65199 10301
0 10303 5 1 1 10302
0 10304 7 1 2 82823 83381
0 10305 5 1 1 10304
0 10306 7 1 2 74189 75817
0 10307 5 1 1 10306
0 10308 7 1 2 10305 10307
0 10309 7 1 2 10303 10308
0 10310 5 1 1 10309
0 10311 7 1 2 57953 10310
0 10312 5 1 1 10311
0 10313 7 1 2 78821 83379
0 10314 5 1 1 10313
0 10315 7 1 2 9587 10314
0 10316 5 1 1 10315
0 10317 7 1 2 64986 10316
0 10318 5 1 1 10317
0 10319 7 1 2 3482 10318
0 10320 5 1 1 10319
0 10321 7 1 2 59293 10320
0 10322 5 1 1 10321
0 10323 7 1 2 10312 10322
0 10324 5 1 1 10323
0 10325 7 1 2 69667 10324
0 10326 5 1 1 10325
0 10327 7 1 2 80642 80183
0 10328 7 3 2 58735 69146
0 10329 7 1 2 76041 83609
0 10330 7 1 2 10327 10329
0 10331 5 1 1 10330
0 10332 7 1 2 10326 10331
0 10333 5 1 1 10332
0 10334 7 1 2 71154 10333
0 10335 5 1 1 10334
0 10336 7 1 2 10285 10335
0 10337 5 1 1 10336
0 10338 7 1 2 61526 10337
0 10339 5 1 1 10338
0 10340 7 1 2 75954 76050
0 10341 5 1 1 10340
0 10342 7 1 2 74663 81923
0 10343 5 1 1 10342
0 10344 7 1 2 10341 10343
0 10345 5 1 1 10344
0 10346 7 1 2 69668 10345
0 10347 5 1 1 10346
0 10348 7 1 2 83522 10347
0 10349 5 1 1 10348
0 10350 7 1 2 60811 10349
0 10351 5 1 1 10350
0 10352 7 1 2 76002 75814
0 10353 5 1 1 10352
0 10354 7 1 2 69669 10353
0 10355 5 1 1 10354
0 10356 7 1 2 83514 10355
0 10357 5 1 1 10356
0 10358 7 1 2 65487 10357
0 10359 5 1 1 10358
0 10360 7 2 2 69670 71359
0 10361 5 1 1 83612
0 10362 7 4 2 63473 82630
0 10363 7 1 2 68752 83614
0 10364 7 1 2 83613 10363
0 10365 5 1 1 10364
0 10366 7 1 2 10359 10365
0 10367 5 1 1 10366
0 10368 7 1 2 64214 10367
0 10369 5 1 1 10368
0 10370 7 1 2 10351 10369
0 10371 5 1 1 10370
0 10372 7 1 2 57954 10371
0 10373 5 1 1 10372
0 10374 7 1 2 79614 79649
0 10375 5 1 1 10374
0 10376 7 2 2 60278 69711
0 10377 5 1 1 83618
0 10378 7 1 2 59294 83619
0 10379 5 1 1 10378
0 10380 7 1 2 10375 10379
0 10381 5 1 1 10380
0 10382 7 1 2 77267 10381
0 10383 5 1 1 10382
0 10384 7 4 2 60812 71471
0 10385 5 3 1 83620
0 10386 7 2 2 69764 83624
0 10387 5 1 1 83627
0 10388 7 1 2 10387 75649
0 10389 5 1 1 10388
0 10390 7 1 2 10383 10389
0 10391 5 1 1 10390
0 10392 7 1 2 69671 10391
0 10393 5 1 1 10392
0 10394 7 1 2 10373 10393
0 10395 5 1 1 10394
0 10396 7 1 2 65200 10395
0 10397 5 1 1 10396
0 10398 7 1 2 57955 82320
0 10399 5 1 1 10398
0 10400 7 1 2 60517 83071
0 10401 5 1 1 10400
0 10402 7 1 2 10399 10401
0 10403 5 1 1 10402
0 10404 7 1 2 59295 10403
0 10405 5 1 1 10404
0 10406 7 1 2 76780 75763
0 10407 5 1 1 10406
0 10408 7 1 2 82322 10407
0 10409 5 1 1 10408
0 10410 7 1 2 71472 10409
0 10411 5 1 1 10410
0 10412 7 1 2 60813 10411
0 10413 7 1 2 10405 10412
0 10414 5 1 1 10413
0 10415 7 2 2 66563 70392
0 10416 7 1 2 64987 83012
0 10417 7 1 2 83629 10416
0 10418 5 1 1 10417
0 10419 7 2 2 68753 66824
0 10420 7 1 2 82819 83631
0 10421 5 1 1 10420
0 10422 7 1 2 65488 10421
0 10423 7 1 2 10418 10422
0 10424 5 1 1 10423
0 10425 7 1 2 69672 10424
0 10426 7 1 2 10414 10425
0 10427 5 1 1 10426
0 10428 7 1 2 10397 10427
0 10429 5 1 1 10428
0 10430 7 1 2 82866 10429
0 10431 5 1 1 10430
0 10432 7 1 2 64215 81990
0 10433 5 1 1 10432
0 10434 7 1 2 83376 10433
0 10435 5 1 1 10434
0 10436 7 1 2 70393 10435
0 10437 5 1 1 10436
0 10438 7 7 2 58736 59489
0 10439 7 1 2 83382 83633
0 10440 5 1 1 10439
0 10441 7 1 2 10437 10440
0 10442 5 1 1 10441
0 10443 7 1 2 58418 10442
0 10444 5 1 1 10443
0 10445 7 7 2 67992 71155
0 10446 5 2 1 83640
0 10447 7 1 2 63165 81991
0 10448 5 1 1 10447
0 10449 7 1 2 83377 10448
0 10450 5 1 1 10449
0 10451 7 1 2 83641 10450
0 10452 5 1 1 10451
0 10453 7 1 2 10444 10452
0 10454 5 1 1 10453
0 10455 7 1 2 61527 10454
0 10456 5 1 1 10455
0 10457 7 4 2 65489 81110
0 10458 7 5 2 58737 82272
0 10459 7 1 2 83649 83653
0 10460 5 1 1 10459
0 10461 7 13 2 63166 63474
0 10462 7 1 2 75732 81383
0 10463 7 2 2 83658 10462
0 10464 5 1 1 83671
0 10465 7 1 2 10460 10464
0 10466 5 1 1 10465
0 10467 7 1 2 58225 10466
0 10468 5 1 1 10467
0 10469 7 1 2 58419 66825
0 10470 7 1 2 83650 10469
0 10471 5 1 1 10470
0 10472 7 1 2 59490 83672
0 10473 5 1 1 10472
0 10474 7 1 2 10471 10473
0 10475 7 1 2 10468 10474
0 10476 5 1 1 10475
0 10477 7 1 2 60279 10476
0 10478 5 1 1 10477
0 10479 7 1 2 66143 74514
0 10480 7 1 2 83370 10479
0 10481 5 1 1 10480
0 10482 7 1 2 10478 10481
0 10483 5 1 1 10482
0 10484 7 1 2 67278 10483
0 10485 5 1 1 10484
0 10486 7 1 2 69733 75764
0 10487 5 1 1 10486
0 10488 7 1 2 83605 10487
0 10489 5 1 1 10488
0 10490 7 1 2 70394 10489
0 10491 5 1 1 10490
0 10492 7 3 2 63993 77268
0 10493 5 2 1 83673
0 10494 7 1 2 70671 83674
0 10495 5 1 1 10494
0 10496 7 1 2 83606 10495
0 10497 5 1 1 10496
0 10498 7 1 2 59491 10497
0 10499 5 1 1 10498
0 10500 7 1 2 10491 10499
0 10501 5 1 1 10500
0 10502 7 1 2 82867 10501
0 10503 5 1 1 10502
0 10504 7 1 2 10485 10503
0 10505 7 1 2 10456 10504
0 10506 5 1 1 10505
0 10507 7 1 2 69673 10506
0 10508 5 1 1 10507
0 10509 7 1 2 75430 76439
0 10510 5 1 1 10509
0 10511 7 7 2 63167 64988
0 10512 5 4 1 83678
0 10513 7 2 2 71156 70159
0 10514 5 1 1 83689
0 10515 7 1 2 83679 83690
0 10516 5 1 1 10515
0 10517 7 1 2 10510 10516
0 10518 5 1 1 10517
0 10519 7 1 2 61528 10518
0 10520 5 1 1 10519
0 10521 7 2 2 81326 78697
0 10522 5 1 1 83691
0 10523 7 1 2 74235 83692
0 10524 5 1 1 10523
0 10525 7 1 2 10520 10524
0 10526 5 1 1 10525
0 10527 7 2 2 66826 67443
0 10528 7 1 2 71103 83693
0 10529 7 1 2 10526 10528
0 10530 5 1 1 10529
0 10531 7 1 2 10508 10530
0 10532 5 1 1 10531
0 10533 7 1 2 68591 10532
0 10534 5 1 1 10533
0 10535 7 1 2 10431 10534
0 10536 7 1 2 10339 10535
0 10537 5 1 1 10536
0 10538 7 1 2 68338 10537
0 10539 5 1 1 10538
0 10540 7 1 2 61906 81809
0 10541 5 1 1 10540
0 10542 7 1 2 9924 10541
0 10543 5 1 1 10542
0 10544 7 1 2 72521 10543
0 10545 5 1 1 10544
0 10546 7 1 2 58226 77611
0 10547 5 1 1 10546
0 10548 7 1 2 79711 10547
0 10549 7 1 2 72371 10548
0 10550 5 1 1 10549
0 10551 7 1 2 75650 10550
0 10552 5 1 1 10551
0 10553 7 1 2 10545 10552
0 10554 5 1 1 10553
0 10555 7 1 2 60814 10554
0 10556 5 1 1 10555
0 10557 7 1 2 75705 8704
0 10558 5 1 1 10557
0 10559 7 1 2 68592 10558
0 10560 5 1 1 10559
0 10561 7 1 2 76009 10560
0 10562 5 1 1 10561
0 10563 7 1 2 67279 10562
0 10564 5 1 1 10563
0 10565 7 3 2 57651 74825
0 10566 7 1 2 61907 75693
0 10567 7 1 2 83695 10566
0 10568 5 1 1 10567
0 10569 7 1 2 82815 10568
0 10570 5 1 1 10569
0 10571 7 1 2 68593 10570
0 10572 5 1 1 10571
0 10573 7 1 2 76020 10572
0 10574 7 1 2 10564 10573
0 10575 5 1 1 10574
0 10576 7 1 2 65201 10575
0 10577 5 1 1 10576
0 10578 7 1 2 67993 75987
0 10579 5 1 1 10578
0 10580 7 1 2 64216 10579
0 10581 7 1 2 10577 10580
0 10582 5 1 1 10581
0 10583 7 1 2 63994 75672
0 10584 5 1 1 10583
0 10585 7 1 2 62328 10584
0 10586 7 1 2 82670 10585
0 10587 5 1 1 10586
0 10588 7 1 2 59492 81988
0 10589 7 1 2 10587 10588
0 10590 5 1 1 10589
0 10591 7 1 2 65490 10590
0 10592 7 1 2 10582 10591
0 10593 5 1 1 10592
0 10594 7 1 2 10556 10593
0 10595 5 1 1 10594
0 10596 7 1 2 69674 10595
0 10597 5 1 1 10596
0 10598 7 2 2 69575 75765
0 10599 7 2 2 70160 73399
0 10600 5 1 1 83700
0 10601 7 2 2 73855 69772
0 10602 7 1 2 64989 73347
0 10603 7 1 2 83702 10602
0 10604 7 1 2 83701 10603
0 10605 7 1 2 83698 10604
0 10606 5 1 1 10605
0 10607 7 1 2 10597 10606
0 10608 5 1 1 10607
0 10609 7 1 2 82893 10608
0 10610 5 1 1 10609
0 10611 7 1 2 59757 10610
0 10612 7 1 2 10539 10611
0 10613 7 1 2 10213 10612
0 10614 5 1 1 10613
0 10615 7 1 2 9340 10614
0 10616 5 1 1 10615
0 10617 7 2 2 64990 77207
0 10618 7 1 2 77378 81810
0 10619 7 1 2 83704 10618
0 10620 5 2 1 10619
0 10621 7 1 2 73205 74424
0 10622 5 1 1 10621
0 10623 7 2 2 74771 82178
0 10624 7 1 2 65491 83708
0 10625 5 1 1 10624
0 10626 7 1 2 10622 10625
0 10627 5 1 1 10626
0 10628 7 1 2 64991 10627
0 10629 5 1 1 10628
0 10630 7 1 2 74447 10629
0 10631 5 2 1 10630
0 10632 7 1 2 64474 83710
0 10633 5 1 1 10632
0 10634 7 1 2 83706 10633
0 10635 5 1 1 10634
0 10636 7 1 2 59296 10635
0 10637 5 1 1 10636
0 10638 7 2 2 74826 74749
0 10639 5 1 1 83712
0 10640 7 1 2 64475 70363
0 10641 7 1 2 83713 10640
0 10642 5 1 1 10641
0 10643 7 1 2 10637 10642
0 10644 5 1 1 10643
0 10645 7 1 2 68594 10644
0 10646 5 1 1 10645
0 10647 7 1 2 77379 81913
0 10648 7 1 2 83632 10647
0 10649 7 1 2 75864 10648
0 10650 5 2 1 10649
0 10651 7 2 2 57652 69872
0 10652 5 3 1 83716
0 10653 7 1 2 78141 83718
0 10654 5 1 1 10653
0 10655 7 1 2 68754 10654
0 10656 5 1 1 10655
0 10657 7 1 2 76280 10656
0 10658 5 1 1 10657
0 10659 7 1 2 74406 10658
0 10660 5 1 1 10659
0 10661 7 4 2 60280 67724
0 10662 5 4 1 83721
0 10663 7 1 2 79514 83725
0 10664 7 1 2 74270 10663
0 10665 5 1 1 10664
0 10666 7 1 2 10660 10665
0 10667 5 1 1 10666
0 10668 7 1 2 65202 10667
0 10669 5 1 1 10668
0 10670 7 1 2 72273 74271
0 10671 5 1 1 10670
0 10672 7 1 2 68755 83709
0 10673 5 1 1 10672
0 10674 7 1 2 10671 10673
0 10675 5 1 1 10674
0 10676 7 1 2 65492 10675
0 10677 5 1 1 10676
0 10678 7 1 2 10669 10677
0 10679 5 2 1 10678
0 10680 7 1 2 64476 83729
0 10681 5 1 1 10680
0 10682 7 1 2 83714 10681
0 10683 5 1 1 10682
0 10684 7 1 2 59297 10683
0 10685 5 1 1 10684
0 10686 7 1 2 10646 10685
0 10687 5 1 1 10686
0 10688 7 1 2 57956 10687
0 10689 5 1 1 10688
0 10690 7 2 2 75848 71638
0 10691 5 2 1 83731
0 10692 7 2 2 83726 83732
0 10693 5 1 1 83735
0 10694 7 1 2 57374 83736
0 10695 5 1 1 10694
0 10696 7 1 2 10695 82080
0 10697 5 2 1 10696
0 10698 7 2 2 65493 67460
0 10699 7 1 2 59983 83739
0 10700 7 2 2 83737 10699
0 10701 7 1 2 67280 79550
0 10702 7 1 2 83741 10701
0 10703 5 1 1 10702
0 10704 7 1 2 64477 70041
0 10705 7 1 2 74445 10704
0 10706 5 1 1 10705
0 10707 7 1 2 10703 10706
0 10708 7 1 2 10689 10707
0 10709 5 1 1 10708
0 10710 7 1 2 71157 10709
0 10711 5 1 1 10710
0 10712 7 1 2 75092 83333
0 10713 5 1 1 10712
0 10714 7 1 2 60518 74272
0 10715 5 1 1 10714
0 10716 7 1 2 10713 10715
0 10717 5 1 1 10716
0 10718 7 1 2 71158 10717
0 10719 5 1 1 10718
0 10720 7 1 2 75319 83218
0 10721 5 1 1 10720
0 10722 7 1 2 82745 83594
0 10723 5 1 1 10722
0 10724 7 1 2 68339 10723
0 10725 5 1 1 10724
0 10726 7 1 2 83499 10725
0 10727 7 1 2 10721 10726
0 10728 5 1 1 10727
0 10729 7 1 2 58227 10728
0 10730 5 1 1 10729
0 10731 7 1 2 67281 83219
0 10732 5 1 1 10731
0 10733 7 1 2 59298 83224
0 10734 5 1 1 10733
0 10735 7 2 2 10732 10734
0 10736 7 3 2 68340 83508
0 10737 5 1 1 83745
0 10738 7 1 2 83743 10737
0 10739 5 1 1 10738
0 10740 7 1 2 59493 10739
0 10741 5 1 1 10740
0 10742 7 3 2 58962 60519
0 10743 7 1 2 83748 69873
0 10744 5 2 1 10743
0 10745 7 2 2 74362 75251
0 10746 5 1 1 83753
0 10747 7 1 2 71869 83754
0 10748 5 1 1 10747
0 10749 7 1 2 83751 10748
0 10750 5 2 1 10749
0 10751 7 1 2 57653 83755
0 10752 5 1 1 10751
0 10753 7 2 2 70768 81689
0 10754 5 1 1 83757
0 10755 7 2 2 10752 10754
0 10756 5 1 1 83759
0 10757 7 1 2 10741 83760
0 10758 5 1 1 10757
0 10759 7 1 2 72522 10758
0 10760 5 1 1 10759
0 10761 7 1 2 10730 10760
0 10762 5 1 1 10761
0 10763 7 1 2 74273 10762
0 10764 5 1 1 10763
0 10765 7 1 2 10719 10764
0 10766 5 1 1 10765
0 10767 7 1 2 60815 10766
0 10768 5 1 1 10767
0 10769 7 1 2 67815 79750
0 10770 5 3 1 10769
0 10771 7 1 2 74092 83761
0 10772 5 2 1 10771
0 10773 7 1 2 59494 75106
0 10774 5 1 1 10773
0 10775 7 1 2 83764 10774
0 10776 5 1 1 10775
0 10777 7 1 2 74274 10776
0 10778 5 1 1 10777
0 10779 7 1 2 57957 79130
0 10780 5 1 1 10779
0 10781 7 1 2 4546 81626
0 10782 5 2 1 10781
0 10783 7 1 2 57958 83766
0 10784 5 1 1 10783
0 10785 7 1 2 73895 75168
0 10786 5 1 1 10785
0 10787 7 1 2 10784 10786
0 10788 5 1 1 10787
0 10789 7 1 2 57654 10788
0 10790 5 1 1 10789
0 10791 7 1 2 10780 10790
0 10792 5 1 1 10791
0 10793 7 2 2 64217 10792
0 10794 5 1 1 83768
0 10795 7 1 2 74407 83769
0 10796 5 1 1 10795
0 10797 7 1 2 10778 10796
0 10798 5 1 1 10797
0 10799 7 1 2 58228 10798
0 10800 5 1 1 10799
0 10801 7 1 2 68070 83140
0 10802 5 1 1 10801
0 10803 7 3 2 67282 10802
0 10804 5 1 1 83770
0 10805 7 1 2 74325 83771
0 10806 5 1 1 10805
0 10807 7 3 2 68595 83308
0 10808 5 1 1 83773
0 10809 7 1 2 71623 83774
0 10810 5 1 1 10809
0 10811 7 1 2 58229 83468
0 10812 5 6 1 10811
0 10813 7 1 2 68429 83776
0 10814 7 1 2 10810 10813
0 10815 7 1 2 10806 10814
0 10816 5 1 1 10815
0 10817 7 1 2 74275 10816
0 10818 5 1 1 10817
0 10819 7 1 2 57959 80724
0 10820 5 1 1 10819
0 10821 7 1 2 70066 10820
0 10822 5 2 1 10821
0 10823 7 1 2 83615 67515
0 10824 7 1 2 83782 10823
0 10825 5 1 1 10824
0 10826 7 1 2 64218 10825
0 10827 7 1 2 10818 10826
0 10828 5 1 1 10827
0 10829 7 2 2 71870 76502
0 10830 5 3 1 83784
0 10831 7 1 2 62329 83786
0 10832 5 1 1 10831
0 10833 7 2 2 81842 10832
0 10834 5 4 1 83789
0 10835 7 2 2 83790 83232
0 10836 5 1 1 83795
0 10837 7 2 2 59299 10836
0 10838 5 1 1 83797
0 10839 7 1 2 60281 83469
0 10840 5 1 1 10839
0 10841 7 1 2 70724 80503
0 10842 5 1 1 10841
0 10843 7 2 2 10840 10842
0 10844 5 1 1 83799
0 10845 7 1 2 83800 83273
0 10846 5 1 1 10845
0 10847 7 1 2 63995 10846
0 10848 5 2 1 10847
0 10849 7 1 2 10838 83801
0 10850 5 1 1 10849
0 10851 7 1 2 74276 10850
0 10852 5 1 1 10851
0 10853 7 1 2 62330 78055
0 10854 5 3 1 10853
0 10855 7 1 2 83321 83803
0 10856 5 1 1 10855
0 10857 7 1 2 58230 10856
0 10858 5 1 1 10857
0 10859 7 2 2 65203 83183
0 10860 5 1 1 83806
0 10861 7 1 2 58231 67561
0 10862 5 1 1 10861
0 10863 7 1 2 10860 10862
0 10864 5 1 1 10863
0 10865 7 1 2 70021 10864
0 10866 5 1 1 10865
0 10867 7 1 2 62331 70037
0 10868 7 1 2 83807 10867
0 10869 5 1 1 10868
0 10870 7 1 2 10866 10869
0 10871 7 1 2 10858 10870
0 10872 5 2 1 10871
0 10873 7 1 2 74408 83808
0 10874 5 1 1 10873
0 10875 7 1 2 59495 10874
0 10876 7 1 2 10852 10875
0 10877 5 1 1 10876
0 10878 7 1 2 65494 10877
0 10879 7 1 2 10828 10878
0 10880 5 1 1 10879
0 10881 7 1 2 62332 69089
0 10882 5 2 1 10881
0 10883 7 6 2 74033 83810
0 10884 5 2 1 83812
0 10885 7 3 2 57655 70868
0 10886 5 2 1 83820
0 10887 7 1 2 83818 83823
0 10888 5 1 1 10887
0 10889 7 1 2 74277 10888
0 10890 5 1 1 10889
0 10891 7 1 2 57656 74778
0 10892 5 1 1 10891
0 10893 7 1 2 10639 10892
0 10894 5 1 1 10893
0 10895 7 1 2 70869 10894
0 10896 5 1 1 10895
0 10897 7 1 2 10890 10896
0 10898 5 1 1 10897
0 10899 7 1 2 69310 73400
0 10900 7 1 2 10898 10899
0 10901 5 1 1 10900
0 10902 7 1 2 10880 10901
0 10903 7 1 2 10800 10902
0 10904 7 1 2 10768 10903
0 10905 5 1 1 10904
0 10906 7 1 2 59758 10905
0 10907 5 1 1 10906
0 10908 7 1 2 10711 10907
0 10909 5 1 1 10908
0 10910 7 1 2 58420 10909
0 10911 5 1 1 10910
0 10912 7 6 2 59759 71159
0 10913 7 1 2 63168 83711
0 10914 5 1 1 10913
0 10915 7 1 2 10914 83707
0 10916 5 1 1 10915
0 10917 7 1 2 59300 10916
0 10918 5 1 1 10917
0 10919 7 1 2 74206 67461
0 10920 7 1 2 81811 10919
0 10921 5 1 1 10920
0 10922 7 1 2 10918 10921
0 10923 5 1 1 10922
0 10924 7 1 2 68596 10923
0 10925 5 1 1 10924
0 10926 7 1 2 63169 83730
0 10927 5 1 1 10926
0 10928 7 1 2 10927 83715
0 10929 5 1 1 10928
0 10930 7 1 2 59301 10929
0 10931 5 1 1 10930
0 10932 7 1 2 10925 10931
0 10933 5 1 1 10932
0 10934 7 1 2 57960 10933
0 10935 5 1 1 10934
0 10936 7 1 2 74207 74278
0 10937 7 1 2 70042 10936
0 10938 5 1 1 10937
0 10939 7 1 2 67283 82797
0 10940 7 1 2 83742 10939
0 10941 5 1 1 10940
0 10942 7 1 2 10938 10941
0 10943 7 1 2 10935 10942
0 10944 5 1 1 10943
0 10945 7 1 2 83825 10944
0 10946 5 1 1 10945
0 10947 7 1 2 61529 10946
0 10948 7 1 2 10911 10947
0 10949 5 1 1 10948
0 10950 7 1 2 57961 76902
0 10951 5 3 1 10950
0 10952 7 1 2 70707 83831
0 10953 7 1 2 80373 10952
0 10954 5 1 1 10953
0 10955 7 1 2 78566 10954
0 10956 5 1 1 10955
0 10957 7 1 2 62333 10956
0 10958 5 1 1 10957
0 10959 7 1 2 58232 83578
0 10960 5 1 1 10959
0 10961 7 1 2 62618 10960
0 10962 5 1 1 10961
0 10963 7 1 2 10958 10962
0 10964 5 1 1 10963
0 10965 7 1 2 60816 10964
0 10966 5 1 1 10965
0 10967 7 2 2 73822 70982
0 10968 7 1 2 62900 83834
0 10969 5 1 1 10968
0 10970 7 1 2 10966 10969
0 10971 5 1 1 10970
0 10972 7 1 2 64219 10971
0 10973 5 1 1 10972
0 10974 7 1 2 64220 77061
0 10975 5 1 1 10974
0 10976 7 1 2 59496 79367
0 10977 5 5 1 10976
0 10978 7 2 2 68477 83836
0 10979 5 1 1 83841
0 10980 7 1 2 63847 83842
0 10981 5 1 1 10980
0 10982 7 1 2 10975 10981
0 10983 5 1 1 10982
0 10984 7 1 2 62334 10983
0 10985 5 1 1 10984
0 10986 7 3 2 60520 70038
0 10987 5 3 1 83843
0 10988 7 1 2 79484 83844
0 10989 5 1 1 10988
0 10990 7 1 2 10985 10989
0 10991 5 1 1 10990
0 10992 7 1 2 76166 10991
0 10993 5 1 1 10992
0 10994 7 1 2 62335 77062
0 10995 5 2 1 10994
0 10996 7 1 2 65495 83846
0 10997 5 1 1 10996
0 10998 7 1 2 60282 10997
0 10999 5 1 1 10998
0 11000 7 1 2 83849 10999
0 11001 5 1 1 11000
0 11002 7 1 2 63996 11001
0 11003 5 1 1 11002
0 11004 7 2 2 62336 69383
0 11005 7 1 2 60817 83851
0 11006 5 1 1 11005
0 11007 7 1 2 11003 11006
0 11008 5 1 1 11007
0 11009 7 1 2 77415 11008
0 11010 5 1 1 11009
0 11011 7 1 2 10993 11010
0 11012 7 1 2 10973 11011
0 11013 5 1 1 11012
0 11014 7 1 2 58421 11013
0 11015 5 1 1 11014
0 11016 7 3 2 62901 72470
0 11017 7 1 2 69813 69917
0 11018 7 1 2 77552 11017
0 11019 7 1 2 83853 11018
0 11020 5 1 1 11019
0 11021 7 1 2 11015 11020
0 11022 5 1 1 11021
0 11023 7 1 2 59760 11022
0 11024 5 1 1 11023
0 11025 7 1 2 74082 74199
0 11026 5 1 1 11025
0 11027 7 1 2 59101 11026
0 11028 5 1 1 11027
0 11029 7 1 2 11028 81210
0 11030 5 1 1 11029
0 11031 7 1 2 57657 11030
0 11032 5 1 1 11031
0 11033 7 1 2 81208 11032
0 11034 5 1 1 11033
0 11035 7 1 2 68756 11034
0 11036 5 1 1 11035
0 11037 7 1 2 81206 11036
0 11038 5 1 1 11037
0 11039 7 1 2 57962 11038
0 11040 5 1 1 11039
0 11041 7 1 2 11040 81204
0 11042 5 1 1 11041
0 11043 7 1 2 64992 11042
0 11044 5 1 1 11043
0 11045 7 1 2 81242 11044
0 11046 5 2 1 11045
0 11047 7 1 2 83856 79637
0 11048 5 1 1 11047
0 11049 7 1 2 78816 83497
0 11050 5 1 1 11049
0 11051 7 1 2 60283 11050
0 11052 5 1 1 11051
0 11053 7 1 2 67843 75236
0 11054 5 1 1 11053
0 11055 7 1 2 83437 76778
0 11056 5 1 1 11055
0 11057 7 1 2 68341 11056
0 11058 5 1 1 11057
0 11059 7 1 2 83116 11058
0 11060 7 1 2 11054 11059
0 11061 7 1 2 11052 11060
0 11062 5 1 1 11061
0 11063 7 1 2 60818 11062
0 11064 5 1 1 11063
0 11065 7 2 2 11064 83495
0 11066 5 1 1 83858
0 11067 7 1 2 59497 11066
0 11068 5 1 1 11067
0 11069 7 2 2 65204 76806
0 11070 5 3 1 83860
0 11071 7 1 2 62902 83862
0 11072 5 1 1 11071
0 11073 7 1 2 59302 11072
0 11074 5 1 1 11073
0 11075 7 4 2 76078 71641
0 11076 5 1 1 83865
0 11077 7 3 2 67725 83866
0 11078 5 1 1 83869
0 11079 7 1 2 57375 81580
0 11080 5 1 1 11079
0 11081 7 4 2 83870 11080
0 11082 5 1 1 83872
0 11083 7 1 2 74363 83873
0 11084 7 1 2 11074 11083
0 11085 5 1 1 11084
0 11086 7 1 2 70395 11085
0 11087 5 1 1 11086
0 11088 7 1 2 67284 80910
0 11089 5 2 1 11088
0 11090 7 1 2 64221 83876
0 11091 7 1 2 11087 11090
0 11092 5 1 1 11091
0 11093 7 1 2 74449 80355
0 11094 5 1 1 11093
0 11095 7 1 2 83186 11094
0 11096 5 1 1 11095
0 11097 7 1 2 62337 11096
0 11098 5 1 1 11097
0 11099 7 2 2 71015 11098
0 11100 5 1 1 83878
0 11101 7 1 2 59498 83879
0 11102 5 1 1 11101
0 11103 7 1 2 65496 11102
0 11104 7 1 2 11092 11103
0 11105 5 1 1 11104
0 11106 7 1 2 83123 69773
0 11107 5 1 1 11106
0 11108 7 1 2 10377 11107
0 11109 5 1 1 11108
0 11110 7 1 2 57963 11109
0 11111 5 1 1 11110
0 11112 7 2 2 68986 74093
0 11113 5 1 1 83880
0 11114 7 1 2 83531 11113
0 11115 5 1 1 11114
0 11116 7 1 2 58233 11115
0 11117 5 1 1 11116
0 11118 7 1 2 11111 11117
0 11119 5 1 1 11118
0 11120 7 1 2 57376 11119
0 11121 5 1 1 11120
0 11122 7 2 2 67285 81615
0 11123 5 2 1 83882
0 11124 7 1 2 83287 83883
0 11125 5 1 1 11124
0 11126 7 1 2 11121 11125
0 11127 5 1 1 11126
0 11128 7 1 2 68342 11127
0 11129 5 1 1 11128
0 11130 7 1 2 70396 67650
0 11131 5 2 1 11130
0 11132 7 1 2 71593 83886
0 11133 5 1 1 11132
0 11134 7 2 2 60819 75237
0 11135 5 1 1 83888
0 11136 7 1 2 77569 11135
0 11137 5 1 1 11136
0 11138 7 1 2 11133 11137
0 11139 5 1 1 11138
0 11140 7 2 2 57964 74364
0 11141 5 2 1 83890
0 11142 7 3 2 67726 72401
0 11143 5 2 1 83894
0 11144 7 1 2 60284 83897
0 11145 5 1 1 11144
0 11146 7 1 2 83892 11145
0 11147 7 1 2 75231 11146
0 11148 5 1 1 11147
0 11149 7 1 2 59303 11148
0 11150 5 1 1 11149
0 11151 7 1 2 76783 11150
0 11152 5 1 1 11151
0 11153 7 1 2 69712 11152
0 11154 5 1 1 11153
0 11155 7 1 2 11139 11154
0 11156 7 1 2 11129 11155
0 11157 7 1 2 11105 11156
0 11158 7 1 2 11068 11157
0 11159 5 1 1 11158
0 11160 7 1 2 76729 11159
0 11161 5 1 1 11160
0 11162 7 1 2 11048 11161
0 11163 7 1 2 11024 11162
0 11164 5 1 1 11163
0 11165 7 1 2 74279 11164
0 11166 5 1 1 11165
0 11167 7 1 2 67727 83453
0 11168 5 1 1 11167
0 11169 7 1 2 75054 11168
0 11170 5 2 1 11169
0 11171 7 1 2 77606 83899
0 11172 5 1 1 11171
0 11173 7 1 2 69754 78786
0 11174 5 1 1 11173
0 11175 7 1 2 63997 11174
0 11176 5 1 1 11175
0 11177 7 1 2 60820 74094
0 11178 5 1 1 11177
0 11179 7 1 2 11176 11178
0 11180 5 1 1 11179
0 11181 7 1 2 70617 11180
0 11182 5 1 1 11181
0 11183 7 1 2 77553 77749
0 11184 5 1 1 11183
0 11185 7 1 2 11182 11184
0 11186 5 1 1 11185
0 11187 7 1 2 63848 11186
0 11188 5 1 1 11187
0 11189 7 1 2 73584 74833
0 11190 5 1 1 11189
0 11191 7 1 2 77612 11190
0 11192 5 1 1 11191
0 11193 7 1 2 79537 11192
0 11194 5 1 1 11193
0 11195 7 1 2 65497 77908
0 11196 5 1 1 11195
0 11197 7 1 2 11194 11196
0 11198 7 1 2 11188 11197
0 11199 5 1 1 11198
0 11200 7 1 2 60285 11199
0 11201 5 1 1 11200
0 11202 7 1 2 11172 11201
0 11203 5 1 1 11202
0 11204 7 1 2 62903 11203
0 11205 5 1 1 11204
0 11206 7 6 2 62164 70894
0 11207 5 3 1 83901
0 11208 7 4 2 63998 79485
0 11209 7 1 2 83902 83910
0 11210 7 1 2 79524 11209
0 11211 5 2 1 11210
0 11212 7 1 2 11205 83914
0 11213 5 1 1 11212
0 11214 7 1 2 76615 11213
0 11215 5 1 1 11214
0 11216 7 1 2 60286 82727
0 11217 5 1 1 11216
0 11218 7 1 2 8591 11217
0 11219 5 1 1 11218
0 11220 7 1 2 71160 11219
0 11221 5 1 1 11220
0 11222 7 5 2 64222 67994
0 11223 5 1 1 83916
0 11224 7 1 2 67651 83917
0 11225 7 1 2 83220 11224
0 11226 5 1 1 11225
0 11227 7 1 2 11221 11226
0 11228 5 1 1 11227
0 11229 7 1 2 65498 11228
0 11230 5 1 1 11229
0 11231 7 6 2 58234 58963
0 11232 5 2 1 83921
0 11233 7 1 2 74178 83922
0 11234 5 1 1 11233
0 11235 7 1 2 70161 72680
0 11236 7 1 2 75281 11235
0 11237 5 1 1 11236
0 11238 7 1 2 11234 11237
0 11239 5 1 1 11238
0 11240 7 1 2 68343 11239
0 11241 5 1 1 11240
0 11242 7 1 2 83403 75138
0 11243 5 1 1 11242
0 11244 7 1 2 11241 11243
0 11245 5 1 1 11244
0 11246 7 1 2 77518 11245
0 11247 5 1 1 11246
0 11248 7 3 2 62338 69783
0 11249 5 5 1 83929
0 11250 7 2 2 68478 83722
0 11251 5 3 1 83937
0 11252 7 1 2 83932 83939
0 11253 5 1 1 11252
0 11254 7 1 2 71096 11253
0 11255 5 1 1 11254
0 11256 7 1 2 79591 83719
0 11257 5 1 1 11256
0 11258 7 1 2 11255 11257
0 11259 5 1 1 11258
0 11260 7 1 2 59499 11259
0 11261 5 1 1 11260
0 11262 7 1 2 11247 11261
0 11263 5 1 1 11262
0 11264 7 1 2 65205 11263
0 11265 5 1 1 11264
0 11266 7 1 2 60821 78927
0 11267 7 1 2 76532 11266
0 11268 7 1 2 77130 11267
0 11269 5 1 1 11268
0 11270 7 1 2 11265 11269
0 11271 7 1 2 11230 11270
0 11272 5 1 1 11271
0 11273 7 1 2 77848 11272
0 11274 5 1 1 11273
0 11275 7 6 2 57965 70162
0 11276 5 21 1 83942
0 11277 7 2 2 83943 79638
0 11278 7 1 2 63170 83969
0 11279 7 1 2 80725 11278
0 11280 5 1 1 11279
0 11281 7 1 2 11274 11280
0 11282 7 1 2 11215 11281
0 11283 5 1 1 11282
0 11284 7 1 2 74409 11283
0 11285 5 1 1 11284
0 11286 7 1 2 66144 11285
0 11287 7 1 2 11166 11286
0 11288 5 1 1 11287
0 11289 7 1 2 70483 11288
0 11290 7 1 2 10949 11289
0 11291 5 1 1 11290
0 11292 7 7 2 60822 67995
0 11293 5 1 1 83971
0 11294 7 1 2 67286 75209
0 11295 5 1 1 11294
0 11296 7 1 2 11293 11295
0 11297 5 1 1 11296
0 11298 7 1 2 75651 11297
0 11299 5 1 1 11298
0 11300 7 2 2 77441 83616
0 11301 7 2 2 60287 81895
0 11302 7 1 2 83978 83980
0 11303 5 1 1 11302
0 11304 7 1 2 11299 11303
0 11305 5 1 1 11304
0 11306 7 1 2 57658 11305
0 11307 5 1 1 11306
0 11308 7 1 2 64993 83385
0 11309 5 1 1 11308
0 11310 7 1 2 11307 11309
0 11311 5 1 1 11310
0 11312 7 1 2 71871 11311
0 11313 5 1 1 11312
0 11314 7 1 2 6441 83972
0 11315 5 2 1 11314
0 11316 7 2 2 67287 76255
0 11317 5 1 1 83984
0 11318 7 1 2 72043 83985
0 11319 5 1 1 11318
0 11320 7 1 2 83982 11319
0 11321 5 2 1 11320
0 11322 7 1 2 83986 75652
0 11323 5 1 1 11322
0 11324 7 1 2 63475 60521
0 11325 7 1 2 68960 11324
0 11326 7 1 2 81896 11325
0 11327 7 1 2 82703 11326
0 11328 5 1 1 11327
0 11329 7 1 2 11323 11328
0 11330 5 1 1 11329
0 11331 7 1 2 68597 11330
0 11332 5 1 1 11331
0 11333 7 1 2 80324 78681
0 11334 5 1 1 11333
0 11335 7 1 2 83319 11334
0 11336 5 1 1 11335
0 11337 7 1 2 68757 11336
0 11338 5 1 1 11337
0 11339 7 1 2 83973 82762
0 11340 5 1 1 11339
0 11341 7 1 2 3158 75307
0 11342 5 1 1 11341
0 11343 7 1 2 60823 72715
0 11344 5 2 1 11343
0 11345 7 1 2 70769 83988
0 11346 7 1 2 11342 11345
0 11347 5 1 1 11346
0 11348 7 1 2 11340 11347
0 11349 7 1 2 11338 11348
0 11350 5 1 1 11349
0 11351 7 1 2 75653 11350
0 11352 5 1 1 11351
0 11353 7 2 2 57966 73742
0 11354 7 1 2 74904 83990
0 11355 7 1 2 82701 11354
0 11356 5 1 1 11355
0 11357 7 1 2 11352 11356
0 11358 7 1 2 11332 11357
0 11359 7 1 2 11313 11358
0 11360 5 1 1 11359
0 11361 7 1 2 71161 11360
0 11362 5 1 1 11361
0 11363 7 1 2 57377 74809
0 11364 7 1 2 68961 11363
0 11365 7 2 2 58738 71473
0 11366 7 1 2 83363 83992
0 11367 7 1 2 11364 11366
0 11368 7 1 2 83436 11367
0 11369 5 1 1 11368
0 11370 7 1 2 11362 11369
0 11371 5 1 1 11370
0 11372 7 1 2 81247 68684
0 11373 7 1 2 11371 11372
0 11374 5 1 1 11373
0 11375 7 1 2 11291 11374
0 11376 7 1 2 10616 11375
0 11377 5 1 1 11376
0 11378 7 1 2 65805 11377
0 11379 5 1 1 11378
0 11380 7 2 2 82798 81017
0 11381 7 25 2 64478 59984
0 11382 5 1 1 83996
0 11383 7 3 2 83997 67920
0 11384 7 1 2 63849 81008
0 11385 7 1 2 84021 11384
0 11386 7 6 2 62051 82093
0 11387 7 3 2 77977 78239
0 11388 7 1 2 84024 84030
0 11389 7 1 2 11385 11388
0 11390 7 1 2 83994 11389
0 11391 5 1 1 11390
0 11392 7 2 2 62339 74450
0 11393 5 3 1 84033
0 11394 7 2 2 67728 72548
0 11395 5 1 1 84038
0 11396 7 1 2 76903 11395
0 11397 5 1 1 11396
0 11398 7 1 2 78454 11397
0 11399 5 1 1 11398
0 11400 7 1 2 84035 11399
0 11401 5 2 1 11400
0 11402 7 1 2 73109 84040
0 11403 5 1 1 11402
0 11404 7 7 2 60288 68223
0 11405 7 1 2 75139 84042
0 11406 5 1 1 11405
0 11407 7 1 2 11403 11406
0 11408 5 1 1 11407
0 11409 7 1 2 62619 11408
0 11410 5 1 1 11409
0 11411 7 2 2 70921 83480
0 11412 7 2 2 71799 73110
0 11413 5 1 1 84051
0 11414 7 1 2 84049 84052
0 11415 5 1 1 11414
0 11416 7 1 2 11410 11415
0 11417 5 1 1 11416
0 11418 7 1 2 66145 11417
0 11419 5 1 1 11418
0 11420 7 1 2 81650 11419
0 11421 5 1 1 11420
0 11422 7 1 2 59500 11421
0 11423 5 1 1 11422
0 11424 7 1 2 11423 81593
0 11425 5 1 1 11424
0 11426 7 1 2 67039 11425
0 11427 5 1 1 11426
0 11428 7 19 2 61530 71162
0 11429 5 2 1 84053
0 11430 7 1 2 82083 84054
0 11431 5 1 1 11430
0 11432 7 1 2 66146 74326
0 11433 7 1 2 81574 11432
0 11434 5 1 1 11433
0 11435 7 1 2 11431 11434
0 11436 5 1 1 11435
0 11437 7 1 2 57378 11436
0 11438 5 1 1 11437
0 11439 7 1 2 72829 69126
0 11440 7 1 2 83179 11439
0 11441 5 1 1 11440
0 11442 7 1 2 11438 11441
0 11443 5 1 1 11442
0 11444 7 1 2 57967 11443
0 11445 5 1 1 11444
0 11446 7 1 2 77450 84050
0 11447 7 1 2 82077 11446
0 11448 5 1 1 11447
0 11449 7 1 2 11445 11448
0 11450 5 1 1 11449
0 11451 7 1 2 60824 11450
0 11452 5 1 1 11451
0 11453 7 3 2 65206 78846
0 11454 5 12 1 84074
0 11455 7 2 2 72716 84075
0 11456 7 1 2 70687 84089
0 11457 5 1 1 11456
0 11458 7 2 2 82154 75299
0 11459 5 1 1 84091
0 11460 7 1 2 57968 84092
0 11461 5 1 1 11460
0 11462 7 1 2 11457 11461
0 11463 5 1 1 11462
0 11464 7 1 2 76426 82376
0 11465 7 1 2 11463 11464
0 11466 5 1 1 11465
0 11467 7 1 2 11452 11466
0 11468 5 1 1 11467
0 11469 7 1 2 66958 11468
0 11470 5 1 1 11469
0 11471 7 1 2 11427 11470
0 11472 5 1 1 11471
0 11473 7 1 2 72560 11472
0 11474 5 1 1 11473
0 11475 7 3 2 67462 72637
0 11476 5 2 1 84093
0 11477 7 1 2 59102 71106
0 11478 5 1 1 11477
0 11479 7 1 2 84096 11478
0 11480 5 1 1 11479
0 11481 7 1 2 58964 11480
0 11482 5 1 1 11481
0 11483 7 1 2 79113 74365
0 11484 5 1 1 11483
0 11485 7 1 2 71945 11484
0 11486 5 1 1 11485
0 11487 7 1 2 11482 11486
0 11488 5 1 1 11487
0 11489 7 1 2 57379 11488
0 11490 5 1 1 11489
0 11491 7 1 2 80045 71946
0 11492 5 1 1 11491
0 11493 7 1 2 11490 11492
0 11494 5 1 1 11493
0 11495 7 1 2 57659 11494
0 11496 5 1 1 11495
0 11497 7 2 2 62052 77131
0 11498 7 3 2 59103 60109
0 11499 7 1 2 67109 84100
0 11500 7 1 2 84098 11499
0 11501 5 1 1 11500
0 11502 7 1 2 11496 11501
0 11503 5 1 1 11502
0 11504 7 1 2 73162 11503
0 11505 5 1 1 11504
0 11506 7 2 2 70163 71947
0 11507 7 1 2 75290 84103
0 11508 5 1 1 11507
0 11509 7 1 2 11505 11508
0 11510 5 1 1 11509
0 11511 7 1 2 57969 11510
0 11512 5 1 1 11511
0 11513 7 1 2 71072 81646
0 11514 5 1 1 11513
0 11515 7 1 2 73287 82174
0 11516 5 2 1 11515
0 11517 7 1 2 77132 84105
0 11518 5 1 1 11517
0 11519 7 1 2 57660 82176
0 11520 5 1 1 11519
0 11521 7 1 2 71872 82127
0 11522 5 1 1 11521
0 11523 7 1 2 80627 11522
0 11524 7 1 2 11520 11523
0 11525 7 1 2 11518 11524
0 11526 5 1 1 11525
0 11527 7 1 2 82013 11526
0 11528 5 1 1 11527
0 11529 7 1 2 11514 11528
0 11530 5 1 1 11529
0 11531 7 1 2 58235 11530
0 11532 5 1 1 11531
0 11533 7 3 2 59104 77133
0 11534 5 1 1 84107
0 11535 7 1 2 76546 11534
0 11536 5 1 1 11535
0 11537 7 1 2 57661 11536
0 11538 5 1 1 11537
0 11539 7 1 2 79718 11538
0 11540 5 1 1 11539
0 11541 7 1 2 84104 11540
0 11542 5 1 1 11541
0 11543 7 1 2 61531 11542
0 11544 7 1 2 11532 11543
0 11545 7 1 2 11512 11544
0 11546 5 1 1 11545
0 11547 7 2 2 71958 67516
0 11548 7 1 2 84041 84110
0 11549 5 1 1 11548
0 11550 7 1 2 83239 83989
0 11551 5 1 1 11550
0 11552 7 1 2 71948 11551
0 11553 5 1 1 11552
0 11554 7 1 2 11549 11553
0 11555 5 1 1 11554
0 11556 7 1 2 63999 11555
0 11557 5 1 1 11556
0 11558 7 1 2 70285 82014
0 11559 5 1 1 11558
0 11560 7 1 2 63850 75140
0 11561 7 1 2 67545 11560
0 11562 5 1 1 11561
0 11563 7 1 2 11559 11562
0 11564 5 1 1 11563
0 11565 7 1 2 75479 11564
0 11566 5 1 1 11565
0 11567 7 3 2 62904 60110
0 11568 7 1 2 67463 84112
0 11569 7 1 2 82006 11568
0 11570 5 1 1 11569
0 11571 7 1 2 11566 11570
0 11572 7 1 2 11557 11571
0 11573 5 1 1 11572
0 11574 7 1 2 62620 11573
0 11575 5 1 1 11574
0 11576 7 1 2 60289 81318
0 11577 5 1 1 11576
0 11578 7 1 2 78436 11577
0 11579 5 1 1 11578
0 11580 7 1 2 71949 11579
0 11581 5 1 1 11580
0 11582 7 4 2 58236 64789
0 11583 7 1 2 72330 84115
0 11584 7 1 2 79209 11583
0 11585 7 1 2 74241 11584
0 11586 5 1 1 11585
0 11587 7 1 2 11581 11586
0 11588 5 1 1 11587
0 11589 7 1 2 62340 11588
0 11590 5 1 1 11589
0 11591 7 4 2 71800 79994
0 11592 7 1 2 84119 82015
0 11593 5 1 1 11592
0 11594 7 1 2 66147 11593
0 11595 7 1 2 11590 11594
0 11596 7 1 2 11575 11595
0 11597 5 1 1 11596
0 11598 7 1 2 59501 11597
0 11599 7 1 2 11546 11598
0 11600 5 1 1 11599
0 11601 7 1 2 71581 81351
0 11602 5 1 1 11601
0 11603 7 8 2 62905 81327
0 11604 5 3 1 84123
0 11605 7 1 2 69320 84124
0 11606 5 1 1 11605
0 11607 7 1 2 11602 11606
0 11608 5 1 1 11607
0 11609 7 1 2 71073 11608
0 11610 5 1 1 11609
0 11611 7 2 2 60111 82094
0 11612 7 1 2 81522 67586
0 11613 7 1 2 84134 11612
0 11614 5 1 1 11613
0 11615 7 1 2 11610 11614
0 11616 5 1 1 11615
0 11617 7 1 2 57380 11616
0 11618 5 1 1 11617
0 11619 7 1 2 76120 8094
0 11620 5 1 1 11619
0 11621 7 1 2 57970 11620
0 11622 5 1 1 11621
0 11623 7 1 2 68921 82016
0 11624 5 1 1 11623
0 11625 7 1 2 11622 11624
0 11626 5 1 1 11625
0 11627 7 1 2 58965 11626
0 11628 5 1 1 11627
0 11629 7 3 2 64994 67996
0 11630 5 1 1 84136
0 11631 7 1 2 67546 84137
0 11632 5 1 1 11631
0 11633 7 1 2 11628 11632
0 11634 5 1 1 11633
0 11635 7 1 2 81424 11634
0 11636 5 1 1 11635
0 11637 7 1 2 11618 11636
0 11638 5 1 1 11637
0 11639 7 1 2 68344 11638
0 11640 5 1 1 11639
0 11641 7 1 2 67890 81425
0 11642 5 1 1 11641
0 11643 7 1 2 64995 81344
0 11644 5 1 1 11643
0 11645 7 1 2 11642 11644
0 11646 5 1 1 11645
0 11647 7 1 2 71950 11646
0 11648 5 1 1 11647
0 11649 7 2 2 58966 67891
0 11650 5 1 1 84139
0 11651 7 2 2 57381 84140
0 11652 5 1 1 84141
0 11653 7 1 2 64996 84142
0 11654 5 1 1 11653
0 11655 7 1 2 82450 11654
0 11656 5 1 1 11655
0 11657 7 1 2 84116 81124
0 11658 7 1 2 11656 11657
0 11659 5 1 1 11658
0 11660 7 1 2 11648 11659
0 11661 7 1 2 11640 11660
0 11662 5 1 1 11661
0 11663 7 1 2 65207 11662
0 11664 5 1 1 11663
0 11665 7 2 2 71390 71074
0 11666 7 1 2 81465 84143
0 11667 5 2 1 11666
0 11668 7 1 2 70079 67547
0 11669 5 1 1 11668
0 11670 7 1 2 67496 11669
0 11671 5 1 1 11670
0 11672 7 1 2 81361 11671
0 11673 5 1 1 11672
0 11674 7 1 2 84145 11673
0 11675 5 1 1 11674
0 11676 7 1 2 68345 11675
0 11677 5 1 1 11676
0 11678 7 1 2 57382 67493
0 11679 5 1 1 11678
0 11680 7 1 2 76121 11679
0 11681 5 1 1 11680
0 11682 7 1 2 71728 11681
0 11683 5 1 1 11682
0 11684 7 1 2 67548 73743
0 11685 5 1 1 11684
0 11686 7 1 2 68987 71951
0 11687 5 2 1 11686
0 11688 7 1 2 11685 84147
0 11689 7 1 2 11683 11688
0 11690 5 1 1 11689
0 11691 7 3 2 58237 59105
0 11692 7 5 2 57662 84149
0 11693 5 2 1 84152
0 11694 7 1 2 61532 84153
0 11695 7 1 2 11690 11694
0 11696 5 1 1 11695
0 11697 7 1 2 11677 11696
0 11698 5 1 1 11697
0 11699 7 1 2 57971 11698
0 11700 5 1 1 11699
0 11701 7 2 2 58238 72325
0 11702 7 7 2 61533 67464
0 11703 7 1 2 84159 84161
0 11704 5 2 1 11703
0 11705 7 1 2 84146 84168
0 11706 5 1 1 11705
0 11707 7 1 2 78632 11706
0 11708 5 1 1 11707
0 11709 7 15 2 60290 66148
0 11710 7 1 2 84170 84144
0 11711 5 1 1 11710
0 11712 7 1 2 84169 11711
0 11713 5 1 1 11712
0 11714 7 1 2 68758 11713
0 11715 5 1 1 11714
0 11716 7 1 2 11708 11715
0 11717 7 1 2 11700 11716
0 11718 5 1 1 11717
0 11719 7 1 2 67844 11718
0 11720 5 1 1 11719
0 11721 7 1 2 11664 11720
0 11722 5 1 1 11721
0 11723 7 1 2 65499 11722
0 11724 5 1 1 11723
0 11725 7 15 2 64223 60522
0 11726 5 8 1 84185
0 11727 7 2 2 84186 81384
0 11728 7 1 2 84208 71952
0 11729 5 1 1 11728
0 11730 7 1 2 81111 80341
0 11731 7 1 2 83356 11730
0 11732 5 1 1 11731
0 11733 7 1 2 11729 11732
0 11734 5 1 1 11733
0 11735 7 1 2 58239 11734
0 11736 5 1 1 11735
0 11737 7 1 2 62621 76547
0 11738 5 2 1 11737
0 11739 7 1 2 84210 76845
0 11740 5 1 1 11739
0 11741 7 1 2 81481 84076
0 11742 5 1 1 11741
0 11743 7 1 2 11740 11742
0 11744 5 1 1 11743
0 11745 7 1 2 71075 11744
0 11746 5 1 1 11745
0 11747 7 1 2 81946 71953
0 11748 5 1 1 11747
0 11749 7 1 2 11746 11748
0 11750 5 1 1 11749
0 11751 7 1 2 68346 11750
0 11752 5 1 1 11751
0 11753 7 1 2 69216 83146
0 11754 5 1 1 11753
0 11755 7 1 2 78698 76118
0 11756 5 1 1 11755
0 11757 7 1 2 11754 11756
0 11758 5 1 1 11757
0 11759 7 1 2 68598 11758
0 11760 5 1 1 11759
0 11761 7 1 2 74515 71954
0 11762 5 1 1 11761
0 11763 7 1 2 76846 67549
0 11764 5 1 1 11763
0 11765 7 1 2 11762 11764
0 11766 5 1 1 11765
0 11767 7 1 2 68759 11766
0 11768 5 1 1 11767
0 11769 7 1 2 77571 82017
0 11770 5 1 1 11769
0 11771 7 1 2 11768 11770
0 11772 7 1 2 11760 11771
0 11773 5 1 1 11772
0 11774 7 1 2 67845 11773
0 11775 5 1 1 11774
0 11776 7 1 2 69335 81914
0 11777 5 1 1 11776
0 11778 7 4 2 64000 61908
0 11779 7 1 2 69242 84212
0 11780 7 1 2 81957 11779
0 11781 5 1 1 11780
0 11782 7 1 2 11777 11781
0 11783 5 1 1 11782
0 11784 7 1 2 76533 11783
0 11785 5 1 1 11784
0 11786 7 1 2 11775 11785
0 11787 7 1 2 11752 11786
0 11788 5 1 1 11787
0 11789 7 1 2 60825 11788
0 11790 5 1 1 11789
0 11791 7 2 2 74327 67465
0 11792 7 1 2 62906 72326
0 11793 7 1 2 84216 11792
0 11794 5 1 1 11793
0 11795 7 1 2 11790 11794
0 11796 5 1 1 11795
0 11797 7 1 2 81328 11796
0 11798 5 1 1 11797
0 11799 7 1 2 11736 11798
0 11800 7 1 2 11724 11799
0 11801 7 1 2 11600 11800
0 11802 5 1 1 11801
0 11803 7 1 2 58851 11802
0 11804 5 1 1 11803
0 11805 7 1 2 61187 11804
0 11806 7 1 2 11474 11805
0 11807 5 1 1 11806
0 11808 7 8 2 66564 69519
0 11809 7 2 2 77341 79769
0 11810 7 1 2 83852 84226
0 11811 5 1 1 11810
0 11812 7 1 2 71391 79136
0 11813 5 1 1 11812
0 11814 7 1 2 11811 11813
0 11815 5 1 1 11814
0 11816 7 1 2 57972 11815
0 11817 5 1 1 11816
0 11818 7 1 2 62341 77085
0 11819 5 1 1 11818
0 11820 7 1 2 83204 11819
0 11821 5 1 1 11820
0 11822 7 1 2 63851 11821
0 11823 5 1 1 11822
0 11824 7 1 2 62342 83206
0 11825 5 1 1 11824
0 11826 7 2 2 62165 78798
0 11827 5 1 1 84228
0 11828 7 1 2 63755 84229
0 11829 5 1 1 11828
0 11830 7 1 2 11825 11829
0 11831 5 1 1 11830
0 11832 7 1 2 65208 11831
0 11833 5 1 1 11832
0 11834 7 1 2 78799 75300
0 11835 5 1 1 11834
0 11836 7 1 2 11833 11835
0 11837 5 1 1 11836
0 11838 7 1 2 60291 11837
0 11839 5 1 1 11838
0 11840 7 1 2 83216 11839
0 11841 7 1 2 11823 11840
0 11842 5 1 1 11841
0 11843 7 1 2 64001 11842
0 11844 5 1 1 11843
0 11845 7 1 2 83192 11844
0 11846 5 1 1 11845
0 11847 7 1 2 71163 11846
0 11848 5 1 1 11847
0 11849 7 1 2 11817 11848
0 11850 5 1 1 11849
0 11851 7 1 2 84218 11850
0 11852 5 1 1 11851
0 11853 7 1 2 83335 10794
0 11854 5 1 1 11853
0 11855 7 1 2 58240 11854
0 11856 5 1 1 11855
0 11857 7 1 2 59502 83809
0 11858 5 1 1 11857
0 11859 7 1 2 69311 83783
0 11860 5 1 1 11859
0 11861 7 1 2 11858 11860
0 11862 5 1 1 11861
0 11863 7 1 2 65500 11862
0 11864 5 1 1 11863
0 11865 7 1 2 83361 11864
0 11866 7 1 2 11856 11865
0 11867 5 1 1 11866
0 11868 7 1 2 72733 11867
0 11869 5 1 1 11868
0 11870 7 1 2 61534 11869
0 11871 7 1 2 11852 11870
0 11872 5 1 1 11871
0 11873 7 2 2 63852 75020
0 11874 5 2 1 84230
0 11875 7 12 2 62343 60826
0 11876 5 6 1 84234
0 11877 7 1 2 65209 84235
0 11878 5 2 1 11877
0 11879 7 1 2 84232 84252
0 11880 5 1 1 11879
0 11881 7 1 2 68479 11880
0 11882 5 1 1 11881
0 11883 7 1 2 68224 83454
0 11884 5 1 1 11883
0 11885 7 1 2 11882 11884
0 11886 5 1 1 11885
0 11887 7 1 2 64224 11886
0 11888 5 1 1 11887
0 11889 7 1 2 75029 79535
0 11890 5 2 1 11889
0 11891 7 2 2 64225 84254
0 11892 5 1 1 84256
0 11893 7 2 2 65210 69918
0 11894 5 1 1 84258
0 11895 7 1 2 4156 78541
0 11896 5 1 1 11895
0 11897 7 1 2 68480 11896
0 11898 5 1 1 11897
0 11899 7 1 2 11894 11898
0 11900 5 1 1 11899
0 11901 7 1 2 84236 11900
0 11902 5 1 1 11901
0 11903 7 1 2 11892 11902
0 11904 5 1 1 11903
0 11905 7 1 2 62622 11904
0 11906 5 1 1 11905
0 11907 7 1 2 11888 11906
0 11908 5 1 1 11907
0 11909 7 1 2 60292 11908
0 11910 5 1 1 11909
0 11911 7 1 2 57663 84233
0 11912 5 1 1 11911
0 11913 7 1 2 77607 83455
0 11914 7 1 2 11912 11913
0 11915 5 1 1 11914
0 11916 7 1 2 11910 11915
0 11917 5 1 1 11916
0 11918 7 1 2 62907 11917
0 11919 5 1 1 11918
0 11920 7 1 2 83915 11919
0 11921 5 1 1 11920
0 11922 7 1 2 72734 11921
0 11923 5 1 1 11922
0 11924 7 9 2 63756 64226
0 11925 7 1 2 84260 72578
0 11926 7 1 2 81849 11925
0 11927 7 2 2 63597 76788
0 11928 7 1 2 77479 84269
0 11929 7 1 2 11926 11928
0 11930 5 1 1 11929
0 11931 7 1 2 66149 11930
0 11932 7 1 2 11923 11931
0 11933 5 1 1 11932
0 11934 7 1 2 66682 11933
0 11935 7 1 2 11872 11934
0 11936 5 1 1 11935
0 11937 7 4 2 63853 81158
0 11938 5 1 1 84271
0 11939 7 1 2 76895 84272
0 11940 5 1 1 11939
0 11941 7 5 2 60523 71251
0 11942 5 3 1 84275
0 11943 7 1 2 59503 80207
0 11944 5 4 1 11943
0 11945 7 1 2 68481 84283
0 11946 5 1 1 11945
0 11947 7 1 2 84280 11946
0 11948 5 1 1 11947
0 11949 7 1 2 62344 11948
0 11950 5 1 1 11949
0 11951 7 1 2 72784 77903
0 11952 7 1 2 11950 11951
0 11953 5 1 1 11952
0 11954 7 1 2 62623 11953
0 11955 5 1 1 11954
0 11956 7 1 2 11940 11955
0 11957 5 1 1 11956
0 11958 7 1 2 66150 11957
0 11959 5 1 1 11958
0 11960 7 1 2 75865 78263
0 11961 5 2 1 11960
0 11962 7 2 2 76167 73585
0 11963 5 3 1 84289
0 11964 7 1 2 84287 84290
0 11965 5 1 1 11964
0 11966 7 11 2 57383 61535
0 11967 5 1 1 84294
0 11968 7 1 2 58967 84295
0 11969 7 1 2 11965 11968
0 11970 5 1 1 11969
0 11971 7 1 2 11959 11970
0 11972 5 1 1 11971
0 11973 7 1 2 60293 11972
0 11974 5 1 1 11973
0 11975 7 1 2 73756 81352
0 11976 5 2 1 11975
0 11977 7 1 2 64227 82729
0 11978 5 1 1 11977
0 11979 7 1 2 58241 11978
0 11980 5 1 1 11979
0 11981 7 1 2 59504 70016
0 11982 5 2 1 11981
0 11983 7 1 2 66151 84307
0 11984 7 1 2 11980 11983
0 11985 5 1 1 11984
0 11986 7 1 2 84305 11985
0 11987 5 1 1 11986
0 11988 7 1 2 62624 11987
0 11989 5 1 1 11988
0 11990 7 1 2 84131 84306
0 11991 5 1 1 11990
0 11992 7 1 2 62345 11991
0 11993 5 1 1 11992
0 11994 7 10 2 60524 61536
0 11995 7 2 2 71392 67729
0 11996 5 3 1 84319
0 11997 7 1 2 78633 84321
0 11998 7 1 2 75320 11997
0 11999 7 1 2 78264 11998
0 12000 5 1 1 11999
0 12001 7 1 2 58242 72523
0 12002 5 1 1 12001
0 12003 7 1 2 81151 81533
0 12004 5 1 1 12003
0 12005 7 1 2 68347 12004
0 12006 5 1 1 12005
0 12007 7 1 2 12002 12006
0 12008 7 1 2 12000 12007
0 12009 5 1 1 12008
0 12010 7 1 2 84309 12009
0 12011 5 1 1 12010
0 12012 7 1 2 11993 12011
0 12013 7 1 2 11989 12012
0 12014 7 1 2 11974 12013
0 12015 5 1 1 12014
0 12016 7 1 2 60827 12015
0 12017 5 1 1 12016
0 12018 7 1 2 76073 78822
0 12019 5 2 1 12018
0 12020 7 6 2 80511 83267
0 12021 5 3 1 84326
0 12022 7 1 2 67869 84332
0 12023 5 1 1 12022
0 12024 7 1 2 84324 12023
0 12025 5 1 1 12024
0 12026 7 1 2 57973 12025
0 12027 5 1 1 12026
0 12028 7 1 2 76088 72701
0 12029 5 1 1 12028
0 12030 7 1 2 62908 79634
0 12031 5 1 1 12030
0 12032 7 1 2 71631 12031
0 12033 5 1 1 12032
0 12034 7 1 2 12029 12033
0 12035 7 1 2 12027 12034
0 12036 5 1 1 12035
0 12037 7 1 2 65501 12036
0 12038 5 1 1 12037
0 12039 7 7 2 57664 70770
0 12040 5 12 1 84335
0 12041 7 1 2 65211 78634
0 12042 5 2 1 12041
0 12043 7 1 2 60828 84354
0 12044 5 2 1 12043
0 12045 7 1 2 68348 84356
0 12046 5 2 1 12045
0 12047 7 1 2 84342 84358
0 12048 5 1 1 12047
0 12049 7 1 2 58243 12048
0 12050 5 1 1 12049
0 12051 7 1 2 69963 79754
0 12052 5 1 1 12051
0 12053 7 1 2 78725 12052
0 12054 5 1 1 12053
0 12055 7 1 2 57974 12054
0 12056 5 1 1 12055
0 12057 7 1 2 78978 76298
0 12058 5 1 1 12057
0 12059 7 1 2 81074 12058
0 12060 5 1 1 12059
0 12061 7 1 2 68349 12060
0 12062 5 1 1 12061
0 12063 7 1 2 64228 12062
0 12064 7 1 2 12056 12063
0 12065 7 1 2 12050 12064
0 12066 7 1 2 12038 12065
0 12067 5 1 1 12066
0 12068 7 1 2 59304 9415
0 12069 5 1 1 12068
0 12070 7 1 2 83802 12069
0 12071 5 1 1 12070
0 12072 7 1 2 65502 12071
0 12073 5 1 1 12072
0 12074 7 1 2 58244 75107
0 12075 5 1 1 12074
0 12076 7 1 2 59505 12075
0 12077 7 1 2 12073 12076
0 12078 5 1 1 12077
0 12079 7 1 2 61537 12078
0 12080 7 1 2 12067 12079
0 12081 5 1 1 12080
0 12082 7 1 2 58245 77913
0 12083 5 2 1 12082
0 12084 7 18 2 73586 84360
0 12085 5 3 1 84362
0 12086 7 3 2 69438 78776
0 12087 7 2 2 63757 84383
0 12088 5 1 1 84386
0 12089 7 1 2 62166 84387
0 12090 5 3 1 12089
0 12091 7 3 2 67730 69384
0 12092 5 1 1 84391
0 12093 7 1 2 84388 12092
0 12094 5 1 1 12093
0 12095 7 1 2 84363 12094
0 12096 5 1 1 12095
0 12097 7 1 2 71393 83835
0 12098 5 1 1 12097
0 12099 7 1 2 12096 12098
0 12100 5 1 1 12099
0 12101 7 1 2 66152 12100
0 12102 5 1 1 12101
0 12103 7 1 2 12081 12102
0 12104 7 1 2 12017 12103
0 12105 5 1 1 12104
0 12106 7 1 2 72686 12105
0 12107 5 1 1 12106
0 12108 7 2 2 80139 83481
0 12109 7 1 2 73357 72112
0 12110 7 1 2 84394 12109
0 12111 5 1 1 12110
0 12112 7 1 2 5636 12111
0 12113 5 1 1 12112
0 12114 7 1 2 66565 82377
0 12115 7 1 2 12113 12114
0 12116 5 1 1 12115
0 12117 7 3 2 60294 73587
0 12118 7 1 2 68482 84396
0 12119 5 1 1 12118
0 12120 7 1 2 77613 12119
0 12121 5 1 1 12120
0 12122 7 1 2 66153 81653
0 12123 7 1 2 72692 12122
0 12124 7 1 2 12121 12123
0 12125 5 1 1 12124
0 12126 7 1 2 12116 12125
0 12127 5 1 1 12126
0 12128 7 1 2 70317 72627
0 12129 7 1 2 12127 12128
0 12130 5 1 1 12129
0 12131 7 1 2 65806 12130
0 12132 7 1 2 12107 12131
0 12133 7 1 2 11936 12132
0 12134 5 1 1 12133
0 12135 7 1 2 63171 12134
0 12136 7 1 2 11807 12135
0 12137 5 1 1 12136
0 12138 7 3 2 66154 73083
0 12139 7 3 2 62909 84399
0 12140 5 2 1 84402
0 12141 7 10 2 63854 77462
0 12142 5 2 1 84407
0 12143 7 2 2 60295 77617
0 12144 5 1 1 84419
0 12145 7 3 2 84408 84420
0 12146 5 2 1 84421
0 12147 7 1 2 72331 84422
0 12148 7 1 2 84403 12147
0 12149 5 1 1 12148
0 12150 7 2 2 61538 80726
0 12151 7 2 2 67997 74683
0 12152 5 2 1 84428
0 12153 7 1 2 64229 84429
0 12154 7 1 2 84426 12153
0 12155 5 1 1 12154
0 12156 7 1 2 12149 12155
0 12157 5 1 1 12156
0 12158 7 1 2 58852 81901
0 12159 7 1 2 12157 12158
0 12160 5 1 1 12159
0 12161 7 1 2 12137 12160
0 12162 5 1 1 12161
0 12163 7 1 2 64479 12162
0 12164 5 1 1 12163
0 12165 7 1 2 71873 80621
0 12166 5 1 1 12165
0 12167 7 1 2 81103 12166
0 12168 5 1 1 12167
0 12169 7 1 2 73650 12168
0 12170 5 1 1 12169
0 12171 7 2 2 73163 73651
0 12172 5 3 1 84432
0 12173 7 1 2 70771 72953
0 12174 5 1 1 12173
0 12175 7 1 2 84434 12174
0 12176 5 1 1 12175
0 12177 7 1 2 69187 12176
0 12178 5 1 1 12177
0 12179 7 1 2 12170 12178
0 12180 5 1 1 12179
0 12181 7 1 2 58246 12180
0 12182 5 1 1 12181
0 12183 7 3 2 70349 73951
0 12184 5 1 1 84437
0 12185 7 2 2 69964 79709
0 12186 5 1 1 84440
0 12187 7 1 2 84438 84441
0 12188 5 1 1 12187
0 12189 7 1 2 12182 12188
0 12190 5 1 1 12189
0 12191 7 1 2 77134 12190
0 12192 5 1 1 12191
0 12193 7 1 2 79045 81092
0 12194 5 1 1 12193
0 12195 7 1 2 12192 12194
0 12196 5 2 1 12195
0 12197 7 5 2 61909 76616
0 12198 7 1 2 84442 84444
0 12199 5 1 1 12198
0 12200 7 2 2 72774 75125
0 12201 7 10 2 62346 63172
0 12202 7 2 2 68483 84451
0 12203 7 2 2 84449 84461
0 12204 7 1 2 70286 73686
0 12205 7 1 2 73371 81915
0 12206 7 1 2 12204 12205
0 12207 7 1 2 84463 12206
0 12208 5 1 1 12207
0 12209 7 1 2 12199 12208
0 12210 5 1 1 12209
0 12211 7 1 2 60112 12210
0 12212 5 1 1 12211
0 12213 7 1 2 81066 81299
0 12214 5 1 1 12213
0 12215 7 1 2 80911 73932
0 12216 5 1 1 12215
0 12217 7 1 2 12214 12216
0 12218 5 3 1 12217
0 12219 7 8 2 65807 66566
0 12220 7 2 2 84465 84468
0 12221 7 6 2 58247 72648
0 12222 5 6 1 84478
0 12223 7 2 2 84479 79178
0 12224 7 1 2 84476 84490
0 12225 5 1 1 12224
0 12226 7 1 2 12212 12225
0 12227 5 1 1 12226
0 12228 7 1 2 58853 12227
0 12229 5 1 1 12228
0 12230 7 2 2 71058 71133
0 12231 7 1 2 76617 84492
0 12232 7 1 2 84477 12231
0 12233 5 1 1 12232
0 12234 7 1 2 12229 12233
0 12235 5 1 1 12234
0 12236 7 1 2 66155 12235
0 12237 5 1 1 12236
0 12238 7 2 2 74530 78475
0 12239 5 1 1 84494
0 12240 7 1 2 76797 84495
0 12241 5 2 1 12240
0 12242 7 8 2 65808 68484
0 12243 7 1 2 70945 84498
0 12244 5 2 1 12243
0 12245 7 1 2 80567 84506
0 12246 5 1 1 12245
0 12247 7 1 2 60829 12246
0 12248 5 1 1 12247
0 12249 7 1 2 68485 72471
0 12250 5 2 1 12249
0 12251 7 1 2 77011 84508
0 12252 5 1 1 12251
0 12253 7 1 2 67731 12252
0 12254 5 1 1 12253
0 12255 7 4 2 62347 65212
0 12256 5 2 1 84510
0 12257 7 1 2 76987 84511
0 12258 5 2 1 12257
0 12259 7 4 2 58422 63758
0 12260 7 2 2 72332 84518
0 12261 5 1 1 84522
0 12262 7 1 2 84516 12261
0 12263 7 1 2 12254 12262
0 12264 5 1 1 12263
0 12265 7 1 2 61188 12264
0 12266 5 1 1 12265
0 12267 7 1 2 12248 12266
0 12268 5 1 1 12267
0 12269 7 1 2 64230 12268
0 12270 5 1 1 12269
0 12271 7 1 2 84496 12270
0 12272 5 1 1 12271
0 12273 7 1 2 76878 12272
0 12274 5 1 1 12273
0 12275 7 3 2 77944 72852
0 12276 5 2 1 84524
0 12277 7 4 2 58423 76168
0 12278 7 1 2 84529 74834
0 12279 7 1 2 84525 12278
0 12280 5 1 1 12279
0 12281 7 2 2 12274 12280
0 12282 5 1 1 84533
0 12283 7 3 2 61539 67921
0 12284 7 1 2 81478 84535
0 12285 7 1 2 12282 12284
0 12286 5 1 1 12285
0 12287 7 1 2 12237 12286
0 12288 5 1 1 12287
0 12289 7 1 2 62053 12288
0 12290 5 1 1 12289
0 12291 7 4 2 69520 77289
0 12292 5 1 1 84538
0 12293 7 1 2 12292 72751
0 12294 5 1 1 12293
0 12295 7 1 2 69919 77706
0 12296 7 1 2 12294 12295
0 12297 5 1 1 12296
0 12298 7 2 2 62625 75899
0 12299 5 3 1 84542
0 12300 7 1 2 78251 72735
0 12301 7 1 2 84543 12300
0 12302 5 1 1 12301
0 12303 7 1 2 12297 12302
0 12304 5 1 1 12303
0 12305 7 1 2 70618 12304
0 12306 5 1 1 12305
0 12307 7 1 2 69920 75357
0 12308 5 1 1 12307
0 12309 7 1 2 67288 71040
0 12310 5 1 1 12309
0 12311 7 5 2 60525 68071
0 12312 5 3 1 84547
0 12313 7 1 2 72785 84548
0 12314 7 1 2 12310 12313
0 12315 5 1 1 12314
0 12316 7 1 2 12308 12315
0 12317 5 1 1 12316
0 12318 7 1 2 72736 12317
0 12319 5 1 1 12318
0 12320 7 1 2 12306 12319
0 12321 5 1 1 12320
0 12322 7 1 2 60296 12321
0 12323 5 1 1 12322
0 12324 7 5 2 60526 75126
0 12325 5 2 1 84555
0 12326 7 1 2 64997 84556
0 12327 5 1 1 12326
0 12328 7 1 2 80383 12327
0 12329 5 1 1 12328
0 12330 7 1 2 64002 72737
0 12331 7 1 2 12329 12330
0 12332 5 1 1 12331
0 12333 7 1 2 12323 12332
0 12334 5 1 1 12333
0 12335 7 1 2 60830 12334
0 12336 5 1 1 12335
0 12337 7 1 2 72738 83212
0 12338 7 1 2 81864 12337
0 12339 5 1 1 12338
0 12340 7 1 2 12336 12339
0 12341 5 1 1 12340
0 12342 7 1 2 73038 12341
0 12343 5 1 1 12342
0 12344 7 4 2 62348 67153
0 12345 5 5 1 84562
0 12346 7 10 2 65809 61910
0 12347 7 1 2 72073 84571
0 12348 7 1 2 84563 12347
0 12349 7 3 2 68486 75000
0 12350 5 1 1 84581
0 12351 7 1 2 74461 12350
0 12352 5 1 1 12351
0 12353 7 2 2 62910 70484
0 12354 7 1 2 12352 84584
0 12355 7 1 2 12348 12354
0 12356 5 1 1 12355
0 12357 7 1 2 12343 12356
0 12358 5 1 1 12357
0 12359 7 1 2 61540 12358
0 12360 5 1 1 12359
0 12361 7 13 2 66156 80413
0 12362 5 1 1 84586
0 12363 7 2 2 78240 84587
0 12364 7 1 2 78457 84599
0 12365 5 1 1 12364
0 12366 7 1 2 57975 70997
0 12367 5 1 1 12366
0 12368 7 1 2 74476 12367
0 12369 5 1 1 12368
0 12370 7 1 2 4128 12369
0 12371 5 1 1 12370
0 12372 7 1 2 78131 12371
0 12373 5 1 1 12372
0 12374 7 1 2 71662 83184
0 12375 5 1 1 12374
0 12376 7 4 2 64003 68225
0 12377 7 1 2 57976 84601
0 12378 5 1 1 12377
0 12379 7 1 2 12375 12378
0 12380 5 1 1 12379
0 12381 7 1 2 65810 12380
0 12382 5 1 1 12381
0 12383 7 1 2 12373 12382
0 12384 5 1 1 12383
0 12385 7 1 2 60527 12384
0 12386 5 1 1 12385
0 12387 7 3 2 68760 73606
0 12388 7 1 2 82140 84605
0 12389 5 1 1 12388
0 12390 7 1 2 62626 70681
0 12391 7 1 2 80135 12390
0 12392 5 1 1 12391
0 12393 7 1 2 75050 12392
0 12394 5 1 1 12393
0 12395 7 1 2 70619 12394
0 12396 5 1 1 12395
0 12397 7 1 2 76336 84246
0 12398 7 1 2 84259 12397
0 12399 5 1 1 12398
0 12400 7 1 2 12396 12399
0 12401 5 1 1 12400
0 12402 7 1 2 65811 12401
0 12403 5 1 1 12402
0 12404 7 1 2 12389 12403
0 12405 7 1 2 12386 12404
0 12406 5 1 1 12405
0 12407 7 1 2 60297 12406
0 12408 5 1 1 12407
0 12409 7 1 2 73197 70129
0 12410 5 1 1 12409
0 12411 7 1 2 68226 78543
0 12412 5 1 1 12411
0 12413 7 1 2 12410 12412
0 12414 5 1 1 12413
0 12415 7 1 2 68761 12414
0 12416 5 1 1 12415
0 12417 7 1 2 65812 77601
0 12418 5 1 1 12417
0 12419 7 1 2 12416 12418
0 12420 5 1 1 12419
0 12421 7 1 2 60831 12420
0 12422 5 1 1 12421
0 12423 7 7 2 62627 74477
0 12424 7 1 2 84608 76995
0 12425 5 1 1 12424
0 12426 7 4 2 64998 80395
0 12427 5 1 1 84615
0 12428 7 2 2 67652 84616
0 12429 5 2 1 84619
0 12430 7 1 2 77764 84620
0 12431 5 1 1 12430
0 12432 7 2 2 59305 80396
0 12433 5 1 1 84623
0 12434 7 3 2 60298 73774
0 12435 5 1 1 84625
0 12436 7 1 2 12433 12435
0 12437 5 1 1 12436
0 12438 7 2 2 62349 76988
0 12439 7 1 2 69365 84628
0 12440 7 1 2 12437 12439
0 12441 5 1 1 12440
0 12442 7 1 2 12431 12441
0 12443 5 1 1 12442
0 12444 7 1 2 68599 12443
0 12445 5 1 1 12444
0 12446 7 1 2 12425 12445
0 12447 7 1 2 12422 12446
0 12448 7 1 2 12408 12447
0 12449 5 1 1 12448
0 12450 7 1 2 61541 12449
0 12451 5 1 1 12450
0 12452 7 1 2 12365 12451
0 12453 5 1 1 12452
0 12454 7 1 2 62911 84219
0 12455 7 1 2 12453 12454
0 12456 5 1 1 12455
0 12457 7 1 2 83532 9758
0 12458 5 1 1 12457
0 12459 7 1 2 58248 12458
0 12460 5 1 1 12459
0 12461 7 1 2 74976 68651
0 12462 5 1 1 12461
0 12463 7 1 2 12460 12462
0 12464 5 1 1 12463
0 12465 7 1 2 60528 12464
0 12466 5 1 1 12465
0 12467 7 1 2 83196 83540
0 12468 5 1 1 12467
0 12469 7 1 2 62912 12468
0 12470 5 1 1 12469
0 12471 7 1 2 81942 74179
0 12472 5 1 1 12471
0 12473 7 1 2 12470 12472
0 12474 5 1 1 12473
0 12475 7 1 2 67846 12474
0 12476 5 1 1 12475
0 12477 7 1 2 78823 74561
0 12478 5 1 1 12477
0 12479 7 1 2 57977 78132
0 12480 5 1 1 12479
0 12481 7 1 2 12478 12480
0 12482 5 1 1 12481
0 12483 7 1 2 62913 12482
0 12484 5 1 1 12483
0 12485 7 1 2 79074 78627
0 12486 5 1 1 12485
0 12487 7 1 2 69188 75044
0 12488 7 1 2 83602 12487
0 12489 5 1 1 12488
0 12490 7 1 2 61189 12489
0 12491 7 1 2 12486 12490
0 12492 7 1 2 12484 12491
0 12493 7 1 2 12476 12492
0 12494 7 1 2 12466 12493
0 12495 5 1 1 12494
0 12496 7 1 2 70318 70245
0 12497 5 1 1 12496
0 12498 7 3 2 62628 70198
0 12499 5 7 1 84630
0 12500 7 1 2 84633 75151
0 12501 5 1 1 12500
0 12502 7 1 2 60529 84582
0 12503 7 1 2 12501 12502
0 12504 5 1 1 12503
0 12505 7 1 2 12497 12504
0 12506 5 1 1 12505
0 12507 7 1 2 63855 12506
0 12508 5 1 1 12507
0 12509 7 3 2 63759 78682
0 12510 7 1 2 77393 84640
0 12511 5 1 1 12510
0 12512 7 1 2 12508 12511
0 12513 5 1 1 12512
0 12514 7 1 2 62350 12513
0 12515 5 1 1 12514
0 12516 7 2 2 62629 76989
0 12517 7 1 2 78444 84643
0 12518 5 1 1 12517
0 12519 7 1 2 65813 12518
0 12520 7 1 2 12515 12519
0 12521 5 1 1 12520
0 12522 7 1 2 61542 12521
0 12523 7 1 2 12495 12522
0 12524 5 1 1 12523
0 12525 7 61 2 61190 66157
0 12526 5 4 1 84645
0 12527 7 1 2 76879 84646
0 12528 7 1 2 76942 12527
0 12529 5 1 1 12528
0 12530 7 1 2 12524 12529
0 12531 5 1 1 12530
0 12532 7 1 2 72739 12531
0 12533 5 1 1 12532
0 12534 7 1 2 12456 12533
0 12535 5 1 1 12534
0 12536 7 1 2 64231 12535
0 12537 5 1 1 12536
0 12538 7 1 2 12360 12537
0 12539 5 1 1 12538
0 12540 7 1 2 66683 12539
0 12541 5 1 1 12540
0 12542 7 2 2 65503 71663
0 12543 5 1 1 84710
0 12544 7 1 2 12543 75308
0 12545 7 1 2 3750 12544
0 12546 5 1 1 12545
0 12547 7 1 2 65213 12546
0 12548 5 1 1 12547
0 12549 7 1 2 60832 79766
0 12550 5 1 1 12549
0 12551 7 1 2 12550 71093
0 12552 7 2 2 12548 12551
0 12553 5 1 1 84712
0 12554 7 1 2 61191 84713
0 12555 5 1 1 12554
0 12556 7 1 2 69979 73288
0 12557 5 1 1 12556
0 12558 7 1 2 81831 12557
0 12559 5 1 1 12558
0 12560 7 1 2 60833 12559
0 12561 5 1 1 12560
0 12562 7 1 2 70319 75412
0 12563 5 1 1 12562
0 12564 7 1 2 68487 12563
0 12565 5 1 1 12564
0 12566 7 1 2 58249 81843
0 12567 5 1 1 12566
0 12568 7 1 2 64004 12567
0 12569 5 1 1 12568
0 12570 7 1 2 12565 12569
0 12571 7 1 2 12561 12570
0 12572 5 1 1 12571
0 12573 7 1 2 62630 12572
0 12574 5 1 1 12573
0 12575 7 1 2 77956 80000
0 12576 5 1 1 12575
0 12577 7 1 2 68488 12576
0 12578 5 2 1 12577
0 12579 7 2 2 63856 75392
0 12580 5 1 1 84716
0 12581 7 1 2 60834 84717
0 12582 5 1 1 12581
0 12583 7 1 2 78437 12582
0 12584 7 1 2 84714 12583
0 12585 5 1 1 12584
0 12586 7 1 2 62351 12585
0 12587 5 1 1 12586
0 12588 7 3 2 62914 75099
0 12589 7 1 2 63857 84718
0 12590 5 1 1 12589
0 12591 7 1 2 65814 12590
0 12592 7 1 2 12587 12591
0 12593 7 1 2 12574 12592
0 12594 5 1 1 12593
0 12595 7 1 2 64232 12594
0 12596 7 1 2 12555 12595
0 12597 5 1 1 12596
0 12598 7 5 2 60299 67154
0 12599 5 3 1 84721
0 12600 7 1 2 77957 84726
0 12601 5 1 1 12600
0 12602 7 1 2 68489 12601
0 12603 5 1 1 12602
0 12604 7 1 2 57978 69792
0 12605 5 4 1 12604
0 12606 7 1 2 73111 84729
0 12607 5 1 1 12606
0 12608 7 1 2 12603 12607
0 12609 5 1 1 12608
0 12610 7 1 2 62352 12609
0 12611 5 1 1 12610
0 12612 7 1 2 72074 84722
0 12613 5 1 1 12612
0 12614 7 1 2 12611 12613
0 12615 5 1 1 12614
0 12616 7 1 2 65815 12615
0 12617 5 2 1 12616
0 12618 7 1 2 78533 84509
0 12619 5 2 1 12618
0 12620 7 1 2 67732 84735
0 12621 5 1 1 12620
0 12622 7 2 2 84517 12621
0 12623 7 1 2 59506 83832
0 12624 5 1 1 12623
0 12625 7 1 2 84737 12624
0 12626 5 1 1 12625
0 12627 7 1 2 61192 12626
0 12628 5 1 1 12627
0 12629 7 1 2 84733 12628
0 12630 5 1 1 12629
0 12631 7 1 2 62915 12630
0 12632 5 1 1 12631
0 12633 7 1 2 73060 84507
0 12634 5 1 1 12633
0 12635 7 1 2 60835 12634
0 12636 5 1 1 12635
0 12637 7 7 2 62167 59507
0 12638 7 1 2 76558 84739
0 12639 5 1 1 12638
0 12640 7 1 2 84738 12639
0 12641 5 1 1 12640
0 12642 7 1 2 61193 12641
0 12643 5 1 1 12642
0 12644 7 1 2 12636 12643
0 12645 5 1 1 12644
0 12646 7 1 2 67155 12645
0 12647 5 1 1 12646
0 12648 7 1 2 84497 12647
0 12649 7 1 2 12632 12648
0 12650 7 1 2 12597 12649
0 12651 5 1 1 12650
0 12652 7 1 2 61543 12651
0 12653 5 1 1 12652
0 12654 7 3 2 70287 69784
0 12655 5 2 1 84746
0 12656 7 2 2 84747 82458
0 12657 5 1 1 84751
0 12658 7 1 2 62353 81319
0 12659 5 1 1 12658
0 12660 7 1 2 78438 12659
0 12661 5 1 1 12660
0 12662 7 1 2 75393 12661
0 12663 5 1 1 12662
0 12664 7 1 2 84237 84719
0 12665 5 1 1 12664
0 12666 7 1 2 12663 12665
0 12667 5 1 1 12666
0 12668 7 1 2 62631 12667
0 12669 5 1 1 12668
0 12670 7 1 2 12657 12669
0 12671 5 1 1 12670
0 12672 7 6 2 66158 72853
0 12673 7 1 2 12671 84753
0 12674 5 1 1 12673
0 12675 7 1 2 12653 12674
0 12676 5 1 1 12675
0 12677 7 1 2 72687 12676
0 12678 5 1 1 12677
0 12679 7 1 2 12541 12678
0 12680 5 1 1 12679
0 12681 7 1 2 77849 12680
0 12682 5 1 1 12681
0 12683 7 2 2 74166 73420
0 12684 7 1 2 71582 82649
0 12685 7 1 2 84759 12684
0 12686 7 1 2 80731 12685
0 12687 5 1 1 12686
0 12688 7 1 2 70485 68705
0 12689 7 1 2 81108 12688
0 12690 5 1 1 12689
0 12691 7 3 2 71801 66959
0 12692 5 2 1 84761
0 12693 7 1 2 67082 84764
0 12694 5 1 1 12693
0 12695 7 1 2 63598 12694
0 12696 5 1 1 12695
0 12697 7 3 2 58854 71065
0 12698 5 4 1 84766
0 12699 7 1 2 12696 84769
0 12700 5 1 1 12699
0 12701 7 1 2 60300 78514
0 12702 7 1 2 12700 12701
0 12703 5 1 1 12702
0 12704 7 1 2 12690 12703
0 12705 5 1 1 12704
0 12706 7 20 2 61194 61544
0 12707 5 1 1 84773
0 12708 7 9 2 60836 84774
0 12709 7 3 2 64233 77416
0 12710 7 1 2 84793 84802
0 12711 7 1 2 12705 12710
0 12712 5 1 1 12711
0 12713 7 1 2 12687 12712
0 12714 5 1 1 12713
0 12715 7 1 2 66684 76618
0 12716 7 1 2 12714 12715
0 12717 5 1 1 12716
0 12718 7 1 2 12682 12717
0 12719 7 1 2 12290 12718
0 12720 7 1 2 12164 12719
0 12721 5 1 1 12720
0 12722 7 1 2 66888 12721
0 12723 5 1 1 12722
0 12724 7 1 2 11391 12723
0 12725 7 1 2 11379 12724
0 12726 7 1 2 8561 12725
0 12727 5 1 1 12726
0 12728 7 1 2 61761 12727
0 12729 5 1 1 12728
0 12730 7 1 2 64846 12729
0 12731 7 1 2 6607 12730
0 12732 5 1 1 12731
0 12733 7 2 2 69965 70719
0 12734 5 3 1 84805
0 12735 7 2 2 83877 84807
0 12736 5 1 1 84810
0 12737 7 2 2 65504 80912
0 12738 5 1 1 84812
0 12739 7 2 2 67156 74366
0 12740 5 1 1 84814
0 12741 7 1 2 58250 12740
0 12742 5 1 1 12741
0 12743 7 1 2 12738 12742
0 12744 7 1 2 84811 12743
0 12745 5 1 1 12744
0 12746 7 1 2 78155 12745
0 12747 5 1 1 12746
0 12748 7 2 2 68350 74013
0 12749 5 1 1 84816
0 12750 7 1 2 60530 77437
0 12751 5 1 1 12750
0 12752 7 1 2 12749 12751
0 12753 5 2 1 12752
0 12754 7 1 2 68762 84818
0 12755 5 1 1 12754
0 12756 7 2 2 70772 73997
0 12757 5 1 1 84820
0 12758 7 1 2 12755 12757
0 12759 5 1 1 12758
0 12760 7 1 2 64999 12759
0 12761 5 1 1 12760
0 12762 7 1 2 78168 12761
0 12763 5 1 1 12762
0 12764 7 1 2 70397 12763
0 12765 5 1 1 12764
0 12766 7 2 2 78833 70978
0 12767 5 2 1 84822
0 12768 7 1 2 59508 84824
0 12769 5 1 1 12768
0 12770 7 2 2 68821 79670
0 12771 5 2 1 84826
0 12772 7 1 2 71574 84828
0 12773 5 1 1 12772
0 12774 7 1 2 12769 12773
0 12775 5 1 1 12774
0 12776 7 1 2 58424 84200
0 12777 5 1 1 12776
0 12778 7 1 2 67289 12777
0 12779 7 1 2 12775 12778
0 12780 5 1 1 12779
0 12781 7 2 2 60531 71583
0 12782 5 1 1 84830
0 12783 7 1 2 69312 84831
0 12784 5 1 1 12783
0 12785 7 1 2 62632 84308
0 12786 5 1 1 12785
0 12787 7 1 2 59509 79223
0 12788 5 2 1 12787
0 12789 7 1 2 84157 84832
0 12790 5 1 1 12789
0 12791 7 1 2 12786 12790
0 12792 5 1 1 12791
0 12793 7 1 2 58425 12792
0 12794 5 1 1 12793
0 12795 7 1 2 12784 12794
0 12796 7 1 2 12780 12795
0 12797 7 1 2 12765 12796
0 12798 5 1 1 12797
0 12799 7 1 2 65505 12798
0 12800 5 1 1 12799
0 12801 7 2 2 65000 72274
0 12802 5 2 1 84834
0 12803 7 1 2 84823 84836
0 12804 5 2 1 12803
0 12805 7 1 2 67998 71474
0 12806 5 3 1 12805
0 12807 7 2 2 82918 84840
0 12808 5 3 1 84843
0 12809 7 1 2 69755 72662
0 12810 7 1 2 84845 12809
0 12811 7 1 2 84838 12810
0 12812 5 1 1 12811
0 12813 7 1 2 12800 12812
0 12814 7 1 2 12747 12813
0 12815 7 1 2 78928 12736
0 12816 5 1 1 12815
0 12817 7 1 2 59510 70946
0 12818 5 1 1 12817
0 12819 7 1 2 78549 76770
0 12820 5 2 1 12819
0 12821 7 1 2 84848 3606
0 12822 7 1 2 12818 12821
0 12823 5 1 1 12822
0 12824 7 1 2 58426 12823
0 12825 5 1 1 12824
0 12826 7 1 2 12816 12825
0 12827 5 1 1 12826
0 12828 7 1 2 60837 12827
0 12829 5 1 1 12828
0 12830 7 1 2 57665 80240
0 12831 5 1 1 12830
0 12832 7 1 2 67290 76828
0 12833 5 1 1 12832
0 12834 7 1 2 12831 12833
0 12835 5 1 1 12834
0 12836 7 1 2 68600 12835
0 12837 5 1 1 12836
0 12838 7 2 2 67291 75866
0 12839 5 2 1 84850
0 12840 7 1 2 68072 84852
0 12841 5 3 1 12840
0 12842 7 1 2 58251 84854
0 12843 5 1 1 12842
0 12844 7 1 2 12837 12843
0 12845 5 2 1 12844
0 12846 7 1 2 69734 84857
0 12847 5 1 1 12846
0 12848 7 5 2 72075 78005
0 12849 7 1 2 71027 84859
0 12850 5 1 1 12849
0 12851 7 4 2 65506 76169
0 12852 5 1 1 84864
0 12853 7 1 2 74932 12852
0 12854 7 1 2 12850 12853
0 12855 5 1 1 12854
0 12856 7 1 2 58427 12855
0 12857 5 1 1 12856
0 12858 7 1 2 12847 12857
0 12859 5 1 1 12858
0 12860 7 1 2 60301 12859
0 12861 5 2 1 12860
0 12862 7 1 2 12829 84868
0 12863 7 1 2 12814 12862
0 12864 5 1 1 12863
0 12865 7 1 2 79312 12864
0 12866 5 1 1 12865
0 12867 7 9 2 62633 63173
0 12868 5 2 1 84870
0 12869 7 9 2 72775 84871
0 12870 5 1 1 84881
0 12871 7 2 2 77634 84882
0 12872 7 2 2 65001 71874
0 12873 5 3 1 84892
0 12874 7 1 2 73289 80169
0 12875 7 1 2 84894 12874
0 12876 7 1 2 84890 12875
0 12877 5 1 1 12876
0 12878 7 1 2 12866 12877
0 12879 5 1 1 12878
0 12880 7 1 2 64480 12879
0 12881 5 1 1 12880
0 12882 7 1 2 64005 73453
0 12883 5 4 1 12882
0 12884 7 1 2 57979 84897
0 12885 5 1 1 12884
0 12886 7 2 2 1375 12885
0 12887 5 2 1 84901
0 12888 7 2 2 71475 84903
0 12889 5 2 1 84905
0 12890 7 4 2 76089 76324
0 12891 5 2 1 84909
0 12892 7 1 2 71252 84913
0 12893 7 1 2 84907 12892
0 12894 5 1 1 12893
0 12895 7 1 2 78360 12894
0 12896 5 1 1 12895
0 12897 7 1 2 71776 73933
0 12898 5 1 1 12897
0 12899 7 7 2 70870 74810
0 12900 5 11 1 84915
0 12901 7 1 2 12898 84922
0 12902 5 1 1 12901
0 12903 7 3 2 71476 82128
0 12904 5 1 1 84933
0 12905 7 1 2 12902 84934
0 12906 5 1 1 12905
0 12907 7 1 2 71164 71777
0 12908 5 1 1 12907
0 12909 7 4 2 70720 74811
0 12910 5 1 1 84936
0 12911 7 1 2 78979 84937
0 12912 5 1 1 12911
0 12913 7 1 2 12908 12912
0 12914 7 1 2 12906 12913
0 12915 5 1 1 12914
0 12916 7 1 2 71875 12915
0 12917 5 1 1 12916
0 12918 7 4 2 70253 4964
0 12919 7 1 2 73896 84940
0 12920 5 1 1 12919
0 12921 7 3 2 81156 84281
0 12922 5 1 1 84944
0 12923 7 2 2 73164 81154
0 12924 7 1 2 84945 84947
0 12925 5 1 1 12924
0 12926 7 1 2 12920 12925
0 12927 7 1 2 12917 12926
0 12928 7 1 2 12896 12927
0 12929 5 1 1 12928
0 12930 7 1 2 58428 12929
0 12931 5 1 1 12930
0 12932 7 1 2 77773 82546
0 12933 7 1 2 78361 12932
0 12934 5 1 1 12933
0 12935 7 2 2 70164 74857
0 12936 5 1 1 84949
0 12937 7 5 2 58252 69814
0 12938 7 1 2 83073 84951
0 12939 7 1 2 84950 12938
0 12940 5 1 1 12939
0 12941 7 1 2 12934 12940
0 12942 7 2 2 12931 12941
0 12943 5 1 1 84956
0 12944 7 1 2 64685 84957
0 12945 5 1 1 12944
0 12946 7 2 2 68351 76904
0 12947 5 4 1 84958
0 12948 7 1 2 84837 72549
0 12949 7 2 2 84960 12948
0 12950 5 1 1 84964
0 12951 7 2 2 67816 84965
0 12952 5 3 1 84966
0 12953 7 1 2 63174 84968
0 12954 5 1 1 12953
0 12955 7 1 2 77417 77572
0 12956 5 1 1 12955
0 12957 7 1 2 84530 83791
0 12958 5 1 1 12957
0 12959 7 1 2 12956 12958
0 12960 7 2 2 12954 12959
0 12961 5 1 1 84971
0 12962 7 1 2 60838 84972
0 12963 5 1 1 12962
0 12964 7 3 2 58429 80879
0 12965 5 21 1 84973
0 12966 7 1 2 84976 72717
0 12967 5 1 1 12966
0 12968 7 4 2 71675 71109
0 12969 5 1 1 84997
0 12970 7 1 2 77044 84998
0 12971 5 1 1 12970
0 12972 7 1 2 63175 71594
0 12973 5 1 1 12972
0 12974 7 1 2 65507 12973
0 12975 7 1 2 12971 12974
0 12976 7 1 2 12967 12975
0 12977 5 1 1 12976
0 12978 7 1 2 64234 12977
0 12979 7 1 2 12963 12978
0 12980 5 1 1 12979
0 12981 7 1 2 84865 72718
0 12982 5 1 1 12981
0 12983 7 5 2 65002 67157
0 12984 5 1 1 85001
0 12985 7 1 2 72143 85002
0 12986 5 1 1 12985
0 12987 7 1 2 12982 12986
0 12988 5 1 1 12987
0 12989 7 1 2 63176 12988
0 12990 5 1 1 12989
0 12991 7 1 2 74531 81833
0 12992 5 2 1 12991
0 12993 7 1 2 84860 80926
0 12994 5 1 1 12993
0 12995 7 1 2 74933 12994
0 12996 5 1 1 12995
0 12997 7 1 2 62354 12996
0 12998 5 1 1 12997
0 12999 7 1 2 85006 12998
0 13000 7 1 2 12990 12999
0 13001 5 1 1 13000
0 13002 7 1 2 84977 13001
0 13003 5 1 1 13002
0 13004 7 1 2 59985 13003
0 13005 7 1 2 12980 13004
0 13006 5 1 1 13005
0 13007 7 1 2 59761 13006
0 13008 7 1 2 12945 13007
0 13009 5 1 1 13008
0 13010 7 2 2 76325 82631
0 13011 5 1 1 85008
0 13012 7 1 2 85009 84480
0 13013 7 1 2 80913 13012
0 13014 5 1 1 13013
0 13015 7 1 2 13009 13014
0 13016 5 1 1 13015
0 13017 7 1 2 69336 13016
0 13018 5 1 1 13017
0 13019 7 1 2 12881 13018
0 13020 5 1 1 13019
0 13021 7 1 2 63476 13020
0 13022 5 1 1 13021
0 13023 7 1 2 82935 81067
0 13024 5 1 1 13023
0 13025 7 1 2 58430 84935
0 13026 5 1 1 13025
0 13027 7 1 2 13024 13026
0 13028 5 1 1 13027
0 13029 7 1 2 59762 13028
0 13030 5 1 1 13029
0 13031 7 1 2 80585 83642
0 13032 5 1 1 13031
0 13033 7 1 2 13030 13032
0 13034 5 1 1 13033
0 13035 7 1 2 80914 13034
0 13036 5 1 1 13035
0 13037 7 2 2 62634 81295
0 13038 5 1 1 85010
0 13039 7 1 2 84941 13038
0 13040 5 1 1 13039
0 13041 7 1 2 71253 81296
0 13042 5 1 1 13041
0 13043 7 1 2 84948 13042
0 13044 5 1 1 13043
0 13045 7 1 2 13040 13044
0 13046 5 1 1 13045
0 13047 7 1 2 76619 13046
0 13048 5 1 1 13047
0 13049 7 1 2 13036 13048
0 13050 5 1 1 13049
0 13051 7 1 2 76026 13050
0 13052 5 1 1 13051
0 13053 7 2 2 59306 68988
0 13054 5 1 1 85012
0 13055 7 2 2 78732 85013
0 13056 5 1 1 85014
0 13057 7 7 2 57980 85015
0 13058 5 3 1 85016
0 13059 7 1 2 70672 85017
0 13060 5 1 1 13059
0 13061 7 2 2 60839 84855
0 13062 5 1 1 85026
0 13063 7 2 2 65508 75321
0 13064 5 1 1 85028
0 13065 7 1 2 60532 85029
0 13066 5 1 1 13065
0 13067 7 1 2 13062 13066
0 13068 5 1 1 13067
0 13069 7 1 2 68763 13068
0 13070 5 1 1 13069
0 13071 7 1 2 67292 82499
0 13072 5 1 1 13071
0 13073 7 1 2 13072 83983
0 13074 7 1 2 13070 13073
0 13075 5 1 1 13074
0 13076 7 1 2 65003 13075
0 13077 5 1 1 13076
0 13078 7 1 2 65509 83500
0 13079 5 1 1 13078
0 13080 7 1 2 57981 75927
0 13081 5 1 1 13080
0 13082 7 1 2 13081 75833
0 13083 5 2 1 13082
0 13084 7 1 2 68601 85030
0 13085 5 1 1 13084
0 13086 7 1 2 60840 80145
0 13087 7 1 2 13085 13086
0 13088 5 1 1 13087
0 13089 7 1 2 13079 13088
0 13090 5 1 1 13089
0 13091 7 1 2 13077 13090
0 13092 5 1 1 13091
0 13093 7 1 2 58253 13092
0 13094 5 1 1 13093
0 13095 7 1 2 13060 13094
0 13096 5 1 1 13095
0 13097 7 1 2 64235 13096
0 13098 5 1 1 13097
0 13099 7 3 2 76376 76392
0 13100 5 2 1 85032
0 13101 7 1 2 67293 85035
0 13102 5 1 1 13101
0 13103 7 1 2 13102 79627
0 13104 5 1 1 13103
0 13105 7 1 2 68352 13104
0 13106 5 2 1 13105
0 13107 7 1 2 82144 82482
0 13108 5 1 1 13107
0 13109 7 1 2 79075 13108
0 13110 5 1 1 13109
0 13111 7 4 2 76170 83887
0 13112 5 4 1 85039
0 13113 7 1 2 65510 83309
0 13114 5 2 1 13113
0 13115 7 1 2 85040 85047
0 13116 7 1 2 13110 13115
0 13117 7 1 2 85037 13116
0 13118 5 1 1 13117
0 13119 7 1 2 59511 13118
0 13120 5 1 1 13119
0 13121 7 1 2 85043 81999
0 13122 5 1 1 13121
0 13123 7 2 2 59512 80490
0 13124 5 2 1 85049
0 13125 7 1 2 78967 76299
0 13126 5 2 1 13125
0 13127 7 1 2 85051 85053
0 13128 5 1 1 13127
0 13129 7 1 2 77927 13128
0 13130 5 1 1 13129
0 13131 7 1 2 63177 64686
0 13132 7 1 2 13130 13131
0 13133 7 1 2 13122 13132
0 13134 7 1 2 13120 13133
0 13135 5 1 1 13134
0 13136 7 1 2 64236 84969
0 13137 5 1 1 13136
0 13138 7 1 2 84849 13137
0 13139 5 2 1 13138
0 13140 7 1 2 60841 85055
0 13141 5 1 1 13140
0 13142 7 1 2 59106 71584
0 13143 5 1 1 13142
0 13144 7 1 2 64237 13143
0 13145 5 1 1 13144
0 13146 7 1 2 84566 13145
0 13147 5 1 1 13146
0 13148 7 1 2 65511 13147
0 13149 5 1 1 13148
0 13150 7 1 2 78539 84238
0 13151 5 1 1 13150
0 13152 7 1 2 58431 13151
0 13153 7 1 2 13149 13152
0 13154 7 1 2 13141 13153
0 13155 5 1 1 13154
0 13156 7 1 2 13135 13155
0 13157 5 1 1 13156
0 13158 7 1 2 84869 13157
0 13159 7 1 2 13098 13158
0 13160 5 1 1 13159
0 13161 7 1 2 72076 79052
0 13162 5 1 1 13161
0 13163 7 2 2 77958 13162
0 13164 5 5 1 85057
0 13165 7 1 2 62355 85059
0 13166 5 1 1 13165
0 13167 7 2 2 13166 84749
0 13168 5 3 1 85064
0 13169 7 1 2 65512 72702
0 13170 5 2 1 13169
0 13171 7 2 2 67158 85069
0 13172 5 1 1 85071
0 13173 7 1 2 85065 13172
0 13174 5 1 1 13173
0 13175 7 6 2 64238 80798
0 13176 5 2 1 85073
0 13177 7 1 2 13174 85074
0 13178 5 1 1 13177
0 13179 7 1 2 59986 13178
0 13180 5 1 1 13179
0 13181 7 1 2 64481 13180
0 13182 7 1 2 13160 13181
0 13183 5 1 1 13182
0 13184 7 11 2 58432 60302
0 13185 5 1 1 85081
0 13186 7 1 2 80202 85082
0 13187 7 1 2 83459 13186
0 13188 5 1 1 13187
0 13189 7 1 2 77838 13188
0 13190 5 1 1 13189
0 13191 7 1 2 82332 13190
0 13192 5 1 1 13191
0 13193 7 5 2 63178 59987
0 13194 7 5 2 64006 64482
0 13195 7 2 2 62635 85097
0 13196 5 2 1 85102
0 13197 7 1 2 85092 85103
0 13198 7 1 2 85060 13197
0 13199 5 1 1 13198
0 13200 7 1 2 13192 13199
0 13201 5 1 1 13200
0 13202 7 1 2 62356 13201
0 13203 5 1 1 13202
0 13204 7 5 2 63179 60303
0 13205 7 2 2 65513 79818
0 13206 5 1 1 85111
0 13207 7 2 2 70288 83998
0 13208 7 1 2 70733 85113
0 13209 5 1 1 13208
0 13210 7 1 2 13206 13209
0 13211 5 1 1 13210
0 13212 7 1 2 85106 13211
0 13213 5 1 1 13212
0 13214 7 1 2 13203 13213
0 13215 5 1 1 13214
0 13216 7 1 2 71254 13215
0 13217 5 1 1 13216
0 13218 7 1 2 64239 12961
0 13219 5 1 1 13218
0 13220 7 3 2 59513 84978
0 13221 7 1 2 83792 85115
0 13222 5 1 1 13221
0 13223 7 1 2 77598 83680
0 13224 5 1 1 13223
0 13225 7 1 2 60842 13224
0 13226 7 1 2 13222 13225
0 13227 7 1 2 13219 13226
0 13228 5 1 1 13227
0 13229 7 3 2 68490 81834
0 13230 5 2 1 85118
0 13231 7 3 2 67294 85121
0 13232 5 1 1 85123
0 13233 7 1 2 84727 85124
0 13234 5 1 1 13233
0 13235 7 19 2 58433 71477
0 13236 5 45 1 85126
0 13237 7 1 2 57666 84728
0 13238 5 2 1 13237
0 13239 7 1 2 85145 85190
0 13240 7 1 2 13234 13239
0 13241 5 1 1 13240
0 13242 7 1 2 71595 72792
0 13243 5 1 1 13242
0 13244 7 1 2 65514 13243
0 13245 7 1 2 13241 13244
0 13246 5 1 1 13245
0 13247 7 1 2 79819 13246
0 13248 7 1 2 13228 13247
0 13249 5 1 1 13248
0 13250 7 1 2 13217 13249
0 13251 7 1 2 13183 13250
0 13252 5 1 1 13251
0 13253 7 1 2 60113 13252
0 13254 5 1 1 13253
0 13255 7 1 2 13052 13254
0 13256 5 1 1 13255
0 13257 7 1 2 74887 13256
0 13258 5 1 1 13257
0 13259 7 1 2 13022 13258
0 13260 5 1 1 13259
0 13261 7 1 2 61195 13260
0 13262 5 1 1 13261
0 13263 7 3 2 58739 76027
0 13264 5 3 1 85192
0 13265 7 4 2 60114 66751
0 13266 5 1 1 85198
0 13267 7 1 2 85195 13266
0 13268 5 1 1 13267
0 13269 7 5 2 62916 76669
0 13270 5 1 1 85202
0 13271 7 4 2 64240 76670
0 13272 5 2 1 85207
0 13273 7 3 2 13270 85211
0 13274 5 3 1 85213
0 13275 7 5 2 75570 85214
0 13276 5 1 1 85219
0 13277 7 2 2 72044 76256
0 13278 7 1 2 68602 85224
0 13279 5 1 1 13278
0 13280 7 2 2 57384 83749
0 13281 5 2 1 85226
0 13282 7 1 2 65515 85227
0 13283 5 1 1 13282
0 13284 7 1 2 81684 13283
0 13285 5 1 1 13284
0 13286 7 1 2 65004 13285
0 13287 5 1 1 13286
0 13288 7 1 2 75867 75210
0 13289 5 1 1 13288
0 13290 7 3 2 69996 74219
0 13291 5 2 1 85230
0 13292 7 1 2 60304 85231
0 13293 5 2 1 13292
0 13294 7 1 2 13289 85235
0 13295 7 1 2 13287 13294
0 13296 7 1 2 13279 13295
0 13297 5 1 1 13296
0 13298 7 1 2 85220 13297
0 13299 5 1 1 13298
0 13300 7 1 2 76620 69713
0 13301 5 1 1 13300
0 13302 7 3 2 58434 78072
0 13303 5 1 1 85237
0 13304 7 1 2 71165 77850
0 13305 5 3 1 13304
0 13306 7 1 2 13303 85240
0 13307 5 1 1 13306
0 13308 7 2 2 68227 72550
0 13309 5 3 1 85243
0 13310 7 1 2 72017 85245
0 13311 7 1 2 13307 13310
0 13312 5 1 1 13311
0 13313 7 1 2 13301 13312
0 13314 7 1 2 13299 13313
0 13315 5 1 1 13314
0 13316 7 1 2 67295 13315
0 13317 5 1 1 13316
0 13318 7 2 2 70773 69815
0 13319 5 1 1 85248
0 13320 7 1 2 73542 85249
0 13321 5 1 1 13320
0 13322 7 1 2 79343 13321
0 13323 5 1 1 13322
0 13324 7 1 2 58435 13323
0 13325 5 1 1 13324
0 13326 7 3 2 63180 72843
0 13327 7 3 2 70774 74120
0 13328 7 1 2 85250 85253
0 13329 5 1 1 13328
0 13330 7 1 2 13325 13329
0 13331 5 1 1 13330
0 13332 7 1 2 68603 13331
0 13333 5 1 1 13332
0 13334 7 3 2 60533 69785
0 13335 5 2 1 85256
0 13336 7 5 2 58436 79334
0 13337 7 1 2 85259 85261
0 13338 5 1 1 13337
0 13339 7 3 2 68764 75571
0 13340 7 1 2 73225 85266
0 13341 7 1 2 83314 13340
0 13342 5 1 1 13341
0 13343 7 1 2 13338 13342
0 13344 7 1 2 13333 13343
0 13345 5 1 1 13344
0 13346 7 1 2 57667 13345
0 13347 5 1 1 13346
0 13348 7 1 2 83787 75674
0 13349 5 1 1 13348
0 13350 7 1 2 85262 13349
0 13351 5 1 1 13350
0 13352 7 1 2 13347 13351
0 13353 5 1 1 13352
0 13354 7 1 2 70398 13353
0 13355 5 1 1 13354
0 13356 7 1 2 79344 79320
0 13357 5 1 1 13356
0 13358 7 1 2 57982 13357
0 13359 5 1 1 13358
0 13360 7 2 2 65516 74638
0 13361 5 1 1 85269
0 13362 7 2 2 69721 13361
0 13363 5 1 1 85271
0 13364 7 1 2 59763 13363
0 13365 5 1 1 13364
0 13366 7 1 2 13359 13365
0 13367 5 1 1 13366
0 13368 7 1 2 59514 13367
0 13369 5 1 1 13368
0 13370 7 1 2 83944 78073
0 13371 5 1 1 13370
0 13372 7 1 2 13369 13371
0 13373 5 1 1 13372
0 13374 7 1 2 58437 13373
0 13375 5 1 1 13374
0 13376 7 1 2 74532 85260
0 13377 5 1 1 13376
0 13378 7 2 2 77309 83289
0 13379 5 1 1 85273
0 13380 7 1 2 59107 85274
0 13381 5 1 1 13380
0 13382 7 1 2 13377 13381
0 13383 5 1 1 13382
0 13384 7 1 2 57668 13383
0 13385 5 1 1 13384
0 13386 7 2 2 70811 84895
0 13387 5 1 1 85275
0 13388 7 1 2 70089 85276
0 13389 5 1 1 13388
0 13390 7 1 2 74533 13389
0 13391 5 1 1 13390
0 13392 7 1 2 13385 13391
0 13393 5 1 1 13392
0 13394 7 1 2 67999 80766
0 13395 5 1 1 13394
0 13396 7 1 2 76671 13395
0 13397 5 7 1 13396
0 13398 7 1 2 13393 85277
0 13399 5 1 1 13398
0 13400 7 1 2 77355 71969
0 13401 5 1 1 13400
0 13402 7 1 2 79672 74534
0 13403 5 2 1 13402
0 13404 7 1 2 13401 85284
0 13405 5 1 1 13404
0 13406 7 1 2 13405 83158
0 13407 5 1 1 13406
0 13408 7 1 2 72018 82735
0 13409 5 1 1 13408
0 13410 7 1 2 85285 13409
0 13411 5 1 1 13410
0 13412 7 1 2 63181 78919
0 13413 5 23 1 13412
0 13414 7 1 2 59764 85286
0 13415 7 1 2 13411 13414
0 13416 5 1 1 13415
0 13417 7 1 2 13407 13416
0 13418 5 1 1 13417
0 13419 7 1 2 68604 13418
0 13420 5 1 1 13419
0 13421 7 1 2 77778 73374
0 13422 7 1 2 79744 13421
0 13423 5 1 1 13422
0 13424 7 1 2 13420 13423
0 13425 7 1 2 13399 13424
0 13426 7 1 2 13375 13425
0 13427 7 1 2 13355 13426
0 13428 7 1 2 13317 13427
0 13429 5 1 1 13428
0 13430 7 1 2 13268 13429
0 13431 5 1 1 13430
0 13432 7 6 2 60115 79873
0 13433 7 1 2 69722 13379
0 13434 5 1 1 13433
0 13435 7 1 2 75322 13434
0 13436 5 1 1 13435
0 13437 7 1 2 67733 84961
0 13438 5 1 1 13437
0 13439 7 1 2 76775 13438
0 13440 5 1 1 13439
0 13441 7 2 2 59515 67734
0 13442 5 1 1 85315
0 13443 7 1 2 65517 13442
0 13444 7 1 2 13440 13443
0 13445 5 1 1 13444
0 13446 7 1 2 57385 80055
0 13447 5 1 1 13446
0 13448 7 1 2 13447 79740
0 13449 5 1 1 13448
0 13450 7 1 2 67296 13449
0 13451 5 1 1 13450
0 13452 7 1 2 12950 78265
0 13453 5 1 1 13452
0 13454 7 1 2 64241 74367
0 13455 5 3 1 13454
0 13456 7 1 2 58254 85317
0 13457 5 1 1 13456
0 13458 7 2 2 60843 13457
0 13459 7 1 2 64242 9228
0 13460 5 1 1 13459
0 13461 7 1 2 67847 13460
0 13462 5 1 1 13461
0 13463 7 1 2 76534 75110
0 13464 5 1 1 13463
0 13465 7 1 2 13462 13464
0 13466 7 1 2 85320 13465
0 13467 7 1 2 13453 13466
0 13468 7 1 2 13451 13467
0 13469 5 1 1 13468
0 13470 7 1 2 13445 13469
0 13471 5 1 1 13470
0 13472 7 1 2 13436 13471
0 13473 5 1 1 13472
0 13474 7 1 2 75506 13473
0 13475 5 1 1 13474
0 13476 7 4 2 65518 73714
0 13477 5 1 1 85322
0 13478 7 1 2 77809 13477
0 13479 5 3 1 13478
0 13480 7 1 2 85119 85326
0 13481 5 1 1 13480
0 13482 7 3 2 60844 77851
0 13483 5 1 1 85329
0 13484 7 1 2 83788 85330
0 13485 5 1 1 13484
0 13486 7 1 2 13485 80852
0 13487 7 1 2 13481 13486
0 13488 5 1 1 13487
0 13489 7 1 2 62357 13488
0 13490 5 1 1 13489
0 13491 7 1 2 64243 72045
0 13492 5 1 1 13491
0 13493 7 1 2 84750 13492
0 13494 5 2 1 13493
0 13495 7 1 2 76730 85332
0 13496 5 1 1 13495
0 13497 7 1 2 13490 13496
0 13498 5 1 1 13497
0 13499 7 1 2 76171 13498
0 13500 5 1 1 13499
0 13501 7 7 2 64007 59765
0 13502 7 3 2 77418 85334
0 13503 5 2 1 85341
0 13504 7 1 2 77839 85344
0 13505 5 1 1 13504
0 13506 7 1 2 85066 13505
0 13507 5 1 1 13506
0 13508 7 9 2 67424 73823
0 13509 5 2 1 85346
0 13510 7 5 2 68073 85347
0 13511 5 1 1 85357
0 13512 7 1 2 72543 75323
0 13513 5 1 1 13512
0 13514 7 1 2 85358 13513
0 13515 5 1 1 13514
0 13516 7 5 2 60305 68074
0 13517 5 2 1 85362
0 13518 7 1 2 78396 85367
0 13519 7 1 2 13515 13518
0 13520 5 1 1 13519
0 13521 7 1 2 13507 13520
0 13522 5 1 1 13521
0 13523 7 1 2 64244 13522
0 13524 5 1 1 13523
0 13525 7 1 2 59516 83249
0 13526 5 1 1 13525
0 13527 7 1 2 64483 13526
0 13528 5 1 1 13527
0 13529 7 2 2 64008 85203
0 13530 7 1 2 1138 85369
0 13531 7 1 2 13528 13530
0 13532 5 1 1 13531
0 13533 7 2 2 65519 80896
0 13534 5 1 1 85371
0 13535 7 1 2 13532 13534
0 13536 5 1 1 13535
0 13537 7 1 2 62636 13536
0 13538 5 1 1 13537
0 13539 7 1 2 13524 13538
0 13540 7 1 2 13500 13539
0 13541 7 1 2 13475 13540
0 13542 5 1 1 13541
0 13543 7 1 2 85309 13542
0 13544 5 1 1 13543
0 13545 7 1 2 13431 13544
0 13546 5 1 1 13545
0 13547 7 1 2 65816 13546
0 13548 5 1 1 13547
0 13549 7 2 2 62637 69211
0 13550 7 2 2 72776 85373
0 13551 7 10 2 83999 82799
0 13552 5 2 1 85377
0 13553 7 1 2 85375 85378
0 13554 7 1 2 85067 13553
0 13555 5 1 1 13554
0 13556 7 1 2 13548 13555
0 13557 5 1 1 13556
0 13558 7 1 2 62054 13557
0 13559 5 1 1 13558
0 13560 7 1 2 13262 13559
0 13561 5 1 1 13560
0 13562 7 1 2 61545 13561
0 13563 5 1 1 13562
0 13564 7 2 2 70620 73607
0 13565 7 1 2 85389 79192
0 13566 5 2 1 13565
0 13567 7 7 2 64245 73608
0 13568 5 1 1 85393
0 13569 7 1 2 71596 85394
0 13570 5 2 1 13569
0 13571 7 4 2 65817 67297
0 13572 5 6 1 85402
0 13573 7 1 2 71255 80445
0 13574 7 1 2 85406 13573
0 13575 5 1 1 13574
0 13576 7 2 2 67159 73609
0 13577 5 3 1 85412
0 13578 7 1 2 85414 74730
0 13579 7 1 2 13575 13578
0 13580 5 1 1 13579
0 13581 7 1 2 70621 13580
0 13582 5 1 1 13581
0 13583 7 1 2 85400 13582
0 13584 5 1 1 13583
0 13585 7 1 2 64484 13584
0 13586 5 1 1 13585
0 13587 7 2 2 85391 13586
0 13588 5 1 1 85417
0 13589 7 2 2 80189 78890
0 13590 7 1 2 79154 85419
0 13591 5 1 1 13590
0 13592 7 1 2 85246 79172
0 13593 5 1 1 13592
0 13594 7 2 2 59766 71478
0 13595 5 6 1 85421
0 13596 7 2 2 85422 78667
0 13597 5 1 1 85429
0 13598 7 1 2 13593 13597
0 13599 7 1 2 13591 13598
0 13600 5 1 1 13599
0 13601 7 1 2 67160 79780
0 13602 5 1 1 13601
0 13603 7 1 2 61196 13602
0 13604 7 1 2 13600 13603
0 13605 5 1 1 13604
0 13606 7 2 2 64485 71256
0 13607 5 5 1 85431
0 13608 7 1 2 67161 85423
0 13609 5 1 1 13608
0 13610 7 1 2 85433 13609
0 13611 5 1 1 13610
0 13612 7 1 2 75244 13611
0 13613 5 1 1 13612
0 13614 7 2 2 64486 84364
0 13615 5 1 1 85438
0 13616 7 1 2 65818 13615
0 13617 7 1 2 13613 13616
0 13618 5 1 1 13617
0 13619 7 1 2 60845 13618
0 13620 7 1 2 13605 13619
0 13621 5 1 1 13620
0 13622 7 1 2 85418 13621
0 13623 5 1 1 13622
0 13624 7 1 2 63182 13623
0 13625 5 1 1 13624
0 13626 7 2 2 72803 84365
0 13627 7 1 2 61197 72551
0 13628 7 1 2 85440 13627
0 13629 5 1 1 13628
0 13630 7 3 2 64246 73775
0 13631 5 1 1 85442
0 13632 7 1 2 80297 85443
0 13633 5 1 1 13632
0 13634 7 1 2 13629 13633
0 13635 5 1 1 13634
0 13636 7 1 2 62358 13635
0 13637 5 1 1 13636
0 13638 7 2 2 62168 65819
0 13639 7 2 2 84261 85445
0 13640 7 3 2 77419 78241
0 13641 5 1 1 85449
0 13642 7 1 2 85447 85450
0 13643 5 1 1 13642
0 13644 7 1 2 13637 13643
0 13645 5 1 1 13644
0 13646 7 1 2 63858 13645
0 13647 5 1 1 13646
0 13648 7 1 2 13647 2668
0 13649 5 1 1 13648
0 13650 7 1 2 60846 13649
0 13651 5 1 1 13650
0 13652 7 1 2 85392 13651
0 13653 5 1 1 13652
0 13654 7 1 2 64487 13653
0 13655 5 1 1 13654
0 13656 7 1 2 13625 13655
0 13657 5 1 1 13656
0 13658 7 1 2 60116 13657
0 13659 5 1 1 13658
0 13660 7 3 2 64790 76621
0 13661 7 1 2 84443 85452
0 13662 5 1 1 13661
0 13663 7 1 2 13659 13662
0 13664 5 1 1 13663
0 13665 7 1 2 66889 13664
0 13666 5 1 1 13665
0 13667 7 1 2 85196 2816
0 13668 5 12 1 13667
0 13669 7 1 2 77135 82739
0 13670 5 1 1 13669
0 13671 7 1 2 75868 82737
0 13672 5 1 1 13671
0 13673 7 1 2 3580 11223
0 13674 7 1 2 13672 13673
0 13675 7 1 2 13670 13674
0 13676 5 1 1 13675
0 13677 7 1 2 63183 13676
0 13678 5 1 1 13677
0 13679 7 1 2 65520 13678
0 13680 5 1 1 13679
0 13681 7 7 2 64247 76172
0 13682 5 4 1 85467
0 13683 7 2 2 84974 85474
0 13684 5 11 1 85478
0 13685 7 1 2 70960 78266
0 13686 5 1 1 13685
0 13687 7 2 2 67298 84336
0 13688 5 1 1 85491
0 13689 7 1 2 13686 13688
0 13690 5 1 1 13689
0 13691 7 1 2 77136 13690
0 13692 5 1 1 13691
0 13693 7 5 2 63184 60847
0 13694 5 2 1 85493
0 13695 7 1 2 79712 85494
0 13696 7 1 2 84361 13695
0 13697 7 1 2 84288 13696
0 13698 7 1 2 13692 13697
0 13699 5 1 1 13698
0 13700 7 1 2 85480 13699
0 13701 7 1 2 13680 13700
0 13702 5 1 1 13701
0 13703 7 1 2 65820 13702
0 13704 5 1 1 13703
0 13705 7 1 2 70961 85287
0 13706 5 1 1 13705
0 13707 7 1 2 58255 85492
0 13708 5 1 1 13707
0 13709 7 1 2 13706 13708
0 13710 5 1 1 13709
0 13711 7 1 2 60848 13710
0 13712 5 1 1 13711
0 13713 7 2 2 68353 73870
0 13714 7 1 2 77707 85500
0 13715 5 1 1 13714
0 13716 7 1 2 13712 13715
0 13717 5 1 1 13716
0 13718 7 1 2 64248 13717
0 13719 5 1 1 13718
0 13720 7 1 2 85044 74208
0 13721 5 1 1 13720
0 13722 7 1 2 13719 13721
0 13723 5 1 1 13722
0 13724 7 1 2 77137 13723
0 13725 5 1 1 13724
0 13726 7 1 2 67299 85247
0 13727 5 1 1 13726
0 13728 7 1 2 76977 13727
0 13729 5 1 1 13728
0 13730 7 1 2 70962 82484
0 13731 5 1 1 13730
0 13732 7 1 2 65214 82142
0 13733 5 1 1 13732
0 13734 7 1 2 13731 13733
0 13735 5 1 1 13734
0 13736 7 1 2 77138 13735
0 13737 5 1 1 13736
0 13738 7 1 2 82487 13737
0 13739 5 1 1 13738
0 13740 7 1 2 63185 13739
0 13741 5 1 1 13740
0 13742 7 1 2 13729 13741
0 13743 5 1 1 13742
0 13744 7 1 2 59517 13743
0 13745 5 1 1 13744
0 13746 7 1 2 67300 84819
0 13747 5 1 1 13746
0 13748 7 1 2 6741 13747
0 13749 5 1 1 13748
0 13750 7 1 2 65521 13749
0 13751 5 1 1 13750
0 13752 7 1 2 83918 80232
0 13753 5 1 1 13752
0 13754 7 1 2 13751 13753
0 13755 5 1 1 13754
0 13756 7 1 2 58256 13755
0 13757 5 1 1 13756
0 13758 7 2 2 60849 80191
0 13759 5 1 1 85502
0 13760 7 1 2 65522 71597
0 13761 5 1 1 13760
0 13762 7 1 2 13759 13761
0 13763 5 1 1 13762
0 13764 7 1 2 75431 13763
0 13765 5 1 1 13764
0 13766 7 1 2 61198 13765
0 13767 7 1 2 13757 13766
0 13768 7 1 2 13745 13767
0 13769 7 1 2 13725 13768
0 13770 5 1 1 13769
0 13771 7 1 2 13704 13770
0 13772 5 1 1 13771
0 13773 7 1 2 73636 73274
0 13774 5 6 1 13773
0 13775 7 4 2 80745 85504
0 13776 5 1 1 85510
0 13777 7 1 2 73024 13776
0 13778 5 2 1 13777
0 13779 7 1 2 76173 85514
0 13780 5 1 1 13779
0 13781 7 1 2 73001 72760
0 13782 5 2 1 13781
0 13783 7 1 2 13780 85516
0 13784 5 1 1 13783
0 13785 7 1 2 58438 13784
0 13786 5 1 1 13785
0 13787 7 1 2 76880 80647
0 13788 5 1 1 13787
0 13789 7 1 2 13786 13788
0 13790 5 1 1 13789
0 13791 7 1 2 70622 13790
0 13792 5 1 1 13791
0 13793 7 1 2 59767 13792
0 13794 7 1 2 13772 13793
0 13795 5 1 1 13794
0 13796 7 1 2 82936 82500
0 13797 5 1 1 13796
0 13798 7 5 2 65523 82916
0 13799 5 1 1 85518
0 13800 7 1 2 65215 85519
0 13801 5 1 1 13800
0 13802 7 1 2 13797 13801
0 13803 5 1 1 13802
0 13804 7 1 2 65821 13803
0 13805 5 1 1 13804
0 13806 7 1 2 61199 85127
0 13807 7 1 2 82471 13806
0 13808 5 1 1 13807
0 13809 7 1 2 13805 13808
0 13810 5 1 1 13809
0 13811 7 1 2 67301 13810
0 13812 5 1 1 13811
0 13813 7 3 2 59518 73241
0 13814 5 1 1 85523
0 13815 7 1 2 79673 85524
0 13816 5 1 1 13815
0 13817 7 1 2 84337 74650
0 13818 5 1 1 13817
0 13819 7 1 2 13816 13818
0 13820 5 1 1 13819
0 13821 7 1 2 85288 13820
0 13822 5 1 1 13821
0 13823 7 1 2 73275 73061
0 13824 5 6 1 13823
0 13825 7 1 2 58439 70963
0 13826 7 1 2 85526 13825
0 13827 5 1 1 13826
0 13828 7 3 2 63186 73687
0 13829 5 7 1 85532
0 13830 7 12 2 58440 65822
0 13831 5 6 1 85542
0 13832 7 1 2 71970 85554
0 13833 7 1 2 85535 13832
0 13834 5 1 1 13833
0 13835 7 1 2 13827 13834
0 13836 5 1 1 13835
0 13837 7 1 2 70399 13836
0 13838 5 1 1 13837
0 13839 7 2 2 58257 70964
0 13840 7 1 2 80640 85560
0 13841 5 1 1 13840
0 13842 7 1 2 13838 13841
0 13843 7 1 2 13822 13842
0 13844 7 1 2 13812 13843
0 13845 5 1 1 13844
0 13846 7 1 2 77139 13845
0 13847 5 1 1 13846
0 13848 7 1 2 69966 77765
0 13849 5 2 1 13848
0 13850 7 3 2 73165 84634
0 13851 5 10 1 85564
0 13852 7 1 2 57669 72490
0 13853 7 1 2 85565 13852
0 13854 5 1 1 13853
0 13855 7 1 2 85562 13854
0 13856 5 2 1 13855
0 13857 7 1 2 59108 85577
0 13858 5 1 1 13857
0 13859 7 1 2 83974 67012
0 13860 5 1 1 13859
0 13861 7 1 2 13858 13860
0 13862 5 1 1 13861
0 13863 7 1 2 82937 13862
0 13864 5 1 1 13863
0 13865 7 1 2 75849 77758
0 13866 5 1 1 13865
0 13867 7 1 2 71257 13866
0 13868 5 2 1 13867
0 13869 7 1 2 60850 85579
0 13870 5 1 1 13869
0 13871 7 1 2 59519 78800
0 13872 5 1 1 13871
0 13873 7 1 2 13870 13872
0 13874 5 1 1 13873
0 13875 7 1 2 58441 13874
0 13876 5 1 1 13875
0 13877 7 1 2 60851 81035
0 13878 5 1 1 13877
0 13879 7 1 2 73206 85520
0 13880 5 1 1 13879
0 13881 7 1 2 13878 13880
0 13882 5 1 1 13881
0 13883 7 1 2 67302 13882
0 13884 5 1 1 13883
0 13885 7 1 2 60852 72649
0 13886 5 2 1 13885
0 13887 7 1 2 59307 85521
0 13888 5 1 1 13887
0 13889 7 1 2 85581 13888
0 13890 5 1 1 13889
0 13891 7 1 2 57983 13890
0 13892 5 1 1 13891
0 13893 7 1 2 13884 13892
0 13894 7 1 2 13876 13893
0 13895 7 1 2 13864 13894
0 13896 5 1 1 13895
0 13897 7 1 2 65823 13896
0 13898 5 1 1 13897
0 13899 7 1 2 84942 80192
0 13900 5 1 1 13899
0 13901 7 1 2 73166 82840
0 13902 7 1 2 85580 13901
0 13903 5 1 1 13902
0 13904 7 1 2 13900 13903
0 13905 5 1 1 13904
0 13906 7 1 2 80553 13905
0 13907 5 1 1 13906
0 13908 7 1 2 64488 13907
0 13909 7 1 2 13898 13908
0 13910 7 1 2 13847 13909
0 13911 5 1 1 13910
0 13912 7 2 2 13795 13911
0 13913 5 1 1 85583
0 13914 7 1 2 85455 85584
0 13915 5 1 1 13914
0 13916 7 4 2 64489 73303
0 13917 5 1 1 85585
0 13918 7 4 2 60306 78476
0 13919 5 4 1 85589
0 13920 7 2 2 79335 85590
0 13921 5 2 1 85597
0 13922 7 1 2 13917 85599
0 13923 5 1 1 13922
0 13924 7 1 2 59520 13923
0 13925 5 1 1 13924
0 13926 7 1 2 78074 73610
0 13927 5 3 1 13926
0 13928 7 1 2 13925 85601
0 13929 5 1 1 13928
0 13930 7 1 2 58442 13929
0 13931 5 1 1 13930
0 13932 7 2 2 65824 77796
0 13933 7 1 2 74121 85604
0 13934 5 1 1 13933
0 13935 7 1 2 13931 13934
0 13936 5 2 1 13935
0 13937 7 1 2 85456 85606
0 13938 5 1 1 13937
0 13939 7 4 2 78477 74977
0 13940 7 1 2 85310 85608
0 13941 7 1 2 80857 13940
0 13942 5 1 1 13941
0 13943 7 1 2 13938 13942
0 13944 5 1 1 13943
0 13945 7 1 2 76955 13944
0 13946 5 1 1 13945
0 13947 7 1 2 13915 13946
0 13948 7 1 2 13666 13947
0 13949 5 1 1 13948
0 13950 7 1 2 83017 13949
0 13951 5 1 1 13950
0 13952 7 1 2 13563 13951
0 13953 5 1 1 13952
0 13954 7 1 2 63599 13953
0 13955 5 1 1 13954
0 13956 7 1 2 76956 85607
0 13957 5 1 1 13956
0 13958 7 1 2 13913 13957
0 13959 5 1 1 13958
0 13960 7 1 2 66752 13959
0 13961 5 1 1 13960
0 13962 7 1 2 75835 76079
0 13963 5 1 1 13962
0 13964 7 1 2 13963 84389
0 13965 5 3 1 13964
0 13966 7 1 2 76174 85612
0 13967 5 1 1 13966
0 13968 7 3 2 59768 76889
0 13969 5 2 1 85615
0 13970 7 1 2 13967 85616
0 13971 5 1 1 13970
0 13972 7 1 2 64490 85420
0 13973 5 1 1 13972
0 13974 7 1 2 64249 13973
0 13975 7 1 2 13971 13974
0 13976 5 1 1 13975
0 13977 7 1 2 85345 73732
0 13978 5 1 1 13977
0 13979 7 1 2 85613 13978
0 13980 5 1 1 13979
0 13981 7 1 2 13980 6463
0 13982 7 1 2 13976 13981
0 13983 5 1 1 13982
0 13984 7 1 2 63187 13983
0 13985 5 1 1 13984
0 13986 7 1 2 85441 85614
0 13987 5 1 1 13986
0 13988 7 8 2 58443 64009
0 13989 7 3 2 62638 85620
0 13990 7 1 2 71394 85628
0 13991 5 1 1 13990
0 13992 7 1 2 13987 13991
0 13993 5 1 1 13992
0 13994 7 1 2 64491 13993
0 13995 5 1 1 13994
0 13996 7 1 2 61200 13995
0 13997 7 1 2 13985 13996
0 13998 5 1 1 13997
0 13999 7 1 2 75245 80989
0 14000 5 1 1 13999
0 14001 7 3 2 63188 84366
0 14002 5 1 1 85631
0 14003 7 1 2 64492 85632
0 14004 5 1 1 14003
0 14005 7 1 2 65825 14004
0 14006 7 1 2 14000 14005
0 14007 5 1 1 14006
0 14008 7 1 2 60853 14007
0 14009 7 1 2 13998 14008
0 14010 5 1 1 14009
0 14011 7 3 2 64010 79155
0 14012 7 5 2 77420 85634
0 14013 7 1 2 85390 85637
0 14014 5 1 1 14013
0 14015 7 1 2 63189 13588
0 14016 5 1 1 14015
0 14017 7 1 2 14014 14016
0 14018 7 1 2 14010 14017
0 14019 5 1 1 14018
0 14020 7 1 2 66890 14019
0 14021 5 1 1 14020
0 14022 7 1 2 13961 14021
0 14023 5 1 1 14022
0 14024 7 1 2 82710 14023
0 14025 5 1 1 14024
0 14026 7 9 2 61201 71395
0 14027 5 8 1 85642
0 14028 7 3 2 67303 85651
0 14029 5 1 1 85659
0 14030 7 2 2 62917 73688
0 14031 5 2 1 85662
0 14032 7 3 2 72887 85664
0 14033 5 3 1 85666
0 14034 7 1 2 14029 85669
0 14035 7 2 2 85068 14034
0 14036 5 1 1 85672
0 14037 7 1 2 85072 85643
0 14038 5 1 1 14037
0 14039 7 1 2 14036 14038
0 14040 5 2 1 14039
0 14041 7 1 2 76069 85674
0 14042 5 1 1 14041
0 14043 7 1 2 85193 85673
0 14044 5 1 1 14043
0 14045 7 1 2 14042 14044
0 14046 5 1 1 14045
0 14047 7 1 2 75507 14046
0 14048 5 1 1 14047
0 14049 7 3 2 64687 76916
0 14050 7 2 2 67304 71166
0 14051 5 26 1 85679
0 14052 7 2 2 67735 85681
0 14053 5 2 1 85707
0 14054 7 1 2 85682 82860
0 14055 5 1 1 14054
0 14056 7 3 2 85709 14055
0 14057 7 1 2 83315 85711
0 14058 5 1 1 14057
0 14059 7 1 2 84952 85027
0 14060 5 1 1 14059
0 14061 7 1 2 14058 14060
0 14062 5 1 1 14061
0 14063 7 1 2 58968 14062
0 14064 5 1 1 14063
0 14065 7 1 2 71167 83987
0 14066 5 1 1 14065
0 14067 7 1 2 14064 14066
0 14068 5 1 1 14067
0 14069 7 1 2 57386 14068
0 14070 5 1 1 14069
0 14071 7 1 2 71729 85031
0 14072 5 1 1 14071
0 14073 7 1 2 80146 14072
0 14074 5 1 1 14073
0 14075 7 1 2 60854 14074
0 14076 5 1 1 14075
0 14077 7 2 2 73215 71642
0 14078 7 1 2 67736 85714
0 14079 5 1 1 14078
0 14080 7 1 2 60307 73871
0 14081 7 1 2 14079 14080
0 14082 5 1 1 14081
0 14083 7 1 2 14076 14082
0 14084 5 1 1 14083
0 14085 7 1 2 71168 14084
0 14086 5 1 1 14085
0 14087 7 1 2 14070 14086
0 14088 5 1 1 14087
0 14089 7 1 2 65826 14088
0 14090 5 1 1 14089
0 14091 7 1 2 76427 73199
0 14092 7 1 2 80915 14091
0 14093 5 1 1 14092
0 14094 7 1 2 14090 14093
0 14095 5 1 1 14094
0 14096 7 1 2 85676 14095
0 14097 5 1 1 14096
0 14098 7 2 2 60855 73084
0 14099 7 1 2 85716 83236
0 14100 5 1 1 14099
0 14101 7 2 2 73637 73025
0 14102 5 11 1 85718
0 14103 7 2 2 70947 85720
0 14104 5 1 1 85731
0 14105 7 1 2 68491 85732
0 14106 5 1 1 14105
0 14107 7 1 2 14100 14106
0 14108 5 1 1 14107
0 14109 7 1 2 58444 14108
0 14110 5 1 1 14109
0 14111 7 1 2 84858 72854
0 14112 5 1 1 14111
0 14113 7 3 2 62918 73652
0 14114 5 2 1 85733
0 14115 7 1 2 67162 85734
0 14116 5 1 1 14115
0 14117 7 1 2 14112 14116
0 14118 5 1 1 14117
0 14119 7 1 2 65524 14118
0 14120 5 1 1 14119
0 14121 7 1 2 14110 14120
0 14122 5 1 1 14121
0 14123 7 1 2 60308 14122
0 14124 5 1 1 14123
0 14125 7 1 2 58445 84158
0 14126 5 1 1 14125
0 14127 7 1 2 68765 85045
0 14128 5 1 1 14127
0 14129 7 1 2 14128 76238
0 14130 5 1 1 14129
0 14131 7 1 2 65005 14130
0 14132 5 1 1 14131
0 14133 7 1 2 78920 14132
0 14134 5 1 1 14133
0 14135 7 1 2 60534 14134
0 14136 5 1 1 14135
0 14137 7 1 2 14126 14136
0 14138 5 1 1 14137
0 14139 7 6 2 61202 69735
0 14140 5 1 1 85738
0 14141 7 1 2 14138 85739
0 14142 5 1 1 14141
0 14143 7 2 2 71802 73085
0 14144 5 1 1 85744
0 14145 7 1 2 62359 85745
0 14146 5 1 1 14145
0 14147 7 1 2 84970 72855
0 14148 5 1 1 14147
0 14149 7 1 2 14146 14148
0 14150 5 1 1 14149
0 14151 7 1 2 58446 14150
0 14152 5 1 1 14151
0 14153 7 1 2 67305 78206
0 14154 5 1 1 14153
0 14155 7 1 2 68075 14154
0 14156 5 2 1 14155
0 14157 7 1 2 57387 85746
0 14158 5 1 1 14157
0 14159 7 1 2 59308 78196
0 14160 5 1 1 14159
0 14161 7 1 2 14158 14160
0 14162 5 1 1 14161
0 14163 7 1 2 71876 14162
0 14164 5 1 1 14163
0 14165 7 1 2 78362 80325
0 14166 5 1 1 14165
0 14167 7 1 2 81061 14166
0 14168 7 1 2 14164 14167
0 14169 5 2 1 14168
0 14170 7 1 2 80476 85748
0 14171 5 1 1 14170
0 14172 7 1 2 14152 14171
0 14173 5 1 1 14172
0 14174 7 1 2 60856 14173
0 14175 5 1 1 14174
0 14176 7 1 2 69756 85498
0 14177 7 3 2 72077 14176
0 14178 7 1 2 80927 85750
0 14179 5 1 1 14178
0 14180 7 1 2 78105 14179
0 14181 5 1 1 14180
0 14182 7 1 2 62360 14181
0 14183 5 1 1 14182
0 14184 7 1 2 58447 85333
0 14185 5 1 1 14184
0 14186 7 1 2 14183 14185
0 14187 5 1 1 14186
0 14188 7 1 2 65827 14187
0 14189 5 1 1 14188
0 14190 7 2 2 61203 72719
0 14191 5 1 1 85753
0 14192 7 1 2 80586 85754
0 14193 5 1 1 14192
0 14194 7 1 2 14189 14193
0 14195 5 1 1 14194
0 14196 7 1 2 76175 14195
0 14197 5 1 1 14196
0 14198 7 4 2 65216 80414
0 14199 7 6 2 58448 65006
0 14200 5 2 1 85759
0 14201 7 1 2 85755 85760
0 14202 5 1 1 14201
0 14203 7 1 2 70357 83250
0 14204 7 1 2 85735 14203
0 14205 5 1 1 14204
0 14206 7 1 2 14202 14205
0 14207 5 1 1 14206
0 14208 7 1 2 64011 14207
0 14209 5 1 1 14208
0 14210 7 2 2 58449 72856
0 14211 5 2 1 85767
0 14212 7 1 2 65525 85768
0 14213 5 1 1 14212
0 14214 7 1 2 14209 14213
0 14215 5 1 1 14214
0 14216 7 1 2 62639 14215
0 14217 5 1 1 14216
0 14218 7 1 2 14197 14217
0 14219 7 1 2 14175 14218
0 14220 7 1 2 14142 14219
0 14221 7 1 2 14124 14220
0 14222 5 1 1 14221
0 14223 7 1 2 66891 14222
0 14224 5 1 1 14223
0 14225 7 10 2 65007 65828
0 14226 5 7 1 85771
0 14227 7 1 2 64250 85772
0 14228 5 1 1 14227
0 14229 7 1 2 73062 14228
0 14230 5 3 1 14229
0 14231 7 1 2 68605 85788
0 14232 5 1 1 14231
0 14233 7 21 2 60309 61204
0 14234 5 6 1 85791
0 14235 7 1 2 74740 82161
0 14236 5 1 1 14235
0 14237 7 1 2 85812 14236
0 14238 5 1 1 14237
0 14239 7 1 2 14232 14238
0 14240 5 1 1 14239
0 14241 7 1 2 65217 14240
0 14242 5 1 1 14241
0 14243 7 1 2 72888 73570
0 14244 7 1 2 75169 14243
0 14245 5 1 1 14244
0 14246 7 1 2 14242 14245
0 14247 5 1 1 14246
0 14248 7 1 2 65526 14247
0 14249 5 1 1 14248
0 14250 7 2 2 58258 85527
0 14251 5 1 1 85818
0 14252 7 1 2 14249 14251
0 14253 5 1 1 14252
0 14254 7 1 2 75324 14253
0 14255 5 1 1 14254
0 14256 7 1 2 79076 85528
0 14257 5 1 1 14256
0 14258 7 5 2 65527 72889
0 14259 5 2 1 85820
0 14260 7 1 2 85781 85821
0 14261 5 1 1 14260
0 14262 7 1 2 14257 14261
0 14263 5 1 1 14262
0 14264 7 1 2 67653 14263
0 14265 5 1 1 14264
0 14266 7 1 2 85529 78756
0 14267 5 1 1 14266
0 14268 7 4 2 59521 85773
0 14269 5 2 1 85827
0 14270 7 1 2 80491 85822
0 14271 7 1 2 85831 14270
0 14272 5 1 1 14271
0 14273 7 1 2 14267 14272
0 14274 5 1 1 14273
0 14275 7 1 2 68354 14274
0 14276 5 1 1 14275
0 14277 7 1 2 14265 14276
0 14278 5 1 1 14277
0 14279 7 1 2 67306 14278
0 14280 5 1 1 14279
0 14281 7 1 2 73026 84621
0 14282 5 1 1 14281
0 14283 7 1 2 81068 14282
0 14284 5 1 1 14283
0 14285 7 7 2 61205 68076
0 14286 5 6 1 85833
0 14287 7 2 2 72524 85840
0 14288 7 1 2 69484 83895
0 14289 5 1 1 14288
0 14290 7 1 2 85846 14289
0 14291 5 1 1 14290
0 14292 7 1 2 78409 76794
0 14293 5 2 1 14292
0 14294 7 1 2 84808 85848
0 14295 7 1 2 14291 14294
0 14296 5 1 1 14295
0 14297 7 1 2 85530 14296
0 14298 5 1 1 14297
0 14299 7 1 2 14284 14298
0 14300 7 1 2 80492 73242
0 14301 5 1 1 14300
0 14302 7 1 2 73611 78757
0 14303 5 1 1 14302
0 14304 7 1 2 14301 14303
0 14305 5 1 1 14304
0 14306 7 1 2 78267 14305
0 14307 5 1 1 14306
0 14308 7 6 2 61206 70400
0 14309 7 1 2 85050 85850
0 14310 5 1 1 14309
0 14311 7 1 2 14307 14310
0 14312 5 1 1 14311
0 14313 7 1 2 68355 14312
0 14314 5 1 1 14313
0 14315 7 1 2 57984 73644
0 14316 5 1 1 14315
0 14317 7 1 2 65829 85270
0 14318 5 1 1 14317
0 14319 7 1 2 58259 85505
0 14320 5 1 1 14319
0 14321 7 1 2 14318 14320
0 14322 7 1 2 14316 14321
0 14323 5 1 1 14322
0 14324 7 1 2 59522 14323
0 14325 5 1 1 14324
0 14326 7 1 2 14314 14325
0 14327 7 1 2 14299 14326
0 14328 7 1 2 14280 14327
0 14329 7 1 2 14255 14328
0 14330 5 1 1 14329
0 14331 7 1 2 79874 14330
0 14332 5 1 1 14331
0 14333 7 1 2 61207 85070
0 14334 7 2 2 64251 79144
0 14335 7 4 2 59988 77421
0 14336 7 1 2 85856 85858
0 14337 7 1 2 14333 14336
0 14338 5 1 1 14337
0 14339 7 1 2 14332 14338
0 14340 5 1 1 14339
0 14341 7 1 2 63190 14340
0 14342 5 1 1 14341
0 14343 7 1 2 72544 85712
0 14344 5 1 1 14343
0 14345 7 1 2 68356 85680
0 14346 5 2 1 14345
0 14347 7 1 2 14344 85862
0 14348 5 1 1 14347
0 14349 7 1 2 65008 14348
0 14350 5 1 1 14349
0 14351 7 1 2 83647 14350
0 14352 5 1 1 14351
0 14353 7 2 2 64688 73304
0 14354 7 1 2 76917 85864
0 14355 7 1 2 14352 14354
0 14356 5 1 1 14355
0 14357 7 1 2 64493 14356
0 14358 7 1 2 14342 14357
0 14359 7 1 2 14224 14358
0 14360 5 1 1 14359
0 14361 7 1 2 68077 80532
0 14362 5 1 1 14361
0 14363 7 1 2 78817 83948
0 14364 5 1 1 14363
0 14365 7 1 2 14362 14364
0 14366 5 1 1 14365
0 14367 7 1 2 85038 14366
0 14368 5 1 1 14367
0 14369 7 1 2 61208 14368
0 14370 5 1 1 14369
0 14371 7 1 2 81293 73216
0 14372 5 1 1 14371
0 14373 7 1 2 73329 85841
0 14374 7 1 2 14372 14373
0 14375 5 1 1 14374
0 14376 7 1 2 14370 14375
0 14377 5 1 1 14376
0 14378 7 1 2 58450 14377
0 14379 5 1 1 14378
0 14380 7 2 2 65830 77310
0 14381 7 2 2 68962 76326
0 14382 5 1 1 85868
0 14383 7 2 2 83074 85869
0 14384 7 1 2 85866 85870
0 14385 5 1 1 14384
0 14386 7 1 2 14379 14385
0 14387 5 1 1 14386
0 14388 7 1 2 71479 14387
0 14389 5 1 1 14388
0 14390 7 2 2 65831 78522
0 14391 5 1 1 85872
0 14392 7 1 2 80568 14391
0 14393 5 1 1 14392
0 14394 7 1 2 58260 14393
0 14395 5 1 1 14394
0 14396 7 3 2 58451 72890
0 14397 5 9 1 85874
0 14398 7 1 2 73571 85875
0 14399 5 1 1 14398
0 14400 7 1 2 14395 14399
0 14401 5 1 1 14400
0 14402 7 1 2 70080 14401
0 14403 5 1 1 14402
0 14404 7 1 2 58452 69816
0 14405 5 1 1 14404
0 14406 7 1 2 80284 14405
0 14407 5 1 1 14406
0 14408 7 1 2 65832 14407
0 14409 5 1 1 14408
0 14410 7 2 2 62919 85877
0 14411 5 2 1 85886
0 14412 7 6 2 85536 85888
0 14413 5 1 1 85890
0 14414 7 5 2 65218 79061
0 14415 5 3 1 85896
0 14416 7 1 2 85891 85897
0 14417 7 1 2 14409 14416
0 14418 5 1 1 14417
0 14419 7 1 2 14403 14418
0 14420 5 1 1 14419
0 14421 7 1 2 65528 14420
0 14422 5 1 1 14421
0 14423 7 1 2 58453 85819
0 14424 5 1 1 14423
0 14425 7 1 2 14422 14424
0 14426 5 1 1 14425
0 14427 7 1 2 75325 14426
0 14428 5 1 1 14427
0 14429 7 1 2 68357 74396
0 14430 5 1 1 14429
0 14431 7 2 2 60857 80038
0 14432 5 1 1 85904
0 14433 7 1 2 14430 14432
0 14434 5 1 1 14433
0 14435 7 1 2 82938 14434
0 14436 5 1 1 14435
0 14437 7 1 2 78937 78169
0 14438 5 4 1 14437
0 14439 7 1 2 65009 85906
0 14440 7 1 2 81094 14439
0 14441 5 1 1 14440
0 14442 7 1 2 14436 14441
0 14443 5 1 1 14442
0 14444 7 1 2 57985 14443
0 14445 5 1 1 14444
0 14446 7 1 2 59309 82939
0 14447 7 1 2 85225 14446
0 14448 5 1 1 14447
0 14449 7 1 2 14445 14448
0 14450 5 1 1 14449
0 14451 7 1 2 68606 14450
0 14452 5 1 1 14451
0 14453 7 2 2 67737 84384
0 14454 7 1 2 82171 85910
0 14455 5 2 1 14454
0 14456 7 1 2 60858 82940
0 14457 7 1 2 85912 14456
0 14458 5 1 1 14457
0 14459 7 1 2 13799 14458
0 14460 5 1 1 14459
0 14461 7 1 2 59310 14460
0 14462 5 1 1 14461
0 14463 7 1 2 85582 14462
0 14464 5 1 1 14463
0 14465 7 1 2 57986 14464
0 14466 5 1 1 14465
0 14467 7 2 2 65219 82941
0 14468 7 1 2 75211 85914
0 14469 5 1 1 14468
0 14470 7 1 2 65010 85522
0 14471 5 1 1 14470
0 14472 7 1 2 14469 14471
0 14473 5 1 1 14472
0 14474 7 1 2 68358 14473
0 14475 5 1 1 14474
0 14476 7 1 2 60859 82172
0 14477 5 2 1 14476
0 14478 7 4 2 67654 82942
0 14479 7 1 2 72046 85918
0 14480 7 1 2 85916 14479
0 14481 5 1 1 14480
0 14482 7 1 2 14475 14481
0 14483 5 1 1 14482
0 14484 7 1 2 67307 14483
0 14485 5 1 1 14484
0 14486 7 1 2 85272 799
0 14487 5 1 1 14486
0 14488 7 1 2 72650 14487
0 14489 5 1 1 14488
0 14490 7 1 2 65833 14489
0 14491 7 1 2 14485 14490
0 14492 7 1 2 14466 14491
0 14493 7 1 2 14452 14492
0 14494 5 1 1 14493
0 14495 7 2 2 62361 75181
0 14496 5 1 1 85922
0 14497 7 3 2 79062 14496
0 14498 5 2 1 85924
0 14499 7 1 2 60860 73217
0 14500 7 1 2 85927 14499
0 14501 5 1 1 14500
0 14502 7 1 2 84481 14501
0 14503 5 1 1 14502
0 14504 7 4 2 68000 83075
0 14505 5 1 1 85929
0 14506 7 1 2 82943 72019
0 14507 7 1 2 85930 14506
0 14508 5 1 1 14507
0 14509 7 1 2 84484 14508
0 14510 5 1 1 14509
0 14511 7 1 2 83785 14510
0 14512 5 1 1 14511
0 14513 7 3 2 57987 68963
0 14514 5 1 1 85933
0 14515 7 2 2 82944 72472
0 14516 7 1 2 85934 85936
0 14517 7 1 2 85925 14516
0 14518 5 1 1 14517
0 14519 7 1 2 61209 14518
0 14520 7 1 2 14512 14519
0 14521 7 1 2 14503 14520
0 14522 5 1 1 14521
0 14523 7 1 2 14494 14522
0 14524 5 1 1 14523
0 14525 7 1 2 14428 14524
0 14526 7 1 2 14389 14525
0 14527 5 1 1 14526
0 14528 7 1 2 66753 14527
0 14529 5 1 1 14528
0 14530 7 1 2 61210 85056
0 14531 5 1 1 14530
0 14532 7 1 2 65834 84367
0 14533 5 2 1 14532
0 14534 7 4 2 65835 85683
0 14535 5 1 1 85940
0 14536 7 1 2 73063 14535
0 14537 5 2 1 14536
0 14538 7 1 2 83793 85944
0 14539 5 1 1 14538
0 14540 7 1 2 85938 14539
0 14541 7 1 2 14531 14540
0 14542 5 1 1 14541
0 14543 7 1 2 60861 14542
0 14544 5 1 1 14543
0 14545 7 2 2 61211 85684
0 14546 7 2 2 65529 85946
0 14547 5 1 1 85948
0 14548 7 1 2 85939 14547
0 14549 5 1 1 14548
0 14550 7 1 2 72720 14549
0 14551 5 1 1 14550
0 14552 7 2 2 70673 85792
0 14553 7 2 2 70022 85950
0 14554 5 1 1 85952
0 14555 7 1 2 62362 85953
0 14556 5 1 1 14555
0 14557 7 3 2 81835 74835
0 14558 5 7 1 85954
0 14559 7 1 2 85941 85955
0 14560 5 1 1 14559
0 14561 7 1 2 85401 14560
0 14562 7 1 2 14556 14561
0 14563 7 1 2 14551 14562
0 14564 7 1 2 14544 14563
0 14565 5 1 1 14564
0 14566 7 1 2 63191 14565
0 14567 5 1 1 14566
0 14568 7 2 2 71396 73612
0 14569 5 1 1 85964
0 14570 7 2 2 64012 85721
0 14571 5 1 1 85966
0 14572 7 2 2 58261 72891
0 14573 5 5 1 85968
0 14574 7 1 2 62640 85970
0 14575 7 1 2 85967 14574
0 14576 5 1 1 14575
0 14577 7 1 2 14569 14576
0 14578 5 1 1 14577
0 14579 7 1 2 85120 14578
0 14580 5 1 1 14579
0 14581 7 2 2 85395 80298
0 14582 5 1 1 85975
0 14583 7 1 2 14580 14582
0 14584 5 1 1 14583
0 14585 7 1 2 62363 14584
0 14586 5 1 1 14585
0 14587 7 3 2 62920 79486
0 14588 5 2 1 85977
0 14589 7 1 2 85413 85978
0 14590 5 1 1 14589
0 14591 7 1 2 80860 73039
0 14592 5 1 1 14591
0 14593 7 5 2 63192 61212
0 14594 5 4 1 85982
0 14595 7 2 2 64252 78995
0 14596 5 1 1 85991
0 14597 7 2 2 85987 85992
0 14598 7 1 2 76176 85407
0 14599 7 1 2 85993 14598
0 14600 5 1 1 14599
0 14601 7 1 2 14592 14600
0 14602 5 2 1 14601
0 14603 7 1 2 83794 85995
0 14604 5 1 1 14603
0 14605 7 3 2 64253 80397
0 14606 5 1 1 85997
0 14607 7 1 2 65011 80299
0 14608 7 1 2 85998 14607
0 14609 5 1 1 14608
0 14610 7 1 2 14604 14609
0 14611 5 1 1 14610
0 14612 7 1 2 60862 14611
0 14613 5 1 1 14612
0 14614 7 1 2 14590 14613
0 14615 7 1 2 14586 14614
0 14616 7 1 2 14567 14615
0 14617 5 1 1 14616
0 14618 7 1 2 66892 14617
0 14619 5 1 1 14618
0 14620 7 1 2 59769 14619
0 14621 7 1 2 14529 14620
0 14622 5 1 1 14621
0 14623 7 1 2 14360 14622
0 14624 5 1 1 14623
0 14625 7 1 2 14097 14624
0 14626 5 1 1 14625
0 14627 7 1 2 64791 14626
0 14628 5 1 1 14627
0 14629 7 1 2 14048 14628
0 14630 5 1 1 14629
0 14631 7 1 2 61546 14630
0 14632 5 1 1 14631
0 14633 7 1 2 14025 14632
0 14634 5 1 1 14633
0 14635 7 1 2 68663 14634
0 14636 5 1 1 14635
0 14637 7 1 2 13955 14636
0 14638 5 1 1 14637
0 14639 7 1 2 61911 14638
0 14640 5 1 1 14639
0 14641 7 1 2 80193 77140
0 14642 5 1 1 14641
0 14643 7 1 2 77696 14642
0 14644 5 1 1 14643
0 14645 7 1 2 60863 14644
0 14646 5 1 1 14645
0 14647 7 1 2 59311 70320
0 14648 7 1 2 76337 14647
0 14649 5 1 1 14648
0 14650 7 1 2 14646 14649
0 14651 5 1 1 14650
0 14652 7 1 2 64254 14651
0 14653 5 1 1 14652
0 14654 7 1 2 77599 84711
0 14655 5 1 1 14654
0 14656 7 3 2 62364 77489
0 14657 5 2 1 86000
0 14658 7 3 2 72333 86001
0 14659 5 1 1 86005
0 14660 7 1 2 67308 14659
0 14661 5 1 1 14660
0 14662 7 1 2 60864 14661
0 14663 5 1 1 14662
0 14664 7 1 2 60535 78468
0 14665 5 1 1 14664
0 14666 7 1 2 77432 14665
0 14667 7 1 2 14663 14666
0 14668 5 1 1 14667
0 14669 7 1 2 59523 14668
0 14670 5 2 1 14669
0 14671 7 1 2 14655 86008
0 14672 7 1 2 14653 14671
0 14673 5 1 1 14672
0 14674 7 1 2 61213 14673
0 14675 5 1 1 14674
0 14676 7 1 2 62365 76522
0 14677 5 2 1 14676
0 14678 7 1 2 81844 86010
0 14679 5 1 1 14678
0 14680 7 1 2 71397 14679
0 14681 5 1 1 14680
0 14682 7 8 2 62921 77583
0 14683 5 2 1 86012
0 14684 7 2 2 64255 76957
0 14685 5 1 1 86022
0 14686 7 1 2 14685 70030
0 14687 5 1 1 14686
0 14688 7 1 2 60536 14687
0 14689 5 1 1 14688
0 14690 7 1 2 71480 14689
0 14691 5 1 1 14690
0 14692 7 1 2 60865 14691
0 14693 5 1 1 14692
0 14694 7 1 2 86020 14693
0 14695 5 1 1 14694
0 14696 7 1 2 62641 14695
0 14697 5 1 1 14696
0 14698 7 1 2 14681 14697
0 14699 5 1 1 14698
0 14700 7 1 2 65836 14699
0 14701 5 1 1 14700
0 14702 7 8 2 65220 73613
0 14703 5 1 1 86024
0 14704 7 1 2 86025 71664
0 14705 5 1 1 14704
0 14706 7 1 2 84734 14705
0 14707 5 1 1 14706
0 14708 7 1 2 71258 14707
0 14709 5 1 1 14708
0 14710 7 1 2 14701 14709
0 14711 7 1 2 14675 14710
0 14712 5 1 1 14711
0 14713 7 1 2 79875 14712
0 14714 5 1 1 14713
0 14715 7 2 2 6248 80687
0 14716 5 2 1 86032
0 14717 7 1 2 67309 86034
0 14718 5 3 1 14717
0 14719 7 1 2 59312 80698
0 14720 5 1 1 14719
0 14721 7 1 2 86036 14720
0 14722 5 1 1 14721
0 14723 7 1 2 65221 14722
0 14724 5 1 1 14723
0 14725 7 1 2 68430 11652
0 14726 7 1 2 14724 14725
0 14727 5 1 1 14726
0 14728 7 1 2 65530 14727
0 14729 5 1 1 14728
0 14730 7 1 2 69967 79759
0 14731 5 1 1 14730
0 14732 7 1 2 14729 14731
0 14733 5 1 1 14732
0 14734 7 8 2 63477 65837
0 14735 7 2 2 77503 86039
0 14736 7 1 2 58262 86047
0 14737 7 1 2 14733 14736
0 14738 5 1 1 14737
0 14739 7 1 2 14714 14738
0 14740 5 1 1 14739
0 14741 7 1 2 58454 14740
0 14742 5 1 1 14741
0 14743 7 3 2 64256 80415
0 14744 5 1 1 86049
0 14745 7 1 2 78903 79876
0 14746 7 1 2 86050 14745
0 14747 7 1 2 80727 14746
0 14748 5 1 1 14747
0 14749 7 1 2 14742 14748
0 14750 5 1 1 14749
0 14751 7 1 2 69521 14750
0 14752 5 1 1 14751
0 14753 7 7 2 66754 70486
0 14754 5 1 1 86052
0 14755 7 1 2 14754 7647
0 14756 5 15 1 14755
0 14757 7 2 2 61214 80996
0 14758 5 2 1 86074
0 14759 7 1 2 77959 72892
0 14760 5 1 1 14759
0 14761 7 3 2 73689 14760
0 14762 7 1 2 74836 86078
0 14763 5 1 1 14762
0 14764 7 1 2 86076 14763
0 14765 5 1 1 14764
0 14766 7 1 2 62922 14765
0 14767 5 1 1 14766
0 14768 7 4 2 62169 84262
0 14769 5 1 1 86081
0 14770 7 6 2 61215 70289
0 14771 7 1 2 68228 86085
0 14772 7 1 2 86082 14771
0 14773 5 1 1 14772
0 14774 7 1 2 14767 14773
0 14775 5 1 1 14774
0 14776 7 1 2 67163 14775
0 14777 5 1 1 14776
0 14778 7 1 2 84526 82459
0 14779 5 1 1 14778
0 14780 7 1 2 14777 14779
0 14781 5 1 1 14780
0 14782 7 1 2 86059 14781
0 14783 5 1 1 14782
0 14784 7 5 2 79877 69522
0 14785 7 1 2 68359 84211
0 14786 5 2 1 14785
0 14787 7 1 2 86096 79764
0 14788 5 2 1 14787
0 14789 7 1 2 59313 86098
0 14790 5 2 1 14789
0 14791 7 1 2 71624 80106
0 14792 5 1 1 14791
0 14793 7 1 2 77650 76539
0 14794 5 1 1 14793
0 14795 7 1 2 14792 14794
0 14796 7 1 2 86100 14795
0 14797 5 1 1 14796
0 14798 7 1 2 61216 14797
0 14799 5 1 1 14798
0 14800 7 1 2 65838 83798
0 14801 5 1 1 14800
0 14802 7 12 2 65012 61217
0 14803 7 1 2 86102 77689
0 14804 5 1 1 14803
0 14805 7 16 2 60310 65839
0 14806 7 4 2 64013 86114
0 14807 5 1 1 86130
0 14808 7 1 2 65222 86131
0 14809 5 1 1 14808
0 14810 7 1 2 14804 14809
0 14811 5 1 1 14810
0 14812 7 1 2 68607 14811
0 14813 5 1 1 14812
0 14814 7 1 2 65013 75358
0 14815 5 1 1 14814
0 14816 7 1 2 85228 14815
0 14817 5 1 1 14816
0 14818 7 1 2 74478 14817
0 14819 5 1 1 14818
0 14820 7 1 2 74694 14807
0 14821 5 1 1 14820
0 14822 7 1 2 14821 83470
0 14823 5 1 1 14822
0 14824 7 1 2 14819 14823
0 14825 7 1 2 14813 14824
0 14826 7 1 2 14801 14825
0 14827 7 1 2 14799 14826
0 14828 5 1 1 14827
0 14829 7 1 2 65531 14828
0 14830 5 1 1 14829
0 14831 7 1 2 70321 75111
0 14832 5 1 1 14831
0 14833 7 1 2 65840 14832
0 14834 5 2 1 14833
0 14835 7 2 2 62642 73290
0 14836 5 3 1 86136
0 14837 7 1 2 72224 86137
0 14838 5 4 1 14837
0 14839 7 1 2 77141 86141
0 14840 5 2 1 14839
0 14841 7 1 2 67164 84343
0 14842 5 2 1 14841
0 14843 7 2 2 70965 86147
0 14844 5 1 1 86149
0 14845 7 1 2 68078 14844
0 14846 7 1 2 86145 14845
0 14847 5 1 1 14846
0 14848 7 1 2 61218 14847
0 14849 5 1 1 14848
0 14850 7 1 2 86134 14849
0 14851 5 1 1 14850
0 14852 7 1 2 58263 14851
0 14853 5 1 1 14852
0 14854 7 2 2 72703 70033
0 14855 5 2 1 86151
0 14856 7 1 2 77658 86153
0 14857 5 1 1 14856
0 14858 7 1 2 60537 14857
0 14859 5 1 1 14858
0 14860 7 1 2 14859 83744
0 14861 5 1 1 14860
0 14862 7 1 2 73243 14861
0 14863 5 1 1 14862
0 14864 7 1 2 74631 84624
0 14865 5 1 1 14864
0 14866 7 2 2 57988 74050
0 14867 5 1 1 86155
0 14868 7 1 2 77142 86156
0 14869 5 1 1 14868
0 14870 7 4 2 60311 73244
0 14871 7 1 2 68766 86157
0 14872 5 3 1 14871
0 14873 7 1 2 14869 86161
0 14874 5 1 1 14873
0 14875 7 1 2 75869 14874
0 14876 5 1 1 14875
0 14877 7 1 2 14865 14876
0 14878 7 1 2 14863 14877
0 14879 7 1 2 14853 14878
0 14880 7 1 2 14830 14879
0 14881 5 1 1 14880
0 14882 7 1 2 59524 14881
0 14883 5 1 1 14882
0 14884 7 1 2 76562 67870
0 14885 5 1 1 14884
0 14886 7 1 2 74328 71639
0 14887 5 1 1 14886
0 14888 7 1 2 14885 14887
0 14889 5 1 1 14888
0 14890 7 1 2 65532 14889
0 14891 5 1 1 14890
0 14892 7 1 2 74329 70120
0 14893 5 1 1 14892
0 14894 7 1 2 14891 14893
0 14895 5 1 1 14894
0 14896 7 1 2 57388 14895
0 14897 5 1 1 14896
0 14898 7 1 2 67871 82260
0 14899 5 1 1 14898
0 14900 7 3 2 59314 74034
0 14901 5 1 1 86164
0 14902 7 1 2 57670 86165
0 14903 5 1 1 14902
0 14904 7 1 2 14899 14903
0 14905 5 1 1 14904
0 14906 7 1 2 65223 14905
0 14907 5 1 1 14906
0 14908 7 1 2 59315 78133
0 14909 5 1 1 14908
0 14910 7 1 2 76433 14909
0 14911 7 1 2 14907 14910
0 14912 7 1 2 14897 14911
0 14913 5 1 1 14912
0 14914 7 1 2 64257 14913
0 14915 5 1 1 14914
0 14916 7 1 2 72721 72402
0 14917 5 1 1 14916
0 14918 7 1 2 68964 14917
0 14919 5 1 1 14918
0 14920 7 1 2 81525 14919
0 14921 5 1 1 14920
0 14922 7 1 2 57389 83246
0 14923 7 1 2 14921 14922
0 14924 5 1 1 14923
0 14925 7 1 2 69908 74106
0 14926 5 1 1 14925
0 14927 7 1 2 64014 74022
0 14928 5 1 1 14927
0 14929 7 1 2 70338 14928
0 14930 5 1 1 14929
0 14931 7 1 2 14926 14930
0 14932 7 1 2 14924 14931
0 14933 7 1 2 14915 14932
0 14934 5 1 1 14933
0 14935 7 1 2 57989 14934
0 14936 5 1 1 14935
0 14937 7 1 2 60538 79604
0 14938 5 3 1 14937
0 14939 7 1 2 86033 79605
0 14940 5 1 1 14939
0 14941 7 3 2 86167 14940
0 14942 7 1 2 69761 86170
0 14943 5 1 1 14942
0 14944 7 1 2 57671 77745
0 14945 5 2 1 14944
0 14946 7 4 2 59109 74095
0 14947 5 1 1 86175
0 14948 7 1 2 74083 14947
0 14949 7 1 2 86173 14948
0 14950 5 1 1 14949
0 14951 7 1 2 65014 14950
0 14952 5 1 1 14951
0 14953 7 1 2 69321 80127
0 14954 5 1 1 14953
0 14955 7 1 2 69736 76563
0 14956 5 1 1 14955
0 14957 7 1 2 14954 14956
0 14958 7 1 2 14952 14957
0 14959 5 1 1 14958
0 14960 7 1 2 57390 14959
0 14961 5 1 1 14960
0 14962 7 2 2 68989 67655
0 14963 5 1 1 86179
0 14964 7 1 2 67102 14963
0 14965 7 1 2 14901 14964
0 14966 5 3 1 14965
0 14967 7 1 2 70290 86181
0 14968 5 1 1 14967
0 14969 7 1 2 68360 76365
0 14970 5 2 1 14969
0 14971 7 1 2 67738 70002
0 14972 5 2 1 14971
0 14973 7 1 2 65224 86186
0 14974 5 1 1 14973
0 14975 7 1 2 86184 14974
0 14976 5 1 1 14975
0 14977 7 1 2 64258 14976
0 14978 5 1 1 14977
0 14979 7 1 2 14968 14978
0 14980 7 1 2 14961 14979
0 14981 5 1 1 14980
0 14982 7 1 2 58264 14981
0 14983 5 1 1 14982
0 14984 7 1 2 14943 14983
0 14985 7 1 2 14936 14984
0 14986 5 1 1 14985
0 14987 7 1 2 65841 14986
0 14988 5 1 1 14987
0 14989 7 2 2 80326 82235
0 14990 5 1 1 86188
0 14991 7 3 2 58265 73614
0 14992 5 2 1 86190
0 14993 7 1 2 86189 86191
0 14994 5 1 1 14993
0 14995 7 3 2 65842 75001
0 14996 5 5 1 86195
0 14997 7 1 2 58969 72932
0 14998 7 2 2 86198 14997
0 14999 5 1 1 86203
0 15000 7 1 2 57391 86204
0 15001 5 1 1 15000
0 15002 7 6 2 65015 73615
0 15003 5 5 1 86205
0 15004 7 1 2 67310 68608
0 15005 7 1 2 86206 15004
0 15006 5 1 1 15005
0 15007 7 1 2 15001 15006
0 15008 5 1 1 15007
0 15009 7 1 2 58266 15008
0 15010 5 1 1 15009
0 15011 7 2 2 72280 86115
0 15012 5 1 1 86216
0 15013 7 1 2 86193 15012
0 15014 5 1 1 15013
0 15015 7 1 2 77442 15014
0 15016 5 1 1 15015
0 15017 7 1 2 15010 15016
0 15018 5 1 1 15017
0 15019 7 1 2 57672 15018
0 15020 5 1 1 15019
0 15021 7 1 2 78904 73616
0 15022 5 1 1 15021
0 15023 7 1 2 15020 15022
0 15024 5 1 1 15023
0 15025 7 1 2 71877 15024
0 15026 5 1 1 15025
0 15027 7 1 2 14994 15026
0 15028 7 1 2 14988 15027
0 15029 7 1 2 14883 15028
0 15030 5 1 1 15029
0 15031 7 1 2 86091 15030
0 15032 5 1 1 15031
0 15033 7 1 2 14783 15032
0 15034 5 1 1 15033
0 15035 7 1 2 63193 15034
0 15036 5 1 1 15035
0 15037 7 1 2 14752 15036
0 15038 5 1 1 15037
0 15039 7 1 2 61547 15038
0 15040 5 1 1 15039
0 15041 7 1 2 74684 84466
0 15042 5 1 1 15041
0 15043 7 1 2 59316 84839
0 15044 5 1 1 15043
0 15045 7 1 2 80905 15044
0 15046 5 1 1 15045
0 15047 7 1 2 57990 15046
0 15048 5 1 1 15047
0 15049 7 1 2 64015 85011
0 15050 5 1 1 15049
0 15051 7 1 2 58267 15050
0 15052 5 1 1 15051
0 15053 7 1 2 83404 81177
0 15054 5 1 1 15053
0 15055 7 1 2 15052 15054
0 15056 7 1 2 15048 15055
0 15057 5 1 1 15056
0 15058 7 1 2 65533 15057
0 15059 5 1 1 15058
0 15060 7 1 2 57392 80248
0 15061 5 1 1 15060
0 15062 7 1 2 76147 78192
0 15063 5 1 1 15062
0 15064 7 1 2 15061 15063
0 15065 5 1 1 15064
0 15066 7 1 2 71878 15065
0 15067 5 1 1 15066
0 15068 7 2 2 80237 80320
0 15069 5 2 1 86218
0 15070 7 1 2 78344 86220
0 15071 5 1 1 15070
0 15072 7 1 2 80241 15071
0 15073 5 1 1 15072
0 15074 7 1 2 15067 15073
0 15075 7 1 2 15059 15074
0 15076 5 1 1 15075
0 15077 7 1 2 59525 15076
0 15078 5 1 1 15077
0 15079 7 1 2 61219 15078
0 15080 5 1 1 15079
0 15081 7 1 2 65534 11100
0 15082 5 1 1 15081
0 15083 7 1 2 65843 15082
0 15084 7 1 2 83859 15083
0 15085 5 1 1 15084
0 15086 7 1 2 59526 15085
0 15087 5 1 1 15086
0 15088 7 1 2 60312 84825
0 15089 5 1 1 15088
0 15090 7 1 2 60539 84835
0 15091 5 1 1 15090
0 15092 7 1 2 15089 15091
0 15093 5 2 1 15092
0 15094 7 1 2 69714 86222
0 15095 5 1 1 15094
0 15096 7 1 2 64259 84813
0 15097 5 1 1 15096
0 15098 7 1 2 15095 15097
0 15099 5 1 1 15098
0 15100 7 1 2 67311 15099
0 15101 5 1 1 15100
0 15102 7 1 2 64260 73463
0 15103 5 1 1 15102
0 15104 7 1 2 86174 15103
0 15105 5 1 1 15104
0 15106 7 1 2 68767 15105
0 15107 5 1 1 15106
0 15108 7 1 2 64261 82472
0 15109 5 1 1 15108
0 15110 7 1 2 15107 15109
0 15111 5 1 1 15110
0 15112 7 1 2 65016 15111
0 15113 5 1 1 15112
0 15114 7 1 2 74143 78692
0 15115 7 1 2 76242 15114
0 15116 5 1 1 15115
0 15117 7 1 2 77741 15116
0 15118 5 1 1 15117
0 15119 7 1 2 68609 15118
0 15120 5 1 1 15119
0 15121 7 2 2 69985 70350
0 15122 5 1 1 86224
0 15123 7 1 2 15120 15122
0 15124 7 1 2 15113 15123
0 15125 5 1 1 15124
0 15126 7 1 2 70401 15125
0 15127 5 1 1 15126
0 15128 7 1 2 78929 70165
0 15129 5 2 1 15128
0 15130 7 1 2 69737 83861
0 15131 5 1 1 15130
0 15132 7 1 2 15131 9459
0 15133 5 1 1 15132
0 15134 7 1 2 59317 15133
0 15135 5 1 1 15134
0 15136 7 1 2 65225 79374
0 15137 5 1 1 15136
0 15138 7 1 2 15135 15137
0 15139 5 1 1 15138
0 15140 7 1 2 57991 15139
0 15141 5 1 1 15140
0 15142 7 1 2 86226 15141
0 15143 7 1 2 15127 15142
0 15144 7 1 2 15101 15143
0 15145 7 1 2 15087 15144
0 15146 5 1 1 15145
0 15147 7 1 2 15080 15146
0 15148 5 2 1 15147
0 15149 7 1 2 15042 86228
0 15150 5 1 1 15149
0 15151 7 1 2 58455 15150
0 15152 5 1 1 15151
0 15153 7 1 2 79046 83857
0 15154 5 1 1 15153
0 15155 7 1 2 15152 15154
0 15156 5 1 1 15155
0 15157 7 1 2 63478 15156
0 15158 5 1 1 15157
0 15159 7 1 2 79869 15158
0 15160 5 1 1 15159
0 15161 7 1 2 73167 83544
0 15162 5 1 1 15161
0 15163 7 1 2 62366 15162
0 15164 5 1 1 15163
0 15165 7 1 2 70199 84392
0 15166 5 1 1 15165
0 15167 7 2 2 68492 75394
0 15168 5 1 1 86230
0 15169 7 1 2 60540 86231
0 15170 5 1 1 15169
0 15171 7 1 2 70254 15170
0 15172 7 1 2 15166 15171
0 15173 7 1 2 15164 15172
0 15174 5 1 1 15173
0 15175 7 1 2 65844 15174
0 15176 5 1 1 15175
0 15177 7 11 2 65535 74330
0 15178 7 5 2 61220 67739
0 15179 5 2 1 86243
0 15180 7 1 2 86232 86244
0 15181 5 1 1 15180
0 15182 7 1 2 15176 15181
0 15183 5 1 1 15182
0 15184 7 1 2 62643 15183
0 15185 5 1 1 15184
0 15186 7 1 2 68361 81947
0 15187 5 1 1 15186
0 15188 7 1 2 67848 81967
0 15189 5 1 1 15188
0 15190 7 1 2 77714 76784
0 15191 7 1 2 15189 15190
0 15192 7 1 2 15187 15191
0 15193 5 1 1 15192
0 15194 7 1 2 60866 15193
0 15195 5 1 1 15194
0 15196 7 1 2 68922 74783
0 15197 5 1 1 15196
0 15198 7 1 2 15195 15197
0 15199 5 1 1 15198
0 15200 7 1 2 61221 15199
0 15201 5 1 1 15200
0 15202 7 1 2 15185 15201
0 15203 5 1 1 15202
0 15204 7 1 2 64262 15203
0 15205 5 1 1 15204
0 15206 7 1 2 83845 79995
0 15207 5 1 1 15206
0 15208 7 1 2 62923 77063
0 15209 5 1 1 15208
0 15210 7 2 2 58268 79368
0 15211 5 3 1 86250
0 15212 7 1 2 70023 86252
0 15213 5 1 1 15212
0 15214 7 1 2 15209 15213
0 15215 5 1 1 15214
0 15216 7 1 2 62367 15215
0 15217 5 1 1 15216
0 15218 7 1 2 15207 15217
0 15219 5 1 1 15218
0 15220 7 1 2 65845 15219
0 15221 5 1 1 15220
0 15222 7 1 2 84617 75141
0 15223 5 2 1 15222
0 15224 7 1 2 15221 86255
0 15225 7 1 2 15205 15224
0 15226 5 1 1 15225
0 15227 7 1 2 73588 15226
0 15228 5 1 1 15227
0 15229 7 1 2 76177 76523
0 15230 5 1 1 15229
0 15231 7 3 2 76450 81667
0 15232 5 1 1 86257
0 15233 7 1 2 58269 15232
0 15234 5 1 1 15233
0 15235 7 1 2 71803 15234
0 15236 5 1 1 15235
0 15237 7 1 2 15230 15236
0 15238 5 1 1 15237
0 15239 7 1 2 62368 15238
0 15240 5 1 1 15239
0 15241 7 1 2 62924 81321
0 15242 5 1 1 15241
0 15243 7 1 2 15240 15242
0 15244 7 1 2 81866 15243
0 15245 5 1 1 15244
0 15246 7 1 2 73040 15245
0 15247 5 1 1 15246
0 15248 7 1 2 65846 84752
0 15249 5 1 1 15248
0 15250 7 1 2 15247 15249
0 15251 7 1 2 15228 15250
0 15252 5 1 1 15251
0 15253 7 1 2 63194 15252
0 15254 5 1 1 15253
0 15255 7 6 2 62925 72857
0 15256 5 7 1 86260
0 15257 7 2 2 82122 86261
0 15258 5 1 1 86273
0 15259 7 1 2 58456 86274
0 15260 5 1 1 15259
0 15261 7 1 2 77028 78511
0 15262 5 1 1 15261
0 15263 7 1 2 65847 77960
0 15264 5 4 1 15263
0 15265 7 1 2 85994 81316
0 15266 7 1 2 86275 15265
0 15267 5 1 1 15266
0 15268 7 1 2 15262 15267
0 15269 5 1 1 15268
0 15270 7 1 2 67165 15269
0 15271 5 1 1 15270
0 15272 7 1 2 77029 77004
0 15273 7 1 2 86262 15272
0 15274 5 1 1 15273
0 15275 7 1 2 15271 15274
0 15276 5 1 1 15275
0 15277 7 1 2 80928 15276
0 15278 5 1 1 15277
0 15279 7 1 2 15260 15278
0 15280 5 1 1 15279
0 15281 7 1 2 62369 15280
0 15282 5 1 1 15281
0 15283 7 2 2 61222 69385
0 15284 7 5 2 58457 63859
0 15285 7 1 2 79193 86281
0 15286 7 1 2 86279 15285
0 15287 5 1 1 15286
0 15288 7 1 2 66799 15287
0 15289 7 1 2 15282 15288
0 15290 7 1 2 15254 15289
0 15291 5 1 1 15290
0 15292 7 1 2 66159 69523
0 15293 7 1 2 15291 15292
0 15294 7 1 2 15160 15293
0 15295 5 1 1 15294
0 15296 7 1 2 15040 15295
0 15297 5 1 1 15296
0 15298 7 1 2 64494 15297
0 15299 5 1 1 15298
0 15300 7 14 2 59527 81036
0 15301 5 1 1 86286
0 15302 7 1 2 75850 86287
0 15303 7 1 2 81346 15302
0 15304 7 1 2 83979 15303
0 15305 5 1 1 15304
0 15306 7 8 2 66160 79878
0 15307 7 1 2 84187 86300
0 15308 7 1 2 84464 15307
0 15309 5 1 1 15308
0 15310 7 1 2 15305 15309
0 15311 5 1 1 15310
0 15312 7 1 2 60313 15311
0 15313 5 1 1 15312
0 15314 7 3 2 65017 70034
0 15315 5 1 1 86308
0 15316 7 10 2 57992 58458
0 15317 7 4 2 86311 72830
0 15318 7 11 2 64689 61548
0 15319 5 1 1 86325
0 15320 7 1 2 78523 86326
0 15321 7 1 2 75806 15320
0 15322 7 1 2 86321 15321
0 15323 7 1 2 86309 15322
0 15324 5 1 1 15323
0 15325 7 1 2 15313 15324
0 15326 5 1 1 15325
0 15327 7 1 2 73245 15326
0 15328 5 1 1 15327
0 15329 7 1 2 65536 85749
0 15330 5 1 1 15329
0 15331 7 2 2 84806 83135
0 15332 5 1 1 86336
0 15333 7 1 2 15330 15332
0 15334 5 1 1 15333
0 15335 7 1 2 74685 15334
0 15336 5 1 1 15335
0 15337 7 1 2 86229 15336
0 15338 5 1 1 15337
0 15339 7 1 2 63195 15338
0 15340 5 1 1 15339
0 15341 7 1 2 74978 4949
0 15342 5 1 1 15341
0 15343 7 1 2 68768 68362
0 15344 5 5 1 15343
0 15345 7 1 2 86338 82148
0 15346 5 1 1 15345
0 15347 7 1 2 65018 76266
0 15348 7 1 2 15346 15347
0 15349 5 1 1 15348
0 15350 7 1 2 15342 15349
0 15351 5 1 1 15350
0 15352 7 1 2 65226 15351
0 15353 5 1 1 15352
0 15354 7 1 2 75225 2804
0 15355 5 1 1 15354
0 15356 7 1 2 57393 15355
0 15357 5 1 1 15356
0 15358 7 1 2 79111 74368
0 15359 5 1 1 15358
0 15360 7 1 2 15357 15359
0 15361 5 1 1 15360
0 15362 7 1 2 57993 15361
0 15363 5 1 1 15362
0 15364 7 1 2 81938 83752
0 15365 5 1 1 15364
0 15366 7 1 2 57394 15365
0 15367 5 1 1 15366
0 15368 7 3 2 57994 69801
0 15369 5 3 1 86343
0 15370 7 1 2 74369 86344
0 15371 5 1 1 15370
0 15372 7 1 2 15367 15371
0 15373 5 1 1 15372
0 15374 7 1 2 57673 15373
0 15375 5 1 1 15374
0 15376 7 1 2 77715 15375
0 15377 7 1 2 15363 15376
0 15378 5 1 1 15377
0 15379 7 1 2 60867 15378
0 15380 5 1 1 15379
0 15381 7 1 2 15353 15380
0 15382 5 1 1 15381
0 15383 7 1 2 61223 15382
0 15384 5 1 1 15383
0 15385 7 2 2 74331 73617
0 15386 5 4 1 86349
0 15387 7 1 2 86116 75087
0 15388 5 1 1 15387
0 15389 7 1 2 86351 15388
0 15390 5 1 1 15389
0 15391 7 1 2 62644 15390
0 15392 5 1 1 15391
0 15393 7 1 2 62926 84626
0 15394 5 1 1 15393
0 15395 7 1 2 15392 15394
0 15396 5 1 1 15395
0 15397 7 1 2 67740 15396
0 15398 5 1 1 15397
0 15399 7 1 2 84247 84390
0 15400 5 1 1 15399
0 15401 7 1 2 76178 15400
0 15402 5 1 1 15401
0 15403 7 1 2 70200 77422
0 15404 5 1 1 15403
0 15405 7 1 2 74870 84239
0 15406 7 1 2 76487 15405
0 15407 5 1 1 15406
0 15408 7 1 2 15404 15407
0 15409 7 1 2 15402 15408
0 15410 5 1 1 15409
0 15411 7 1 2 65848 15410
0 15412 5 1 1 15411
0 15413 7 1 2 15398 15412
0 15414 7 1 2 15384 15413
0 15415 5 1 1 15414
0 15416 7 1 2 58459 15415
0 15417 5 1 1 15416
0 15418 7 1 2 80453 82441
0 15419 7 1 2 75238 15418
0 15420 5 1 1 15419
0 15421 7 1 2 15417 15420
0 15422 5 1 1 15421
0 15423 7 1 2 64263 15422
0 15424 5 1 1 15423
0 15425 7 1 2 58460 69386
0 15426 5 3 1 15425
0 15427 7 1 2 62370 74925
0 15428 7 1 2 86233 15427
0 15429 5 1 1 15428
0 15430 7 1 2 86355 15429
0 15431 5 1 1 15430
0 15432 7 1 2 68493 15431
0 15433 5 1 1 15432
0 15434 7 1 2 81845 83850
0 15435 5 1 1 15434
0 15436 7 1 2 58461 15435
0 15437 5 1 1 15436
0 15438 7 1 2 15433 15437
0 15439 5 1 1 15438
0 15440 7 1 2 65849 15439
0 15441 5 1 1 15440
0 15442 7 1 2 80554 86234
0 15443 5 1 1 15442
0 15444 7 1 2 15441 15443
0 15445 5 1 1 15444
0 15446 7 1 2 64016 15445
0 15447 5 1 1 15446
0 15448 7 1 2 58462 73041
0 15449 7 1 2 82007 15448
0 15450 5 1 1 15449
0 15451 7 1 2 15447 15450
0 15452 5 1 1 15451
0 15453 7 1 2 62645 15452
0 15454 5 1 1 15453
0 15455 7 1 2 72078 73042
0 15456 5 1 1 15455
0 15457 7 2 2 71676 86276
0 15458 5 1 1 86358
0 15459 7 1 2 62170 72893
0 15460 7 1 2 86359 15459
0 15461 5 2 1 15460
0 15462 7 1 2 15456 86360
0 15463 5 1 1 15462
0 15464 7 1 2 62371 15463
0 15465 5 1 1 15464
0 15466 7 3 2 78524 85793
0 15467 5 1 1 86362
0 15468 7 2 2 63860 86363
0 15469 5 1 1 86365
0 15470 7 1 2 15465 15469
0 15471 5 1 1 15470
0 15472 7 1 2 58463 15471
0 15473 5 1 1 15472
0 15474 7 1 2 15454 15473
0 15475 5 1 1 15474
0 15476 7 1 2 62927 15475
0 15477 5 1 1 15476
0 15478 7 4 2 59528 80416
0 15479 5 4 1 86367
0 15480 7 1 2 86361 86371
0 15481 5 1 1 15480
0 15482 7 1 2 67166 15481
0 15483 5 1 1 15482
0 15484 7 2 2 74926 86086
0 15485 5 1 1 86375
0 15486 7 1 2 80929 86376
0 15487 5 1 1 15486
0 15488 7 1 2 15483 15487
0 15489 5 1 1 15488
0 15490 7 1 2 62372 15489
0 15491 5 1 1 15490
0 15492 7 1 2 70734 86364
0 15493 5 1 1 15492
0 15494 7 1 2 15491 15493
0 15495 5 1 1 15494
0 15496 7 1 2 58464 15495
0 15497 5 1 1 15496
0 15498 7 1 2 66161 15497
0 15499 7 1 2 15477 15498
0 15500 7 1 2 15424 15499
0 15501 7 1 2 15340 15500
0 15502 5 1 1 15501
0 15503 7 1 2 59529 83796
0 15504 5 1 1 15503
0 15505 7 1 2 67849 84333
0 15506 5 1 1 15505
0 15507 7 1 2 64264 77659
0 15508 7 1 2 84325 15507
0 15509 7 1 2 15506 15508
0 15510 5 1 1 15509
0 15511 7 1 2 65537 15510
0 15512 7 1 2 15504 15511
0 15513 5 1 1 15512
0 15514 7 1 2 59530 9405
0 15515 5 1 1 15514
0 15516 7 1 2 80107 83221
0 15517 5 2 1 15516
0 15518 7 1 2 12782 86377
0 15519 7 1 2 15515 15518
0 15520 5 1 1 15519
0 15521 7 1 2 60868 15520
0 15522 5 1 1 15521
0 15523 7 1 2 69189 86176
0 15524 5 1 1 15523
0 15525 7 1 2 15522 15524
0 15526 7 1 2 15513 15525
0 15527 5 1 1 15526
0 15528 7 1 2 65850 15527
0 15529 5 1 1 15528
0 15530 7 1 2 78635 74743
0 15531 5 1 1 15530
0 15532 7 1 2 68769 85652
0 15533 7 1 2 86199 15532
0 15534 5 1 1 15533
0 15535 7 1 2 15531 15534
0 15536 5 1 1 15535
0 15537 7 1 2 73401 15536
0 15538 5 1 1 15537
0 15539 7 1 2 85969 72958
0 15540 5 1 1 15539
0 15541 7 1 2 15538 15540
0 15542 5 1 1 15541
0 15543 7 1 2 68363 15542
0 15544 5 1 1 15543
0 15545 7 1 2 71481 86099
0 15546 5 1 1 15545
0 15547 7 1 2 70056 83762
0 15548 5 1 1 15547
0 15549 7 1 2 15546 15548
0 15550 5 1 1 15549
0 15551 7 1 2 65538 15550
0 15552 5 1 1 15551
0 15553 7 1 2 81171 81958
0 15554 5 1 1 15553
0 15555 7 4 2 57995 71169
0 15556 5 1 1 86379
0 15557 7 1 2 15554 15556
0 15558 7 1 2 15552 15557
0 15559 5 1 1 15558
0 15560 7 1 2 61224 15559
0 15561 5 1 1 15560
0 15562 7 1 2 15544 15561
0 15563 7 1 2 15529 15562
0 15564 5 1 1 15563
0 15565 7 1 2 59318 15564
0 15566 5 1 1 15565
0 15567 7 1 2 74479 10844
0 15568 5 1 1 15567
0 15569 7 1 2 62928 12910
0 15570 5 3 1 15569
0 15571 7 1 2 71879 86383
0 15572 5 1 1 15571
0 15573 7 1 2 57996 70775
0 15574 5 2 1 15573
0 15575 7 1 2 62929 86386
0 15576 5 1 1 15575
0 15577 7 1 2 78312 15576
0 15578 5 1 1 15577
0 15579 7 2 2 71598 15578
0 15580 5 1 1 86388
0 15581 7 1 2 15572 86389
0 15582 5 2 1 15581
0 15583 7 1 2 61225 86390
0 15584 5 1 1 15583
0 15585 7 1 2 15568 15584
0 15586 5 1 1 15585
0 15587 7 1 2 65539 15586
0 15588 5 1 1 15587
0 15589 7 3 2 61226 71730
0 15590 7 1 2 77690 86392
0 15591 5 1 1 15590
0 15592 7 1 2 65851 76564
0 15593 7 1 2 75108 15592
0 15594 5 1 1 15593
0 15595 7 1 2 15591 15594
0 15596 5 1 1 15595
0 15597 7 1 2 65540 15596
0 15598 5 1 1 15597
0 15599 7 1 2 73246 69322
0 15600 5 2 1 15599
0 15601 7 1 2 61227 81523
0 15602 5 1 1 15601
0 15603 7 1 2 86395 15602
0 15604 5 1 1 15603
0 15605 7 1 2 80194 15604
0 15606 5 1 1 15605
0 15607 7 1 2 65852 74516
0 15608 7 1 2 75311 15607
0 15609 5 1 1 15608
0 15610 7 1 2 15606 15609
0 15611 7 1 2 15598 15610
0 15612 5 1 1 15611
0 15613 7 1 2 57395 15612
0 15614 5 1 1 15613
0 15615 7 1 2 71880 78219
0 15616 5 1 1 15615
0 15617 7 2 2 73897 78313
0 15618 5 1 1 86397
0 15619 7 1 2 15616 15618
0 15620 5 2 1 15619
0 15621 7 1 2 61228 86399
0 15622 5 1 1 15621
0 15623 7 1 2 86135 15622
0 15624 5 1 1 15623
0 15625 7 1 2 58270 15624
0 15626 5 1 1 15625
0 15627 7 4 2 60541 73247
0 15628 5 1 1 86401
0 15629 7 1 2 68990 67850
0 15630 5 1 1 15629
0 15631 7 1 2 77660 15630
0 15632 5 1 1 15631
0 15633 7 1 2 86402 15632
0 15634 5 1 1 15633
0 15635 7 1 2 15626 15634
0 15636 7 1 2 15614 15635
0 15637 7 1 2 15588 15636
0 15638 5 1 1 15637
0 15639 7 1 2 59531 15638
0 15640 5 1 1 15639
0 15641 7 1 2 65541 71632
0 15642 5 1 1 15641
0 15643 7 1 2 84359 15642
0 15644 5 1 1 15643
0 15645 7 1 2 64265 15644
0 15646 5 1 1 15645
0 15647 7 5 2 65019 70291
0 15648 7 1 2 68610 86405
0 15649 5 1 1 15648
0 15650 7 1 2 74103 15649
0 15651 5 1 1 15650
0 15652 7 1 2 67851 15651
0 15653 5 1 1 15652
0 15654 7 1 2 70292 77651
0 15655 5 1 1 15654
0 15656 7 1 2 60869 7212
0 15657 5 1 1 15656
0 15658 7 1 2 57997 74144
0 15659 7 1 2 15657 15658
0 15660 5 1 1 15659
0 15661 7 1 2 15655 15660
0 15662 7 1 2 15653 15661
0 15663 7 1 2 15646 15662
0 15664 5 1 1 15663
0 15665 7 1 2 65853 15664
0 15666 5 1 1 15665
0 15667 7 1 2 80398 77753
0 15668 5 1 1 15667
0 15669 7 1 2 76327 78843
0 15670 7 1 2 86393 15669
0 15671 5 1 1 15670
0 15672 7 1 2 86162 15671
0 15673 5 1 1 15672
0 15674 7 1 2 75870 15673
0 15675 5 1 1 15674
0 15676 7 1 2 15668 15675
0 15677 7 1 2 15666 15676
0 15678 5 1 1 15677
0 15679 7 1 2 58271 15678
0 15680 5 1 1 15679
0 15681 7 1 2 77519 73305
0 15682 7 1 2 86171 15681
0 15683 5 1 1 15682
0 15684 7 1 2 15680 15683
0 15685 7 1 2 15640 15684
0 15686 7 1 2 15566 15685
0 15687 5 1 1 15686
0 15688 7 1 2 58465 15687
0 15689 5 1 1 15688
0 15690 7 1 2 73799 68925
0 15691 5 1 1 15690
0 15692 7 1 2 57674 15691
0 15693 5 1 1 15692
0 15694 7 1 2 60870 69886
0 15695 5 4 1 15694
0 15696 7 1 2 59319 86410
0 15697 5 1 1 15696
0 15698 7 1 2 15693 15697
0 15699 5 1 1 15698
0 15700 7 1 2 74014 15699
0 15701 5 1 1 15700
0 15702 7 1 2 83405 86406
0 15703 5 1 1 15702
0 15704 7 1 2 15701 15703
0 15705 5 1 1 15704
0 15706 7 1 2 57998 15705
0 15707 5 1 1 15706
0 15708 7 1 2 81227 15707
0 15709 5 1 1 15708
0 15710 7 1 2 68611 15709
0 15711 5 1 1 15710
0 15712 7 1 2 73872 83738
0 15713 5 1 1 15712
0 15714 7 1 2 63861 74370
0 15715 5 1 1 15714
0 15716 7 1 2 65542 15715
0 15717 5 1 1 15716
0 15718 7 1 2 76247 15717
0 15719 5 1 1 15718
0 15720 7 1 2 68001 15719
0 15721 5 1 1 15720
0 15722 7 1 2 15713 15721
0 15723 5 1 1 15722
0 15724 7 1 2 63196 15723
0 15725 5 1 1 15724
0 15726 7 1 2 60314 80233
0 15727 5 1 1 15726
0 15728 7 1 2 74200 15727
0 15729 5 1 1 15728
0 15730 7 1 2 59320 77443
0 15731 7 1 2 15729 15730
0 15732 5 1 1 15731
0 15733 7 1 2 15725 15732
0 15734 7 1 2 15711 15733
0 15735 5 1 1 15734
0 15736 7 1 2 79047 15735
0 15737 5 1 1 15736
0 15738 7 1 2 61549 15737
0 15739 7 1 2 15689 15738
0 15740 5 1 1 15739
0 15741 7 1 2 63479 15740
0 15742 7 1 2 15502 15741
0 15743 5 1 1 15742
0 15744 7 1 2 79870 15743
0 15745 5 1 1 15744
0 15746 7 1 2 64266 12553
0 15747 5 1 1 15746
0 15748 7 2 2 71654 71780
0 15749 5 1 1 86414
0 15750 7 1 2 84866 86415
0 15751 5 1 1 15750
0 15752 7 1 2 61229 15751
0 15753 7 1 2 86009 15752
0 15754 7 1 2 15747 15753
0 15755 5 1 1 15754
0 15756 7 2 2 62646 69980
0 15757 5 2 1 86416
0 15758 7 1 2 12580 86418
0 15759 5 1 1 15758
0 15760 7 1 2 64267 15759
0 15761 5 1 1 15760
0 15762 7 5 2 62930 75395
0 15763 5 1 1 86420
0 15764 7 1 2 63862 86421
0 15765 5 1 1 15764
0 15766 7 1 2 15761 15765
0 15767 5 1 1 15766
0 15768 7 1 2 60871 15767
0 15769 5 1 1 15768
0 15770 7 1 2 70910 84715
0 15771 5 1 1 15770
0 15772 7 1 2 73589 15771
0 15773 5 1 1 15772
0 15774 7 2 2 60872 81850
0 15775 5 1 1 86425
0 15776 7 1 2 4868 15775
0 15777 5 1 1 15776
0 15778 7 1 2 68494 15777
0 15779 5 1 1 15778
0 15780 7 1 2 15773 15779
0 15781 7 1 2 15769 15780
0 15782 5 1 1 15781
0 15783 7 1 2 62373 15782
0 15784 5 1 1 15783
0 15785 7 1 2 65543 75406
0 15786 5 3 1 15785
0 15787 7 1 2 63863 86427
0 15788 5 1 1 15787
0 15789 7 1 2 83572 15788
0 15790 5 1 1 15789
0 15791 7 1 2 60542 15790
0 15792 5 1 1 15791
0 15793 7 2 2 64017 74979
0 15794 5 3 1 86430
0 15795 7 1 2 70255 86432
0 15796 7 1 2 15792 15795
0 15797 5 1 1 15796
0 15798 7 1 2 64268 15797
0 15799 5 1 1 15798
0 15800 7 1 2 60873 86422
0 15801 5 1 1 15800
0 15802 7 1 2 15799 15801
0 15803 5 1 1 15802
0 15804 7 1 2 62647 15803
0 15805 5 1 1 15804
0 15806 7 1 2 73590 84120
0 15807 5 1 1 15806
0 15808 7 1 2 65854 15807
0 15809 7 1 2 15805 15808
0 15810 7 1 2 15784 15809
0 15811 5 1 1 15810
0 15812 7 1 2 63197 15811
0 15813 7 1 2 15755 15812
0 15814 5 1 1 15813
0 15815 7 1 2 84534 15814
0 15816 5 1 1 15815
0 15817 7 1 2 61550 15816
0 15818 5 1 1 15817
0 15819 7 2 2 63198 84647
0 15820 7 5 2 64018 77978
0 15821 5 3 1 86437
0 15822 7 2 2 77423 86438
0 15823 5 2 1 86445
0 15824 7 1 2 67167 78030
0 15825 5 1 1 15824
0 15826 7 1 2 71398 77945
0 15827 5 1 1 15826
0 15828 7 1 2 15825 15827
0 15829 5 1 1 15828
0 15830 7 1 2 80930 15829
0 15831 5 1 1 15830
0 15832 7 1 2 86447 15831
0 15833 5 1 1 15832
0 15834 7 1 2 62374 15833
0 15835 5 1 1 15834
0 15836 7 1 2 77909 84121
0 15837 5 1 1 15836
0 15838 7 1 2 15835 15837
0 15839 5 1 1 15838
0 15840 7 1 2 86435 15839
0 15841 5 1 1 15840
0 15842 7 1 2 66800 15841
0 15843 7 1 2 15818 15842
0 15844 5 1 1 15843
0 15845 7 1 2 59770 15844
0 15846 7 1 2 15745 15845
0 15847 5 1 1 15846
0 15848 7 1 2 15328 15847
0 15849 5 1 1 15848
0 15850 7 1 2 69524 15849
0 15851 5 1 1 15850
0 15852 7 1 2 15299 15851
0 15853 5 1 1 15852
0 15854 7 1 2 67466 15853
0 15855 5 1 1 15854
0 15856 7 2 2 14640 15855
0 15857 5 1 1 86449
0 15858 7 60 2 65855 61551
0 15859 5 6 1 86451
0 15860 7 2 2 63864 67040
0 15861 5 2 1 86517
0 15862 7 1 2 86452 86518
0 15863 5 1 1 15862
0 15864 7 5 2 66567 84648
0 15865 7 2 2 70904 72105
0 15866 7 1 2 86521 86526
0 15867 5 1 1 15866
0 15868 7 1 2 15863 15867
0 15869 5 1 1 15868
0 15870 7 1 2 62648 15869
0 15871 5 1 1 15870
0 15872 7 1 2 74436 81024
0 15873 5 1 1 15872
0 15874 7 6 2 62931 66960
0 15875 5 3 1 86528
0 15876 7 1 2 63865 86529
0 15877 5 1 1 15876
0 15878 7 1 2 15873 15877
0 15879 5 1 1 15878
0 15880 7 1 2 86453 15879
0 15881 5 1 1 15880
0 15882 7 1 2 15871 15881
0 15883 5 1 1 15882
0 15884 7 1 2 63600 15883
0 15885 5 1 1 15884
0 15886 7 1 2 75002 2435
0 15887 5 3 1 15886
0 15888 7 3 2 61912 86537
0 15889 7 1 2 70450 86454
0 15890 7 1 2 86540 15889
0 15891 5 1 1 15890
0 15892 7 1 2 15885 15891
0 15893 5 1 1 15892
0 15894 7 1 2 77852 15893
0 15895 5 1 1 15894
0 15896 7 1 2 58272 75940
0 15897 5 1 1 15896
0 15898 7 6 2 63199 63866
0 15899 7 2 2 86543 79930
0 15900 7 25 2 65856 66162
0 15901 5 1 1 86551
0 15902 7 1 2 86552 66961
0 15903 7 1 2 86549 15902
0 15904 7 1 2 15897 15903
0 15905 5 1 1 15904
0 15906 7 1 2 15895 15905
0 15907 5 1 1 15906
0 15908 7 1 2 64269 15907
0 15909 5 1 1 15908
0 15910 7 10 2 62932 59771
0 15911 7 2 2 86455 86576
0 15912 5 1 1 86586
0 15913 7 1 2 70487 86587
0 15914 7 1 2 86541 15913
0 15915 5 1 1 15914
0 15916 7 3 2 60874 72894
0 15917 7 4 2 78996 86588
0 15918 7 4 2 64495 84171
0 15919 5 1 1 86595
0 15920 7 1 2 86596 84539
0 15921 7 1 2 86591 15920
0 15922 5 1 1 15921
0 15923 7 1 2 15915 15922
0 15924 5 1 1 15923
0 15925 7 1 2 63200 15924
0 15926 5 1 1 15925
0 15927 7 1 2 15909 15926
0 15928 5 1 1 15927
0 15929 7 1 2 66893 15928
0 15930 5 1 1 15929
0 15931 7 4 2 63201 77891
0 15932 7 3 2 61552 73360
0 15933 7 2 2 61913 79970
0 15934 7 2 2 86603 86606
0 15935 7 1 2 86599 86608
0 15936 5 1 1 15935
0 15937 7 6 2 66163 66568
0 15938 7 2 2 65857 86610
0 15939 7 1 2 74980 86616
0 15940 7 4 2 64792 80457
0 15941 7 1 2 86618 79036
0 15942 7 1 2 15939 15941
0 15943 5 1 1 15942
0 15944 7 1 2 15936 15943
0 15945 5 1 1 15944
0 15946 7 1 2 62933 15945
0 15947 5 1 1 15946
0 15948 7 3 2 65858 77892
0 15949 5 1 1 86622
0 15950 7 1 2 59532 85794
0 15951 5 3 1 15950
0 15952 7 1 2 15949 86625
0 15953 5 2 1 15952
0 15954 7 2 2 66569 81385
0 15955 7 1 2 85677 79187
0 15956 7 1 2 86630 15955
0 15957 7 1 2 86628 15956
0 15958 5 1 1 15957
0 15959 7 1 2 15947 15958
0 15960 5 1 1 15959
0 15961 7 1 2 62649 15960
0 15962 5 1 1 15961
0 15963 7 4 2 60315 85495
0 15964 5 1 1 86632
0 15965 7 1 2 86609 86633
0 15966 5 1 1 15965
0 15967 7 2 2 79297 86617
0 15968 7 6 2 63867 59772
0 15969 7 3 2 58466 86638
0 15970 7 1 2 79231 86644
0 15971 7 1 2 86636 15970
0 15972 5 1 1 15971
0 15973 7 1 2 15966 15972
0 15974 5 1 1 15973
0 15975 7 1 2 71399 15974
0 15976 5 1 1 15975
0 15977 7 1 2 15962 15976
0 15978 7 1 2 15930 15977
0 15979 5 1 1 15978
0 15980 7 1 2 62055 15979
0 15981 5 1 1 15980
0 15982 7 8 2 61553 80417
0 15983 7 3 2 67517 86647
0 15984 7 3 2 84872 77394
0 15985 7 1 2 86658 79232
0 15986 7 2 2 86655 15985
0 15987 7 17 2 64496 64690
0 15988 5 3 1 86663
0 15989 7 3 2 72106 86664
0 15990 7 1 2 84263 86683
0 15991 7 1 2 86661 15990
0 15992 5 1 1 15991
0 15993 7 1 2 15981 15992
0 15994 5 1 1 15993
0 15995 7 1 2 70983 15994
0 15996 5 1 1 15995
0 15997 7 1 2 86450 15996
0 15998 5 1 1 15997
0 15999 7 1 2 61762 15998
0 16000 5 1 1 15999
0 16001 7 1 2 85685 86006
0 16002 5 1 1 16001
0 16003 7 1 2 84380 16002
0 16004 5 1 1 16003
0 16005 7 1 2 65859 16004
0 16006 5 1 1 16005
0 16007 7 1 2 64270 80953
0 16008 5 1 1 16007
0 16009 7 1 2 60316 75246
0 16010 5 1 1 16009
0 16011 7 1 2 73579 16010
0 16012 5 1 1 16011
0 16013 7 1 2 61230 16012
0 16014 7 1 2 16008 16013
0 16015 5 1 1 16014
0 16016 7 1 2 16006 16015
0 16017 5 1 1 16016
0 16018 7 1 2 66164 16017
0 16019 5 1 1 16018
0 16020 7 1 2 86456 78387
0 16021 5 1 1 16020
0 16022 7 1 2 16019 16021
0 16023 5 1 1 16022
0 16024 7 1 2 58467 16023
0 16025 5 1 1 16024
0 16026 7 4 2 64271 84649
0 16027 5 3 1 86686
0 16028 7 4 2 59533 86457
0 16029 5 9 1 86693
0 16030 7 1 2 86690 86697
0 16031 5 9 1 16030
0 16032 7 1 2 84938 86706
0 16033 5 1 1 16032
0 16034 7 21 2 63202 65860
0 16035 5 11 1 86715
0 16036 7 1 2 86716 81546
0 16037 5 1 1 16036
0 16038 7 1 2 16033 16037
0 16039 5 1 1 16038
0 16040 7 1 2 57396 16039
0 16041 5 1 1 16040
0 16042 7 2 2 66165 78314
0 16043 7 1 2 86717 86747
0 16044 5 1 1 16043
0 16045 7 1 2 16041 16044
0 16046 5 1 1 16045
0 16047 7 1 2 72241 16046
0 16048 5 1 1 16047
0 16049 7 3 2 66166 86718
0 16050 7 1 2 67168 77726
0 16051 5 1 1 16050
0 16052 7 1 2 86749 16051
0 16053 5 1 1 16052
0 16054 7 1 2 68002 86707
0 16055 7 1 2 78363 16054
0 16056 5 1 1 16055
0 16057 7 1 2 16053 16056
0 16058 5 1 1 16057
0 16059 7 1 2 71881 16058
0 16060 5 1 1 16059
0 16061 7 1 2 76090 86708
0 16062 7 1 2 78230 16061
0 16063 5 1 1 16062
0 16064 7 3 2 64019 75271
0 16065 5 1 1 86752
0 16066 7 1 2 62375 86753
0 16067 5 1 1 16066
0 16068 7 1 2 57999 86750
0 16069 7 1 2 16067 16068
0 16070 5 1 1 16069
0 16071 7 1 2 16063 16070
0 16072 7 1 2 16060 16071
0 16073 7 1 2 16048 16072
0 16074 5 1 1 16073
0 16075 7 1 2 58273 16074
0 16076 5 1 1 16075
0 16077 7 1 2 57675 72525
0 16078 7 1 2 75282 16077
0 16079 5 1 1 16078
0 16080 7 1 2 79713 16079
0 16081 5 1 1 16080
0 16082 7 1 2 71882 16081
0 16083 5 1 1 16082
0 16084 7 3 2 59321 73757
0 16085 5 1 1 86755
0 16086 7 3 2 59534 70776
0 16087 5 1 1 86758
0 16088 7 1 2 73280 16087
0 16089 5 1 1 16088
0 16090 7 1 2 82236 16089
0 16091 5 1 1 16090
0 16092 7 1 2 16085 16091
0 16093 7 1 2 16083 16092
0 16094 5 1 1 16093
0 16095 7 1 2 86751 16094
0 16096 5 1 1 16095
0 16097 7 1 2 60875 16096
0 16098 7 1 2 16076 16097
0 16099 7 1 2 16025 16098
0 16100 5 1 1 16099
0 16101 7 2 2 58274 69802
0 16102 5 2 1 86761
0 16103 7 1 2 69911 86763
0 16104 5 1 1 16103
0 16105 7 1 2 58000 16104
0 16106 5 1 1 16105
0 16107 7 2 2 69097 69807
0 16108 5 2 1 86765
0 16109 7 1 2 58275 86767
0 16110 5 1 1 16109
0 16111 7 1 2 16106 16110
0 16112 5 1 1 16111
0 16113 7 1 2 57676 16112
0 16114 5 1 1 16113
0 16115 7 1 2 68079 77532
0 16116 5 1 1 16115
0 16117 7 2 2 67312 16116
0 16118 5 2 1 86769
0 16119 7 2 2 58276 86770
0 16120 5 1 1 86773
0 16121 7 3 2 16114 16120
0 16122 5 1 1 86775
0 16123 7 1 2 63203 86776
0 16124 5 1 1 16123
0 16125 7 1 2 58468 80699
0 16126 5 1 1 16125
0 16127 7 1 2 16124 16126
0 16128 5 1 1 16127
0 16129 7 1 2 61554 16128
0 16130 5 1 1 16129
0 16131 7 3 2 68229 84979
0 16132 5 1 1 86778
0 16133 7 1 2 66167 16132
0 16134 5 1 1 16133
0 16135 7 1 2 59535 16134
0 16136 7 1 2 16130 16135
0 16137 5 1 1 16136
0 16138 7 1 2 67313 74035
0 16139 5 1 1 16138
0 16140 7 1 2 64020 80691
0 16141 5 1 1 16140
0 16142 7 2 2 57677 16141
0 16143 5 1 1 86781
0 16144 7 1 2 16139 16143
0 16145 5 1 1 16144
0 16146 7 1 2 57397 16145
0 16147 5 1 1 16146
0 16148 7 1 2 67901 16147
0 16149 5 1 1 16148
0 16150 7 1 2 81248 16149
0 16151 5 1 1 16150
0 16152 7 1 2 67314 83813
0 16153 5 1 1 16152
0 16154 7 2 2 68080 16153
0 16155 5 1 1 86783
0 16156 7 1 2 82868 16155
0 16157 5 1 1 16156
0 16158 7 2 2 66168 73976
0 16159 5 1 1 86785
0 16160 7 1 2 81267 16159
0 16161 5 1 1 16160
0 16162 7 1 2 67315 16161
0 16163 7 1 2 11076 16162
0 16164 5 1 1 16163
0 16165 7 1 2 61555 85023
0 16166 5 1 1 16165
0 16167 7 1 2 58277 81189
0 16168 7 1 2 16166 16167
0 16169 5 1 1 16168
0 16170 7 1 2 16164 16169
0 16171 7 1 2 16157 16170
0 16172 7 1 2 16151 16171
0 16173 5 1 1 16172
0 16174 7 1 2 64272 16173
0 16175 5 1 1 16174
0 16176 7 1 2 65861 16175
0 16177 7 1 2 16137 16176
0 16178 5 1 1 16177
0 16179 7 1 2 81190 86777
0 16180 5 1 1 16179
0 16181 7 1 2 59536 15168
0 16182 5 2 1 16181
0 16183 7 1 2 81152 86787
0 16184 5 1 1 16183
0 16185 7 5 2 60317 71259
0 16186 5 1 1 86789
0 16187 7 2 2 68495 86790
0 16188 5 2 1 86794
0 16189 7 1 2 81185 86796
0 16190 7 1 2 16184 16189
0 16191 5 1 1 16190
0 16192 7 8 2 63204 61556
0 16193 5 3 1 86798
0 16194 7 1 2 16191 86806
0 16195 7 1 2 16180 16194
0 16196 5 1 1 16195
0 16197 7 1 2 67316 69803
0 16198 5 3 1 16197
0 16199 7 1 2 62171 86809
0 16200 5 1 1 16199
0 16201 7 1 2 86782 16200
0 16202 5 1 1 16201
0 16203 7 2 2 86771 16202
0 16204 5 1 1 86812
0 16205 7 1 2 62934 86813
0 16206 5 2 1 16205
0 16207 7 1 2 85018 81426
0 16208 5 1 1 16207
0 16209 7 1 2 82891 16208
0 16210 5 1 1 16209
0 16211 7 1 2 59537 16210
0 16212 7 1 2 86814 16211
0 16213 5 1 1 16212
0 16214 7 1 2 61231 16213
0 16215 7 1 2 16196 16214
0 16216 5 1 1 16215
0 16217 7 1 2 65227 16216
0 16218 7 1 2 16178 16217
0 16219 5 1 1 16218
0 16220 7 1 2 84154 68612
0 16221 5 1 1 16220
0 16222 7 1 2 63205 16221
0 16223 5 1 1 16222
0 16224 7 1 2 67317 16223
0 16225 5 1 1 16224
0 16226 7 1 2 85289 76807
0 16227 5 1 1 16226
0 16228 7 1 2 16225 16227
0 16229 5 1 1 16228
0 16230 7 1 2 69387 16229
0 16231 5 1 1 16230
0 16232 7 2 2 58278 83772
0 16233 7 3 2 65020 86816
0 16234 5 1 1 86818
0 16235 7 1 2 63206 86819
0 16236 5 1 1 16235
0 16237 7 1 2 16231 16236
0 16238 5 1 1 16237
0 16239 7 1 2 61557 16238
0 16240 5 1 1 16239
0 16241 7 2 2 58469 81441
0 16242 5 3 1 86821
0 16243 7 1 2 59322 82869
0 16244 5 1 1 16243
0 16245 7 1 2 86823 16244
0 16246 5 1 1 16245
0 16247 7 1 2 62650 16246
0 16248 5 1 1 16247
0 16249 7 3 2 62172 66169
0 16250 7 5 2 63207 63760
0 16251 7 2 2 86826 86829
0 16252 5 1 1 86834
0 16253 7 1 2 74962 86835
0 16254 5 1 1 16253
0 16255 7 1 2 59538 16254
0 16256 7 1 2 16248 16255
0 16257 7 1 2 16240 16256
0 16258 5 1 1 16257
0 16259 7 7 2 57398 66170
0 16260 7 2 2 58970 86836
0 16261 7 1 2 63208 86843
0 16262 5 1 1 16261
0 16263 7 1 2 86824 16262
0 16264 5 1 1 16263
0 16265 7 1 2 67892 16264
0 16266 5 1 1 16265
0 16267 7 7 2 57399 58470
0 16268 7 4 2 58971 86845
0 16269 7 1 2 81347 86852
0 16270 7 1 2 82749 16269
0 16271 5 1 1 16270
0 16272 7 1 2 64273 16271
0 16273 7 1 2 16266 16272
0 16274 5 1 1 16273
0 16275 7 1 2 16258 16274
0 16276 5 1 1 16275
0 16277 7 1 2 77005 82674
0 16278 5 2 1 16277
0 16279 7 1 2 83681 81329
0 16280 5 1 1 16279
0 16281 7 1 2 86856 16280
0 16282 5 1 1 16281
0 16283 7 1 2 83775 16282
0 16284 5 1 1 16283
0 16285 7 1 2 71599 77929
0 16286 5 1 1 16285
0 16287 7 2 2 66171 72793
0 16288 5 1 1 86858
0 16289 7 1 2 16288 86857
0 16290 5 1 1 16289
0 16291 7 1 2 16286 16290
0 16292 5 1 1 16291
0 16293 7 4 2 58471 82675
0 16294 5 1 1 86860
0 16295 7 1 2 74963 86861
0 16296 5 1 1 16295
0 16297 7 1 2 69774 86786
0 16298 5 1 1 16297
0 16299 7 1 2 16296 16298
0 16300 5 1 1 16299
0 16301 7 1 2 58279 16300
0 16302 5 1 1 16301
0 16303 7 1 2 65862 16302
0 16304 7 1 2 16292 16303
0 16305 7 1 2 16284 16304
0 16306 7 1 2 16276 16305
0 16307 5 1 1 16306
0 16308 7 1 2 62651 84284
0 16309 5 1 1 16308
0 16310 7 1 2 62935 73814
0 16311 5 1 1 16310
0 16312 7 1 2 16309 16311
0 16313 5 2 1 16312
0 16314 7 1 2 58472 86864
0 16315 5 1 1 16314
0 16316 7 1 2 71260 10804
0 16317 5 1 1 16316
0 16318 7 1 2 63209 71482
0 16319 7 1 2 16317 16318
0 16320 5 1 1 16319
0 16321 7 1 2 16315 16320
0 16322 5 1 1 16321
0 16323 7 1 2 65021 16322
0 16324 5 1 1 16323
0 16325 7 1 2 58280 83583
0 16326 5 1 1 16325
0 16327 7 1 2 78170 16326
0 16328 5 1 1 16327
0 16329 7 1 2 68652 16328
0 16330 5 1 1 16329
0 16331 7 3 2 58473 84188
0 16332 5 1 1 86866
0 16333 7 1 2 60318 86867
0 16334 5 1 1 16333
0 16335 7 1 2 82906 16334
0 16336 5 1 1 16335
0 16337 7 3 2 77480 79210
0 16338 5 4 1 86869
0 16339 7 1 2 16336 86872
0 16340 5 1 1 16339
0 16341 7 1 2 16330 16340
0 16342 7 1 2 16324 16341
0 16343 5 1 1 16342
0 16344 7 1 2 66172 16343
0 16345 5 1 1 16344
0 16346 7 3 2 70922 69798
0 16347 5 7 1 86876
0 16348 7 1 2 82844 86879
0 16349 5 1 1 16348
0 16350 7 1 2 86037 16349
0 16351 5 1 1 16350
0 16352 7 2 2 71483 16351
0 16353 5 1 1 86886
0 16354 7 1 2 81249 86887
0 16355 5 1 1 16354
0 16356 7 1 2 61232 16355
0 16357 7 1 2 16345 16356
0 16358 5 1 1 16357
0 16359 7 1 2 16307 16358
0 16360 5 1 1 16359
0 16361 7 1 2 65544 16360
0 16362 7 1 2 16219 16361
0 16363 5 1 1 16362
0 16364 7 1 2 16100 16363
0 16365 5 1 1 16364
0 16366 7 1 2 59323 77185
0 16367 5 1 1 16366
0 16368 7 1 2 72388 80227
0 16369 5 5 1 16368
0 16370 7 1 2 16367 86888
0 16371 5 1 1 16370
0 16372 7 1 2 58001 16371
0 16373 5 1 1 16372
0 16374 7 1 2 16373 83149
0 16375 5 2 1 16374
0 16376 7 1 2 71484 86893
0 16377 5 1 1 16376
0 16378 7 1 2 67169 77172
0 16379 7 1 2 78898 16378
0 16380 5 1 1 16379
0 16381 7 1 2 71170 16380
0 16382 5 1 1 16381
0 16383 7 1 2 61233 16382
0 16384 7 1 2 16377 16383
0 16385 5 1 1 16384
0 16386 7 5 2 65863 71261
0 16387 5 2 1 86895
0 16388 7 1 2 86900 81250
0 16389 7 1 2 78943 16388
0 16390 7 1 2 16385 16389
0 16391 5 1 1 16390
0 16392 7 1 2 85468 83237
0 16393 5 1 1 16392
0 16394 7 1 2 80861 76896
0 16395 5 1 1 16394
0 16396 7 1 2 16393 16395
0 16397 5 1 1 16396
0 16398 7 1 2 65864 16397
0 16399 5 1 1 16398
0 16400 7 4 2 62652 77342
0 16401 7 2 2 85591 86902
0 16402 5 1 1 86906
0 16403 7 1 2 16399 16402
0 16404 5 1 1 16403
0 16405 7 1 2 58474 16404
0 16406 5 1 1 16405
0 16407 7 1 2 70402 81634
0 16408 5 1 1 16407
0 16409 7 1 2 58281 85957
0 16410 5 1 1 16409
0 16411 7 1 2 75170 70098
0 16412 5 5 1 16411
0 16413 7 2 2 16410 86908
0 16414 5 4 1 86913
0 16415 7 1 2 67318 86915
0 16416 5 1 1 16415
0 16417 7 9 2 59324 71585
0 16418 5 3 1 86919
0 16419 7 1 2 16416 86928
0 16420 7 1 2 16408 16419
0 16421 5 1 1 16420
0 16422 7 1 2 61234 78156
0 16423 7 1 2 16421 16422
0 16424 5 1 1 16423
0 16425 7 1 2 16406 16424
0 16426 5 1 1 16425
0 16427 7 1 2 66173 16426
0 16428 5 1 1 16427
0 16429 7 1 2 85083 85947
0 16430 5 1 1 16429
0 16431 7 1 2 85116 84499
0 16432 5 1 1 16431
0 16433 7 1 2 16430 16432
0 16434 5 1 1 16433
0 16435 7 1 2 66174 16434
0 16436 5 1 1 16435
0 16437 7 11 2 59539 60319
0 16438 5 2 1 86931
0 16439 7 8 2 61558 85543
0 16440 7 1 2 86932 86944
0 16441 5 1 1 16440
0 16442 7 1 2 16436 16441
0 16443 5 1 1 16442
0 16444 7 1 2 65228 16443
0 16445 5 1 1 16444
0 16446 7 3 2 60543 86553
0 16447 7 2 2 63210 72986
0 16448 7 1 2 86952 86955
0 16449 5 1 1 16448
0 16450 7 1 2 16445 16449
0 16451 5 1 1 16450
0 16452 7 1 2 65545 16451
0 16453 5 1 1 16452
0 16454 7 1 2 81186 78445
0 16455 7 1 2 84609 16454
0 16456 5 1 1 16455
0 16457 7 1 2 16453 16456
0 16458 5 1 1 16457
0 16459 7 1 2 67741 16458
0 16460 5 1 1 16459
0 16461 7 1 2 16428 16460
0 16462 7 1 2 16391 16461
0 16463 7 1 2 16365 16462
0 16464 5 1 1 16463
0 16465 7 1 2 59989 16464
0 16466 5 1 1 16465
0 16467 7 4 2 71171 82637
0 16468 5 1 1 86957
0 16469 7 1 2 66175 86958
0 16470 7 1 2 80753 16469
0 16471 5 1 1 16470
0 16472 7 1 2 16466 16471
0 16473 5 1 1 16472
0 16474 7 1 2 61914 16473
0 16475 5 1 1 16474
0 16476 7 1 2 64274 2593
0 16477 5 1 1 16476
0 16478 7 1 2 79408 77645
0 16479 5 1 1 16478
0 16480 7 1 2 62936 16479
0 16481 5 1 1 16480
0 16482 7 1 2 16477 16481
0 16483 5 1 1 16482
0 16484 7 1 2 61559 16483
0 16485 5 1 1 16484
0 16486 7 1 2 84450 84209
0 16487 5 1 1 16486
0 16488 7 1 2 16485 16487
0 16489 5 1 1 16488
0 16490 7 1 2 61235 16489
0 16491 5 1 1 16490
0 16492 7 3 2 71400 86458
0 16493 5 1 1 86961
0 16494 7 1 2 67170 86962
0 16495 5 1 1 16494
0 16496 7 1 2 16491 16495
0 16497 5 1 1 16496
0 16498 7 1 2 63211 16497
0 16499 5 1 1 16498
0 16500 7 1 2 79487 84650
0 16501 5 3 1 16500
0 16502 7 1 2 86511 86964
0 16503 5 1 1 16502
0 16504 7 1 2 63212 16503
0 16505 5 1 1 16504
0 16506 7 3 2 75432 84775
0 16507 5 1 1 86967
0 16508 7 1 2 16505 16507
0 16509 5 1 1 16508
0 16510 7 1 2 67171 16509
0 16511 5 1 1 16510
0 16512 7 3 2 65865 72794
0 16513 5 2 1 86970
0 16514 7 1 2 61560 86971
0 16515 5 1 1 16514
0 16516 7 1 2 16511 16515
0 16517 5 1 1 16516
0 16518 7 1 2 62937 16517
0 16519 5 1 1 16518
0 16520 7 4 2 63213 64021
0 16521 7 3 2 62653 86975
0 16522 5 1 1 86979
0 16523 7 2 2 59540 84776
0 16524 7 1 2 86980 86982
0 16525 5 1 1 16524
0 16526 7 1 2 16519 16525
0 16527 5 1 1 16526
0 16528 7 1 2 16527 75064
0 16529 5 1 1 16528
0 16530 7 1 2 16499 16529
0 16531 5 1 1 16530
0 16532 7 1 2 75733 16531
0 16533 5 1 1 16532
0 16534 7 1 2 16475 16533
0 16535 5 1 1 16534
0 16536 7 1 2 59773 16535
0 16537 5 1 1 16536
0 16538 7 1 2 73002 82638
0 16539 5 1 1 16538
0 16540 7 4 2 63214 72895
0 16541 5 4 1 86984
0 16542 7 11 2 58475 59990
0 16543 5 1 1 86992
0 16544 7 1 2 67172 16543
0 16545 7 1 2 2077 16544
0 16546 7 1 2 86988 16545
0 16547 5 1 1 16546
0 16548 7 1 2 16539 16547
0 16549 5 1 1 16548
0 16550 7 1 2 62938 16549
0 16551 5 1 1 16550
0 16552 7 1 2 61236 77504
0 16553 7 1 2 85629 16552
0 16554 5 1 1 16553
0 16555 7 1 2 16551 16554
0 16556 5 1 1 16555
0 16557 7 1 2 75065 16556
0 16558 5 1 1 16557
0 16559 7 4 2 65866 74180
0 16560 5 1 1 87003
0 16561 7 1 2 87004 83746
0 16562 5 1 1 16561
0 16563 7 1 2 74220 82456
0 16564 5 1 1 16563
0 16565 7 4 2 65546 70403
0 16566 5 1 1 87007
0 16567 7 1 2 71646 87008
0 16568 5 1 1 16567
0 16569 7 1 2 76239 16568
0 16570 7 1 2 16564 16569
0 16571 5 1 1 16570
0 16572 7 1 2 61237 16571
0 16573 5 1 1 16572
0 16574 7 1 2 16562 16573
0 16575 5 1 1 16574
0 16576 7 1 2 71731 16575
0 16577 5 1 1 16576
0 16578 7 1 2 61238 76348
0 16579 5 1 1 16578
0 16580 7 1 2 69190 86403
0 16581 5 1 1 16580
0 16582 7 1 2 16579 16581
0 16583 5 1 1 16582
0 16584 7 1 2 74036 16583
0 16585 5 1 1 16584
0 16586 7 1 2 61239 2904
0 16587 5 1 1 16586
0 16588 7 1 2 73248 69117
0 16589 7 1 2 76781 16588
0 16590 5 1 1 16589
0 16591 7 1 2 16587 16590
0 16592 7 1 2 16585 16591
0 16593 7 1 2 16577 16592
0 16594 5 1 1 16593
0 16595 7 1 2 63215 16594
0 16596 5 1 1 16595
0 16597 7 10 2 62939 58476
0 16598 5 2 1 87011
0 16599 7 4 2 64022 80418
0 16600 5 2 1 87023
0 16601 7 1 2 87012 87024
0 16602 5 1 1 16601
0 16603 7 1 2 62940 80555
0 16604 5 3 1 16603
0 16605 7 1 2 70166 86719
0 16606 5 2 1 16605
0 16607 7 1 2 87029 87032
0 16608 5 1 1 16607
0 16609 7 1 2 74882 16608
0 16610 5 1 1 16609
0 16611 7 1 2 16602 16610
0 16612 7 1 2 16596 16611
0 16613 5 1 1 16612
0 16614 7 1 2 59541 16613
0 16615 5 1 1 16614
0 16616 7 2 2 61240 76338
0 16617 5 2 1 87034
0 16618 7 1 2 68364 72959
0 16619 7 1 2 87036 16618
0 16620 5 1 1 16619
0 16621 7 1 2 67852 86026
0 16622 5 1 1 16621
0 16623 7 1 2 16620 16622
0 16624 5 1 1 16623
0 16625 7 1 2 59325 16624
0 16626 5 1 1 16625
0 16627 7 1 2 73249 83747
0 16628 5 1 1 16627
0 16629 7 1 2 16626 16628
0 16630 5 1 1 16629
0 16631 7 1 2 77779 16630
0 16632 5 1 1 16631
0 16633 7 1 2 78478 85621
0 16634 5 1 1 16633
0 16635 7 1 2 70404 86720
0 16636 5 1 1 16635
0 16637 7 1 2 16634 16636
0 16638 5 1 1 16637
0 16639 7 1 2 68365 16638
0 16640 5 1 1 16639
0 16641 7 1 2 69968 86721
0 16642 7 1 2 67853 16641
0 16643 5 1 1 16642
0 16644 7 1 2 16640 16643
0 16645 5 1 1 16644
0 16646 7 1 2 65547 16645
0 16647 5 1 1 16646
0 16648 7 1 2 58477 87027
0 16649 5 2 1 16648
0 16650 7 1 2 63216 78997
0 16651 5 2 1 16650
0 16652 7 1 2 81287 87040
0 16653 7 1 2 87038 16652
0 16654 5 1 1 16653
0 16655 7 1 2 16647 16654
0 16656 5 1 1 16655
0 16657 7 1 2 64275 16656
0 16658 5 1 1 16657
0 16659 7 1 2 16632 16658
0 16660 5 1 1 16659
0 16661 7 1 2 57400 16660
0 16662 5 1 1 16661
0 16663 7 1 2 61241 78108
0 16664 7 1 2 85355 16663
0 16665 5 1 1 16664
0 16666 7 1 2 16662 16665
0 16667 5 1 1 16666
0 16668 7 1 2 71732 16667
0 16669 5 1 1 16668
0 16670 7 1 2 69451 74705
0 16671 5 1 1 16670
0 16672 7 1 2 70057 73003
0 16673 5 1 1 16672
0 16674 7 1 2 16671 16673
0 16675 5 1 1 16674
0 16676 7 1 2 63217 16675
0 16677 5 1 1 16676
0 16678 7 3 2 58478 77584
0 16679 7 1 2 85756 87042
0 16680 5 1 1 16679
0 16681 7 1 2 16677 16680
0 16682 5 1 1 16681
0 16683 7 1 2 58002 16682
0 16684 5 1 1 16683
0 16685 7 3 2 58972 85774
0 16686 5 1 1 87045
0 16687 7 1 2 77780 87046
0 16688 5 1 1 16687
0 16689 7 1 2 75433 78949
0 16690 5 1 1 16689
0 16691 7 1 2 16688 16690
0 16692 5 1 1 16691
0 16693 7 1 2 75303 16692
0 16694 5 1 1 16693
0 16695 7 3 2 58479 73618
0 16696 5 1 1 87048
0 16697 7 1 2 87049 81519
0 16698 5 1 1 16697
0 16699 7 1 2 16694 16698
0 16700 5 1 1 16699
0 16701 7 1 2 60544 16700
0 16702 5 1 1 16701
0 16703 7 1 2 69997 86722
0 16704 7 1 2 79375 16703
0 16705 5 1 1 16704
0 16706 7 1 2 16702 16705
0 16707 7 1 2 16684 16706
0 16708 5 1 1 16707
0 16709 7 1 2 68366 16708
0 16710 5 1 1 16709
0 16711 7 1 2 75434 87025
0 16712 5 1 1 16711
0 16713 7 2 2 59326 73306
0 16714 5 2 1 87051
0 16715 7 1 2 62941 87053
0 16716 5 1 1 16715
0 16717 7 1 2 72933 85533
0 16718 7 1 2 16716 16717
0 16719 5 1 1 16718
0 16720 7 1 2 16712 16719
0 16721 5 1 1 16720
0 16722 7 1 2 65229 16721
0 16723 5 1 1 16722
0 16724 7 3 2 80419 75435
0 16725 5 1 1 87055
0 16726 7 1 2 72529 87056
0 16727 5 1 1 16726
0 16728 7 1 2 16723 16727
0 16729 5 1 1 16728
0 16730 7 1 2 67854 16729
0 16731 5 1 1 16730
0 16732 7 1 2 63218 6916
0 16733 5 1 1 16732
0 16734 7 3 2 59327 80420
0 16735 5 2 1 87058
0 16736 7 2 2 57401 84189
0 16737 7 1 2 87059 87063
0 16738 7 1 2 16733 16737
0 16739 5 1 1 16738
0 16740 7 1 2 16731 16739
0 16741 5 1 1 16740
0 16742 7 1 2 68991 16741
0 16743 5 1 1 16742
0 16744 7 1 2 77781 74646
0 16745 5 1 1 16744
0 16746 7 1 2 87033 6184
0 16747 5 1 1 16746
0 16748 7 1 2 58003 16747
0 16749 5 1 1 16748
0 16750 7 1 2 78982 74190
0 16751 5 1 1 16750
0 16752 7 1 2 16749 16751
0 16753 5 1 1 16752
0 16754 7 1 2 64276 16753
0 16755 5 1 1 16754
0 16756 7 1 2 16745 16755
0 16757 5 1 1 16756
0 16758 7 1 2 67656 16757
0 16759 5 1 1 16758
0 16760 7 1 2 85644 86312
0 16761 5 1 1 16760
0 16762 7 2 2 72858 87013
0 16763 5 1 1 87065
0 16764 7 1 2 83390 74700
0 16765 7 1 2 77143 16764
0 16766 5 1 1 16765
0 16767 7 1 2 16763 16766
0 16768 5 1 1 16767
0 16769 7 4 2 72267 78645
0 16770 5 2 1 87067
0 16771 7 1 2 65230 87071
0 16772 7 1 2 16768 16771
0 16773 5 1 1 16772
0 16774 7 1 2 16761 16773
0 16775 5 1 1 16774
0 16776 7 1 2 73168 16775
0 16777 5 1 1 16776
0 16778 7 2 2 63219 70241
0 16779 5 2 1 87073
0 16780 7 1 2 84980 73004
0 16781 7 1 2 87075 16780
0 16782 5 1 1 16781
0 16783 7 1 2 16777 16782
0 16784 7 1 2 16759 16783
0 16785 7 1 2 16743 16784
0 16786 7 1 2 16710 16785
0 16787 7 1 2 16669 16786
0 16788 7 1 2 16615 16787
0 16789 5 1 1 16788
0 16790 7 1 2 64691 16789
0 16791 5 1 1 16790
0 16792 7 1 2 16558 16791
0 16793 5 1 1 16792
0 16794 7 1 2 66570 16793
0 16795 5 1 1 16794
0 16796 7 1 2 1209 86810
0 16797 7 1 2 69098 16796
0 16798 5 1 1 16797
0 16799 7 1 2 57678 16798
0 16800 5 1 1 16799
0 16801 7 1 2 86772 16800
0 16802 5 1 1 16801
0 16803 7 1 2 59542 16802
0 16804 5 1 1 16803
0 16805 7 1 2 75171 82442
0 16806 5 1 1 16805
0 16807 7 1 2 16804 16806
0 16808 5 1 1 16807
0 16809 7 1 2 58282 16808
0 16810 5 1 1 16809
0 16811 7 1 2 59543 85019
0 16812 5 1 1 16811
0 16813 7 1 2 16810 16812
0 16814 5 1 1 16813
0 16815 7 1 2 65231 16814
0 16816 5 1 1 16815
0 16817 7 1 2 59544 86820
0 16818 5 1 1 16817
0 16819 7 1 2 16816 16818
0 16820 5 1 1 16819
0 16821 7 1 2 85544 83364
0 16822 7 1 2 16820 16821
0 16823 5 1 1 16822
0 16824 7 1 2 61561 16823
0 16825 7 1 2 16795 16824
0 16826 5 1 1 16825
0 16827 7 1 2 61242 82856
0 16828 5 1 1 16827
0 16829 7 1 2 78268 87005
0 16830 5 1 1 16829
0 16831 7 1 2 74741 78960
0 16832 5 2 1 16831
0 16833 7 1 2 73873 87077
0 16834 5 1 1 16833
0 16835 7 1 2 16830 16834
0 16836 7 1 2 16828 16835
0 16837 5 1 1 16836
0 16838 7 1 2 75871 16837
0 16839 5 1 1 16838
0 16840 7 2 2 73064 78961
0 16841 5 1 1 87079
0 16842 7 1 2 87080 84430
0 16843 5 1 1 16842
0 16844 7 1 2 87009 16843
0 16845 5 1 1 16844
0 16846 7 1 2 73065 16560
0 16847 5 2 1 16846
0 16848 7 1 2 76148 87081
0 16849 5 1 1 16848
0 16850 7 1 2 85525 72820
0 16851 5 1 1 16850
0 16852 7 1 2 16849 16851
0 16853 7 1 2 16845 16852
0 16854 7 1 2 16839 16853
0 16855 5 1 1 16854
0 16856 7 1 2 71733 16855
0 16857 5 1 1 16856
0 16858 7 1 2 69023 79681
0 16859 5 4 1 16858
0 16860 7 1 2 74858 87083
0 16861 5 2 1 16860
0 16862 7 1 2 87087 82085
0 16863 5 1 1 16862
0 16864 7 1 2 57402 16863
0 16865 5 1 1 16864
0 16866 7 1 2 67657 73402
0 16867 5 3 1 16866
0 16868 7 1 2 16865 87089
0 16869 5 1 1 16868
0 16870 7 1 2 71485 16869
0 16871 5 1 1 16870
0 16872 7 1 2 71172 84560
0 16873 5 1 1 16872
0 16874 7 1 2 16871 16873
0 16875 5 1 1 16874
0 16876 7 1 2 73169 16875
0 16877 5 1 1 16876
0 16878 7 1 2 57403 86138
0 16879 5 1 1 16878
0 16880 7 4 2 62654 75182
0 16881 5 5 1 87092
0 16882 7 1 2 70966 87096
0 16883 5 1 1 16882
0 16884 7 1 2 16879 16883
0 16885 5 1 1 16884
0 16886 7 1 2 84943 16885
0 16887 5 1 1 16886
0 16888 7 1 2 71262 78378
0 16889 7 1 2 8463 16888
0 16890 5 1 1 16889
0 16891 7 1 2 70167 84946
0 16892 7 1 2 16890 16891
0 16893 5 1 1 16892
0 16894 7 1 2 84939 79386
0 16895 5 1 1 16894
0 16896 7 1 2 71173 70934
0 16897 5 1 1 16896
0 16898 7 1 2 16895 16897
0 16899 5 1 1 16898
0 16900 7 1 2 84898 16899
0 16901 5 1 1 16900
0 16902 7 1 2 61243 16901
0 16903 7 1 2 16893 16902
0 16904 7 1 2 16887 16903
0 16905 7 1 2 16877 16904
0 16906 5 1 1 16905
0 16907 7 1 2 60876 86391
0 16908 5 1 1 16907
0 16909 7 1 2 69738 86400
0 16910 5 1 1 16909
0 16911 7 2 2 59545 79538
0 16912 5 1 1 87101
0 16913 7 1 2 16910 16912
0 16914 7 1 2 16908 16913
0 16915 5 1 1 16914
0 16916 7 1 2 59328 16915
0 16917 5 1 1 16916
0 16918 7 1 2 64277 15580
0 16919 5 1 1 16918
0 16920 7 2 2 68496 73758
0 16921 5 1 1 87103
0 16922 7 1 2 62376 87104
0 16923 5 1 1 16922
0 16924 7 1 2 16919 16923
0 16925 5 1 1 16924
0 16926 7 1 2 65548 16925
0 16927 5 1 1 16926
0 16928 7 1 2 78220 83621
0 16929 5 1 1 16928
0 16930 7 1 2 69739 86384
0 16931 5 1 1 16930
0 16932 7 1 2 16929 16931
0 16933 5 1 1 16932
0 16934 7 1 2 71883 16933
0 16935 5 1 1 16934
0 16936 7 1 2 86398 83622
0 16937 5 1 1 16936
0 16938 7 1 2 65867 16937
0 16939 7 1 2 16935 16938
0 16940 7 1 2 16927 16939
0 16941 7 1 2 16917 16940
0 16942 5 1 1 16941
0 16943 7 1 2 16906 16942
0 16944 5 1 1 16943
0 16945 7 1 2 16857 16944
0 16946 5 1 1 16945
0 16947 7 1 2 75955 16946
0 16948 5 1 1 16947
0 16949 7 4 2 61915 73307
0 16950 7 2 2 87105 82273
0 16951 7 1 2 87109 80218
0 16952 5 1 1 16951
0 16953 7 1 2 67173 79996
0 16954 7 1 2 75734 16953
0 16955 7 1 2 86075 16954
0 16956 5 1 1 16955
0 16957 7 1 2 16952 16956
0 16958 5 1 1 16957
0 16959 7 1 2 70623 16958
0 16960 5 1 1 16959
0 16961 7 1 2 59329 87110
0 16962 5 1 1 16961
0 16963 7 1 2 69921 86263
0 16964 7 1 2 77213 16963
0 16965 5 1 1 16964
0 16966 7 1 2 16962 16965
0 16967 5 1 1 16966
0 16968 7 1 2 62655 16967
0 16969 5 1 1 16968
0 16970 7 1 2 58480 16969
0 16971 7 1 2 16960 16970
0 16972 7 1 2 16948 16971
0 16973 5 1 1 16972
0 16974 7 1 2 75735 4287
0 16975 5 1 1 16974
0 16976 7 2 2 71884 77144
0 16977 5 1 1 87111
0 16978 7 1 2 67420 87112
0 16979 5 1 1 16978
0 16980 7 1 2 59330 74859
0 16981 5 8 1 16980
0 16982 7 1 2 14990 87113
0 16983 7 1 2 16979 16982
0 16984 5 1 1 16983
0 16985 7 1 2 79048 83365
0 16986 7 1 2 16984 16985
0 16987 5 1 1 16986
0 16988 7 1 2 63220 16987
0 16989 7 1 2 16975 16988
0 16990 5 1 1 16989
0 16991 7 1 2 16973 16990
0 16992 5 1 1 16991
0 16993 7 3 2 79114 80512
0 16994 5 1 1 87121
0 16995 7 1 2 73250 16994
0 16996 5 1 1 16995
0 16997 7 1 2 86027 69127
0 16998 5 1 1 16997
0 16999 7 1 2 16996 16998
0 17000 5 1 1 16999
0 17001 7 1 2 57404 17000
0 17002 5 1 1 17001
0 17003 7 1 2 80046 73251
0 17004 5 1 1 17003
0 17005 7 1 2 17002 17004
0 17006 5 1 1 17005
0 17007 7 1 2 57679 17006
0 17008 5 1 1 17007
0 17009 7 1 2 73952 83485
0 17010 5 1 1 17009
0 17011 7 1 2 17008 17010
0 17012 5 1 1 17011
0 17013 7 1 2 83643 75956
0 17014 7 1 2 17012 17013
0 17015 5 1 1 17014
0 17016 7 1 2 66176 17015
0 17017 7 1 2 16992 17016
0 17018 5 1 1 17017
0 17019 7 1 2 64497 17018
0 17020 7 1 2 16826 17019
0 17021 5 1 1 17020
0 17022 7 1 2 65868 80539
0 17023 5 1 1 17022
0 17024 7 1 2 17023 80618
0 17025 5 1 1 17024
0 17026 7 1 2 59991 81112
0 17027 7 1 2 84482 17026
0 17028 7 1 2 17025 17027
0 17029 5 1 1 17028
0 17030 7 1 2 63480 17029
0 17031 7 1 2 17021 17030
0 17032 7 1 2 16537 17031
0 17033 5 1 1 17032
0 17034 7 3 2 63868 72473
0 17035 5 2 1 87124
0 17036 7 1 2 77012 87127
0 17037 5 3 1 17036
0 17038 7 1 2 85342 87129
0 17039 5 1 1 17038
0 17040 7 2 2 70674 68653
0 17041 7 1 2 77230 87132
0 17042 5 1 1 17041
0 17043 7 1 2 17039 17042
0 17044 5 1 1 17043
0 17045 7 8 2 59992 61244
0 17046 5 3 1 87134
0 17047 7 3 2 64278 87135
0 17048 5 1 1 87145
0 17049 7 1 2 17044 87146
0 17050 5 1 1 17049
0 17051 7 1 2 82945 68654
0 17052 5 1 1 17051
0 17053 7 1 2 85128 86873
0 17054 5 1 1 17053
0 17055 7 1 2 17052 17054
0 17056 5 1 1 17055
0 17057 7 1 2 65549 17056
0 17058 5 1 1 17057
0 17059 7 1 2 84485 17058
0 17060 5 1 1 17059
0 17061 7 1 2 60545 17060
0 17062 5 1 1 17061
0 17063 7 1 2 72651 87125
0 17064 5 1 1 17063
0 17065 7 1 2 17062 17064
0 17066 5 1 1 17065
0 17067 7 1 2 64692 17066
0 17068 5 1 1 17067
0 17069 7 7 2 59993 60877
0 17070 7 1 2 80799 87148
0 17071 7 1 2 78065 17070
0 17072 5 1 1 17071
0 17073 7 1 2 17068 17072
0 17074 5 1 1 17073
0 17075 7 1 2 59774 17074
0 17076 5 1 1 17075
0 17077 7 1 2 73591 76798
0 17078 5 1 1 17077
0 17079 7 1 2 78269 17078
0 17080 5 1 1 17079
0 17081 7 1 2 71263 77925
0 17082 7 1 2 17080 17081
0 17083 5 1 1 17082
0 17084 7 1 2 60546 78051
0 17085 7 1 2 17083 17084
0 17086 5 1 1 17085
0 17087 7 1 2 78110 17086
0 17088 5 1 1 17087
0 17089 7 1 2 63221 17088
0 17090 5 1 1 17089
0 17091 7 2 2 62942 78112
0 17092 5 1 1 87155
0 17093 7 2 2 67174 87156
0 17094 5 1 1 87157
0 17095 7 1 2 17090 17094
0 17096 5 1 1 17095
0 17097 7 1 2 84000 17096
0 17098 5 1 1 17097
0 17099 7 1 2 86959 87133
0 17100 5 1 1 17099
0 17101 7 1 2 17098 17100
0 17102 7 1 2 17076 17101
0 17103 5 1 1 17102
0 17104 7 1 2 65869 17103
0 17105 5 1 1 17104
0 17106 7 1 2 17050 17105
0 17107 5 1 1 17106
0 17108 7 1 2 61562 17107
0 17109 5 1 1 17108
0 17110 7 3 2 63222 84001
0 17111 5 1 1 87159
0 17112 7 3 2 58481 79820
0 17113 5 5 1 87162
0 17114 7 1 2 17111 87165
0 17115 5 5 1 17114
0 17116 7 1 2 76179 87170
0 17117 5 1 1 17116
0 17118 7 2 2 84883 79849
0 17119 5 1 1 87175
0 17120 7 1 2 17117 17119
0 17121 5 1 1 17120
0 17122 7 1 2 66177 17121
0 17123 5 1 1 17122
0 17124 7 11 2 64279 61563
0 17125 5 3 1 87177
0 17126 7 1 2 85335 87178
0 17127 7 1 2 85859 17126
0 17128 5 1 1 17127
0 17129 7 1 2 17123 17128
0 17130 5 1 1 17129
0 17131 7 1 2 72474 17130
0 17132 5 1 1 17131
0 17133 7 2 2 62656 79255
0 17134 7 2 2 63223 69922
0 17135 7 1 2 78446 81386
0 17136 7 1 2 87193 17135
0 17137 7 1 2 87191 17136
0 17138 5 1 1 17137
0 17139 7 1 2 17132 17138
0 17140 5 1 1 17139
0 17141 7 1 2 61245 17140
0 17142 5 1 1 17141
0 17143 7 18 2 60878 84651
0 17144 5 6 1 87195
0 17145 7 2 2 71804 87196
0 17146 5 4 1 87219
0 17147 7 4 2 65232 86459
0 17148 7 2 2 65550 87225
0 17149 5 1 1 87229
0 17150 7 1 2 87221 17149
0 17151 5 1 1 17150
0 17152 7 1 2 59546 17151
0 17153 5 1 1 17152
0 17154 7 10 2 65233 66178
0 17155 5 2 1 87231
0 17156 7 1 2 85740 87232
0 17157 5 1 1 17156
0 17158 7 1 2 17153 17157
0 17159 5 1 1 17158
0 17160 7 1 2 84981 84002
0 17161 5 1 1 17160
0 17162 7 1 2 87166 17161
0 17163 5 1 1 17162
0 17164 7 1 2 17159 17163
0 17165 5 1 1 17164
0 17166 7 1 2 58482 78024
0 17167 5 2 1 17166
0 17168 7 1 2 59994 86460
0 17169 7 1 2 85343 17168
0 17170 7 1 2 87243 17169
0 17171 5 1 1 17170
0 17172 7 1 2 17165 17171
0 17173 7 1 2 17142 17172
0 17174 5 1 1 17173
0 17175 7 1 2 70624 17174
0 17176 5 1 1 17175
0 17177 7 1 2 78534 87128
0 17178 5 1 1 17177
0 17179 7 1 2 67175 17178
0 17180 5 1 1 17179
0 17181 7 1 2 71264 74451
0 17182 5 1 1 17181
0 17183 7 4 2 60547 86874
0 17184 5 2 1 87245
0 17185 7 1 2 64280 87246
0 17186 5 1 1 17185
0 17187 7 1 2 17182 17186
0 17188 5 1 1 17187
0 17189 7 1 2 65551 17188
0 17190 5 1 1 17189
0 17191 7 1 2 17180 17190
0 17192 5 1 1 17191
0 17193 7 1 2 87171 17192
0 17194 5 1 1 17193
0 17195 7 2 2 63869 80842
0 17196 7 1 2 81753 87251
0 17197 5 1 1 17196
0 17198 7 1 2 75373 73963
0 17199 7 1 2 68655 17198
0 17200 5 1 1 17199
0 17201 7 1 2 17197 17200
0 17202 5 1 1 17201
0 17203 7 1 2 69740 17202
0 17204 5 1 1 17203
0 17205 7 1 2 17194 17204
0 17206 5 1 1 17205
0 17207 7 1 2 84652 17206
0 17208 5 1 1 17207
0 17209 7 1 2 17176 17208
0 17210 7 1 2 17109 17209
0 17211 5 1 1 17210
0 17212 7 1 2 60320 17211
0 17213 5 1 1 17212
0 17214 7 22 2 64498 61564
0 17215 5 2 1 87253
0 17216 7 1 2 71486 78430
0 17217 5 1 1 17216
0 17218 7 1 2 71265 83411
0 17219 5 1 1 17218
0 17220 7 3 2 68822 71266
0 17221 5 1 1 87277
0 17222 7 1 2 65022 17221
0 17223 7 1 2 17219 17222
0 17224 5 1 1 17223
0 17225 7 2 2 17217 17224
0 17226 7 1 2 70067 77930
0 17227 7 1 2 10808 17226
0 17228 5 1 1 17227
0 17229 7 1 2 59547 17228
0 17230 5 1 1 17229
0 17231 7 1 2 87280 17230
0 17232 5 1 1 17231
0 17233 7 1 2 65552 17232
0 17234 5 1 1 17233
0 17235 7 1 2 70405 77186
0 17236 5 1 1 17235
0 17237 7 1 2 78830 17236
0 17238 5 1 1 17237
0 17239 7 1 2 59548 17238
0 17240 5 1 1 17239
0 17241 7 1 2 17234 17240
0 17242 5 2 1 17241
0 17243 7 1 2 87254 87282
0 17244 5 1 1 17243
0 17245 7 5 2 62943 77893
0 17246 5 1 1 87284
0 17247 7 1 2 72296 87285
0 17248 5 1 1 17247
0 17249 7 1 2 60879 73715
0 17250 5 1 1 17249
0 17251 7 1 2 17248 17250
0 17252 5 1 1 17251
0 17253 7 1 2 64023 17252
0 17254 5 1 1 17253
0 17255 7 1 2 79156 77053
0 17256 5 1 1 17255
0 17257 7 1 2 17254 17256
0 17258 5 1 1 17257
0 17259 7 1 2 62657 17258
0 17260 5 1 1 17259
0 17261 7 1 2 75152 2554
0 17262 5 1 1 17261
0 17263 7 1 2 69414 17262
0 17264 5 1 1 17263
0 17265 7 1 2 68613 86142
0 17266 5 1 1 17265
0 17267 7 1 2 57680 82169
0 17268 5 1 1 17267
0 17269 7 2 2 68992 79104
0 17270 5 2 1 87289
0 17271 7 1 2 85359 87291
0 17272 7 1 2 17268 17271
0 17273 7 1 2 17266 17272
0 17274 5 1 1 17273
0 17275 7 1 2 60880 17274
0 17276 5 1 1 17275
0 17277 7 1 2 17264 17276
0 17278 5 2 1 17277
0 17279 7 1 2 79157 87293
0 17280 5 1 1 17279
0 17281 7 1 2 17260 17280
0 17282 5 1 1 17281
0 17283 7 1 2 66179 17282
0 17284 5 1 1 17283
0 17285 7 1 2 61246 17284
0 17286 7 1 2 17244 17285
0 17287 5 1 1 17286
0 17288 7 1 2 78388 87255
0 17289 5 1 1 17288
0 17290 7 1 2 76799 82517
0 17291 7 1 2 85618 17290
0 17292 5 1 1 17291
0 17293 7 1 2 17289 17292
0 17294 5 1 1 17293
0 17295 7 1 2 60881 17294
0 17296 5 1 1 17295
0 17297 7 1 2 79158 81494
0 17298 7 1 2 78431 17297
0 17299 5 1 1 17298
0 17300 7 2 2 63870 82548
0 17301 5 2 1 87295
0 17302 7 2 2 68497 82194
0 17303 5 3 1 87299
0 17304 7 1 2 87297 87301
0 17305 5 1 1 17304
0 17306 7 1 2 79294 17305
0 17307 5 1 1 17306
0 17308 7 2 2 61565 69415
0 17309 7 1 2 85323 87304
0 17310 5 1 1 17309
0 17311 7 1 2 17307 17310
0 17312 5 1 1 17311
0 17313 7 1 2 62658 17312
0 17314 5 1 1 17313
0 17315 7 1 2 65870 17314
0 17316 7 1 2 17299 17315
0 17317 7 1 2 17296 17316
0 17318 5 1 1 17317
0 17319 7 1 2 63224 17318
0 17320 7 1 2 17287 17319
0 17321 5 1 1 17320
0 17322 7 3 2 62377 82195
0 17323 5 1 1 87306
0 17324 7 1 2 85448 87307
0 17325 5 1 1 17324
0 17326 7 2 2 59775 70625
0 17327 7 1 2 86983 87309
0 17328 5 1 1 17327
0 17329 7 1 2 17325 17328
0 17330 5 1 1 17329
0 17331 7 1 2 71805 17330
0 17332 5 1 1 17331
0 17333 7 2 2 64281 73496
0 17334 5 4 1 87311
0 17335 7 2 2 81251 87312
0 17336 5 1 1 87317
0 17337 7 1 2 17332 17336
0 17338 5 1 1 17337
0 17339 7 1 2 80862 17338
0 17340 5 1 1 17339
0 17341 7 4 2 64282 73361
0 17342 5 1 1 87319
0 17343 7 1 2 81427 87320
0 17344 7 1 2 86894 17343
0 17345 5 1 1 17344
0 17346 7 1 2 17340 17345
0 17347 5 1 1 17346
0 17348 7 1 2 60882 17347
0 17349 5 1 1 17348
0 17350 7 1 2 70626 87318
0 17351 5 1 1 17350
0 17352 7 3 2 64499 86554
0 17353 5 1 1 87323
0 17354 7 2 2 84462 87324
0 17355 5 1 1 87326
0 17356 7 1 2 17351 17355
0 17357 5 1 1 17356
0 17358 7 1 2 60883 17357
0 17359 5 1 1 17358
0 17360 7 2 2 63225 77356
0 17361 7 4 2 65553 84653
0 17362 5 1 1 87330
0 17363 7 1 2 87328 87331
0 17364 5 1 1 17363
0 17365 7 1 2 17359 17364
0 17366 5 1 1 17365
0 17367 7 1 2 71806 17366
0 17368 5 1 1 17367
0 17369 7 1 2 64283 87327
0 17370 5 1 1 17369
0 17371 7 1 2 17368 17370
0 17372 5 1 1 17371
0 17373 7 1 2 76180 17372
0 17374 5 1 1 17373
0 17375 7 1 2 82590 82220
0 17376 5 14 1 17375
0 17377 7 2 2 61247 87334
0 17378 5 1 1 87348
0 17379 7 3 2 59549 87256
0 17380 5 2 1 87350
0 17381 7 1 2 17378 87353
0 17382 5 1 1 17381
0 17383 7 2 2 73066 17382
0 17384 7 2 2 65554 87355
0 17385 7 1 2 85003 81851
0 17386 7 1 2 87357 17385
0 17387 5 1 1 17386
0 17388 7 1 2 59995 17387
0 17389 7 1 2 17374 17388
0 17390 7 1 2 17349 17389
0 17391 7 1 2 17321 17390
0 17392 5 1 1 17391
0 17393 7 1 2 78185 78373
0 17394 5 1 1 17393
0 17395 7 2 2 70812 75797
0 17396 5 1 1 87359
0 17397 7 1 2 67319 17396
0 17398 5 1 1 17397
0 17399 7 1 2 68770 75917
0 17400 5 1 1 17399
0 17401 7 1 2 82849 17400
0 17402 7 1 2 17398 17401
0 17403 5 1 1 17402
0 17404 7 1 2 71487 17403
0 17405 5 1 1 17404
0 17406 7 1 2 17394 17405
0 17407 5 1 1 17406
0 17408 7 1 2 65023 17407
0 17409 5 1 1 17408
0 17410 7 1 2 71174 76808
0 17411 5 1 1 17410
0 17412 7 1 2 71488 68656
0 17413 5 1 1 17412
0 17414 7 1 2 17411 17413
0 17415 7 1 2 17409 17414
0 17416 5 1 1 17415
0 17417 7 1 2 61566 17416
0 17418 5 1 1 17417
0 17419 7 1 2 86865 81567
0 17420 5 1 1 17419
0 17421 7 1 2 71600 81330
0 17422 5 1 1 17421
0 17423 7 1 2 68081 71665
0 17424 5 2 1 17423
0 17425 7 1 2 87361 84291
0 17426 5 1 1 17425
0 17427 7 1 2 71267 17426
0 17428 5 1 1 17427
0 17429 7 1 2 61567 17428
0 17430 5 1 1 17429
0 17431 7 1 2 17422 17430
0 17432 5 1 1 17431
0 17433 7 1 2 65234 17432
0 17434 5 1 1 17433
0 17435 7 1 2 17420 17434
0 17436 7 1 2 17418 17435
0 17437 5 1 1 17436
0 17438 7 1 2 65555 17437
0 17439 5 1 1 17438
0 17440 7 1 2 82857 81442
0 17441 5 1 1 17440
0 17442 7 1 2 82505 17441
0 17443 5 1 1 17442
0 17444 7 1 2 71657 17443
0 17445 5 1 1 17444
0 17446 7 2 2 69505 81387
0 17447 7 1 2 75796 87363
0 17448 5 1 1 17447
0 17449 7 3 2 70813 75721
0 17450 5 1 1 87365
0 17451 7 1 2 75798 87366
0 17452 5 3 1 17451
0 17453 7 3 2 61568 71489
0 17454 7 1 2 82845 87371
0 17455 7 1 2 87368 17454
0 17456 5 1 1 17455
0 17457 7 1 2 17448 17456
0 17458 7 1 2 17445 17457
0 17459 7 1 2 57405 74037
0 17460 5 1 1 17459
0 17461 7 3 2 59110 76565
0 17462 5 2 1 87374
0 17463 7 1 2 17460 87377
0 17464 5 1 1 17463
0 17465 7 1 2 57681 17464
0 17466 5 1 1 17465
0 17467 7 1 2 58004 83591
0 17468 5 1 1 17467
0 17469 7 2 2 64284 17468
0 17470 7 1 2 17466 87379
0 17471 5 1 1 17470
0 17472 7 1 2 73592 81388
0 17473 7 1 2 17471 17472
0 17474 5 1 1 17473
0 17475 7 4 2 67658 74221
0 17476 5 3 1 87381
0 17477 7 1 2 78380 87382
0 17478 5 1 1 17477
0 17479 7 1 2 71268 17478
0 17480 5 1 1 17479
0 17481 7 1 2 61569 17480
0 17482 5 1 1 17481
0 17483 7 1 2 76809 82507
0 17484 5 1 1 17483
0 17485 7 1 2 17482 17484
0 17486 5 1 1 17485
0 17487 7 1 2 67320 17486
0 17488 5 1 1 17487
0 17489 7 1 2 17474 17488
0 17490 7 1 2 17458 17489
0 17491 7 1 2 17439 17490
0 17492 5 1 1 17491
0 17493 7 1 2 58483 17492
0 17494 5 1 1 17493
0 17495 7 2 2 72281 81331
0 17496 7 1 2 80493 87388
0 17497 5 1 1 17496
0 17498 7 1 2 74122 81353
0 17499 5 1 1 17498
0 17500 7 1 2 6892 17499
0 17501 5 1 1 17500
0 17502 7 1 2 78758 17501
0 17503 5 1 1 17502
0 17504 7 1 2 17497 17503
0 17505 5 1 1 17504
0 17506 7 1 2 59111 17505
0 17507 5 1 1 17506
0 17508 7 3 2 59331 76503
0 17509 5 2 1 87390
0 17510 7 2 2 78410 87391
0 17511 5 2 1 87395
0 17512 7 1 2 81366 87396
0 17513 5 1 1 17512
0 17514 7 1 2 17507 17513
0 17515 5 1 1 17514
0 17516 7 1 2 57682 17515
0 17517 5 1 1 17516
0 17518 7 1 2 79131 87389
0 17519 5 1 1 17518
0 17520 7 1 2 17517 17519
0 17521 5 1 1 17520
0 17522 7 1 2 58005 17521
0 17523 5 1 1 17522
0 17524 7 1 2 83406 78824
0 17525 7 1 2 87364 17524
0 17526 5 1 1 17525
0 17527 7 1 2 17523 17526
0 17528 5 1 1 17527
0 17529 7 1 2 58283 17528
0 17530 5 1 1 17529
0 17531 7 1 2 61248 17530
0 17532 7 1 2 17494 17531
0 17533 5 1 1 17532
0 17534 7 1 2 74535 80047
0 17535 5 1 1 17534
0 17536 7 1 2 68993 82478
0 17537 5 1 1 17536
0 17538 7 1 2 73815 17537
0 17539 5 1 1 17538
0 17540 7 1 2 57683 74145
0 17541 7 1 2 17539 17540
0 17542 5 1 1 17541
0 17543 7 1 2 17535 17542
0 17544 5 1 1 17543
0 17545 7 1 2 57406 17544
0 17546 5 1 1 17545
0 17547 7 2 2 65024 67013
0 17548 5 1 1 87399
0 17549 7 1 2 83733 17548
0 17550 5 1 1 17549
0 17551 7 1 2 74536 17550
0 17552 5 1 1 17551
0 17553 7 1 2 17546 17552
0 17554 5 1 1 17553
0 17555 7 1 2 85290 17554
0 17556 5 1 1 17555
0 17557 7 1 2 59332 80108
0 17558 5 1 1 17557
0 17559 7 1 2 71490 67855
0 17560 5 2 1 17559
0 17561 7 1 2 17558 87401
0 17562 5 1 1 17561
0 17563 7 1 2 60884 17562
0 17564 5 1 1 17563
0 17565 7 1 2 78818 72508
0 17566 5 1 1 17565
0 17567 7 1 2 65556 79714
0 17568 7 1 2 17566 17567
0 17569 5 1 1 17568
0 17570 7 1 2 17564 17569
0 17571 5 2 1 17570
0 17572 7 1 2 58484 87403
0 17573 5 1 1 17572
0 17574 7 1 2 71175 83409
0 17575 5 1 1 17574
0 17576 7 1 2 17573 17575
0 17577 5 1 1 17576
0 17578 7 1 2 69416 17577
0 17579 5 1 1 17578
0 17580 7 1 2 63226 13319
0 17581 5 1 1 17580
0 17582 7 1 2 78905 17581
0 17583 5 1 1 17582
0 17584 7 2 2 58485 70406
0 17585 5 2 1 87405
0 17586 7 2 2 67742 76307
0 17587 5 2 1 87409
0 17588 7 1 2 57407 87411
0 17589 5 1 1 17588
0 17590 7 2 2 83447 17589
0 17591 7 1 2 64285 78424
0 17592 7 1 2 87413 17591
0 17593 5 1 1 17592
0 17594 7 1 2 87406 17593
0 17595 5 1 1 17594
0 17596 7 1 2 17583 17595
0 17597 5 1 1 17596
0 17598 7 1 2 60885 17597
0 17599 5 1 1 17598
0 17600 7 1 2 85129 76810
0 17601 5 1 1 17600
0 17602 7 1 2 74332 82946
0 17603 7 1 2 79596 17602
0 17604 5 1 1 17603
0 17605 7 1 2 17601 17604
0 17606 5 1 1 17605
0 17607 7 1 2 60886 17606
0 17608 5 1 1 17607
0 17609 7 2 2 65557 75436
0 17610 7 1 2 4338 87415
0 17611 5 1 1 17610
0 17612 7 1 2 17608 17611
0 17613 5 1 1 17612
0 17614 7 1 2 67321 17613
0 17615 5 1 1 17614
0 17616 7 1 2 61570 17615
0 17617 7 1 2 17599 17616
0 17618 7 1 2 17579 17617
0 17619 7 1 2 17556 17618
0 17620 5 1 1 17619
0 17621 7 1 2 78031 78115
0 17622 5 1 1 17621
0 17623 7 4 2 62944 74123
0 17624 5 2 1 87417
0 17625 7 1 2 65235 87418
0 17626 5 1 1 17625
0 17627 7 1 2 78106 17626
0 17628 5 1 1 17627
0 17629 7 1 2 62378 17628
0 17630 5 1 1 17629
0 17631 7 1 2 17092 17630
0 17632 5 1 1 17631
0 17633 7 1 2 67176 17632
0 17634 5 1 1 17633
0 17635 7 1 2 17622 17634
0 17636 5 1 1 17635
0 17637 7 1 2 68498 17636
0 17638 5 1 1 17637
0 17639 7 1 2 62379 87158
0 17640 5 1 1 17639
0 17641 7 1 2 66180 17640
0 17642 7 1 2 17638 17641
0 17643 5 1 1 17642
0 17644 7 1 2 17620 17643
0 17645 5 1 1 17644
0 17646 7 1 2 65871 17645
0 17647 5 1 1 17646
0 17648 7 1 2 59776 17647
0 17649 7 1 2 17533 17648
0 17650 5 1 1 17649
0 17651 7 1 2 78335 81252
0 17652 5 1 1 17651
0 17653 7 2 2 74812 82602
0 17654 5 1 1 87423
0 17655 7 1 2 17652 17654
0 17656 5 1 1 17655
0 17657 7 1 2 60887 17656
0 17658 5 1 1 17657
0 17659 7 1 2 66181 78397
0 17660 5 1 1 17659
0 17661 7 1 2 17658 17660
0 17662 5 1 1 17661
0 17663 7 1 2 59333 17662
0 17664 5 1 1 17663
0 17665 7 5 2 64500 72020
0 17666 7 5 2 58973 66182
0 17667 7 1 2 73998 87430
0 17668 7 1 2 87425 17667
0 17669 5 1 1 17668
0 17670 7 1 2 17664 17669
0 17671 5 1 1 17670
0 17672 7 1 2 73653 17671
0 17673 5 1 1 17672
0 17674 7 1 2 57408 80556
0 17675 7 1 2 79398 17674
0 17676 7 1 2 86748 17675
0 17677 5 1 1 17676
0 17678 7 1 2 17673 17677
0 17679 5 1 1 17678
0 17680 7 1 2 71885 17679
0 17681 5 1 1 17680
0 17682 7 2 2 57409 82196
0 17683 5 2 1 87435
0 17684 7 1 2 81268 87437
0 17685 5 2 1 17684
0 17686 7 1 2 72282 87439
0 17687 5 1 1 17686
0 17688 7 8 2 63227 82197
0 17689 5 2 1 87441
0 17690 7 1 2 78968 87442
0 17691 5 1 1 17690
0 17692 7 1 2 17687 17691
0 17693 5 1 1 17692
0 17694 7 1 2 73654 17693
0 17695 5 1 1 17694
0 17696 7 6 2 64501 84654
0 17697 5 3 1 87451
0 17698 7 1 2 80635 87452
0 17699 5 1 1 17698
0 17700 7 1 2 17695 17699
0 17701 5 1 1 17700
0 17702 7 1 2 75872 17701
0 17703 5 1 1 17702
0 17704 7 8 2 57410 65872
0 17705 5 2 1 87460
0 17706 7 1 2 82870 87461
0 17707 7 1 2 79404 17706
0 17708 5 1 1 17707
0 17709 7 1 2 17703 17708
0 17710 5 1 1 17709
0 17711 7 1 2 71734 17710
0 17712 5 1 1 17711
0 17713 7 2 2 74124 86723
0 17714 5 1 1 87470
0 17715 7 2 2 68994 82198
0 17716 5 1 1 87472
0 17717 7 1 2 87471 87473
0 17718 5 1 1 17717
0 17719 7 7 2 61571 73655
0 17720 5 1 1 87474
0 17721 7 1 2 60888 87475
0 17722 5 1 1 17721
0 17723 7 1 2 87457 17722
0 17724 5 2 1 17723
0 17725 7 1 2 58486 70081
0 17726 7 1 2 87481 17725
0 17727 5 1 1 17726
0 17728 7 7 2 65558 86555
0 17729 5 1 1 87483
0 17730 7 1 2 80897 87484
0 17731 5 1 1 17730
0 17732 7 1 2 17727 17731
0 17733 5 1 1 17732
0 17734 7 1 2 57684 17733
0 17735 5 1 1 17734
0 17736 7 1 2 17718 17735
0 17737 5 1 1 17736
0 17738 7 1 2 72242 17737
0 17739 5 1 1 17738
0 17740 7 2 2 68614 82199
0 17741 5 1 1 87490
0 17742 7 1 2 80557 87491
0 17743 7 1 2 76278 17742
0 17744 5 1 1 17743
0 17745 7 1 2 17739 17744
0 17746 7 1 2 17712 17745
0 17747 7 1 2 17681 17746
0 17748 5 1 1 17747
0 17749 7 1 2 58006 17748
0 17750 5 1 1 17749
0 17751 7 2 2 73543 84655
0 17752 5 1 1 87492
0 17753 7 1 2 76811 87493
0 17754 5 1 1 17753
0 17755 7 14 2 59777 65873
0 17756 5 1 1 87494
0 17757 7 1 2 72896 17756
0 17758 7 1 2 80612 17757
0 17759 5 1 1 17758
0 17760 7 1 2 13814 17759
0 17761 5 1 1 17760
0 17762 7 1 2 61572 17761
0 17763 5 1 1 17762
0 17764 7 1 2 87458 17763
0 17765 5 1 1 17764
0 17766 7 1 2 57411 17765
0 17767 5 1 1 17766
0 17768 7 1 2 57685 87482
0 17769 5 1 1 17768
0 17770 7 1 2 17767 17769
0 17771 5 1 1 17770
0 17772 7 1 2 70777 17771
0 17773 5 1 1 17772
0 17774 7 1 2 17754 17773
0 17775 5 1 1 17774
0 17776 7 1 2 58487 17775
0 17777 5 1 1 17776
0 17778 7 1 2 68995 73252
0 17779 5 2 1 17778
0 17780 7 1 2 61249 79620
0 17781 5 2 1 17780
0 17782 7 1 2 57686 73330
0 17783 7 1 2 87510 17782
0 17784 5 1 1 17783
0 17785 7 1 2 87508 17784
0 17786 5 1 1 17785
0 17787 7 4 2 64502 87233
0 17788 5 2 1 87512
0 17789 7 1 2 73226 87513
0 17790 7 1 2 17786 17789
0 17791 5 1 1 17790
0 17792 7 1 2 17777 17791
0 17793 5 1 1 17792
0 17794 7 1 2 58007 17793
0 17795 5 1 1 17794
0 17796 7 1 2 86103 86853
0 17797 5 1 1 17796
0 17798 7 1 2 17714 17797
0 17799 5 1 1 17798
0 17800 7 1 2 65236 17799
0 17801 5 1 1 17800
0 17802 7 2 2 63228 73656
0 17803 5 1 1 87518
0 17804 7 1 2 65025 87519
0 17805 5 1 1 17804
0 17806 7 1 2 80569 17805
0 17807 5 1 1 17806
0 17808 7 1 2 68615 17807
0 17809 5 1 1 17808
0 17810 7 3 2 58974 73977
0 17811 7 1 2 73657 87520
0 17812 5 1 1 17811
0 17813 7 1 2 17809 17812
0 17814 5 1 1 17813
0 17815 7 1 2 65559 17814
0 17816 5 1 1 17815
0 17817 7 1 2 17801 17816
0 17818 5 1 1 17817
0 17819 7 1 2 67659 17818
0 17820 5 1 1 17819
0 17821 7 2 2 73207 73308
0 17822 5 1 1 87523
0 17823 7 1 2 78157 77145
0 17824 7 1 2 87524 17823
0 17825 5 1 1 17824
0 17826 7 1 2 17820 17825
0 17827 5 1 1 17826
0 17828 7 1 2 82200 17827
0 17829 5 1 1 17828
0 17830 7 2 2 67014 70082
0 17831 7 1 2 59112 74537
0 17832 7 1 2 86945 17831
0 17833 7 1 2 87525 17832
0 17834 5 1 1 17833
0 17835 7 1 2 17829 17834
0 17836 7 1 2 17795 17835
0 17837 5 1 1 17836
0 17838 7 1 2 59334 17837
0 17839 5 1 1 17838
0 17840 7 1 2 17750 17839
0 17841 5 1 1 17840
0 17842 7 1 2 58284 17841
0 17843 5 1 1 17842
0 17844 7 1 2 64693 17843
0 17845 7 1 2 17650 17844
0 17846 5 1 1 17845
0 17847 7 1 2 17392 17846
0 17848 5 1 1 17847
0 17849 7 16 2 64694 66183
0 17850 5 3 1 87527
0 17851 7 1 2 70068 77935
0 17852 5 1 1 17851
0 17853 7 1 2 59550 17852
0 17854 5 1 1 17853
0 17855 7 1 2 87281 17854
0 17856 5 1 1 17855
0 17857 7 1 2 87528 17856
0 17858 5 1 1 17857
0 17859 7 13 2 59996 61573
0 17860 5 8 1 87546
0 17861 7 2 2 80384 76826
0 17862 5 1 1 87567
0 17863 7 1 2 64286 17862
0 17864 5 1 1 17863
0 17865 7 1 2 69840 70627
0 17866 5 2 1 17865
0 17867 7 1 2 77319 87569
0 17868 5 1 1 17867
0 17869 7 1 2 85686 17868
0 17870 5 1 1 17869
0 17871 7 1 2 17864 17870
0 17872 5 1 1 17871
0 17873 7 1 2 87547 17872
0 17874 5 1 1 17873
0 17875 7 1 2 17858 17874
0 17876 5 1 1 17875
0 17877 7 1 2 61250 17876
0 17878 5 1 1 17877
0 17879 7 1 2 65237 16122
0 17880 5 1 1 17879
0 17881 7 1 2 61574 16234
0 17882 7 1 2 17880 17881
0 17883 5 1 1 17882
0 17884 7 1 2 70370 84853
0 17885 5 1 1 17884
0 17886 7 1 2 75283 17885
0 17887 5 1 1 17886
0 17888 7 2 2 62945 75900
0 17889 5 1 1 87571
0 17890 7 1 2 75921 87572
0 17891 5 2 1 17890
0 17892 7 1 2 58008 87573
0 17893 5 1 1 17892
0 17894 7 1 2 83092 17893
0 17895 7 1 2 17887 17894
0 17896 5 1 1 17895
0 17897 7 1 2 66184 17896
0 17898 5 1 1 17897
0 17899 7 1 2 64287 17898
0 17900 5 1 1 17899
0 17901 7 9 2 64695 65874
0 17902 7 1 2 59335 83833
0 17903 5 1 1 17902
0 17904 7 1 2 78252 84039
0 17905 5 1 1 17904
0 17906 7 1 2 84036 81869
0 17907 7 1 2 17905 17906
0 17908 7 1 2 17903 17907
0 17909 5 1 1 17908
0 17910 7 1 2 87575 17909
0 17911 7 1 2 17900 17910
0 17912 7 1 2 17883 17911
0 17913 5 1 1 17912
0 17914 7 1 2 17878 17913
0 17915 5 1 1 17914
0 17916 7 1 2 65560 17915
0 17917 5 1 1 17916
0 17918 7 1 2 80921 9530
0 17919 5 1 1 17918
0 17920 7 1 2 77979 17919
0 17921 5 1 1 17920
0 17922 7 2 2 76181 70628
0 17923 7 1 2 77967 87584
0 17924 5 1 1 17923
0 17925 7 1 2 17921 17924
0 17926 5 1 1 17925
0 17927 7 1 2 60321 17926
0 17928 5 1 1 17927
0 17929 7 2 2 67177 78142
0 17930 7 1 2 79775 87586
0 17931 5 1 1 17930
0 17932 7 1 2 17928 17931
0 17933 5 1 1 17932
0 17934 7 1 2 86461 17933
0 17935 5 1 1 17934
0 17936 7 1 2 67178 77190
0 17937 5 2 1 17936
0 17938 7 1 2 87179 87588
0 17939 5 1 1 17938
0 17940 7 1 2 85469 84172
0 17941 5 2 1 17940
0 17942 7 1 2 82390 87590
0 17943 5 1 1 17942
0 17944 7 1 2 60889 75247
0 17945 7 1 2 17943 17944
0 17946 5 1 1 17945
0 17947 7 1 2 82391 84132
0 17948 5 1 1 17947
0 17949 7 1 2 67179 17948
0 17950 5 1 1 17949
0 17951 7 1 2 17946 17950
0 17952 7 1 2 17939 17951
0 17953 5 1 1 17952
0 17954 7 1 2 61251 77064
0 17955 7 1 2 17953 17954
0 17956 5 1 1 17955
0 17957 7 1 2 17935 17956
0 17958 5 1 1 17957
0 17959 7 1 2 59997 17958
0 17960 5 1 1 17959
0 17961 7 4 2 61252 67322
0 17962 5 2 1 87592
0 17963 7 1 2 87383 87593
0 17964 5 1 1 17963
0 17965 7 1 2 80195 73253
0 17966 5 1 1 17965
0 17967 7 1 2 17964 17966
0 17968 5 1 1 17967
0 17969 7 1 2 68996 17968
0 17970 5 1 1 17969
0 17971 7 1 2 70083 85851
0 17972 5 1 1 17971
0 17973 7 1 2 58009 73254
0 17974 5 1 1 17973
0 17975 7 1 2 17972 17974
0 17976 5 1 1 17975
0 17977 7 1 2 70967 17976
0 17978 5 1 1 17977
0 17979 7 1 2 65875 85905
0 17980 5 1 1 17979
0 17981 7 1 2 17978 17980
0 17982 7 1 2 17970 17981
0 17983 5 1 1 17982
0 17984 7 1 2 59551 17983
0 17985 5 1 1 17984
0 17986 7 2 2 81856 72217
0 17987 5 2 1 87598
0 17988 7 1 2 58010 87600
0 17989 5 1 1 17988
0 17990 7 1 2 58285 75928
0 17991 5 1 1 17990
0 17992 7 1 2 17989 17991
0 17993 5 1 1 17992
0 17994 7 1 2 85531 17993
0 17995 5 1 1 17994
0 17996 7 1 2 70407 75873
0 17997 5 1 1 17996
0 17998 7 1 2 76182 17997
0 17999 5 1 1 17998
0 18000 7 1 2 71735 87082
0 18001 5 1 1 18000
0 18002 7 1 2 87509 73601
0 18003 7 1 2 18001 18002
0 18004 5 1 1 18003
0 18005 7 1 2 17999 18004
0 18006 5 1 1 18005
0 18007 7 1 2 73658 75252
0 18008 7 1 2 85503 18007
0 18009 5 1 1 18008
0 18010 7 1 2 18006 18009
0 18011 7 1 2 17995 18010
0 18012 7 1 2 17985 18011
0 18013 5 1 1 18012
0 18014 7 1 2 87529 18013
0 18015 5 1 1 18014
0 18016 7 1 2 17960 18015
0 18017 7 1 2 17917 18016
0 18018 5 1 1 18017
0 18019 7 1 2 76731 18018
0 18020 5 1 1 18019
0 18021 7 1 2 17848 18020
0 18022 7 1 2 17213 18021
0 18023 5 1 1 18022
0 18024 7 1 2 61916 18023
0 18025 5 1 1 18024
0 18026 7 4 2 72079 71269
0 18027 7 6 2 59998 65876
0 18028 7 2 2 82650 87606
0 18029 5 1 1 87612
0 18030 7 4 2 74653 82095
0 18031 7 1 2 67180 70629
0 18032 7 1 2 87614 18031
0 18033 5 1 1 18032
0 18034 7 1 2 18029 18033
0 18035 5 1 1 18034
0 18036 7 1 2 64503 18035
0 18037 5 1 1 18036
0 18038 7 2 2 61575 79256
0 18039 5 1 1 87618
0 18040 7 2 2 84572 87619
0 18041 5 1 1 87620
0 18042 7 1 2 18037 18041
0 18043 5 1 1 18042
0 18044 7 1 2 63229 18043
0 18045 5 1 1 18044
0 18046 7 10 2 64504 87548
0 18047 5 4 1 87622
0 18048 7 7 2 59778 87530
0 18049 5 2 1 87636
0 18050 7 1 2 87632 87643
0 18051 5 5 1 18050
0 18052 7 2 2 58488 87645
0 18053 5 2 1 87650
0 18054 7 1 2 84573 87651
0 18055 5 1 1 18054
0 18056 7 1 2 18045 18055
0 18057 5 1 1 18056
0 18058 7 1 2 71401 18057
0 18059 5 1 1 18058
0 18060 7 3 2 66185 87172
0 18061 7 1 2 61917 84610
0 18062 7 1 2 87654 18061
0 18063 5 1 1 18062
0 18064 7 1 2 18059 18063
0 18065 5 1 1 18064
0 18066 7 1 2 87602 18065
0 18067 5 1 1 18066
0 18068 7 1 2 58740 18067
0 18069 7 1 2 18025 18068
0 18070 5 1 1 18069
0 18071 7 1 2 17033 18070
0 18072 5 1 1 18071
0 18073 7 7 2 65877 82651
0 18074 7 1 2 82312 87657
0 18075 5 1 1 18074
0 18076 7 1 2 62659 73776
0 18077 7 1 2 70630 18076
0 18078 5 1 1 18077
0 18079 7 1 2 74695 18078
0 18080 5 1 1 18079
0 18081 7 5 2 66571 86327
0 18082 7 1 2 77894 87664
0 18083 7 1 2 18080 18082
0 18084 5 1 1 18083
0 18085 7 1 2 18075 18084
0 18086 5 1 1 18085
0 18087 7 1 2 63481 18086
0 18088 5 1 1 18087
0 18089 7 4 2 58286 73659
0 18090 5 1 1 87669
0 18091 7 1 2 79431 82652
0 18092 7 1 2 87670 18091
0 18093 5 1 1 18092
0 18094 7 1 2 18088 18093
0 18095 5 1 1 18094
0 18096 7 1 2 77853 18095
0 18097 5 1 1 18096
0 18098 7 5 2 64696 75508
0 18099 7 3 2 66572 86462
0 18100 7 1 2 83060 87678
0 18101 7 1 2 87673 18100
0 18102 7 1 2 82733 18101
0 18103 5 1 1 18102
0 18104 7 1 2 18097 18103
0 18105 5 1 1 18104
0 18106 7 1 2 70201 18105
0 18107 5 1 1 18106
0 18108 7 1 2 69525 18107
0 18109 7 1 2 18072 18108
0 18110 5 1 1 18109
0 18111 7 1 2 66755 87283
0 18112 5 1 1 18111
0 18113 7 3 2 62660 79879
0 18114 7 1 2 72080 86013
0 18115 7 1 2 87681 18114
0 18116 5 1 1 18115
0 18117 7 1 2 18112 18116
0 18118 5 1 1 18117
0 18119 7 1 2 61253 18118
0 18120 5 1 1 18119
0 18121 7 6 2 65878 66756
0 18122 7 1 2 59113 80537
0 18123 5 1 1 18122
0 18124 7 1 2 65238 79581
0 18125 5 1 1 18124
0 18126 7 1 2 83625 18125
0 18127 7 1 2 18123 18126
0 18128 5 1 1 18127
0 18129 7 1 2 57687 18128
0 18130 5 1 1 18129
0 18131 7 1 2 72021 86177
0 18132 5 1 1 18131
0 18133 7 1 2 71491 77039
0 18134 7 1 2 77065 18133
0 18135 5 1 1 18134
0 18136 7 1 2 18132 18135
0 18137 7 1 2 18130 18136
0 18138 5 1 1 18137
0 18139 7 1 2 67323 18138
0 18140 5 1 1 18139
0 18141 7 1 2 69417 87404
0 18142 5 1 1 18141
0 18143 7 1 2 76374 77066
0 18144 5 1 1 18143
0 18145 7 1 2 60890 87400
0 18146 5 1 1 18145
0 18147 7 3 2 63871 72190
0 18148 5 3 1 87690
0 18149 7 1 2 87693 77193
0 18150 5 1 1 18149
0 18151 7 1 2 18146 18150
0 18152 7 1 2 18144 18151
0 18153 5 1 1 18152
0 18154 7 1 2 78270 18153
0 18155 5 1 1 18154
0 18156 7 1 2 65561 76972
0 18157 5 1 1 18156
0 18158 7 1 2 77716 18157
0 18159 5 1 1 18158
0 18160 7 1 2 86933 18159
0 18161 5 1 1 18160
0 18162 7 1 2 82000 79017
0 18163 5 1 1 18162
0 18164 7 1 2 71492 78713
0 18165 5 1 1 18164
0 18166 7 1 2 18163 18165
0 18167 5 1 1 18166
0 18168 7 1 2 75326 18167
0 18169 5 1 1 18168
0 18170 7 1 2 18161 18169
0 18171 7 1 2 58011 83528
0 18172 5 1 1 18171
0 18173 7 1 2 83628 18172
0 18174 5 1 1 18173
0 18175 7 1 2 68367 81178
0 18176 7 1 2 18174 18175
0 18177 5 1 1 18176
0 18178 7 1 2 68003 77922
0 18179 5 1 1 18178
0 18180 7 1 2 64288 77538
0 18181 7 1 2 18179 18180
0 18182 5 1 1 18181
0 18183 7 1 2 60891 70408
0 18184 7 1 2 18182 18183
0 18185 5 1 1 18184
0 18186 7 1 2 18177 18185
0 18187 7 1 2 18170 18186
0 18188 7 1 2 18155 18187
0 18189 7 1 2 18142 18188
0 18190 7 1 2 18140 18189
0 18191 5 1 1 18190
0 18192 7 1 2 87684 18191
0 18193 5 1 1 18192
0 18194 7 3 2 64289 85795
0 18195 5 3 1 87696
0 18196 7 2 2 65879 79502
0 18197 5 3 1 87702
0 18198 7 2 2 77946 87704
0 18199 5 1 1 87707
0 18200 7 1 2 87699 18199
0 18201 5 1 1 18200
0 18202 7 1 2 62946 18201
0 18203 5 1 1 18202
0 18204 7 1 2 84527 18203
0 18205 5 1 1 18204
0 18206 7 1 2 67181 18205
0 18207 5 1 1 18206
0 18208 7 5 2 60548 80421
0 18209 7 1 2 87286 87709
0 18210 5 2 1 18209
0 18211 7 1 2 18207 87714
0 18212 5 1 1 18211
0 18213 7 1 2 79880 70631
0 18214 7 1 2 18212 18213
0 18215 5 1 1 18214
0 18216 7 1 2 18193 18215
0 18217 7 1 2 18120 18216
0 18218 5 1 1 18217
0 18219 7 1 2 63230 18218
0 18220 5 1 1 18219
0 18221 7 1 2 77067 87589
0 18222 5 1 1 18221
0 18223 7 1 2 87568 77320
0 18224 5 2 1 18223
0 18225 7 1 2 65562 87716
0 18226 5 1 1 18225
0 18227 7 1 2 61254 18226
0 18228 7 1 2 18222 18227
0 18229 5 1 1 18228
0 18230 7 1 2 75932 75100
0 18231 5 1 1 18230
0 18232 7 1 2 65880 18231
0 18233 7 1 2 70012 86538
0 18234 5 1 1 18233
0 18235 7 1 2 18234 78439
0 18236 7 1 2 18232 18235
0 18237 5 1 1 18236
0 18238 7 1 2 58489 18237
0 18239 7 1 2 18229 18238
0 18240 5 1 1 18239
0 18241 7 1 2 58012 77198
0 18242 5 1 1 18241
0 18243 7 1 2 3422 18242
0 18244 5 1 1 18243
0 18245 7 1 2 74686 18244
0 18246 5 1 1 18245
0 18247 7 1 2 18240 18246
0 18248 5 1 1 18247
0 18249 7 1 2 64290 18248
0 18250 5 1 1 18249
0 18251 7 1 2 77947 80558
0 18252 5 1 1 18251
0 18253 7 1 2 73561 71994
0 18254 7 1 2 80300 18253
0 18255 5 1 1 18254
0 18256 7 1 2 18252 18255
0 18257 5 1 1 18256
0 18258 7 1 2 59552 18257
0 18259 5 1 1 18258
0 18260 7 2 2 65881 77968
0 18261 5 1 1 87718
0 18262 7 1 2 76183 87719
0 18263 5 1 1 18262
0 18264 7 1 2 65239 85949
0 18265 5 1 1 18264
0 18266 7 1 2 85517 18265
0 18267 7 1 2 18263 18266
0 18268 5 1 1 18267
0 18269 7 1 2 85084 18268
0 18270 5 1 1 18269
0 18271 7 1 2 18259 18270
0 18272 5 1 1 18271
0 18273 7 1 2 70632 18272
0 18274 5 1 1 18273
0 18275 7 1 2 80570 85736
0 18276 5 3 1 18275
0 18277 7 3 2 65563 87720
0 18278 5 1 1 87723
0 18279 7 1 2 77317 87724
0 18280 5 1 1 18279
0 18281 7 8 2 62947 65882
0 18282 5 3 1 87726
0 18283 7 1 2 73067 87734
0 18284 5 3 1 18283
0 18285 7 1 2 58490 77068
0 18286 7 1 2 87737 18285
0 18287 5 1 1 18286
0 18288 7 1 2 18280 18287
0 18289 5 1 1 18288
0 18290 7 1 2 67182 18289
0 18291 5 1 1 18290
0 18292 7 2 2 61255 77311
0 18293 7 1 2 75142 86282
0 18294 7 1 2 87740 18293
0 18295 5 1 1 18294
0 18296 7 1 2 18291 18295
0 18297 7 1 2 18274 18296
0 18298 7 1 2 18250 18297
0 18299 5 1 1 18298
0 18300 7 1 2 66757 18299
0 18301 5 1 1 18300
0 18302 7 1 2 18220 18301
0 18303 5 1 1 18302
0 18304 7 1 2 61576 18303
0 18305 5 1 1 18304
0 18306 7 1 2 64291 87130
0 18307 5 1 1 18306
0 18308 7 3 2 64292 72491
0 18309 5 2 1 87742
0 18310 7 1 2 70633 87745
0 18311 7 1 2 77969 18310
0 18312 5 2 1 18311
0 18313 7 1 2 18307 87747
0 18314 5 1 1 18313
0 18315 7 1 2 60322 18314
0 18316 5 1 1 18315
0 18317 7 1 2 64293 76997
0 18318 5 1 1 18317
0 18319 7 1 2 18316 18318
0 18320 5 1 1 18319
0 18321 7 1 2 62948 18320
0 18322 5 1 1 18321
0 18323 7 1 2 78158 77069
0 18324 5 1 1 18323
0 18325 7 1 2 18322 18324
0 18326 5 1 1 18325
0 18327 7 1 2 64024 18326
0 18328 5 1 1 18327
0 18329 7 1 2 72795 77054
0 18330 5 1 1 18329
0 18331 7 1 2 18328 18330
0 18332 5 1 1 18331
0 18333 7 1 2 62661 18332
0 18334 5 1 1 18333
0 18335 7 3 2 65564 70814
0 18336 5 1 1 87749
0 18337 7 1 2 64294 87750
0 18338 7 1 2 70746 18337
0 18339 5 1 1 18338
0 18340 7 1 2 87748 18339
0 18341 5 1 1 18340
0 18342 7 1 2 60323 18341
0 18343 5 1 1 18342
0 18344 7 1 2 64295 87294
0 18345 5 1 1 18344
0 18346 7 1 2 18343 18345
0 18347 5 1 1 18346
0 18348 7 1 2 63231 18347
0 18349 5 1 1 18348
0 18350 7 1 2 18334 18349
0 18351 5 1 1 18350
0 18352 7 1 2 61256 18351
0 18353 5 1 1 18352
0 18354 7 1 2 75437 72761
0 18355 5 1 1 18354
0 18356 7 1 2 1782 18355
0 18357 5 1 1 18356
0 18358 7 1 2 70634 18357
0 18359 5 1 1 18358
0 18360 7 1 2 74015 76990
0 18361 5 1 1 18360
0 18362 7 1 2 18359 18361
0 18363 5 1 1 18362
0 18364 7 1 2 60324 18363
0 18365 5 1 1 18364
0 18366 7 1 2 83682 78125
0 18367 5 1 1 18366
0 18368 7 1 2 18365 18367
0 18369 5 1 1 18368
0 18370 7 1 2 61257 18369
0 18371 5 1 1 18370
0 18372 7 1 2 86724 81003
0 18373 5 1 1 18372
0 18374 7 1 2 18371 18373
0 18375 5 1 1 18374
0 18376 7 1 2 76184 18375
0 18377 5 1 1 18376
0 18378 7 1 2 80863 87244
0 18379 5 1 1 18378
0 18380 7 1 2 72796 72762
0 18381 5 1 1 18380
0 18382 7 1 2 18379 18381
0 18383 5 1 1 18382
0 18384 7 1 2 74837 18383
0 18385 5 1 1 18384
0 18386 7 4 2 64025 72081
0 18387 5 2 1 87752
0 18388 7 5 2 62662 80800
0 18389 7 1 2 87753 87758
0 18390 5 1 1 18389
0 18391 7 1 2 18385 18390
0 18392 5 1 1 18391
0 18393 7 1 2 65883 18392
0 18394 5 1 1 18393
0 18395 7 1 2 18377 18394
0 18396 7 1 2 18353 18395
0 18397 5 1 1 18396
0 18398 7 1 2 18397 82188
0 18399 5 1 1 18398
0 18400 7 1 2 18305 18399
0 18401 5 1 1 18400
0 18402 7 1 2 64505 18401
0 18403 5 1 1 18402
0 18404 7 1 2 63232 78037
0 18405 5 1 1 18404
0 18406 7 1 2 76881 78020
0 18407 5 1 1 18406
0 18408 7 1 2 18405 18407
0 18409 5 1 1 18408
0 18410 7 1 2 70635 18409
0 18411 5 1 1 18410
0 18412 7 2 2 63233 78041
0 18413 5 2 1 87763
0 18414 7 1 2 78066 87764
0 18415 5 1 1 18414
0 18416 7 1 2 18411 18415
0 18417 5 1 1 18416
0 18418 7 1 2 60325 18417
0 18419 5 1 1 18418
0 18420 7 1 2 78664 78143
0 18421 5 1 1 18420
0 18422 7 1 2 64296 78434
0 18423 5 1 1 18422
0 18424 7 1 2 18421 18423
0 18425 5 1 1 18424
0 18426 7 1 2 63234 18425
0 18427 5 1 1 18426
0 18428 7 1 2 18419 18427
0 18429 5 1 1 18428
0 18430 7 1 2 86463 18429
0 18431 5 1 1 18430
0 18432 7 1 2 63235 87717
0 18433 5 1 1 18432
0 18434 7 1 2 76882 77318
0 18435 5 1 1 18434
0 18436 7 1 2 18433 18435
0 18437 5 1 1 18436
0 18438 7 1 2 65565 18437
0 18439 5 1 1 18438
0 18440 7 1 2 63236 77188
0 18441 5 1 1 18440
0 18442 7 1 2 18439 18441
0 18443 5 1 1 18442
0 18444 7 1 2 87180 18443
0 18445 5 1 1 18444
0 18446 7 5 2 65240 81495
0 18447 5 1 1 87767
0 18448 7 2 2 66186 78021
0 18449 5 1 1 87772
0 18450 7 1 2 18447 18449
0 18451 5 1 1 18450
0 18452 7 1 2 85107 18451
0 18453 5 1 1 18452
0 18454 7 3 2 76978 87181
0 18455 5 1 1 87774
0 18456 7 1 2 71807 87775
0 18457 5 1 1 18456
0 18458 7 1 2 18453 18457
0 18459 5 1 1 18458
0 18460 7 1 2 76185 18459
0 18461 5 1 1 18460
0 18462 7 2 2 69741 69841
0 18463 5 1 1 87777
0 18464 7 1 2 74934 18463
0 18465 5 1 1 18464
0 18466 7 4 2 61577 84982
0 18467 7 1 2 18465 87779
0 18468 5 1 1 18467
0 18469 7 5 2 62949 86544
0 18470 7 3 2 60549 81389
0 18471 7 1 2 84723 87788
0 18472 7 1 2 87783 18471
0 18473 5 1 1 18472
0 18474 7 1 2 18468 18473
0 18475 7 1 2 18461 18474
0 18476 5 1 1 18475
0 18477 7 1 2 70636 18476
0 18478 5 1 1 18477
0 18479 7 1 2 86981 82378
0 18480 5 1 1 18479
0 18481 7 1 2 80864 82894
0 18482 5 1 1 18481
0 18483 7 1 2 63237 81376
0 18484 5 1 1 18483
0 18485 7 1 2 18482 18484
0 18486 5 1 1 18485
0 18487 7 1 2 64297 18486
0 18488 5 1 1 18487
0 18489 7 1 2 18480 18488
0 18490 5 1 1 18489
0 18491 7 1 2 77070 18490
0 18492 5 1 1 18491
0 18493 7 1 2 76991 86799
0 18494 7 1 2 76186 18493
0 18495 7 1 2 77312 18494
0 18496 5 1 1 18495
0 18497 7 1 2 18492 18496
0 18498 7 1 2 18478 18497
0 18499 7 1 2 18445 18498
0 18500 5 1 1 18499
0 18501 7 1 2 61258 18500
0 18502 5 1 1 18501
0 18503 7 1 2 18431 18502
0 18504 5 1 1 18503
0 18505 7 1 2 59779 18504
0 18506 5 1 1 18505
0 18507 7 6 2 60892 68230
0 18508 5 4 1 87791
0 18509 7 1 2 73777 87792
0 18510 5 1 1 18509
0 18511 7 1 2 80405 18510
0 18512 5 1 1 18511
0 18513 7 1 2 68499 18512
0 18514 5 1 1 18513
0 18515 7 2 2 60326 84512
0 18516 5 1 1 87801
0 18517 7 1 2 77321 18516
0 18518 5 1 1 18517
0 18519 7 1 2 73619 18518
0 18520 5 1 1 18519
0 18521 7 1 2 18514 18520
0 18522 5 1 1 18521
0 18523 7 3 2 80801 81332
0 18524 5 3 1 87803
0 18525 7 1 2 67183 87804
0 18526 7 1 2 18522 18525
0 18527 5 1 1 18526
0 18528 7 1 2 18506 18527
0 18529 5 1 1 18528
0 18530 7 1 2 66758 18529
0 18531 5 1 1 18530
0 18532 7 1 2 18403 18531
0 18533 5 1 1 18532
0 18534 7 1 2 61918 18533
0 18535 5 1 1 18534
0 18536 7 1 2 69564 18535
0 18537 5 1 1 18536
0 18538 7 7 2 66404 62056
0 18539 7 1 2 67946 87809
0 18540 7 1 2 18537 18539
0 18541 7 1 2 18110 18540
0 18542 5 2 1 18541
0 18543 7 1 2 60171 87816
0 18544 7 1 2 16000 18543
0 18545 5 1 1 18544
0 18546 7 1 2 63657 18545
0 18547 7 1 2 12732 18546
0 18548 5 1 1 18547
0 18549 7 1 2 61763 15857
0 18550 5 1 1 18549
0 18551 7 1 2 18550 87817
0 18552 5 1 1 18551
0 18553 7 1 2 64847 18552
0 18554 5 1 1 18553
0 18555 7 2 2 65884 79881
0 18556 7 4 2 64506 75438
0 18557 5 1 1 87820
0 18558 7 1 2 71270 77797
0 18559 5 1 1 18558
0 18560 7 1 2 18557 18559
0 18561 5 7 1 18560
0 18562 7 1 2 87818 87824
0 18563 5 1 1 18562
0 18564 7 2 2 85075 79567
0 18565 5 1 1 87831
0 18566 7 1 2 61259 87832
0 18567 5 1 1 18566
0 18568 7 1 2 18563 18567
0 18569 5 1 1 18568
0 18570 7 1 2 70488 18569
0 18571 5 1 1 18570
0 18572 7 6 2 60117 61260
0 18573 7 2 2 64697 87833
0 18574 5 1 1 87839
0 18575 7 2 2 79960 80679
0 18576 7 1 2 87840 87841
0 18577 5 1 1 18576
0 18578 7 1 2 18571 18577
0 18579 5 1 1 18578
0 18580 7 1 2 64848 18579
0 18581 5 1 1 18580
0 18582 7 6 2 63238 66759
0 18583 7 3 2 62950 79159
0 18584 5 1 1 87849
0 18585 7 2 2 87843 87850
0 18586 7 5 2 64793 60172
0 18587 7 6 2 63601 87854
0 18588 5 1 1 87859
0 18589 7 2 2 61261 87860
0 18590 7 1 2 87852 87865
0 18591 5 1 1 18590
0 18592 7 1 2 18581 18591
0 18593 5 1 1 18592
0 18594 7 1 2 86542 18593
0 18595 5 1 1 18594
0 18596 7 3 2 77854 79882
0 18597 7 2 2 66573 87867
0 18598 7 6 2 64794 64849
0 18599 7 1 2 69937 87872
0 18600 7 1 2 86623 18599
0 18601 7 1 2 87870 18600
0 18602 5 1 1 18601
0 18603 7 1 2 18595 18602
0 18604 5 1 1 18603
0 18605 7 1 2 61578 18604
0 18606 5 1 1 18605
0 18607 7 1 2 80001 3825
0 18608 5 1 1 18607
0 18609 7 1 2 75933 18608
0 18610 5 1 1 18609
0 18611 7 1 2 17246 18610
0 18612 5 1 1 18611
0 18613 7 1 2 65885 18612
0 18614 5 1 1 18613
0 18615 7 4 2 60327 80422
0 18616 7 1 2 77451 87878
0 18617 5 1 1 18616
0 18618 7 1 2 18614 18617
0 18619 5 1 1 18618
0 18620 7 5 2 79821 76918
0 18621 5 1 1 87882
0 18622 7 1 2 75509 66894
0 18623 5 1 1 18622
0 18624 7 1 2 18621 18623
0 18625 5 5 1 18624
0 18626 7 1 2 18619 87887
0 18627 5 1 1 18626
0 18628 7 1 2 87057 79446
0 18629 5 1 1 18628
0 18630 7 3 2 72859 70905
0 18631 5 1 1 87892
0 18632 7 1 2 77798 87893
0 18633 5 1 1 18632
0 18634 7 1 2 18629 18633
0 18635 5 1 1 18634
0 18636 7 1 2 60328 87682
0 18637 7 1 2 18635 18636
0 18638 5 1 1 18637
0 18639 7 1 2 18627 18638
0 18640 5 1 1 18639
0 18641 7 4 2 64850 66187
0 18642 7 1 2 87895 84220
0 18643 7 1 2 18640 18642
0 18644 5 1 1 18643
0 18645 7 1 2 18606 18644
0 18646 5 1 1 18645
0 18647 7 1 2 62057 18646
0 18648 5 1 1 18647
0 18649 7 6 2 64851 60329
0 18650 7 2 2 79298 87899
0 18651 7 1 2 63761 79160
0 18652 7 1 2 87905 18651
0 18653 7 1 2 86662 18652
0 18654 5 1 1 18653
0 18655 7 1 2 18648 18654
0 18656 5 1 1 18655
0 18657 7 1 2 70984 18656
0 18658 5 1 1 18657
0 18659 7 2 2 60173 61579
0 18660 7 8 2 63482 64507
0 18661 5 2 1 87909
0 18662 7 5 2 87910 83422
0 18663 7 2 2 79299 87919
0 18664 7 3 2 87907 87924
0 18665 5 1 1 87926
0 18666 7 1 2 67952 87927
0 18667 7 1 2 85675 18666
0 18668 5 1 1 18667
0 18669 7 1 2 18658 18668
0 18670 5 1 1 18669
0 18671 7 1 2 61764 18670
0 18672 5 1 1 18671
0 18673 7 1 2 18554 18672
0 18674 5 1 1 18673
0 18675 7 1 2 58906 18674
0 18676 5 1 1 18675
0 18677 7 3 2 78938 78506
0 18678 5 14 1 87929
0 18679 7 2 2 62173 78283
0 18680 5 2 1 87946
0 18681 7 3 2 58013 87948
0 18682 7 1 2 83811 87950
0 18683 5 3 1 18682
0 18684 7 1 2 69675 87953
0 18685 5 1 1 18684
0 18686 7 1 2 85229 83209
0 18687 5 1 1 18686
0 18688 7 1 2 60330 18687
0 18689 5 1 1 18688
0 18690 7 1 2 67583 4808
0 18691 5 1 1 18690
0 18692 7 1 2 18689 18691
0 18693 5 1 1 18692
0 18694 7 1 2 58014 18693
0 18695 5 1 1 18694
0 18696 7 1 2 69199 84514
0 18697 7 1 2 78061 18696
0 18698 7 1 2 78636 18697
0 18699 5 1 1 18698
0 18700 7 1 2 18695 18699
0 18701 5 1 1 18700
0 18702 7 1 2 63872 18701
0 18703 5 1 1 18702
0 18704 7 1 2 62663 10756
0 18705 5 1 1 18704
0 18706 7 1 2 74860 79081
0 18707 5 1 1 18706
0 18708 7 2 2 65026 71017
0 18709 5 1 1 87956
0 18710 7 1 2 68616 87957
0 18711 5 1 1 18710
0 18712 7 1 2 18707 18711
0 18713 5 1 1 18712
0 18714 7 1 2 62380 18713
0 18715 5 1 1 18714
0 18716 7 4 2 62174 58015
0 18717 7 1 2 71677 74579
0 18718 7 1 2 87958 18717
0 18719 5 1 1 18718
0 18720 7 1 2 18715 18719
0 18721 7 1 2 18705 18720
0 18722 7 1 2 18703 18721
0 18723 5 1 1 18722
0 18724 7 1 2 60893 18723
0 18725 5 1 1 18724
0 18726 7 5 2 62175 65241
0 18727 7 1 2 79281 87962
0 18728 5 1 1 18727
0 18729 7 1 2 80513 83266
0 18730 5 1 1 18729
0 18731 7 1 2 62381 18730
0 18732 7 1 2 18728 18731
0 18733 5 1 1 18732
0 18734 7 1 2 78777 84644
0 18735 7 1 2 18733 18734
0 18736 5 1 1 18735
0 18737 7 1 2 18725 18736
0 18738 5 1 1 18737
0 18739 7 1 2 69268 18738
0 18740 5 1 1 18739
0 18741 7 1 2 18685 18740
0 18742 5 1 1 18741
0 18743 7 1 2 87674 18742
0 18744 5 1 1 18743
0 18745 7 4 2 59780 70489
0 18746 7 2 2 62058 87967
0 18747 7 1 2 86993 87971
0 18748 7 1 2 87954 18747
0 18749 5 1 1 18748
0 18750 7 1 2 18744 18749
0 18751 5 1 1 18750
0 18752 7 1 2 66188 18751
0 18753 5 1 1 18752
0 18754 7 1 2 60550 82237
0 18755 5 1 1 18754
0 18756 7 1 2 72722 87963
0 18757 5 1 1 18756
0 18758 7 1 2 18755 18757
0 18759 5 1 1 18758
0 18760 7 1 2 60894 18759
0 18761 5 1 1 18760
0 18762 7 1 2 71028 77194
0 18763 5 1 1 18762
0 18764 7 1 2 18761 18763
0 18765 5 1 1 18764
0 18766 7 1 2 58016 18765
0 18767 5 1 1 18766
0 18768 7 3 2 65027 70589
0 18769 5 1 1 87973
0 18770 7 1 2 78783 87974
0 18771 5 1 1 18770
0 18772 7 1 2 18767 18771
0 18773 5 1 1 18772
0 18774 7 1 2 63873 18773
0 18775 5 1 1 18774
0 18776 7 2 2 62382 87959
0 18777 5 1 1 87976
0 18778 7 1 2 69842 87977
0 18779 5 3 1 18778
0 18780 7 4 2 57688 62664
0 18781 5 2 1 87981
0 18782 7 1 2 83756 87982
0 18783 5 1 1 18782
0 18784 7 1 2 87978 18783
0 18785 5 1 1 18784
0 18786 7 1 2 60895 18785
0 18787 5 1 1 18786
0 18788 7 2 2 59114 78279
0 18789 5 11 1 87987
0 18790 7 1 2 84344 80514
0 18791 7 2 2 87989 18790
0 18792 7 1 2 3794 11827
0 18793 5 1 1 18792
0 18794 7 1 2 71886 18793
0 18795 7 1 2 88000 18794
0 18796 5 1 1 18795
0 18797 7 1 2 18787 18796
0 18798 7 1 2 18775 18797
0 18799 5 1 1 18798
0 18800 7 1 2 69269 18799
0 18801 5 1 1 18800
0 18802 7 1 2 76874 80131
0 18803 5 1 1 18802
0 18804 7 1 2 68695 18803
0 18805 5 1 1 18804
0 18806 7 1 2 62176 18805
0 18807 5 1 1 18806
0 18808 7 1 2 76339 79682
0 18809 7 1 2 69576 73803
0 18810 7 1 2 18808 18809
0 18811 5 1 1 18810
0 18812 7 1 2 18807 18811
0 18813 5 1 1 18812
0 18814 7 1 2 69024 18813
0 18815 5 1 1 18814
0 18816 7 1 2 58017 78280
0 18817 5 1 1 18816
0 18818 7 1 2 69351 18817
0 18819 5 1 1 18818
0 18820 7 1 2 18815 18819
0 18821 7 1 2 18801 18820
0 18822 5 1 1 18821
0 18823 7 1 2 77855 86328
0 18824 7 1 2 18822 18823
0 18825 5 1 1 18824
0 18826 7 1 2 18753 18825
0 18827 5 1 1 18826
0 18828 7 1 2 63483 18827
0 18829 5 1 1 18828
0 18830 7 1 2 87655 87955
0 18831 5 1 1 18830
0 18832 7 17 2 61580 77856
0 18833 7 3 2 57689 77116
0 18834 5 4 1 88019
0 18835 7 3 2 74569 88020
0 18836 5 3 1 88026
0 18837 7 2 2 88002 88029
0 18838 7 1 2 59999 88032
0 18839 5 1 1 18838
0 18840 7 1 2 18831 18839
0 18841 5 1 1 18840
0 18842 7 1 2 79834 18841
0 18843 5 1 1 18842
0 18844 7 1 2 18829 18843
0 18845 5 1 1 18844
0 18846 7 1 2 61262 18845
0 18847 5 1 1 18846
0 18848 7 4 2 76622 79883
0 18849 5 3 1 88034
0 18850 7 1 2 85387 88038
0 18851 5 10 1 18850
0 18852 7 1 2 70490 88041
0 18853 5 2 1 18852
0 18854 7 2 2 63484 60118
0 18855 7 2 2 75510 88053
0 18856 5 1 1 88055
0 18857 7 2 2 64698 88056
0 18858 5 1 1 88057
0 18859 7 3 2 58855 88058
0 18860 5 1 1 88059
0 18861 7 1 2 88051 18860
0 18862 5 1 1 18861
0 18863 7 1 2 83018 79359
0 18864 7 1 2 78705 18863
0 18865 7 1 2 18862 18864
0 18866 5 1 1 18865
0 18867 7 1 2 18847 18866
0 18868 5 1 1 18867
0 18869 7 1 2 64852 18868
0 18870 5 1 1 18869
0 18871 7 1 2 61263 88033
0 18872 5 1 1 18871
0 18873 7 2 2 71678 70293
0 18874 5 2 1 88062
0 18875 7 1 2 65886 88064
0 18876 5 2 1 18875
0 18877 7 1 2 62383 88066
0 18878 5 1 1 18877
0 18879 7 1 2 15458 18878
0 18880 5 1 1 18879
0 18881 7 1 2 62177 18880
0 18882 5 1 1 18881
0 18883 7 2 2 61264 69025
0 18884 5 4 1 88068
0 18885 7 1 2 62384 88069
0 18886 5 1 1 18885
0 18887 7 1 2 65887 79369
0 18888 5 2 1 18887
0 18889 7 1 2 77661 88074
0 18890 5 1 1 18889
0 18891 7 1 2 18886 18890
0 18892 7 1 2 18882 18891
0 18893 5 1 1 18892
0 18894 7 1 2 87443 18893
0 18895 5 1 1 18894
0 18896 7 1 2 18872 18895
0 18897 5 1 1 18896
0 18898 7 2 2 62059 18897
0 18899 7 5 2 64795 79233
0 18900 7 1 2 64699 60174
0 18901 7 3 2 88078 18900
0 18902 5 1 1 88083
0 18903 7 1 2 88076 88084
0 18904 5 1 1 18903
0 18905 7 1 2 18870 18904
0 18906 5 1 1 18905
0 18907 7 1 2 63658 18906
0 18908 5 1 1 18907
0 18909 7 5 2 63602 58907
0 18910 7 6 2 87873 88086
0 18911 5 1 1 88091
0 18912 7 3 2 66760 88092
0 18913 5 1 1 88097
0 18914 7 1 2 88077 88098
0 18915 5 1 1 18914
0 18916 7 1 2 18908 18915
0 18917 5 1 1 18916
0 18918 7 1 2 66574 18917
0 18919 5 1 1 18918
0 18920 7 4 2 86060 88003
0 18921 7 1 2 80504 7149
0 18922 5 1 1 18921
0 18923 7 1 2 74371 84417
0 18924 5 1 1 18923
0 18925 7 1 2 83274 18924
0 18926 7 1 2 18922 18925
0 18927 5 1 1 18926
0 18928 7 1 2 88100 18927
0 18929 5 1 1 18928
0 18930 7 1 2 64796 88042
0 18931 5 1 1 18930
0 18932 7 1 2 18858 18931
0 18933 5 1 1 18932
0 18934 7 1 2 63603 18933
0 18935 5 1 1 18934
0 18936 7 3 2 64797 79198
0 18937 7 1 2 87844 88104
0 18938 5 1 1 18937
0 18939 7 1 2 18935 18938
0 18940 5 6 1 18939
0 18941 7 2 2 78284 69887
0 18942 5 1 1 88113
0 18943 7 1 2 78340 88114
0 18944 5 1 1 18943
0 18945 7 1 2 60551 18944
0 18946 5 1 1 18945
0 18947 7 1 2 80163 9388
0 18948 5 1 1 18947
0 18949 7 1 2 65242 18948
0 18950 5 1 1 18949
0 18951 7 1 2 71041 74585
0 18952 5 1 1 18951
0 18953 7 1 2 18950 18952
0 18954 7 1 2 18946 18953
0 18955 5 1 1 18954
0 18956 7 1 2 66189 18955
0 18957 7 1 2 88107 18956
0 18958 5 1 1 18957
0 18959 7 1 2 18929 18958
0 18960 5 1 1 18959
0 18961 7 1 2 60896 18960
0 18962 5 1 1 18961
0 18963 7 1 2 68823 88101
0 18964 5 1 1 18963
0 18965 7 2 2 63762 66190
0 18966 7 1 2 62178 88115
0 18967 7 1 2 88108 18966
0 18968 5 1 1 18967
0 18969 7 1 2 18964 18968
0 18970 5 1 1 18969
0 18971 7 1 2 77662 18970
0 18972 5 1 1 18971
0 18973 7 1 2 67817 88102
0 18974 5 1 1 18973
0 18975 7 1 2 18972 18974
0 18976 5 1 1 18975
0 18977 7 1 2 65566 18976
0 18978 5 1 1 18977
0 18979 7 1 2 18962 18978
0 18980 5 1 1 18979
0 18981 7 20 2 63659 64853
0 18982 5 4 1 88117
0 18983 7 14 2 66685 88118
0 18984 7 1 2 72967 88141
0 18985 7 1 2 18980 18984
0 18986 5 1 1 18985
0 18987 7 1 2 18919 18986
0 18988 5 1 1 18987
0 18989 7 1 2 64026 18988
0 18990 5 1 1 18989
0 18991 7 2 2 62060 88030
0 18992 7 1 2 88099 88155
0 18993 5 1 1 18992
0 18994 7 1 2 64854 79971
0 18995 5 1 1 18994
0 18996 7 1 2 18902 18995
0 18997 5 2 1 18996
0 18998 7 1 2 88156 88157
0 18999 5 1 1 18998
0 19000 7 3 2 60552 83300
0 19001 5 1 1 88159
0 19002 7 1 2 75291 88160
0 19003 5 1 1 19002
0 19004 7 2 2 67743 77089
0 19005 5 4 1 88162
0 19006 7 1 2 65243 88163
0 19007 5 1 1 19006
0 19008 7 1 2 62665 19007
0 19009 7 1 2 19003 19008
0 19010 5 1 1 19009
0 19011 7 1 2 58018 75292
0 19012 5 2 1 19011
0 19013 7 2 2 69243 74167
0 19014 7 1 2 64855 66761
0 19015 7 1 2 73411 19014
0 19016 7 1 2 88170 19015
0 19017 7 1 2 88168 19016
0 19018 7 1 2 19010 19017
0 19019 5 1 1 19018
0 19020 7 1 2 18999 19019
0 19021 5 1 1 19020
0 19022 7 1 2 63660 19021
0 19023 5 1 1 19022
0 19024 7 1 2 18993 19023
0 19025 5 1 1 19024
0 19026 7 1 2 88004 19025
0 19027 5 1 1 19026
0 19028 7 2 2 71887 72198
0 19029 5 2 1 88172
0 19030 7 1 2 87951 88173
0 19031 5 1 1 19030
0 19032 7 5 2 62061 19031
0 19033 7 1 2 79950 88176
0 19034 5 1 1 19033
0 19035 7 1 2 67922 88177
0 19036 5 1 1 19035
0 19037 7 2 2 65244 71770
0 19038 5 1 1 88181
0 19039 7 7 2 72723 77146
0 19040 5 1 1 88183
0 19041 7 1 2 57690 68824
0 19042 5 1 1 19041
0 19043 7 2 2 19040 19042
0 19044 5 4 1 88190
0 19045 7 1 2 60553 88191
0 19046 5 1 1 19045
0 19047 7 1 2 65245 78364
0 19048 5 1 1 19047
0 19049 7 1 2 63874 19048
0 19050 7 1 2 19046 19049
0 19051 5 1 1 19050
0 19052 7 1 2 19038 19051
0 19053 5 1 1 19052
0 19054 7 2 2 62666 63604
0 19055 7 1 2 80020 88196
0 19056 7 1 2 19053 19055
0 19057 5 1 1 19056
0 19058 7 1 2 19036 19057
0 19059 5 1 1 19058
0 19060 7 1 2 66762 19059
0 19061 5 1 1 19060
0 19062 7 1 2 19034 19061
0 19063 5 1 1 19062
0 19064 7 1 2 75511 19063
0 19065 5 1 1 19064
0 19066 7 1 2 70491 88035
0 19067 7 1 2 88178 19066
0 19068 5 1 1 19067
0 19069 7 1 2 19065 19068
0 19070 5 1 1 19069
0 19071 7 1 2 64856 19070
0 19072 5 1 1 19071
0 19073 7 4 2 64700 87855
0 19074 7 2 2 87920 88198
0 19075 5 1 1 88202
0 19076 7 1 2 88179 88203
0 19077 5 1 1 19076
0 19078 7 1 2 19072 19077
0 19079 5 1 1 19078
0 19080 7 1 2 63661 19079
0 19081 5 1 1 19080
0 19082 7 2 2 58908 87874
0 19083 7 4 2 87921 88204
0 19084 5 1 1 88206
0 19085 7 3 2 64701 88207
0 19086 5 1 1 88210
0 19087 7 1 2 88211 88180
0 19088 5 1 1 19087
0 19089 7 1 2 19081 19088
0 19090 5 1 1 19089
0 19091 7 1 2 66191 19090
0 19092 5 1 1 19091
0 19093 7 1 2 19027 19092
0 19094 5 1 1 19093
0 19095 7 1 2 60897 19094
0 19096 5 1 1 19095
0 19097 7 4 2 59336 64857
0 19098 7 1 2 82871 69244
0 19099 7 1 2 88213 19098
0 19100 7 1 2 63662 64702
0 19101 7 1 2 73544 19100
0 19102 7 1 2 79241 19101
0 19103 7 1 2 19099 19102
0 19104 7 1 2 78458 19103
0 19105 5 1 1 19104
0 19106 7 1 2 66575 19105
0 19107 7 1 2 19096 19106
0 19108 5 1 1 19107
0 19109 7 1 2 72144 74598
0 19110 5 1 1 19109
0 19111 7 2 2 71679 74871
0 19112 5 1 1 88217
0 19113 7 1 2 65567 88218
0 19114 5 1 1 19113
0 19115 7 1 2 19110 19114
0 19116 5 1 1 19115
0 19117 7 1 2 62179 19116
0 19118 5 1 1 19117
0 19119 7 5 2 65028 72145
0 19120 5 1 1 88219
0 19121 7 1 2 77490 88220
0 19122 5 1 1 19121
0 19123 7 4 2 72082 83251
0 19124 7 1 2 62667 88224
0 19125 5 1 1 19124
0 19126 7 1 2 19122 19125
0 19127 7 1 2 19118 19126
0 19128 5 1 1 19127
0 19129 7 1 2 62385 19128
0 19130 5 1 1 19129
0 19131 7 1 2 68825 88225
0 19132 5 1 1 19131
0 19133 7 1 2 63875 77305
0 19134 7 1 2 80071 19133
0 19135 5 2 1 19134
0 19136 7 1 2 19132 88228
0 19137 5 1 1 19136
0 19138 7 1 2 62668 19137
0 19139 5 1 1 19138
0 19140 7 1 2 19130 19139
0 19141 5 1 1 19140
0 19142 7 2 2 88005 19141
0 19143 7 1 2 85199 88230
0 19144 5 1 1 19143
0 19145 7 1 2 85871 86301
0 19146 5 1 1 19145
0 19147 7 1 2 68771 67856
0 19148 5 2 1 19147
0 19149 7 2 2 77663 88232
0 19150 5 1 1 88234
0 19151 7 17 2 60898 61581
0 19152 7 2 2 66827 88236
0 19153 7 1 2 88235 88253
0 19154 5 1 1 19153
0 19155 7 1 2 70168 86302
0 19156 7 1 2 74572 19155
0 19157 5 1 1 19156
0 19158 7 1 2 19154 19157
0 19159 5 1 1 19158
0 19160 7 1 2 65029 19159
0 19161 5 1 1 19160
0 19162 7 1 2 19146 19161
0 19163 5 1 1 19162
0 19164 7 1 2 65246 19163
0 19165 5 1 1 19164
0 19166 7 5 2 65030 74813
0 19167 5 2 1 88255
0 19168 7 1 2 84557 88260
0 19169 5 1 1 19168
0 19170 7 1 2 78567 2335
0 19171 5 1 1 19170
0 19172 7 1 2 62180 74872
0 19173 7 1 2 19171 19172
0 19174 5 1 1 19173
0 19175 7 1 2 19169 19174
0 19176 5 1 1 19175
0 19177 7 15 2 58741 61582
0 19178 5 5 1 88262
0 19179 7 1 2 82362 88263
0 19180 7 1 2 19176 19179
0 19181 5 1 1 19180
0 19182 7 1 2 19165 19181
0 19183 5 1 1 19182
0 19184 7 1 2 64798 77857
0 19185 7 1 2 19183 19184
0 19186 5 1 1 19185
0 19187 7 1 2 19144 19186
0 19188 5 1 1 19187
0 19189 7 1 2 63605 19188
0 19190 5 1 1 19189
0 19191 7 5 2 79961 79300
0 19192 7 1 2 88282 88231
0 19193 5 1 1 19192
0 19194 7 1 2 19190 19193
0 19195 5 1 1 19194
0 19196 7 1 2 66686 19195
0 19197 5 1 1 19196
0 19198 7 1 2 85093 87335
0 19199 5 1 1 19198
0 19200 7 1 2 87652 19199
0 19201 5 1 1 19200
0 19202 7 1 2 58742 19201
0 19203 5 1 1 19202
0 19204 7 4 2 66192 76919
0 19205 7 1 2 79257 88287
0 19206 5 1 1 19205
0 19207 7 1 2 19203 19206
0 19208 5 1 1 19207
0 19209 7 2 2 62062 77071
0 19210 7 1 2 67923 88291
0 19211 7 1 2 19208 19210
0 19212 5 1 1 19211
0 19213 7 1 2 64858 19212
0 19214 7 1 2 19197 19213
0 19215 5 1 1 19214
0 19216 7 2 2 88103 88292
0 19217 5 1 1 88293
0 19218 7 1 2 60175 19217
0 19219 5 1 1 19218
0 19220 7 1 2 63663 19219
0 19221 7 1 2 19215 19220
0 19222 5 1 1 19221
0 19223 7 20 2 58909 60176
0 19224 5 4 1 88295
0 19225 7 26 2 88137 88315
0 19226 5 1 1 88319
0 19227 7 2 2 83019 88320
0 19228 7 1 2 77072 88345
0 19229 5 1 1 19228
0 19230 7 22 2 64859 66687
0 19231 7 12 2 63664 88347
0 19232 7 1 2 61583 86337
0 19233 5 1 1 19232
0 19234 7 1 2 75127 81466
0 19235 7 1 2 77727 19234
0 19236 5 1 1 19235
0 19237 7 1 2 19233 19236
0 19238 5 1 1 19237
0 19239 7 1 2 65568 19238
0 19240 5 1 1 19239
0 19241 7 1 2 74333 72191
0 19242 5 1 1 19241
0 19243 7 1 2 69767 19242
0 19244 5 1 1 19243
0 19245 7 1 2 62181 19244
0 19246 5 1 1 19245
0 19247 7 1 2 78285 74964
0 19248 5 1 1 19247
0 19249 7 1 2 19246 19248
0 19250 5 1 1 19249
0 19251 7 1 2 63876 19250
0 19252 5 1 1 19251
0 19253 7 1 2 74334 83460
0 19254 5 1 1 19253
0 19255 7 1 2 19252 19254
0 19256 5 1 1 19255
0 19257 7 1 2 81390 19256
0 19258 5 1 1 19257
0 19259 7 1 2 19240 19258
0 19260 5 1 1 19259
0 19261 7 1 2 88369 19260
0 19262 5 1 1 19261
0 19263 7 1 2 19229 19262
0 19264 5 1 1 19263
0 19265 7 1 2 88109 19264
0 19266 5 1 1 19265
0 19267 7 12 2 58910 64860
0 19268 7 1 2 88381 88294
0 19269 5 1 1 19268
0 19270 7 1 2 61919 19269
0 19271 7 1 2 19266 19270
0 19272 7 1 2 19222 19271
0 19273 5 1 1 19272
0 19274 7 1 2 61265 19273
0 19275 7 1 2 19108 19274
0 19276 5 1 1 19275
0 19277 7 1 2 18990 19276
0 19278 5 1 1 19277
0 19279 7 1 2 66405 19278
0 19280 5 1 1 19279
0 19281 7 9 2 61266 61765
0 19282 7 7 2 61920 86061
0 19283 7 1 2 79755 88402
0 19284 5 1 1 19283
0 19285 7 1 2 69526 74006
0 19286 7 1 2 81729 19285
0 19287 5 1 1 19286
0 19288 7 1 2 19284 19287
0 19289 5 1 1 19288
0 19290 7 2 2 82538 19289
0 19291 7 2 2 71123 72667
0 19292 5 1 1 88411
0 19293 7 1 2 88409 88412
0 19294 5 1 1 19293
0 19295 7 4 2 64508 68004
0 19296 7 1 2 88410 88413
0 19297 5 1 1 19296
0 19298 7 1 2 60331 83900
0 19299 5 1 1 19298
0 19300 7 1 2 77664 75021
0 19301 5 1 1 19300
0 19302 7 1 2 19299 19301
0 19303 5 1 1 19302
0 19304 7 1 2 68826 19303
0 19305 5 1 1 19304
0 19306 7 1 2 76905 75407
0 19307 5 1 1 19306
0 19308 7 1 2 77665 19307
0 19309 5 1 1 19308
0 19310 7 1 2 73291 86417
0 19311 5 1 1 19310
0 19312 7 2 2 19309 19311
0 19313 5 1 1 88417
0 19314 7 1 2 65569 19313
0 19315 5 1 1 19314
0 19316 7 2 2 74023 84564
0 19317 5 2 1 88419
0 19318 7 1 2 68082 88421
0 19319 5 2 1 19318
0 19320 7 1 2 15749 88423
0 19321 5 1 1 19320
0 19322 7 1 2 60899 19321
0 19323 5 1 1 19322
0 19324 7 1 2 19315 19323
0 19325 7 1 2 19305 19324
0 19326 5 1 1 19325
0 19327 7 1 2 79238 71066
0 19328 7 1 2 10086 19327
0 19329 7 1 2 79871 19328
0 19330 7 1 2 19326 19329
0 19331 5 1 1 19330
0 19332 7 1 2 57412 78198
0 19333 5 1 1 19332
0 19334 7 1 2 62669 75491
0 19335 5 1 1 19334
0 19336 7 2 2 70923 79282
0 19337 5 1 1 88425
0 19338 7 1 2 19335 19337
0 19339 7 1 2 19333 19338
0 19340 5 6 1 19339
0 19341 7 1 2 59337 88427
0 19342 5 2 1 19341
0 19343 7 2 2 57691 87097
0 19344 5 1 1 88435
0 19345 7 1 2 64027 88436
0 19346 5 1 1 19345
0 19347 7 1 2 88433 19346
0 19348 5 1 1 19347
0 19349 7 1 2 71808 19348
0 19350 5 1 1 19349
0 19351 7 1 2 79286 74586
0 19352 5 1 1 19351
0 19353 7 3 2 62670 71888
0 19354 5 1 1 88437
0 19355 7 1 2 76455 88438
0 19356 5 1 1 19355
0 19357 7 1 2 19352 19356
0 19358 5 1 1 19357
0 19359 7 1 2 57692 19358
0 19360 5 2 1 19359
0 19361 7 1 2 62386 87098
0 19362 5 1 1 19361
0 19363 7 1 2 58019 76451
0 19364 5 1 1 19363
0 19365 7 1 2 19362 19364
0 19366 5 1 1 19365
0 19367 7 1 2 74587 19366
0 19368 5 2 1 19367
0 19369 7 1 2 62182 75480
0 19370 5 2 1 19369
0 19371 7 1 2 71889 88444
0 19372 5 1 1 19371
0 19373 7 1 2 76316 19372
0 19374 5 1 1 19373
0 19375 7 1 2 88442 19374
0 19376 7 1 2 88440 19375
0 19377 5 1 1 19376
0 19378 7 1 2 64028 19377
0 19379 5 1 1 19378
0 19380 7 1 2 19350 19379
0 19381 5 1 1 19380
0 19382 7 1 2 66962 19381
0 19383 5 1 1 19382
0 19384 7 3 2 77173 71781
0 19385 5 1 1 88446
0 19386 7 1 2 88424 19385
0 19387 5 1 1 19386
0 19388 7 1 2 67041 19387
0 19389 5 1 1 19388
0 19390 7 1 2 60900 19389
0 19391 7 1 2 19383 19390
0 19392 5 1 1 19391
0 19393 7 1 2 75408 83579
0 19394 5 1 1 19393
0 19395 7 1 2 62387 19394
0 19396 5 1 1 19395
0 19397 7 1 2 64029 84730
0 19398 5 1 1 19397
0 19399 7 1 2 19396 19398
0 19400 5 1 1 19399
0 19401 7 1 2 68827 19400
0 19402 5 1 1 19401
0 19403 7 1 2 88418 19402
0 19404 5 1 1 19403
0 19405 7 1 2 67042 19404
0 19406 5 1 1 19405
0 19407 7 1 2 77208 76789
0 19408 7 1 2 78459 19407
0 19409 5 1 1 19408
0 19410 7 1 2 65570 19409
0 19411 7 1 2 19406 19410
0 19412 5 1 1 19411
0 19413 7 3 2 64703 79234
0 19414 7 1 2 19412 88449
0 19415 7 1 2 19392 19414
0 19416 5 1 1 19415
0 19417 7 1 2 19331 19416
0 19418 5 1 1 19417
0 19419 7 1 2 66193 19418
0 19420 5 1 1 19419
0 19421 7 2 2 82443 81496
0 19422 5 1 1 88452
0 19423 7 1 2 67112 88453
0 19424 5 1 1 19423
0 19425 7 4 2 60119 82653
0 19426 7 1 2 73112 88454
0 19427 5 1 1 19426
0 19428 7 1 2 19424 19427
0 19429 5 1 1 19428
0 19430 7 1 2 57413 19429
0 19431 5 1 1 19430
0 19432 7 1 2 81391 81482
0 19433 7 1 2 84762 19432
0 19434 5 1 1 19433
0 19435 7 1 2 19431 19434
0 19436 5 1 1 19435
0 19437 7 1 2 63606 19436
0 19438 5 1 1 19437
0 19439 7 2 2 57414 82654
0 19440 7 1 2 71959 77386
0 19441 7 1 2 88458 19440
0 19442 5 1 1 19441
0 19443 7 1 2 19438 19442
0 19444 5 1 1 19443
0 19445 7 1 2 66763 19444
0 19446 5 1 1 19445
0 19447 7 1 2 61921 81392
0 19448 7 1 2 80345 19447
0 19449 7 1 2 82766 19448
0 19450 5 1 1 19449
0 19451 7 1 2 19446 19450
0 19452 5 1 1 19451
0 19453 7 1 2 71736 19452
0 19454 5 1 1 19453
0 19455 7 1 2 75736 76790
0 19456 7 1 2 87768 19455
0 19457 7 1 2 71368 76100
0 19458 7 1 2 19456 19457
0 19459 5 1 1 19458
0 19460 7 1 2 19454 19459
0 19461 7 1 2 19420 19460
0 19462 5 1 1 19461
0 19463 7 1 2 59781 19462
0 19464 5 1 1 19463
0 19465 7 1 2 19297 19464
0 19466 5 1 1 19465
0 19467 7 1 2 58491 19466
0 19468 5 1 1 19467
0 19469 7 1 2 19294 19468
0 19470 5 1 1 19469
0 19471 7 1 2 66688 19470
0 19472 5 1 1 19471
0 19473 7 9 2 66576 79972
0 19474 7 1 2 76403 88460
0 19475 5 1 1 19474
0 19476 7 1 2 68932 83558
0 19477 5 1 1 19476
0 19478 7 1 2 19475 19477
0 19479 5 1 1 19478
0 19480 7 2 2 76623 83020
0 19481 7 1 2 19479 88469
0 19482 5 1 1 19481
0 19483 7 1 2 19472 19482
0 19484 5 1 1 19483
0 19485 7 1 2 64861 19484
0 19486 5 1 1 19485
0 19487 7 1 2 66963 76404
0 19488 5 1 1 19487
0 19489 7 1 2 68942 19488
0 19490 5 1 1 19489
0 19491 7 1 2 63607 19490
0 19492 5 1 1 19491
0 19493 7 1 2 70451 68933
0 19494 5 1 1 19493
0 19495 7 1 2 19492 19494
0 19496 5 1 1 19495
0 19497 7 1 2 66764 19496
0 19498 5 1 1 19497
0 19499 7 1 2 83383 82355
0 19500 5 1 1 19499
0 19501 7 1 2 19498 19500
0 19502 5 1 1 19501
0 19503 7 2 2 83021 19502
0 19504 7 3 2 60177 76624
0 19505 7 1 2 88471 88473
0 19506 5 1 1 19505
0 19507 7 1 2 19486 19506
0 19508 5 1 1 19507
0 19509 7 1 2 63665 19508
0 19510 5 1 1 19509
0 19511 7 1 2 76625 88382
0 19512 7 1 2 88472 19511
0 19513 5 1 1 19512
0 19514 7 2 2 74024 75262
0 19515 5 1 1 88476
0 19516 7 1 2 60554 88477
0 19517 5 1 1 19516
0 19518 7 1 2 80688 75158
0 19519 7 1 2 19517 19518
0 19520 5 1 1 19519
0 19521 7 1 2 19354 19520
0 19522 5 1 1 19521
0 19523 7 1 2 79347 19522
0 19524 5 1 1 19523
0 19525 7 5 2 65571 77147
0 19526 5 1 1 88478
0 19527 7 1 2 72006 79654
0 19528 7 1 2 88479 19527
0 19529 5 1 1 19528
0 19530 7 1 2 19524 19529
0 19531 5 1 1 19530
0 19532 7 1 2 57693 19531
0 19533 5 1 1 19532
0 19534 7 1 2 80312 88184
0 19535 5 1 1 19534
0 19536 7 1 2 64030 84090
0 19537 5 1 1 19536
0 19538 7 1 2 82746 19537
0 19539 5 1 1 19538
0 19540 7 3 2 78315 87952
0 19541 5 3 1 88483
0 19542 7 1 2 59338 88484
0 19543 5 2 1 19542
0 19544 7 1 2 63877 88489
0 19545 7 1 2 19539 19544
0 19546 5 1 1 19545
0 19547 7 1 2 19535 19546
0 19548 5 1 1 19547
0 19549 7 1 2 60901 19548
0 19550 5 1 1 19549
0 19551 7 3 2 65572 78345
0 19552 7 1 2 84558 88491
0 19553 5 1 1 19552
0 19554 7 1 2 19550 19553
0 19555 5 1 1 19554
0 19556 7 1 2 59782 19555
0 19557 5 1 1 19556
0 19558 7 1 2 19533 19557
0 19559 5 1 1 19558
0 19560 7 1 2 63239 19559
0 19561 5 1 1 19560
0 19562 7 2 2 59115 88192
0 19563 5 1 1 88494
0 19564 7 2 2 69323 67594
0 19565 5 2 1 88496
0 19566 7 1 2 19563 88498
0 19567 5 1 1 19566
0 19568 7 1 2 64031 19567
0 19569 5 1 1 19568
0 19570 7 2 2 62671 18769
0 19571 5 4 1 88500
0 19572 7 1 2 64032 88501
0 19573 5 1 1 19572
0 19574 7 2 2 88490 19573
0 19575 7 1 2 63878 88506
0 19576 5 1 1 19575
0 19577 7 1 2 19569 19576
0 19578 5 1 1 19577
0 19579 7 1 2 60902 19578
0 19580 5 1 1 19579
0 19581 7 1 2 75128 88492
0 19582 5 1 1 19581
0 19583 7 1 2 19580 19582
0 19584 5 1 1 19583
0 19585 7 1 2 60555 19584
0 19586 5 1 1 19585
0 19587 7 1 2 63879 88193
0 19588 5 1 1 19587
0 19589 7 1 2 87985 19588
0 19590 5 1 1 19589
0 19591 7 1 2 71890 73113
0 19592 7 1 2 19590 19591
0 19593 5 1 1 19592
0 19594 7 1 2 19586 19593
0 19595 5 1 1 19594
0 19596 7 1 2 77817 19595
0 19597 5 1 1 19596
0 19598 7 1 2 19561 19597
0 19599 5 1 1 19598
0 19600 7 3 2 63666 69527
0 19601 7 3 2 88508 88348
0 19602 7 1 2 19599 88511
0 19603 5 1 1 19602
0 19604 7 1 2 69528 88321
0 19605 5 1 1 19604
0 19606 7 6 2 67924 88119
0 19607 5 2 1 88514
0 19608 7 1 2 19605 88520
0 19609 5 18 1 19608
0 19610 7 10 2 62063 88522
0 19611 7 1 2 70202 77858
0 19612 7 1 2 88540 19611
0 19613 5 1 1 19612
0 19614 7 1 2 19603 19613
0 19615 5 1 1 19614
0 19616 7 1 2 61584 19615
0 19617 5 1 1 19616
0 19618 7 13 2 66194 75512
0 19619 7 1 2 72047 88541
0 19620 5 1 1 19619
0 19621 7 2 2 57694 79283
0 19622 5 1 1 88563
0 19623 7 1 2 81939 19622
0 19624 5 1 1 19623
0 19625 7 2 2 62183 19624
0 19626 5 1 1 88565
0 19627 7 1 2 78286 78336
0 19628 5 2 1 19627
0 19629 7 4 2 62388 58020
0 19630 5 1 1 88569
0 19631 7 1 2 88567 19630
0 19632 7 1 2 19626 19631
0 19633 5 2 1 19632
0 19634 7 1 2 74588 88573
0 19635 5 1 1 19634
0 19636 7 1 2 5175 19344
0 19637 5 1 1 19636
0 19638 7 1 2 71809 19637
0 19639 5 1 1 19638
0 19640 7 1 2 74873 76456
0 19641 7 1 2 86139 19640
0 19642 5 1 1 19641
0 19643 7 1 2 19642 87979
0 19644 7 1 2 19639 19643
0 19645 7 1 2 19635 19644
0 19646 5 1 1 19645
0 19647 7 4 2 64862 60903
0 19648 7 3 2 66689 88575
0 19649 7 4 2 63667 88579
0 19650 7 1 2 69529 88582
0 19651 7 1 2 19646 19650
0 19652 5 1 1 19651
0 19653 7 1 2 19620 19652
0 19654 5 1 1 19653
0 19655 7 1 2 64033 19654
0 19656 5 1 1 19655
0 19657 7 3 2 63763 72022
0 19658 5 2 1 88586
0 19659 7 1 2 81018 88587
0 19660 5 1 1 19659
0 19661 7 1 2 72283 88428
0 19662 5 1 1 19661
0 19663 7 1 2 19660 19662
0 19664 5 1 1 19663
0 19665 7 1 2 71810 88512
0 19666 7 1 2 19664 19665
0 19667 5 1 1 19666
0 19668 7 1 2 19656 19667
0 19669 5 1 1 19668
0 19670 7 1 2 88550 19669
0 19671 5 1 1 19670
0 19672 7 1 2 19617 19671
0 19673 5 1 1 19672
0 19674 7 1 2 66577 19673
0 19675 5 1 1 19674
0 19676 7 19 2 62064 88322
0 19677 7 3 2 58492 87257
0 19678 5 4 1 88610
0 19679 7 2 2 63240 87336
0 19680 5 4 1 88617
0 19681 7 1 2 88613 88619
0 19682 5 1 1 19681
0 19683 7 2 2 60904 19682
0 19684 5 1 1 88623
0 19685 7 1 2 88591 88624
0 19686 5 1 1 19685
0 19687 7 2 2 60556 76958
0 19688 5 1 1 88625
0 19689 7 1 2 88169 88626
0 19690 5 1 1 19689
0 19691 7 1 2 58021 75783
0 19692 5 4 1 19691
0 19693 7 1 2 60332 88627
0 19694 5 1 1 19693
0 19695 7 1 2 83079 84731
0 19696 5 1 1 19695
0 19697 7 1 2 19694 19696
0 19698 5 1 1 19697
0 19699 7 1 2 64034 19698
0 19700 5 1 1 19699
0 19701 7 1 2 19690 19700
0 19702 5 1 1 19701
0 19703 7 1 2 65573 19702
0 19704 5 1 1 19703
0 19705 7 1 2 83187 5768
0 19706 5 1 1 19705
0 19707 7 1 2 60905 19706
0 19708 5 1 1 19707
0 19709 7 1 2 72146 77177
0 19710 5 2 1 19709
0 19711 7 1 2 19708 88631
0 19712 7 1 2 19704 19711
0 19713 5 1 1 19712
0 19714 7 1 2 87444 19713
0 19715 5 1 1 19714
0 19716 7 1 2 68828 75003
0 19717 7 1 2 86428 19716
0 19718 5 2 1 19717
0 19719 7 2 2 64035 80356
0 19720 5 1 1 88635
0 19721 7 1 2 88633 19720
0 19722 5 1 1 19721
0 19723 7 1 2 62389 19722
0 19724 5 1 1 19723
0 19725 7 1 2 70778 83210
0 19726 5 1 1 19725
0 19727 7 1 2 76906 74981
0 19728 7 1 2 19726 19727
0 19729 5 1 1 19728
0 19730 7 1 2 62672 79539
0 19731 5 1 1 19730
0 19732 7 1 2 78795 19731
0 19733 7 1 2 19729 19732
0 19734 7 1 2 19724 19733
0 19735 5 1 1 19734
0 19736 7 1 2 88006 19735
0 19737 5 1 1 19736
0 19738 7 1 2 85098 82872
0 19739 5 1 1 19738
0 19740 7 3 2 61585 69388
0 19741 7 1 2 77859 88637
0 19742 5 1 1 19741
0 19743 7 1 2 19739 19742
0 19744 5 1 1 19743
0 19745 7 2 2 65574 72275
0 19746 5 1 1 88640
0 19747 7 2 2 77030 77463
0 19748 5 1 1 88642
0 19749 7 1 2 19746 19748
0 19750 7 1 2 19744 19749
0 19751 5 1 1 19750
0 19752 7 1 2 19737 19751
0 19753 7 1 2 19715 19752
0 19754 5 1 1 19753
0 19755 7 1 2 19754 88370
0 19756 5 1 1 19755
0 19757 7 1 2 19686 19756
0 19758 5 1 1 19757
0 19759 7 1 2 72740 19758
0 19760 5 1 1 19759
0 19761 7 1 2 19675 19760
0 19762 5 1 1 19761
0 19763 7 1 2 66895 19762
0 19764 5 1 1 19763
0 19765 7 1 2 19513 19764
0 19766 7 1 2 19510 19765
0 19767 5 1 1 19766
0 19768 7 1 2 88393 19767
0 19769 5 1 1 19768
0 19770 7 9 2 60000 61766
0 19771 5 3 1 88644
0 19772 7 15 2 64704 66406
0 19773 5 1 1 88656
0 19774 7 1 2 59339 88657
0 19775 5 2 1 19774
0 19776 7 1 2 88653 88671
0 19777 5 1 1 19776
0 19778 7 1 2 58743 19777
0 19779 5 1 1 19778
0 19780 7 3 2 60001 66407
0 19781 7 1 2 75807 88673
0 19782 5 2 1 19781
0 19783 7 1 2 19779 88676
0 19784 5 3 1 19783
0 19785 7 1 2 61922 88678
0 19786 5 1 1 19785
0 19787 7 1 2 62673 83863
0 19788 5 2 1 19787
0 19789 7 29 2 61767 66578
0 19790 7 2 2 66765 88683
0 19791 7 1 2 88681 88712
0 19792 5 1 1 19791
0 19793 7 1 2 19786 19792
0 19794 5 1 1 19793
0 19795 7 1 2 64799 19794
0 19796 5 1 1 19795
0 19797 7 11 2 61768 61923
0 19798 7 2 2 85200 88714
0 19799 5 1 1 88725
0 19800 7 1 2 19796 19799
0 19801 5 1 1 19800
0 19802 7 1 2 63608 19801
0 19803 5 1 1 19802
0 19804 7 2 2 88715 88283
0 19805 5 1 1 88727
0 19806 7 1 2 19803 19805
0 19807 5 1 1 19806
0 19808 7 1 2 88383 19807
0 19809 5 1 1 19808
0 19810 7 6 2 65247 61769
0 19811 7 4 2 60002 88729
0 19812 5 5 1 88735
0 19813 7 1 2 88672 88739
0 19814 5 1 1 19813
0 19815 7 1 2 58744 19814
0 19816 5 1 1 19815
0 19817 7 1 2 88677 19816
0 19818 5 1 1 19817
0 19819 7 1 2 76812 19818
0 19820 5 1 1 19819
0 19821 7 1 2 58022 88679
0 19822 5 1 1 19821
0 19823 7 1 2 19820 19822
0 19824 5 1 1 19823
0 19825 7 1 2 64863 70492
0 19826 7 1 2 19824 19825
0 19827 5 1 1 19826
0 19828 7 8 2 60120 64864
0 19829 7 1 2 58856 88744
0 19830 5 1 1 19829
0 19831 7 1 2 18588 19830
0 19832 5 10 1 19831
0 19833 7 4 2 61770 88752
0 19834 7 1 2 66766 88682
0 19835 7 1 2 88762 19834
0 19836 5 1 1 19835
0 19837 7 1 2 66579 19836
0 19838 7 1 2 19827 19837
0 19839 5 1 1 19838
0 19840 7 1 2 88680 88753
0 19841 5 1 1 19840
0 19842 7 6 2 60178 61771
0 19843 7 1 2 86053 88766
0 19844 5 1 1 19843
0 19845 7 1 2 61924 19844
0 19846 7 1 2 19841 19845
0 19847 5 1 1 19846
0 19848 7 1 2 63668 19847
0 19849 7 1 2 19839 19848
0 19850 5 1 1 19849
0 19851 7 1 2 19809 19850
0 19852 5 1 1 19851
0 19853 7 1 2 62065 19852
0 19854 5 1 1 19853
0 19855 7 1 2 57695 76457
0 19856 7 1 2 83344 19855
0 19857 5 1 1 19856
0 19858 7 1 2 60557 88566
0 19859 5 1 1 19858
0 19860 7 1 2 19857 19859
0 19861 5 1 1 19860
0 19862 7 1 2 59116 19861
0 19863 5 1 1 19862
0 19864 7 1 2 57696 86346
0 19865 5 1 1 19864
0 19866 7 1 2 59117 78199
0 19867 5 1 1 19866
0 19868 7 1 2 19865 19867
0 19869 5 1 1 19868
0 19870 7 1 2 57415 19869
0 19871 5 1 1 19870
0 19872 7 6 2 62184 67744
0 19873 5 3 1 88772
0 19874 7 1 2 68368 79284
0 19875 5 1 1 19874
0 19876 7 1 2 81940 19875
0 19877 5 1 1 19876
0 19878 7 1 2 88773 19877
0 19879 5 1 1 19878
0 19880 7 2 2 62674 68369
0 19881 5 1 1 88781
0 19882 7 1 2 83727 88782
0 19883 5 1 1 19882
0 19884 7 1 2 19879 19883
0 19885 7 1 2 19871 19884
0 19886 5 1 1 19885
0 19887 7 1 2 65248 19886
0 19888 5 1 1 19887
0 19889 7 1 2 19863 19888
0 19890 5 1 1 19889
0 19891 7 1 2 59340 19890
0 19892 5 1 1 19891
0 19893 7 1 2 74589 74612
0 19894 5 1 1 19893
0 19895 7 1 2 65249 79699
0 19896 5 1 1 19895
0 19897 7 1 2 19894 19896
0 19898 5 1 1 19897
0 19899 7 1 2 87099 19898
0 19900 5 1 1 19899
0 19901 7 3 2 59118 81483
0 19902 7 1 2 74335 88783
0 19903 5 1 1 19902
0 19904 7 1 2 19900 19903
0 19905 7 1 2 19892 19904
0 19906 5 1 1 19905
0 19907 7 1 2 64705 88684
0 19908 7 1 2 19906 19907
0 19909 5 1 1 19908
0 19910 7 1 2 7759 19881
0 19911 5 1 1 19910
0 19912 7 1 2 65250 19911
0 19913 5 1 1 19912
0 19914 7 1 2 68829 79692
0 19915 5 1 1 19914
0 19916 7 1 2 59341 87986
0 19917 7 1 2 87570 19916
0 19918 5 1 1 19917
0 19919 7 1 2 59119 19918
0 19920 5 1 1 19919
0 19921 7 1 2 19915 19920
0 19922 7 1 2 19913 19921
0 19923 5 1 1 19922
0 19924 7 1 2 72243 19923
0 19925 5 1 1 19924
0 19926 7 1 2 11459 19925
0 19927 5 1 1 19926
0 19928 7 2 2 66408 75957
0 19929 7 1 2 67324 88786
0 19930 7 1 2 19927 19929
0 19931 5 1 1 19930
0 19932 7 1 2 19909 19931
0 19933 5 1 1 19932
0 19934 7 1 2 63485 19933
0 19935 5 1 1 19934
0 19936 7 1 2 79693 88658
0 19937 5 1 1 19936
0 19938 7 1 2 88740 19937
0 19939 5 1 1 19938
0 19940 7 1 2 68830 19939
0 19941 5 1 1 19940
0 19942 7 1 2 70779 88659
0 19943 7 1 2 70637 19942
0 19944 5 1 1 19943
0 19945 7 1 2 88654 19773
0 19946 5 6 1 19945
0 19947 7 1 2 68772 2605
0 19948 7 1 2 7526 19947
0 19949 7 1 2 88788 19948
0 19950 5 1 1 19949
0 19951 7 1 2 19944 19950
0 19952 5 1 1 19951
0 19953 7 1 2 60333 19952
0 19954 5 1 1 19953
0 19955 7 1 2 67660 88660
0 19956 5 1 1 19955
0 19957 7 1 2 88741 19956
0 19958 5 1 1 19957
0 19959 7 1 2 62675 19958
0 19960 5 1 1 19959
0 19961 7 1 2 78062 88645
0 19962 7 1 2 70110 19961
0 19963 5 1 1 19962
0 19964 7 1 2 19960 19963
0 19965 7 1 2 19954 19964
0 19966 7 1 2 19941 19965
0 19967 5 1 1 19966
0 19968 7 1 2 59342 19967
0 19969 5 1 1 19968
0 19970 7 2 2 82155 88646
0 19971 5 1 1 88794
0 19972 7 1 2 83185 88661
0 19973 5 1 1 19972
0 19974 7 1 2 19971 19973
0 19975 5 1 1 19974
0 19976 7 1 2 65251 19975
0 19977 5 1 1 19976
0 19978 7 1 2 66409 82162
0 19979 5 1 1 19978
0 19980 7 1 2 82742 88789
0 19981 7 1 2 19979 19980
0 19982 5 1 1 19981
0 19983 7 1 2 19977 19982
0 19984 5 1 1 19983
0 19985 7 1 2 68370 19984
0 19986 5 1 1 19985
0 19987 7 1 2 67857 88795
0 19988 5 1 1 19987
0 19989 7 5 2 65252 66410
0 19990 7 3 2 64706 88796
0 19991 5 1 1 88801
0 19992 7 1 2 88784 88802
0 19993 5 1 1 19992
0 19994 7 1 2 19988 19993
0 19995 7 1 2 19986 19994
0 19996 7 1 2 19969 19995
0 19997 5 1 1 19996
0 19998 7 1 2 75681 19997
0 19999 5 1 1 19998
0 20000 7 1 2 19935 19999
0 20001 5 1 1 20000
0 20002 7 1 2 64800 20001
0 20003 5 1 1 20002
0 20004 7 1 2 82156 86143
0 20005 5 1 1 20004
0 20006 7 2 2 65253 8403
0 20007 5 2 1 88804
0 20008 7 1 2 59343 88805
0 20009 5 1 1 20008
0 20010 7 7 2 68083 68231
0 20011 5 4 1 88808
0 20012 7 1 2 82743 88815
0 20013 5 1 1 20012
0 20014 7 1 2 20009 20013
0 20015 7 1 2 20005 20014
0 20016 5 2 1 20015
0 20017 7 1 2 88726 88819
0 20018 5 1 1 20017
0 20019 7 1 2 20003 20018
0 20020 5 1 1 20019
0 20021 7 1 2 63609 20020
0 20022 5 1 1 20021
0 20023 7 1 2 88728 88820
0 20024 5 1 1 20023
0 20025 7 1 2 61772 75327
0 20026 7 1 2 85457 20025
0 20027 5 1 1 20026
0 20028 7 5 2 66411 79884
0 20029 7 2 2 62390 59120
0 20030 5 1 1 88826
0 20031 7 1 2 69138 88827
0 20032 7 1 2 88821 20031
0 20033 5 1 1 20032
0 20034 7 1 2 20027 20033
0 20035 5 1 1 20034
0 20036 7 1 2 60558 20035
0 20037 5 1 1 20036
0 20038 7 1 2 79701 71098
0 20039 7 1 2 88822 20038
0 20040 5 1 1 20039
0 20041 7 1 2 20037 20040
0 20042 5 1 1 20041
0 20043 7 1 2 63610 20042
0 20044 5 1 1 20043
0 20045 7 3 2 60559 61773
0 20046 7 1 2 88284 88828
0 20047 7 1 2 75328 20046
0 20048 5 1 1 20047
0 20049 7 1 2 20044 20048
0 20050 5 1 1 20049
0 20051 7 1 2 72448 20050
0 20052 5 1 1 20051
0 20053 7 2 2 65254 88685
0 20054 7 4 2 66767 69530
0 20055 7 1 2 88833 88785
0 20056 7 1 2 88831 20055
0 20057 5 1 1 20056
0 20058 7 1 2 20052 20057
0 20059 5 1 1 20058
0 20060 7 1 2 68617 20059
0 20061 5 1 1 20060
0 20062 7 1 2 20024 20061
0 20063 7 1 2 20022 20062
0 20064 5 1 1 20063
0 20065 7 1 2 88142 20064
0 20066 5 1 1 20065
0 20067 7 1 2 19854 20066
0 20068 5 1 1 20067
0 20069 7 1 2 65575 20068
0 20070 5 1 1 20069
0 20071 7 2 2 67661 67444
0 20072 7 1 2 68773 72319
0 20073 7 1 2 88837 20072
0 20074 5 1 1 20073
0 20075 7 1 2 72184 20074
0 20076 5 1 1 20075
0 20077 7 1 2 77269 20076
0 20078 5 1 1 20077
0 20079 7 1 2 83694 84111
0 20080 7 1 2 71658 20079
0 20081 5 1 1 20080
0 20082 7 1 2 20078 20081
0 20083 5 1 1 20082
0 20084 7 1 2 65255 20083
0 20085 5 1 1 20084
0 20086 7 1 2 72284 78587
0 20087 7 1 2 81768 20086
0 20088 5 1 1 20087
0 20089 7 1 2 20085 20088
0 20090 5 1 1 20089
0 20091 7 1 2 65031 20090
0 20092 5 1 1 20091
0 20093 7 2 2 60906 81769
0 20094 5 1 1 88839
0 20095 7 1 2 86097 88233
0 20096 5 1 1 20095
0 20097 7 1 2 59344 20096
0 20098 5 1 1 20097
0 20099 7 1 2 87090 20098
0 20100 5 1 1 20099
0 20101 7 1 2 88840 20100
0 20102 5 1 1 20101
0 20103 7 2 2 66768 74242
0 20104 7 1 2 65256 79760
0 20105 5 1 1 20104
0 20106 7 1 2 86101 20105
0 20107 5 1 1 20106
0 20108 7 1 2 88841 20107
0 20109 5 1 1 20108
0 20110 7 1 2 74419 84217
0 20111 5 1 1 20110
0 20112 7 1 2 20109 20111
0 20113 5 1 1 20112
0 20114 7 1 2 70493 20113
0 20115 5 1 1 20114
0 20116 7 1 2 20102 20115
0 20117 7 1 2 20092 20116
0 20118 5 1 1 20117
0 20119 7 1 2 61774 20118
0 20120 5 1 1 20119
0 20121 7 4 2 61925 79885
0 20122 7 5 2 64801 66412
0 20123 7 1 2 77766 72561
0 20124 7 1 2 88847 20123
0 20125 7 1 2 88843 20124
0 20126 7 1 2 82089 20125
0 20127 5 1 1 20126
0 20128 7 1 2 20120 20127
0 20129 5 1 1 20128
0 20130 7 1 2 64865 20129
0 20131 5 1 1 20130
0 20132 7 7 2 61775 62066
0 20133 7 2 2 75737 88852
0 20134 7 2 2 69139 88859
0 20135 7 1 2 60179 74336
0 20136 7 1 2 79235 20135
0 20137 7 1 2 88861 20136
0 20138 5 1 1 20137
0 20139 7 1 2 20131 20138
0 20140 5 1 1 20139
0 20141 7 1 2 63669 20140
0 20142 5 1 1 20141
0 20143 7 4 2 64866 65032
0 20144 7 1 2 63486 65257
0 20145 7 1 2 88087 20144
0 20146 7 1 2 88863 20145
0 20147 7 1 2 88862 20146
0 20148 5 1 1 20147
0 20149 7 1 2 20142 20148
0 20150 7 1 2 20070 20149
0 20151 5 1 1 20150
0 20152 7 1 2 66195 20151
0 20153 5 1 1 20152
0 20154 7 12 2 61776 79886
0 20155 5 1 1 88867
0 20156 7 2 2 3251 71963
0 20157 7 3 2 57416 64802
0 20158 5 1 1 88881
0 20159 7 1 2 63611 20158
0 20160 7 1 2 88879 20159
0 20161 5 1 1 20160
0 20162 7 1 2 84770 20161
0 20163 5 1 1 20162
0 20164 7 1 2 78287 20163
0 20165 5 1 1 20164
0 20166 7 1 2 72754 81578
0 20167 5 1 1 20166
0 20168 7 1 2 59121 76458
0 20169 5 1 1 20168
0 20170 7 1 2 72741 20169
0 20171 5 1 1 20170
0 20172 7 1 2 20167 20171
0 20173 7 1 2 20165 20172
0 20174 5 1 1 20173
0 20175 7 1 2 62676 20174
0 20176 5 1 1 20175
0 20177 7 1 2 68232 77090
0 20178 7 1 2 72742 20177
0 20179 5 1 1 20178
0 20180 7 1 2 20176 20179
0 20181 5 1 1 20180
0 20182 7 1 2 88868 20181
0 20183 5 1 1 20182
0 20184 7 2 2 86347 80693
0 20185 5 1 1 88884
0 20186 7 1 2 62391 88885
0 20187 5 1 1 20186
0 20188 7 3 2 59122 76504
0 20189 5 2 1 88886
0 20190 7 1 2 87093 88889
0 20191 5 1 1 20190
0 20192 7 1 2 20187 20191
0 20193 5 1 1 20192
0 20194 7 4 2 66413 86062
0 20195 7 1 2 61926 88891
0 20196 7 1 2 20193 20195
0 20197 5 1 1 20196
0 20198 7 1 2 20183 20197
0 20199 5 1 1 20198
0 20200 7 1 2 60560 20199
0 20201 5 1 1 20200
0 20202 7 24 2 66414 61927
0 20203 7 1 2 77091 88895
0 20204 7 1 2 84409 20203
0 20205 7 1 2 86063 20204
0 20206 5 1 1 20205
0 20207 7 1 2 20201 20206
0 20208 5 1 1 20207
0 20209 7 9 2 61586 66690
0 20210 7 1 2 73114 88120
0 20211 7 1 2 88919 20210
0 20212 7 1 2 20208 20211
0 20213 5 1 1 20212
0 20214 7 1 2 20153 20213
0 20215 5 1 1 20214
0 20216 7 1 2 76732 20215
0 20217 5 1 1 20216
0 20218 7 1 2 75112 72688
0 20219 5 1 1 20218
0 20220 7 3 2 62677 69026
0 20221 5 1 1 88928
0 20222 7 3 2 75263 88929
0 20223 5 1 1 88931
0 20224 7 1 2 72743 20223
0 20225 5 1 1 20224
0 20226 7 1 2 70090 80505
0 20227 5 1 1 20226
0 20228 7 3 2 75232 20227
0 20229 5 2 1 88934
0 20230 7 1 2 57697 88937
0 20231 5 1 1 20230
0 20232 7 3 2 62392 65033
0 20233 7 1 2 78825 88939
0 20234 5 1 1 20233
0 20235 7 1 2 83438 20234
0 20236 7 1 2 20231 20235
0 20237 5 1 1 20236
0 20238 7 1 2 63880 20237
0 20239 5 1 1 20238
0 20240 7 1 2 69843 88570
0 20241 5 1 1 20240
0 20242 7 1 2 62393 88935
0 20243 5 1 1 20242
0 20244 7 2 2 63764 69844
0 20245 5 1 1 88942
0 20246 7 1 2 74522 20245
0 20247 5 3 1 20246
0 20248 7 7 2 83268 88944
0 20249 5 1 1 88947
0 20250 7 1 2 57698 20249
0 20251 5 1 1 20250
0 20252 7 1 2 59123 20251
0 20253 7 1 2 20243 20252
0 20254 5 1 1 20253
0 20255 7 1 2 20241 20254
0 20256 7 1 2 20239 20255
0 20257 5 1 1 20256
0 20258 7 1 2 84221 20257
0 20259 5 1 1 20258
0 20260 7 1 2 20225 20259
0 20261 5 1 1 20260
0 20262 7 1 2 59345 20261
0 20263 5 1 1 20262
0 20264 7 1 2 83188 6996
0 20265 5 5 1 20264
0 20266 7 1 2 65034 88954
0 20267 5 1 1 20266
0 20268 7 1 2 64036 74570
0 20269 5 1 1 20268
0 20270 7 1 2 20267 20269
0 20271 5 1 1 20270
0 20272 7 1 2 66964 20271
0 20273 5 1 1 20272
0 20274 7 1 2 77148 67043
0 20275 5 1 1 20274
0 20276 7 1 2 20273 20275
0 20277 5 1 1 20276
0 20278 7 1 2 65258 20277
0 20279 5 1 1 20278
0 20280 7 2 2 58023 66965
0 20281 7 1 2 65035 81370
0 20282 5 1 1 20281
0 20283 7 1 2 69768 20282
0 20284 5 1 1 20283
0 20285 7 1 2 88959 20284
0 20286 5 1 1 20285
0 20287 7 1 2 8755 20286
0 20288 7 1 2 20279 20287
0 20289 5 1 1 20288
0 20290 7 1 2 63612 20289
0 20291 5 1 1 20290
0 20292 7 1 2 64037 84077
0 20293 5 1 1 20292
0 20294 7 1 2 84767 20293
0 20295 5 1 1 20294
0 20296 7 1 2 20291 20295
0 20297 5 1 1 20296
0 20298 7 1 2 68371 20297
0 20299 5 1 1 20298
0 20300 7 6 2 77209 72107
0 20301 5 1 1 88961
0 20302 7 1 2 59346 88962
0 20303 5 1 1 20302
0 20304 7 1 2 72504 20303
0 20305 5 1 1 20304
0 20306 7 1 2 63613 20305
0 20307 5 1 1 20306
0 20308 7 1 2 70452 72449
0 20309 5 1 1 20308
0 20310 7 1 2 20307 20309
0 20311 5 1 1 20310
0 20312 7 1 2 68618 20311
0 20313 5 1 1 20312
0 20314 7 1 2 79839 67113
0 20315 5 1 1 20314
0 20316 7 1 2 67083 20315
0 20317 5 1 1 20316
0 20318 7 1 2 63614 20317
0 20319 5 1 1 20318
0 20320 7 1 2 84771 20319
0 20321 5 1 1 20320
0 20322 7 1 2 68774 20321
0 20323 5 1 1 20322
0 20324 7 1 2 20313 20323
0 20325 5 1 1 20324
0 20326 7 1 2 67858 20325
0 20327 5 1 1 20326
0 20328 7 1 2 70590 82901
0 20329 7 1 2 88963 20328
0 20330 5 1 1 20329
0 20331 7 1 2 20327 20330
0 20332 7 1 2 20299 20331
0 20333 7 1 2 20263 20332
0 20334 5 1 1 20333
0 20335 7 1 2 66691 20334
0 20336 5 1 1 20335
0 20337 7 1 2 20219 20336
0 20338 5 1 1 20337
0 20339 7 5 2 61777 75513
0 20340 7 1 2 20338 88967
0 20341 5 1 1 20340
0 20342 7 1 2 57699 20185
0 20343 5 1 1 20342
0 20344 7 1 2 80706 20343
0 20345 5 2 1 20344
0 20346 7 1 2 60561 88972
0 20347 5 1 1 20346
0 20348 7 1 2 60562 83874
0 20349 5 1 1 20348
0 20350 7 1 2 63881 80360
0 20351 5 1 1 20350
0 20352 7 1 2 77728 20351
0 20353 5 2 1 20352
0 20354 7 1 2 70708 76813
0 20355 5 1 1 20354
0 20356 7 1 2 65259 20355
0 20357 7 1 2 88974 20356
0 20358 5 1 1 20357
0 20359 7 1 2 59347 20358
0 20360 7 1 2 20349 20359
0 20361 5 1 1 20360
0 20362 7 1 2 20347 20361
0 20363 5 1 1 20362
0 20364 7 3 2 66692 20363
0 20365 7 3 2 58493 64803
0 20366 7 3 2 82718 88979
0 20367 7 1 2 88896 88982
0 20368 7 1 2 88976 20367
0 20369 5 1 1 20368
0 20370 7 1 2 20341 20369
0 20371 5 1 1 20370
0 20372 7 1 2 64867 20371
0 20373 5 1 1 20372
0 20374 7 1 2 75113 84222
0 20375 5 1 1 20374
0 20376 7 1 2 72752 20375
0 20377 5 2 1 20376
0 20378 7 2 2 88985 88853
0 20379 7 4 2 64509 60180
0 20380 7 2 2 63241 88989
0 20381 7 1 2 88987 88993
0 20382 5 1 1 20381
0 20383 7 1 2 20373 20382
0 20384 5 1 1 20383
0 20385 7 1 2 63670 20384
0 20386 5 1 1 20385
0 20387 7 3 2 66415 67953
0 20388 7 2 2 88474 88995
0 20389 5 1 1 88998
0 20390 7 1 2 81223 88349
0 20391 7 4 2 64510 88686
0 20392 7 1 2 88955 89000
0 20393 7 1 2 20390 20392
0 20394 5 1 1 20393
0 20395 7 1 2 20389 20394
0 20396 5 1 1 20395
0 20397 7 1 2 63671 20396
0 20398 5 1 1 20397
0 20399 7 6 2 66416 76626
0 20400 7 2 2 67954 88384
0 20401 7 1 2 89004 89010
0 20402 5 1 1 20401
0 20403 7 1 2 20398 20402
0 20404 5 1 1 20403
0 20405 7 1 2 69531 20404
0 20406 5 1 1 20405
0 20407 7 3 2 58494 67925
0 20408 7 4 2 63672 59783
0 20409 7 2 2 89012 89015
0 20410 7 5 2 64868 66417
0 20411 7 2 2 67955 89021
0 20412 7 1 2 89019 89026
0 20413 5 1 1 20412
0 20414 7 1 2 20406 20413
0 20415 5 1 1 20414
0 20416 7 1 2 69418 20415
0 20417 5 1 1 20416
0 20418 7 1 2 75514 88385
0 20419 7 1 2 88988 20418
0 20420 5 1 1 20419
0 20421 7 1 2 20417 20420
0 20422 7 1 2 20386 20421
0 20423 5 1 1 20422
0 20424 7 1 2 66896 20423
0 20425 5 1 1 20424
0 20426 7 2 2 64038 78748
0 20427 5 3 1 89028
0 20428 7 1 2 84515 74463
0 20429 5 1 1 20428
0 20430 7 1 2 60334 20429
0 20431 5 1 1 20430
0 20432 7 1 2 77322 20431
0 20433 5 1 1 20432
0 20434 7 1 2 89030 20433
0 20435 5 1 1 20434
0 20436 7 1 2 69389 76945
0 20437 5 1 1 20436
0 20438 7 1 2 65036 87369
0 20439 5 1 1 20438
0 20440 7 1 2 73208 70998
0 20441 5 1 1 20440
0 20442 7 1 2 20439 20441
0 20443 5 1 1 20442
0 20444 7 1 2 64039 20443
0 20445 5 1 1 20444
0 20446 7 1 2 20437 20445
0 20447 7 1 2 20435 20446
0 20448 5 1 1 20447
0 20449 7 1 2 58024 20448
0 20450 5 1 1 20449
0 20451 7 1 2 59124 88938
0 20452 5 1 1 20451
0 20453 7 1 2 68775 75073
0 20454 5 1 1 20453
0 20455 7 1 2 62394 20454
0 20456 7 1 2 20452 20455
0 20457 5 1 1 20456
0 20458 7 1 2 63882 88936
0 20459 5 1 1 20458
0 20460 7 1 2 62185 88945
0 20461 5 2 1 20460
0 20462 7 1 2 69442 79063
0 20463 5 1 1 20462
0 20464 7 1 2 59125 70730
0 20465 7 1 2 20463 20464
0 20466 7 1 2 89033 20465
0 20467 5 1 1 20466
0 20468 7 1 2 20459 20467
0 20469 5 1 1 20468
0 20470 7 1 2 83233 82754
0 20471 5 1 1 20470
0 20472 7 1 2 57700 20471
0 20473 7 1 2 20469 20472
0 20474 5 1 1 20473
0 20475 7 1 2 20457 20474
0 20476 5 1 1 20475
0 20477 7 1 2 59348 18709
0 20478 7 1 2 20476 20477
0 20479 5 1 1 20478
0 20480 7 1 2 89031 20479
0 20481 5 1 1 20480
0 20482 7 1 2 20450 20481
0 20483 5 1 1 20482
0 20484 7 1 2 72755 20483
0 20485 5 1 1 20484
0 20486 7 1 2 59349 83471
0 20487 5 1 1 20486
0 20488 7 1 2 86146 20487
0 20489 5 1 1 20488
0 20490 7 2 2 61928 20489
0 20491 7 1 2 70494 89035
0 20492 5 1 1 20491
0 20493 7 1 2 20485 20492
0 20494 5 1 1 20493
0 20495 7 1 2 66769 20494
0 20496 5 1 1 20495
0 20497 7 1 2 82064 89036
0 20498 5 1 1 20497
0 20499 7 1 2 66693 20498
0 20500 7 1 2 20496 20499
0 20501 5 1 1 20500
0 20502 7 1 2 75114 88461
0 20503 5 1 1 20502
0 20504 7 5 2 77016 83551
0 20505 5 4 1 89037
0 20506 7 1 2 62067 89042
0 20507 7 1 2 20503 20506
0 20508 5 1 1 20507
0 20509 7 1 2 63673 20508
0 20510 7 1 2 20501 20509
0 20511 5 1 1 20510
0 20512 7 1 2 19226 20511
0 20513 5 1 1 20512
0 20514 7 18 2 61778 76627
0 20515 5 2 1 89046
0 20516 7 1 2 66770 88986
0 20517 5 1 1 20516
0 20518 7 2 2 69532 75654
0 20519 5 1 1 89066
0 20520 7 1 2 20517 20519
0 20521 5 1 1 20520
0 20522 7 1 2 62068 20521
0 20523 5 1 1 20522
0 20524 7 1 2 88138 20523
0 20525 5 1 1 20524
0 20526 7 1 2 89047 20525
0 20527 7 1 2 20513 20526
0 20528 5 1 1 20527
0 20529 7 1 2 69533 88977
0 20530 5 1 1 20529
0 20531 7 2 2 62069 69419
0 20532 7 1 2 67926 89068
0 20533 5 1 1 20532
0 20534 7 1 2 20530 20533
0 20535 5 1 1 20534
0 20536 7 1 2 66828 20535
0 20537 5 1 1 20536
0 20538 7 1 2 86054 88978
0 20539 5 1 1 20538
0 20540 7 1 2 20537 20539
0 20541 5 1 1 20540
0 20542 7 1 2 61929 20541
0 20543 5 1 1 20542
0 20544 7 1 2 62395 77533
0 20545 5 2 1 20544
0 20546 7 2 2 71680 68197
0 20547 5 1 1 89072
0 20548 7 1 2 89070 20547
0 20549 5 4 1 20548
0 20550 7 1 2 58025 89074
0 20551 5 1 1 20550
0 20552 7 1 2 69888 87983
0 20553 7 1 2 75284 20552
0 20554 5 1 1 20553
0 20555 7 1 2 20551 20554
0 20556 5 1 1 20555
0 20557 7 1 2 59350 20556
0 20558 5 1 1 20557
0 20559 7 1 2 88495 88956
0 20560 5 1 1 20559
0 20561 7 1 2 20558 20560
0 20562 5 1 1 20561
0 20563 7 1 2 65260 20562
0 20564 5 1 1 20563
0 20565 7 1 2 78346 83509
0 20566 5 1 1 20565
0 20567 7 1 2 83230 77724
0 20568 5 1 1 20567
0 20569 7 1 2 20566 20568
0 20570 5 1 1 20569
0 20571 7 1 2 68965 20570
0 20572 5 1 1 20571
0 20573 7 1 2 20564 20572
0 20574 5 1 1 20573
0 20575 7 1 2 83699 20574
0 20576 5 1 1 20575
0 20577 7 1 2 88121 20576
0 20578 7 1 2 20543 20577
0 20579 5 1 1 20578
0 20580 7 1 2 88403 89069
0 20581 5 1 1 20580
0 20582 7 1 2 88139 20581
0 20583 5 1 1 20582
0 20584 7 18 2 66418 75515
0 20585 7 1 2 88316 89078
0 20586 7 1 2 20583 20585
0 20587 7 1 2 20579 20586
0 20588 5 1 1 20587
0 20589 7 1 2 20528 20588
0 20590 7 1 2 20425 20589
0 20591 5 1 1 20590
0 20592 7 1 2 65576 20591
0 20593 5 1 1 20592
0 20594 7 15 2 62070 88386
0 20595 5 2 1 89096
0 20596 7 31 2 60181 62071
0 20597 5 1 1 89113
0 20598 7 1 2 88580 19150
0 20599 5 1 1 20598
0 20600 7 1 2 20597 20599
0 20601 5 1 1 20600
0 20602 7 1 2 63674 20601
0 20603 5 1 1 20602
0 20604 7 1 2 89111 20603
0 20605 5 1 1 20604
0 20606 7 1 2 65261 20605
0 20607 5 1 1 20606
0 20608 7 1 2 58026 88583
0 20609 7 1 2 77181 20608
0 20610 5 1 1 20609
0 20611 7 1 2 20607 20610
0 20612 5 1 1 20611
0 20613 7 1 2 66966 20612
0 20614 5 1 1 20613
0 20615 7 1 2 76505 80196
0 20616 5 1 1 20615
0 20617 7 2 2 70968 68776
0 20618 5 1 1 89144
0 20619 7 1 2 65037 89145
0 20620 5 1 1 20619
0 20621 7 1 2 20616 20620
0 20622 5 1 1 20621
0 20623 7 2 2 67518 20622
0 20624 7 1 2 63675 88745
0 20625 7 1 2 89146 20624
0 20626 5 1 1 20625
0 20627 7 1 2 20614 20626
0 20628 5 1 1 20627
0 20629 7 1 2 63615 20628
0 20630 5 1 1 20629
0 20631 7 6 2 58857 63676
0 20632 7 4 2 64869 89148
0 20633 7 1 2 64804 89147
0 20634 5 1 1 20633
0 20635 7 1 2 84097 20634
0 20636 5 1 1 20635
0 20637 7 1 2 89154 20636
0 20638 5 1 1 20637
0 20639 7 1 2 20630 20638
0 20640 5 1 1 20639
0 20641 7 1 2 88968 20640
0 20642 5 1 1 20641
0 20643 7 7 2 59784 64870
0 20644 7 5 2 63677 89158
0 20645 7 1 2 72309 88897
0 20646 7 1 2 86619 20645
0 20647 7 1 2 89165 20646
0 20648 7 1 2 88973 20647
0 20649 5 1 1 20648
0 20650 7 1 2 20642 20649
0 20651 5 1 1 20650
0 20652 7 1 2 59351 20651
0 20653 5 1 1 20652
0 20654 7 5 2 76628 88898
0 20655 5 3 1 89170
0 20656 7 1 2 86035 89171
0 20657 5 1 1 20656
0 20658 7 3 2 57701 64511
0 20659 7 2 2 73856 89178
0 20660 7 6 2 63242 58975
0 20661 5 1 1 89183
0 20662 7 1 2 88687 89184
0 20663 7 1 2 89181 20662
0 20664 5 1 1 20663
0 20665 7 1 2 20657 20664
0 20666 5 1 1 20665
0 20667 7 1 2 69534 73403
0 20668 7 1 2 88584 20667
0 20669 7 1 2 20666 20668
0 20670 5 1 1 20669
0 20671 7 1 2 20653 20670
0 20672 5 1 1 20671
0 20673 7 1 2 66897 20672
0 20674 5 1 1 20673
0 20675 7 4 2 87883 88688
0 20676 7 1 2 59352 89189
0 20677 5 1 1 20676
0 20678 7 3 2 68997 79568
0 20679 7 1 2 73978 88899
0 20680 7 1 2 89193 20679
0 20681 5 1 1 20680
0 20682 7 1 2 20677 20681
0 20683 5 1 1 20682
0 20684 7 1 2 65262 20683
0 20685 5 1 1 20684
0 20686 7 1 2 85379 88900
0 20687 5 1 1 20686
0 20688 7 1 2 57417 89190
0 20689 5 1 1 20688
0 20690 7 1 2 20687 20689
0 20691 5 1 1 20690
0 20692 7 1 2 71737 20691
0 20693 5 1 1 20692
0 20694 7 4 2 63243 79551
0 20695 5 1 1 89196
0 20696 7 2 2 88787 89197
0 20697 7 1 2 57418 89200
0 20698 5 1 1 20697
0 20699 7 6 2 58976 59785
0 20700 5 1 1 89202
0 20701 7 2 2 88689 89203
0 20702 7 1 2 82639 83416
0 20703 7 1 2 89208 20702
0 20704 5 1 1 20703
0 20705 7 1 2 20698 20704
0 20706 7 1 2 20693 20705
0 20707 5 1 1 20706
0 20708 7 1 2 59353 20707
0 20709 5 1 1 20708
0 20710 7 1 2 20685 20709
0 20711 5 1 1 20710
0 20712 7 1 2 77767 20711
0 20713 5 1 1 20712
0 20714 7 1 2 61779 74420
0 20715 7 2 2 84445 20714
0 20716 7 1 2 79077 89210
0 20717 5 1 1 20716
0 20718 7 1 2 20713 20717
0 20719 5 1 1 20718
0 20720 7 1 2 68372 20719
0 20721 5 1 1 20720
0 20722 7 1 2 13054 73412
0 20723 5 1 1 20722
0 20724 7 1 2 57419 20723
0 20725 5 1 1 20724
0 20726 7 2 2 64040 80515
0 20727 5 2 1 89212
0 20728 7 1 2 58027 89214
0 20729 5 1 1 20728
0 20730 7 1 2 20725 20729
0 20731 5 1 1 20730
0 20732 7 1 2 20731 89201
0 20733 5 1 1 20732
0 20734 7 1 2 68084 76548
0 20735 5 1 1 20734
0 20736 7 1 2 67325 89191
0 20737 7 1 2 20735 20736
0 20738 5 1 1 20737
0 20739 7 1 2 20733 20738
0 20740 5 1 1 20739
0 20741 7 1 2 60907 20740
0 20742 5 1 1 20741
0 20743 7 1 2 76506 89211
0 20744 5 1 1 20743
0 20745 7 1 2 20742 20744
0 20746 5 1 1 20745
0 20747 7 1 2 67662 20746
0 20748 5 1 1 20747
0 20749 7 1 2 76446 83340
0 20750 5 1 1 20749
0 20751 7 1 2 75655 20750
0 20752 5 1 1 20751
0 20753 7 1 2 72389 77768
0 20754 7 1 2 82056 20753
0 20755 5 1 1 20754
0 20756 7 1 2 20752 20755
0 20757 5 1 1 20756
0 20758 7 1 2 89048 20757
0 20759 5 1 1 20758
0 20760 7 3 2 60908 88901
0 20761 7 1 2 80643 89216
0 20762 7 1 2 89194 20761
0 20763 5 1 1 20762
0 20764 7 1 2 20759 20763
0 20765 5 1 1 20764
0 20766 7 1 2 59354 20765
0 20767 5 1 1 20766
0 20768 7 1 2 20748 20767
0 20769 7 1 2 20721 20768
0 20770 5 1 1 20769
0 20771 7 1 2 69270 20770
0 20772 5 1 1 20771
0 20773 7 21 2 59786 61780
0 20774 7 4 2 58495 89219
0 20775 5 7 1 89240
0 20776 7 21 2 64512 66419
0 20777 7 2 2 73999 89251
0 20778 7 1 2 60909 89272
0 20779 5 1 1 20778
0 20780 7 1 2 89244 20779
0 20781 5 1 1 20780
0 20782 7 1 2 80695 20781
0 20783 5 1 1 20782
0 20784 7 2 2 77769 89079
0 20785 5 1 1 89274
0 20786 7 1 2 59126 89275
0 20787 5 1 1 20786
0 20788 7 3 2 76629 88730
0 20789 5 1 1 89276
0 20790 7 1 2 79064 89277
0 20791 5 1 1 20790
0 20792 7 1 2 20787 20791
0 20793 5 1 1 20792
0 20794 7 1 2 57702 20793
0 20795 5 1 1 20794
0 20796 7 1 2 20783 20795
0 20797 5 1 1 20796
0 20798 7 1 2 59355 20797
0 20799 5 1 1 20798
0 20800 7 2 2 74016 89252
0 20801 7 2 2 77770 89279
0 20802 5 1 1 89281
0 20803 7 1 2 80636 89220
0 20804 5 1 1 20803
0 20805 7 1 2 20802 20804
0 20806 5 1 1 20805
0 20807 7 1 2 57703 20806
0 20808 5 1 1 20807
0 20809 7 1 2 20785 20789
0 20810 5 1 1 20809
0 20811 7 1 2 59356 20810
0 20812 5 1 1 20811
0 20813 7 1 2 20808 20812
0 20814 5 1 1 20813
0 20815 7 1 2 77529 20814
0 20816 5 1 1 20815
0 20817 7 1 2 80686 89282
0 20818 5 1 1 20817
0 20819 7 1 2 20816 20818
0 20820 7 1 2 20799 20819
0 20821 5 1 1 20820
0 20822 7 1 2 74410 20821
0 20823 5 1 1 20822
0 20824 7 4 2 66580 76630
0 20825 7 1 2 69969 66829
0 20826 7 1 2 88854 20825
0 20827 7 1 2 89283 20826
0 20828 5 1 1 20827
0 20829 7 1 2 20823 20828
0 20830 5 1 1 20829
0 20831 7 1 2 70495 20830
0 20832 5 1 1 20831
0 20833 7 2 2 76920 81880
0 20834 7 4 2 62072 88690
0 20835 7 6 2 59787 65263
0 20836 7 1 2 72327 89293
0 20837 7 1 2 89289 20836
0 20838 7 1 2 89287 20837
0 20839 5 1 1 20838
0 20840 7 1 2 20832 20839
0 20841 7 1 2 20772 20840
0 20842 5 1 1 20841
0 20843 7 1 2 64871 20842
0 20844 5 1 1 20843
0 20845 7 1 2 69970 67467
0 20846 7 1 2 88767 20845
0 20847 7 3 2 58496 79236
0 20848 7 3 2 64805 79822
0 20849 7 1 2 89299 89302
0 20850 7 1 2 20846 20849
0 20851 5 1 1 20850
0 20852 7 1 2 20844 20851
0 20853 5 1 1 20852
0 20854 7 1 2 63678 20853
0 20855 5 1 1 20854
0 20856 7 1 2 69971 87875
0 20857 7 1 2 89221 20856
0 20858 7 2 2 58911 67468
0 20859 7 2 2 66771 80458
0 20860 7 1 2 89305 89307
0 20861 7 1 2 20857 20860
0 20862 5 1 1 20861
0 20863 7 1 2 20855 20862
0 20864 7 1 2 20674 20863
0 20865 7 1 2 20593 20864
0 20866 5 1 1 20865
0 20867 7 1 2 61587 20866
0 20868 5 1 1 20867
0 20869 7 5 2 66420 66581
0 20870 7 7 2 62073 89309
0 20871 7 6 2 82800 87623
0 20872 5 1 1 89321
0 20873 7 1 2 57420 89322
0 20874 5 1 1 20873
0 20875 7 3 2 66196 77860
0 20876 7 1 2 68373 89327
0 20877 5 1 1 20876
0 20878 7 2 2 86846 82549
0 20879 5 1 1 89330
0 20880 7 1 2 20877 20879
0 20881 5 1 1 20880
0 20882 7 1 2 66898 20881
0 20883 5 1 1 20882
0 20884 7 1 2 20874 20883
0 20885 5 1 1 20884
0 20886 7 1 2 70496 20885
0 20887 5 1 1 20886
0 20888 7 4 2 58858 76058
0 20889 7 3 2 83659 89332
0 20890 7 4 2 64513 89336
0 20891 5 1 1 89339
0 20892 7 1 2 84296 89340
0 20893 5 1 1 20892
0 20894 7 1 2 20887 20893
0 20895 5 1 1 20894
0 20896 7 1 2 64872 20895
0 20897 5 1 1 20896
0 20898 7 2 2 64806 86665
0 20899 7 3 2 87908 89343
0 20900 7 2 2 83423 74502
0 20901 7 1 2 89345 89348
0 20902 5 1 1 20901
0 20903 7 1 2 20897 20902
0 20904 5 1 1 20903
0 20905 7 1 2 63679 20904
0 20906 5 1 1 20905
0 20907 7 1 2 84297 88212
0 20908 5 1 1 20907
0 20909 7 1 2 20906 20908
0 20910 5 1 1 20909
0 20911 7 1 2 71738 20910
0 20912 5 1 1 20911
0 20913 7 2 2 86329 88208
0 20914 5 1 1 89350
0 20915 7 11 2 61588 76631
0 20916 5 3 1 89352
0 20917 7 1 2 76733 86837
0 20918 5 1 1 20917
0 20919 7 1 2 89363 20918
0 20920 5 1 1 20919
0 20921 7 1 2 66899 20920
0 20922 5 1 1 20921
0 20923 7 1 2 20872 20922
0 20924 5 1 1 20923
0 20925 7 1 2 70497 20924
0 20926 5 1 1 20925
0 20927 7 2 2 86800 79206
0 20928 5 1 1 89366
0 20929 7 1 2 20926 20928
0 20930 5 1 1 20929
0 20931 7 1 2 64873 20930
0 20932 5 1 1 20931
0 20933 7 1 2 18665 20932
0 20934 5 1 1 20933
0 20935 7 1 2 63680 20934
0 20936 5 1 1 20935
0 20937 7 1 2 20914 20936
0 20938 5 1 1 20937
0 20939 7 1 2 81581 20938
0 20940 5 1 1 20939
0 20941 7 4 2 79887 70498
0 20942 7 2 2 67859 77861
0 20943 7 3 2 66197 88122
0 20944 7 1 2 89372 89374
0 20945 7 1 2 89368 20944
0 20946 5 1 1 20945
0 20947 7 1 2 20940 20946
0 20948 7 1 2 20912 20947
0 20949 5 1 1 20948
0 20950 7 1 2 65264 20949
0 20951 5 1 1 20950
0 20952 7 1 2 58028 89351
0 20953 5 1 1 20952
0 20954 7 1 2 58029 89323
0 20955 5 1 1 20954
0 20956 7 1 2 67818 86339
0 20957 5 3 1 20956
0 20958 7 3 2 77862 81568
0 20959 7 1 2 89377 89380
0 20960 5 1 1 20959
0 20961 7 9 2 58497 82550
0 20962 5 4 1 89383
0 20963 7 1 2 58030 89384
0 20964 5 1 1 20963
0 20965 7 1 2 20960 20964
0 20966 5 1 1 20965
0 20967 7 1 2 66900 20966
0 20968 5 1 1 20967
0 20969 7 1 2 20955 20968
0 20970 5 1 1 20969
0 20971 7 1 2 70499 20970
0 20972 5 1 1 20971
0 20973 7 1 2 58031 89367
0 20974 5 1 1 20973
0 20975 7 1 2 20972 20974
0 20976 5 1 1 20975
0 20977 7 1 2 64874 20976
0 20978 5 1 1 20977
0 20979 7 1 2 83424 76096
0 20980 7 1 2 89346 20979
0 20981 5 1 1 20980
0 20982 7 1 2 20978 20981
0 20983 5 1 1 20982
0 20984 7 1 2 63681 20983
0 20985 5 1 1 20984
0 20986 7 1 2 20953 20985
0 20987 7 1 2 20951 20986
0 20988 5 1 1 20987
0 20989 7 1 2 89314 20988
0 20990 5 1 1 20989
0 20991 7 1 2 70500 87888
0 20992 5 1 1 20991
0 20993 7 2 2 86994 79179
0 20994 7 1 2 76108 89396
0 20995 5 1 1 20994
0 20996 7 1 2 20992 20995
0 20997 5 1 1 20996
0 20998 7 3 2 61589 88716
0 20999 7 1 2 88143 89398
0 21000 7 1 2 77701 20999
0 21001 7 1 2 20997 21000
0 21002 5 1 1 21001
0 21003 7 1 2 20990 21002
0 21004 5 1 1 21003
0 21005 7 1 2 73170 21004
0 21006 5 1 1 21005
0 21007 7 5 2 61781 70501
0 21008 7 5 2 62186 63244
0 21009 5 1 1 89406
0 21010 7 2 2 64514 89407
0 21011 7 2 2 89401 89411
0 21012 5 1 1 89413
0 21013 7 4 2 69786 72192
0 21014 5 2 1 89415
0 21015 7 1 2 89414 89416
0 21016 5 1 1 21015
0 21017 7 2 2 76632 88848
0 21018 7 1 2 76999 89421
0 21019 5 1 1 21018
0 21020 7 1 2 21012 21019
0 21021 5 1 1 21020
0 21022 7 1 2 78288 21021
0 21023 5 1 1 21022
0 21024 7 1 2 67745 70502
0 21025 7 1 2 88969 21024
0 21026 5 1 1 21025
0 21027 7 7 2 59788 66421
0 21028 7 1 2 68198 89423
0 21029 7 1 2 86620 21028
0 21030 5 1 1 21029
0 21031 7 1 2 21026 21030
0 21032 5 1 1 21031
0 21033 7 1 2 69027 21032
0 21034 5 1 1 21033
0 21035 7 5 2 63245 80658
0 21036 7 1 2 67604 89430
0 21037 7 1 2 89402 21036
0 21038 5 1 1 21037
0 21039 7 1 2 21034 21038
0 21040 7 1 2 21023 21039
0 21041 5 1 1 21040
0 21042 7 1 2 62678 21041
0 21043 5 1 1 21042
0 21044 7 1 2 21016 21043
0 21045 5 1 1 21044
0 21046 7 1 2 61930 21045
0 21047 5 1 1 21046
0 21048 7 3 2 64807 61782
0 21049 7 2 2 66582 89435
0 21050 7 1 2 86550 77554
0 21051 7 1 2 89438 21050
0 21052 5 1 1 21051
0 21053 7 1 2 21047 21052
0 21054 5 1 1 21053
0 21055 7 1 2 66901 21054
0 21056 5 1 1 21055
0 21057 7 2 2 86545 89253
0 21058 5 1 1 89440
0 21059 7 1 2 62187 89441
0 21060 5 1 1 21059
0 21061 7 2 2 61783 67746
0 21062 7 1 2 76633 89442
0 21063 5 1 1 21062
0 21064 7 1 2 21060 21063
0 21065 5 1 1 21064
0 21066 7 1 2 69028 21065
0 21067 5 1 1 21066
0 21068 7 8 2 58498 61784
0 21069 7 2 2 86639 89444
0 21070 7 1 2 67605 89452
0 21071 5 1 1 21070
0 21072 7 6 2 62188 58499
0 21073 7 1 2 89222 89454
0 21074 5 1 1 21073
0 21075 7 1 2 21058 21074
0 21076 5 1 1 21075
0 21077 7 1 2 78289 21076
0 21078 5 1 1 21077
0 21079 7 1 2 21071 21078
0 21080 7 1 2 21067 21079
0 21081 5 1 1 21080
0 21082 7 1 2 62679 21081
0 21083 5 1 1 21082
0 21084 7 2 2 62396 89049
0 21085 7 1 2 89073 89460
0 21086 5 1 1 21085
0 21087 7 1 2 21083 21086
0 21088 5 1 1 21087
0 21089 7 1 2 88404 21088
0 21090 5 1 1 21089
0 21091 7 1 2 63765 88691
0 21092 7 1 2 86645 21091
0 21093 7 1 2 81019 88834
0 21094 7 1 2 21092 21093
0 21095 5 1 1 21094
0 21096 7 1 2 21090 21095
0 21097 7 1 2 21056 21096
0 21098 5 1 1 21097
0 21099 7 1 2 78242 72310
0 21100 7 1 2 89375 21099
0 21101 7 1 2 21098 21100
0 21102 5 1 1 21101
0 21103 7 1 2 21006 21102
0 21104 7 1 2 20868 21103
0 21105 7 1 2 20217 21104
0 21106 5 1 1 21105
0 21107 7 1 2 65888 21106
0 21108 5 1 1 21107
0 21109 7 1 2 19769 21108
0 21110 7 1 2 19280 21109
0 21111 5 1 1 21110
0 21112 7 1 2 87932 21111
0 21113 5 1 1 21112
0 21114 7 1 2 65265 69793
0 21115 5 7 1 21114
0 21116 7 3 2 61931 87834
0 21117 7 1 2 74538 89469
0 21118 5 2 1 21117
0 21119 7 6 2 64808 65889
0 21120 7 2 2 66583 84368
0 21121 7 1 2 89474 89480
0 21122 5 1 1 21121
0 21123 7 1 2 89472 21122
0 21124 5 1 1 21123
0 21125 7 1 2 89462 21124
0 21126 5 1 1 21125
0 21127 7 2 2 72023 74452
0 21128 5 1 1 89482
0 21129 7 1 2 78535 21128
0 21130 5 1 1 21129
0 21131 7 1 2 76187 21130
0 21132 5 1 1 21131
0 21133 7 1 2 86235 77895
0 21134 5 1 1 21133
0 21135 7 1 2 21132 21134
0 21136 5 2 1 21135
0 21137 7 1 2 61267 89484
0 21138 5 1 1 21137
0 21139 7 1 2 86439 78552
0 21140 5 1 1 21139
0 21141 7 1 2 21138 21140
0 21142 5 1 1 21141
0 21143 7 1 2 66967 21142
0 21144 5 1 1 21143
0 21145 7 1 2 21126 21144
0 21146 5 1 1 21145
0 21147 7 1 2 59789 21146
0 21148 5 1 1 21147
0 21149 7 1 2 65890 72631
0 21150 7 1 2 82542 89463
0 21151 7 1 2 21149 21150
0 21152 5 1 1 21151
0 21153 7 1 2 21148 21152
0 21154 5 1 1 21153
0 21155 7 1 2 61785 21154
0 21156 5 1 1 21155
0 21157 7 1 2 76188 68939
0 21158 5 1 1 21157
0 21159 7 1 2 67184 86530
0 21160 5 1 1 21159
0 21161 7 1 2 21158 21160
0 21162 5 1 1 21161
0 21163 7 1 2 71811 21162
0 21164 5 1 1 21163
0 21165 7 3 2 64809 81897
0 21166 5 1 1 89486
0 21167 7 1 2 76883 89487
0 21168 5 1 1 21167
0 21169 7 1 2 21164 21168
0 21170 5 1 1 21169
0 21171 7 3 2 66422 79161
0 21172 7 1 2 61268 89489
0 21173 7 1 2 21170 21172
0 21174 5 1 1 21173
0 21175 7 1 2 66198 21174
0 21176 7 1 2 21156 21175
0 21177 5 1 1 21176
0 21178 7 1 2 74967 75078
0 21179 5 1 1 21178
0 21180 7 2 2 73828 21179
0 21181 7 5 2 65577 61786
0 21182 7 1 2 66968 89494
0 21183 7 1 2 89492 21182
0 21184 5 1 1 21183
0 21185 7 1 2 76189 77970
0 21186 5 1 1 21185
0 21187 7 1 2 78025 21186
0 21188 5 1 1 21187
0 21189 7 1 2 67044 89254
0 21190 7 1 2 21188 21189
0 21191 5 1 1 21190
0 21192 7 1 2 21184 21191
0 21193 5 1 1 21192
0 21194 7 1 2 65891 21193
0 21195 5 1 1 21194
0 21196 7 13 2 61269 66423
0 21197 7 1 2 71371 89499
0 21198 7 1 2 85687 21197
0 21199 7 1 2 83397 21198
0 21200 5 1 1 21199
0 21201 7 1 2 61590 21200
0 21202 7 1 2 21195 21201
0 21203 5 1 1 21202
0 21204 7 1 2 58500 21203
0 21205 7 1 2 21177 21204
0 21206 5 1 1 21205
0 21207 7 1 2 72897 87708
0 21208 5 1 1 21207
0 21209 7 1 2 73620 69506
0 21210 5 4 1 21209
0 21211 7 1 2 21208 89512
0 21212 5 1 1 21211
0 21213 7 1 2 66199 21212
0 21214 5 1 1 21213
0 21215 7 3 2 73660 81443
0 21216 5 1 1 89516
0 21217 7 1 2 65578 89517
0 21218 5 3 1 21217
0 21219 7 1 2 21214 89519
0 21220 5 1 1 21219
0 21221 7 1 2 64515 21220
0 21222 5 1 1 21221
0 21223 7 3 2 64298 82551
0 21224 5 3 1 89522
0 21225 7 1 2 71812 73255
0 21226 5 3 1 21225
0 21227 7 2 2 86211 89528
0 21228 5 3 1 89531
0 21229 7 1 2 89523 89533
0 21230 5 1 1 21229
0 21231 7 1 2 21222 21230
0 21232 5 1 1 21231
0 21233 7 2 2 60121 80865
0 21234 7 1 2 88902 89536
0 21235 7 1 2 21232 21234
0 21236 5 1 1 21235
0 21237 7 1 2 21206 21236
0 21238 5 1 1 21237
0 21239 7 1 2 62074 21238
0 21240 5 1 1 21239
0 21241 7 1 2 77452 87754
0 21242 5 1 1 21241
0 21243 7 1 2 78558 21242
0 21244 5 1 1 21243
0 21245 7 1 2 61270 21244
0 21246 5 1 1 21245
0 21247 7 4 2 72083 84369
0 21248 5 1 1 89538
0 21249 7 1 2 86196 89539
0 21250 5 1 1 21249
0 21251 7 1 2 21246 21250
0 21252 5 2 1 21251
0 21253 7 1 2 66969 89542
0 21254 5 1 1 21253
0 21255 7 3 2 61271 72024
0 21256 5 1 1 89544
0 21257 7 1 2 65892 84748
0 21258 5 1 1 21257
0 21259 7 1 2 21256 21258
0 21260 5 2 1 21259
0 21261 7 1 2 85688 89547
0 21262 5 1 1 21261
0 21263 7 1 2 84370 86117
0 21264 5 2 1 21263
0 21265 7 2 2 21262 89549
0 21266 5 1 1 89551
0 21267 7 1 2 15485 89552
0 21268 5 1 1 21267
0 21269 7 1 2 67045 21268
0 21270 5 1 1 21269
0 21271 7 1 2 21254 21270
0 21272 5 1 1 21271
0 21273 7 1 2 66200 21272
0 21274 5 1 1 21273
0 21275 7 1 2 87476 72454
0 21276 5 1 1 21275
0 21277 7 1 2 21274 21276
0 21278 5 1 1 21277
0 21279 7 1 2 66424 21278
0 21280 5 1 1 21279
0 21281 7 1 2 62951 86079
0 21282 5 1 1 21281
0 21283 7 1 2 84528 21282
0 21284 5 1 1 21283
0 21285 7 1 2 67185 21284
0 21286 5 1 1 21285
0 21287 7 1 2 87715 21286
0 21288 5 4 1 21287
0 21289 7 2 2 82676 88692
0 21290 7 2 2 89553 89557
0 21291 5 1 1 89559
0 21292 7 1 2 60122 89560
0 21293 5 1 1 21292
0 21294 7 1 2 64516 21293
0 21295 7 1 2 21280 21294
0 21296 5 1 1 21295
0 21297 7 2 2 64299 86531
0 21298 5 1 1 89561
0 21299 7 1 2 68943 21298
0 21300 5 1 1 21299
0 21301 7 1 2 71813 71271
0 21302 7 1 2 21300 21301
0 21303 5 1 1 21302
0 21304 7 1 2 60910 89562
0 21305 5 1 1 21304
0 21306 7 1 2 21303 21305
0 21307 5 1 1 21306
0 21308 7 1 2 66201 21307
0 21309 5 1 1 21308
0 21310 7 1 2 81497 72501
0 21311 5 1 1 21310
0 21312 7 1 2 21309 21311
0 21313 5 1 1 21312
0 21314 7 1 2 67186 21313
0 21315 5 1 1 21314
0 21316 7 3 2 62952 81393
0 21317 7 1 2 77901 89563
0 21318 5 1 1 21317
0 21319 7 1 2 8375 21318
0 21320 5 1 1 21319
0 21321 7 1 2 71272 67046
0 21322 7 1 2 21320 21321
0 21323 5 1 1 21322
0 21324 7 1 2 21315 21323
0 21325 5 1 1 21324
0 21326 7 1 2 89500 21325
0 21327 5 1 1 21326
0 21328 7 7 2 60123 61591
0 21329 7 2 2 88903 89566
0 21330 7 1 2 78038 89573
0 21331 5 1 1 21330
0 21332 7 25 2 66202 61787
0 21333 7 4 2 66584 89575
0 21334 7 1 2 74125 69140
0 21335 7 1 2 89464 21334
0 21336 7 1 2 89600 21335
0 21337 5 1 1 21336
0 21338 7 1 2 21331 21337
0 21339 5 1 1 21338
0 21340 7 1 2 65893 21339
0 21341 5 1 1 21340
0 21342 7 1 2 59790 21341
0 21343 7 1 2 21327 21342
0 21344 5 1 1 21343
0 21345 7 1 2 21296 21344
0 21346 5 1 1 21345
0 21347 7 9 2 66203 88904
0 21348 7 1 2 85376 89604
0 21349 7 1 2 89548 21348
0 21350 5 1 1 21349
0 21351 7 1 2 21346 21350
0 21352 5 1 1 21351
0 21353 7 1 2 62075 21352
0 21354 5 1 1 21353
0 21355 7 1 2 65579 81846
0 21356 5 4 1 21355
0 21357 7 3 2 72968 88920
0 21358 7 1 2 89436 89617
0 21359 7 1 2 85638 21358
0 21360 7 1 2 89613 21359
0 21361 5 1 1 21360
0 21362 7 1 2 21354 21361
0 21363 5 1 1 21362
0 21364 7 1 2 63246 21363
0 21365 5 1 1 21364
0 21366 7 1 2 21240 21365
0 21367 5 1 1 21366
0 21368 7 1 2 62397 21367
0 21369 5 1 1 21368
0 21370 7 2 2 85722 89576
0 21371 5 2 1 89620
0 21372 7 9 2 65894 89577
0 21373 5 2 1 89624
0 21374 7 27 2 61592 66425
0 21375 7 2 2 72860 89635
0 21376 5 1 1 89662
0 21377 7 1 2 89633 21376
0 21378 5 4 1 21377
0 21379 7 2 2 60911 89664
0 21380 7 1 2 71814 89668
0 21381 5 1 1 21380
0 21382 7 1 2 89622 21381
0 21383 5 1 1 21382
0 21384 7 1 2 76190 21383
0 21385 5 1 1 21384
0 21386 7 3 2 64300 61788
0 21387 7 2 2 66204 89670
0 21388 7 1 2 85511 89673
0 21389 5 1 1 21388
0 21390 7 1 2 21385 21389
0 21391 5 1 1 21390
0 21392 7 1 2 76634 21391
0 21393 5 1 1 21392
0 21394 7 1 2 58501 85617
0 21395 5 4 1 21394
0 21396 7 4 2 73309 89578
0 21397 5 2 1 89679
0 21398 7 4 2 66426 84777
0 21399 7 1 2 77948 89685
0 21400 5 1 1 21399
0 21401 7 1 2 89683 21400
0 21402 5 3 1 21401
0 21403 7 1 2 80778 89689
0 21404 7 1 2 89675 21403
0 21405 5 1 1 21404
0 21406 7 1 2 21393 21405
0 21407 5 1 1 21406
0 21408 7 1 2 60335 21407
0 21409 5 1 1 21408
0 21410 7 9 2 65580 86464
0 21411 5 2 1 89692
0 21412 7 1 2 87222 89701
0 21413 5 2 1 21412
0 21414 7 3 2 61789 73829
0 21415 7 1 2 58502 89705
0 21416 7 1 2 89703 21415
0 21417 5 1 1 21416
0 21418 7 1 2 21409 21417
0 21419 5 1 1 21418
0 21420 7 1 2 67047 21419
0 21421 5 1 1 21420
0 21422 7 2 2 59357 88226
0 21423 5 1 1 89708
0 21424 7 2 2 70662 71094
0 21425 5 1 1 89710
0 21426 7 1 2 60336 21425
0 21427 5 1 1 21426
0 21428 7 1 2 21423 21427
0 21429 5 1 1 21428
0 21430 7 1 2 73716 21429
0 21431 5 1 1 21430
0 21432 7 1 2 77980 78561
0 21433 5 1 1 21432
0 21434 7 1 2 21248 21433
0 21435 5 1 1 21434
0 21436 7 1 2 59791 21435
0 21437 5 1 1 21436
0 21438 7 1 2 21431 21437
0 21439 5 1 1 21438
0 21440 7 1 2 65895 21439
0 21441 5 1 1 21440
0 21442 7 6 2 59553 76191
0 21443 7 1 2 72084 89712
0 21444 5 1 1 21443
0 21445 7 1 2 69507 83201
0 21446 5 1 1 21445
0 21447 7 1 2 21444 21446
0 21448 5 1 1 21447
0 21449 7 1 2 73497 21448
0 21450 5 1 1 21449
0 21451 7 1 2 21441 21450
0 21452 5 1 1 21451
0 21453 7 1 2 66205 21452
0 21454 5 1 1 21453
0 21455 7 1 2 59358 86465
0 21456 7 2 2 79540 21455
0 21457 5 1 1 89718
0 21458 7 1 2 73830 89719
0 21459 5 1 1 21458
0 21460 7 1 2 21454 21459
0 21461 5 1 1 21460
0 21462 7 1 2 61790 21461
0 21463 5 1 1 21462
0 21464 7 1 2 86903 73362
0 21465 5 1 1 21464
0 21466 7 1 2 87313 73521
0 21467 5 4 1 21466
0 21468 7 1 2 77920 87596
0 21469 7 1 2 89720 21468
0 21470 5 1 1 21469
0 21471 7 1 2 21465 21470
0 21472 5 1 1 21471
0 21473 7 1 2 72085 21472
0 21474 5 1 1 21473
0 21475 7 1 2 73043 80199
0 21476 5 1 1 21475
0 21477 7 2 2 70203 78562
0 21478 5 1 1 89724
0 21479 7 1 2 73005 89725
0 21480 5 1 1 21479
0 21481 7 1 2 21476 21480
0 21482 5 1 1 21481
0 21483 7 1 2 64517 21482
0 21484 5 1 1 21483
0 21485 7 1 2 21474 21484
0 21486 5 1 1 21485
0 21487 7 3 2 66427 82677
0 21488 7 1 2 21486 89726
0 21489 5 1 1 21488
0 21490 7 1 2 58503 21489
0 21491 7 1 2 21463 21490
0 21492 5 1 1 21491
0 21493 7 3 2 59792 89636
0 21494 7 1 2 72940 78563
0 21495 5 1 1 21494
0 21496 7 1 2 73593 78435
0 21497 5 1 1 21496
0 21498 7 1 2 21495 21497
0 21499 5 1 1 21498
0 21500 7 1 2 89729 21499
0 21501 5 1 1 21500
0 21502 7 6 2 64518 89637
0 21503 5 1 1 89732
0 21504 7 1 2 69723 70691
0 21505 5 1 1 21504
0 21506 7 1 2 89733 21505
0 21507 5 1 1 21506
0 21508 7 1 2 89711 21507
0 21509 5 1 1 21508
0 21510 7 5 2 59793 89579
0 21511 5 6 1 89738
0 21512 7 1 2 21503 89743
0 21513 5 3 1 21512
0 21514 7 1 2 59554 89749
0 21515 7 1 2 21509 21514
0 21516 5 1 1 21515
0 21517 7 1 2 21501 21516
0 21518 5 1 1 21517
0 21519 7 1 2 65896 21518
0 21520 5 1 1 21519
0 21521 7 1 2 73847 89638
0 21522 7 1 2 6826 21521
0 21523 5 1 1 21522
0 21524 7 1 2 21520 21523
0 21525 5 1 1 21524
0 21526 7 1 2 60337 21525
0 21527 5 1 1 21526
0 21528 7 5 2 73661 82405
0 21529 7 1 2 61791 89752
0 21530 7 1 2 89709 21529
0 21531 5 1 1 21530
0 21532 7 1 2 63247 21531
0 21533 7 1 2 21527 21532
0 21534 5 1 1 21533
0 21535 7 1 2 66970 21534
0 21536 7 1 2 21492 21535
0 21537 5 1 1 21536
0 21538 7 1 2 21421 21537
0 21539 5 1 1 21538
0 21540 7 1 2 62076 21539
0 21541 5 1 1 21540
0 21542 7 1 2 21369 21541
0 21543 5 1 1 21542
0 21544 7 1 2 63616 21543
0 21545 5 1 1 21544
0 21546 7 2 2 89399 89554
0 21547 7 1 2 71372 89757
0 21548 5 1 1 21547
0 21549 7 2 2 59555 79323
0 21550 7 2 2 61932 89690
0 21551 7 1 2 89759 89761
0 21552 5 1 1 21551
0 21553 7 2 2 72025 86466
0 21554 5 3 1 89763
0 21555 7 1 2 87223 89765
0 21556 5 1 1 21555
0 21557 7 1 2 59556 21556
0 21558 5 1 1 21557
0 21559 7 1 2 66206 21266
0 21560 5 1 1 21559
0 21561 7 1 2 21558 21560
0 21562 5 1 1 21561
0 21563 7 1 2 88905 21562
0 21564 5 1 1 21563
0 21565 7 1 2 21291 21564
0 21566 5 1 1 21565
0 21567 7 1 2 64519 21566
0 21568 5 1 1 21567
0 21569 7 5 2 78479 81394
0 21570 5 2 1 89768
0 21571 7 1 2 87287 89769
0 21572 5 1 1 21571
0 21573 7 3 2 61593 71273
0 21574 5 1 1 89775
0 21575 7 1 2 74731 89532
0 21576 5 1 1 21575
0 21577 7 1 2 89776 21576
0 21578 5 1 1 21577
0 21579 7 1 2 21572 21578
0 21580 5 1 1 21579
0 21581 7 1 2 59794 21580
0 21582 5 1 1 21581
0 21583 7 1 2 59795 77949
0 21584 5 1 1 21583
0 21585 7 1 2 79583 21584
0 21586 5 1 1 21585
0 21587 7 1 2 62953 21586
0 21588 5 1 1 21587
0 21589 7 1 2 78094 21588
0 21590 5 1 1 21589
0 21591 7 1 2 66207 21590
0 21592 5 1 1 21591
0 21593 7 1 2 72844 81498
0 21594 5 2 1 21593
0 21595 7 1 2 61272 89778
0 21596 7 1 2 21592 21595
0 21597 5 1 1 21596
0 21598 7 1 2 82552 78035
0 21599 5 1 1 21598
0 21600 7 1 2 84122 81367
0 21601 5 1 1 21600
0 21602 7 1 2 65897 21601
0 21603 7 1 2 21599 21602
0 21604 5 1 1 21603
0 21605 7 1 2 67187 21604
0 21606 7 1 2 21597 21605
0 21607 5 1 1 21606
0 21608 7 1 2 21582 21607
0 21609 5 1 1 21608
0 21610 7 1 2 88906 21609
0 21611 5 1 1 21610
0 21612 7 1 2 21568 21611
0 21613 5 1 1 21612
0 21614 7 1 2 62398 21613
0 21615 5 1 1 21614
0 21616 7 1 2 21552 21615
0 21617 5 1 1 21616
0 21618 7 1 2 64810 21617
0 21619 5 1 1 21618
0 21620 7 1 2 21548 21619
0 21621 5 2 1 21620
0 21622 7 1 2 63248 89780
0 21623 5 1 1 21622
0 21624 7 3 2 73292 89465
0 21625 5 1 1 89782
0 21626 7 2 2 73044 89783
0 21627 5 1 1 89785
0 21628 7 1 2 60912 89786
0 21629 5 1 1 21628
0 21630 7 5 2 64301 86118
0 21631 5 2 1 89787
0 21632 7 1 2 76192 89788
0 21633 5 1 1 21632
0 21634 7 1 2 21629 21633
0 21635 5 1 1 21634
0 21636 7 1 2 66208 21635
0 21637 5 1 1 21636
0 21638 7 1 2 74126 86467
0 21639 5 2 1 21638
0 21640 7 1 2 21637 89794
0 21641 5 1 1 21640
0 21642 7 1 2 59796 21641
0 21643 5 1 1 21642
0 21644 7 2 2 85324 86556
0 21645 5 1 1 89796
0 21646 7 1 2 60338 89797
0 21647 5 1 1 21646
0 21648 7 1 2 21643 21647
0 21649 5 1 1 21648
0 21650 7 1 2 61792 21649
0 21651 5 1 1 21650
0 21652 7 1 2 61793 84173
0 21653 7 2 2 85512 21652
0 21654 7 1 2 59797 89798
0 21655 5 1 1 21654
0 21656 7 4 2 62399 61594
0 21657 7 1 2 89255 89800
0 21658 7 1 2 89534 21657
0 21659 5 1 1 21658
0 21660 7 1 2 21655 21659
0 21661 5 1 1 21660
0 21662 7 1 2 85689 21661
0 21663 5 1 1 21662
0 21664 7 1 2 86512 87224
0 21665 5 1 1 21664
0 21666 7 2 2 62400 64520
0 21667 7 1 2 85470 89804
0 21668 7 1 2 21665 21667
0 21669 5 1 1 21668
0 21670 7 6 2 64521 60339
0 21671 7 2 2 59557 89806
0 21672 5 1 1 89812
0 21673 7 5 2 60340 76193
0 21674 5 1 1 89814
0 21675 7 1 2 78075 89815
0 21676 5 1 1 21675
0 21677 7 1 2 21672 21676
0 21678 5 1 1 21677
0 21679 7 2 2 71815 80423
0 21680 7 1 2 61595 89819
0 21681 7 1 2 21678 21680
0 21682 5 1 1 21681
0 21683 7 1 2 21669 21682
0 21684 5 1 1 21683
0 21685 7 1 2 66428 21684
0 21686 5 1 1 21685
0 21687 7 1 2 21663 21686
0 21688 7 1 2 21651 21687
0 21689 5 1 1 21688
0 21690 7 1 2 58504 21689
0 21691 5 1 1 21690
0 21692 7 1 2 87358 88940
0 21693 5 1 1 21692
0 21694 7 4 2 59798 82678
0 21695 5 5 1 89821
0 21696 7 1 2 17323 89825
0 21697 5 1 1 21696
0 21698 7 1 2 73045 21697
0 21699 5 1 1 21698
0 21700 7 1 2 82591 15919
0 21701 5 8 1 21700
0 21702 7 1 2 62401 73006
0 21703 7 1 2 89830 21702
0 21704 5 1 1 21703
0 21705 7 1 2 21699 21704
0 21706 5 1 1 21705
0 21707 7 1 2 72763 21706
0 21708 5 1 1 21707
0 21709 7 1 2 21693 21708
0 21710 5 1 1 21709
0 21711 7 1 2 66429 21710
0 21712 5 1 1 21711
0 21713 7 1 2 89680 89760
0 21714 5 1 1 21713
0 21715 7 1 2 21712 21714
0 21716 5 1 1 21715
0 21717 7 1 2 80866 21716
0 21718 5 1 1 21717
0 21719 7 1 2 21691 21718
0 21720 5 1 1 21719
0 21721 7 2 2 71067 21720
0 21722 5 1 1 89838
0 21723 7 1 2 21623 21722
0 21724 5 1 1 21723
0 21725 7 1 2 68664 21724
0 21726 5 1 1 21725
0 21727 7 1 2 21545 21726
0 21728 5 1 1 21727
0 21729 7 1 2 66772 21728
0 21730 5 1 1 21729
0 21731 7 1 2 63617 89781
0 21732 5 1 1 21731
0 21733 7 1 2 88105 89758
0 21734 5 1 1 21733
0 21735 7 1 2 21732 21734
0 21736 5 1 1 21735
0 21737 7 1 2 63249 21736
0 21738 5 1 1 21737
0 21739 7 1 2 63618 89839
0 21740 5 1 1 21739
0 21741 7 1 2 21738 21740
0 21742 5 1 1 21741
0 21743 7 1 2 74247 21742
0 21744 5 1 1 21743
0 21745 7 2 2 21730 21744
0 21746 5 1 1 89840
0 21747 7 1 2 64875 21746
0 21748 5 1 1 21747
0 21749 7 3 2 62077 88717
0 21750 7 1 2 87928 89842
0 21751 7 1 2 89555 21750
0 21752 5 1 1 21751
0 21753 7 1 2 21748 21752
0 21754 5 1 1 21753
0 21755 7 1 2 58912 21754
0 21756 5 1 1 21755
0 21757 7 1 2 60182 89841
0 21758 5 1 1 21757
0 21759 7 4 2 62954 75439
0 21760 5 3 1 89845
0 21761 7 1 2 82907 89849
0 21762 5 3 1 21761
0 21763 7 1 2 69390 89734
0 21764 5 1 1 21763
0 21765 7 1 2 63883 89739
0 21766 5 1 1 21765
0 21767 7 1 2 21764 21766
0 21768 5 1 1 21767
0 21769 7 1 2 89852 21768
0 21770 5 1 1 21769
0 21771 7 6 2 60563 66430
0 21772 7 2 2 82679 89855
0 21773 7 3 2 80802 78076
0 21774 7 1 2 89861 89863
0 21775 5 1 1 21774
0 21776 7 1 2 66209 80659
0 21777 5 1 1 21776
0 21778 7 1 2 89826 21777
0 21779 5 1 1 21778
0 21780 7 6 2 59558 61794
0 21781 7 5 2 81037 89866
0 21782 5 1 1 89872
0 21783 7 1 2 21779 89873
0 21784 5 1 1 21783
0 21785 7 1 2 21775 21784
0 21786 7 1 2 21770 21785
0 21787 5 1 1 21786
0 21788 7 1 2 64041 21787
0 21789 5 1 1 21788
0 21790 7 10 2 61596 61795
0 21791 7 2 2 77939 89877
0 21792 7 1 2 86283 79324
0 21793 7 1 2 89887 21792
0 21794 5 1 1 21793
0 21795 7 1 2 65581 21794
0 21796 7 1 2 21789 21795
0 21797 5 1 1 21796
0 21798 7 2 2 63884 66210
0 21799 7 2 2 59799 88731
0 21800 7 1 2 89889 89891
0 21801 5 1 1 21800
0 21802 7 1 2 74965 89735
0 21803 5 1 1 21802
0 21804 7 1 2 21801 21803
0 21805 5 1 1 21804
0 21806 7 1 2 89853 21805
0 21807 5 1 1 21806
0 21808 7 1 2 84055 89278
0 21809 5 1 1 21808
0 21810 7 20 2 66211 66431
0 21811 7 1 2 70688 89893
0 21812 7 1 2 80680 21811
0 21813 5 1 1 21812
0 21814 7 1 2 21809 21813
0 21815 5 1 1 21814
0 21816 7 1 2 60341 21815
0 21817 5 1 1 21816
0 21818 7 6 2 58505 89580
0 21819 5 1 1 89913
0 21820 7 2 2 79639 89914
0 21821 5 1 1 89919
0 21822 7 1 2 74453 89920
0 21823 5 1 1 21822
0 21824 7 4 2 71402 89639
0 21825 7 6 2 63250 60564
0 21826 5 3 1 89925
0 21827 7 1 2 72668 89926
0 21828 7 1 2 89921 21827
0 21829 5 1 1 21828
0 21830 7 1 2 60913 21829
0 21831 7 1 2 21823 21830
0 21832 7 1 2 21817 21831
0 21833 7 1 2 21807 21832
0 21834 5 1 1 21833
0 21835 7 1 2 65898 21834
0 21836 7 1 2 21797 21835
0 21837 5 1 1 21836
0 21838 7 1 2 85622 86087
0 21839 7 3 2 82406 89867
0 21840 7 1 2 79773 89934
0 21841 7 1 2 21838 21840
0 21842 5 1 1 21841
0 21843 7 3 2 21837 21842
0 21844 5 1 1 89937
0 21845 7 1 2 64811 21844
0 21846 5 1 1 21845
0 21847 7 2 2 69757 79409
0 21848 5 2 1 89940
0 21849 7 1 2 77708 89942
0 21850 5 2 1 21849
0 21851 7 1 2 79413 75074
0 21852 5 1 1 21851
0 21853 7 1 2 89944 21852
0 21854 5 3 1 21853
0 21855 7 1 2 64522 88849
0 21856 7 1 2 89946 21855
0 21857 5 1 1 21856
0 21858 7 1 2 58506 21857
0 21859 5 1 1 21858
0 21860 7 2 2 61597 21859
0 21861 7 3 2 59800 88850
0 21862 7 1 2 89947 89951
0 21863 5 1 1 21862
0 21864 7 2 2 61796 89614
0 21865 7 2 2 85635 84113
0 21866 7 1 2 89954 89956
0 21867 5 1 1 21866
0 21868 7 1 2 63251 21867
0 21869 7 1 2 21863 21868
0 21870 5 2 1 21869
0 21871 7 1 2 89949 89958
0 21872 5 1 1 21871
0 21873 7 1 2 69889 75143
0 21874 5 1 1 21873
0 21875 7 1 2 83548 21874
0 21876 5 1 1 21875
0 21877 7 1 2 59559 21876
0 21878 5 1 1 21877
0 21879 7 1 2 59359 87778
0 21880 5 1 1 21879
0 21881 7 1 2 21878 21880
0 21882 5 1 1 21881
0 21883 7 3 2 89581 21882
0 21884 7 1 2 85453 89960
0 21885 5 1 1 21884
0 21886 7 1 2 21872 21885
0 21887 5 1 1 21886
0 21888 7 1 2 61273 21887
0 21889 5 1 1 21888
0 21890 7 1 2 80803 75101
0 21891 7 1 2 89490 21890
0 21892 5 1 1 21891
0 21893 7 3 2 59560 77863
0 21894 7 1 2 77717 7736
0 21895 5 2 1 21894
0 21896 7 1 2 61797 89966
0 21897 7 1 2 89963 21896
0 21898 5 1 1 21897
0 21899 7 1 2 21892 21898
0 21900 5 1 1 21899
0 21901 7 1 2 66212 21900
0 21902 5 1 1 21901
0 21903 7 7 2 59801 72652
0 21904 7 2 2 61798 82680
0 21905 7 1 2 69972 89975
0 21906 7 1 2 89968 21905
0 21907 5 1 1 21906
0 21908 7 1 2 21902 21907
0 21909 5 1 1 21908
0 21910 7 1 2 65582 21909
0 21911 5 1 1 21910
0 21912 7 2 2 72147 69923
0 21913 7 1 2 87014 89740
0 21914 7 1 2 89977 21913
0 21915 5 1 1 21914
0 21916 7 1 2 21911 21915
0 21917 5 1 1 21916
0 21918 7 3 2 65899 21917
0 21919 5 1 1 89979
0 21920 7 1 2 64812 89980
0 21921 5 1 1 21920
0 21922 7 1 2 21889 21921
0 21923 5 1 1 21922
0 21924 7 1 2 62680 21923
0 21925 5 1 1 21924
0 21926 7 1 2 21846 21925
0 21927 5 1 1 21926
0 21928 7 1 2 61933 21927
0 21929 5 1 1 21928
0 21930 7 2 2 71403 70735
0 21931 7 5 2 82096 88394
0 21932 7 1 2 80221 78390
0 21933 7 1 2 89984 21932
0 21934 7 1 2 89982 21933
0 21935 5 1 1 21934
0 21936 7 1 2 58859 21935
0 21937 7 1 2 21929 21936
0 21938 5 1 1 21937
0 21939 7 1 2 76635 89961
0 21940 5 1 1 21939
0 21941 7 2 2 66432 76672
0 21942 7 1 2 61598 89989
0 21943 7 1 2 89948 21942
0 21944 5 1 1 21943
0 21945 7 1 2 21940 21944
0 21946 5 1 1 21945
0 21947 7 1 2 61274 75572
0 21948 7 1 2 21946 21947
0 21949 5 1 1 21948
0 21950 7 1 2 21919 21949
0 21951 5 1 1 21950
0 21952 7 1 2 62681 21951
0 21953 5 1 1 21952
0 21954 7 1 2 89938 21953
0 21955 5 1 1 21954
0 21956 7 1 2 67048 21955
0 21957 5 1 1 21956
0 21958 7 1 2 62955 79695
0 21959 7 2 2 61275 89927
0 21960 5 1 1 89991
0 21961 7 8 2 65583 89894
0 21962 7 1 2 89992 89993
0 21963 7 1 2 21958 21962
0 21964 5 1 1 21963
0 21965 7 4 2 81253 89223
0 21966 5 2 1 90001
0 21967 7 5 2 59561 78983
0 21968 5 6 1 90007
0 21969 7 1 2 79355 90008
0 21970 7 1 2 90002 21969
0 21971 5 1 1 21970
0 21972 7 1 2 21964 21971
0 21973 5 1 1 21972
0 21974 7 1 2 59127 21973
0 21975 5 1 1 21974
0 21976 7 2 2 78077 87015
0 21977 5 1 1 90018
0 21978 7 1 2 85241 21977
0 21979 5 4 1 21978
0 21980 7 10 2 61276 89640
0 21981 7 1 2 73115 90024
0 21982 5 2 1 21981
0 21983 7 1 2 70169 89625
0 21984 5 1 1 21983
0 21985 7 1 2 90034 21984
0 21986 5 1 1 21985
0 21987 7 1 2 90020 21986
0 21988 5 1 1 21987
0 21989 7 2 2 61277 89582
0 21990 7 1 2 86288 79348
0 21991 7 1 2 90036 21990
0 21992 5 1 1 21991
0 21993 7 1 2 21988 21992
0 21994 5 1 1 21993
0 21995 7 1 2 85257 21994
0 21996 5 1 1 21995
0 21997 7 3 2 64042 72026
0 21998 5 4 1 90038
0 21999 7 1 2 72294 90041
0 22000 5 3 1 21999
0 22001 7 1 2 85545 81428
0 22002 7 1 2 89706 22001
0 22003 7 1 2 90045 22002
0 22004 5 1 1 22003
0 22005 7 1 2 21996 22004
0 22006 5 1 1 22005
0 22007 7 1 2 62682 22006
0 22008 5 1 1 22007
0 22009 7 1 2 21975 22008
0 22010 5 1 1 22009
0 22011 7 1 2 64813 22010
0 22012 5 1 1 22011
0 22013 7 2 2 87784 75057
0 22014 7 2 2 88395 88237
0 22015 7 1 2 79918 90050
0 22016 7 1 2 90048 22015
0 22017 5 1 1 22016
0 22018 7 1 2 22012 22017
0 22019 5 1 1 22018
0 22020 7 1 2 66585 22019
0 22021 5 1 1 22020
0 22022 7 1 2 63619 22021
0 22023 7 1 2 21957 22022
0 22024 5 1 1 22023
0 22025 7 1 2 66773 22024
0 22026 7 1 2 21938 22025
0 22027 5 1 1 22026
0 22028 7 1 2 62683 89981
0 22029 5 1 1 22028
0 22030 7 1 2 22029 89939
0 22031 5 1 1 22030
0 22032 7 1 2 69535 22031
0 22033 5 1 1 22032
0 22034 7 10 2 62684 61278
0 22035 7 1 2 88983 89962
0 22036 5 1 1 22035
0 22037 7 1 2 63620 89959
0 22038 5 1 1 22037
0 22039 7 1 2 75516 70453
0 22040 7 1 2 86014 22039
0 22041 7 1 2 89955 22040
0 22042 5 1 1 22041
0 22043 7 1 2 22038 22042
0 22044 5 1 1 22043
0 22045 7 1 2 89950 22044
0 22046 5 1 1 22045
0 22047 7 1 2 22036 22046
0 22048 5 1 1 22047
0 22049 7 1 2 90052 22048
0 22050 5 1 1 22049
0 22051 7 1 2 22033 22050
0 22052 5 1 1 22051
0 22053 7 1 2 61934 22052
0 22054 5 1 1 22053
0 22055 7 2 2 80804 89985
0 22056 7 4 2 62685 69536
0 22057 7 1 2 80660 84031
0 22058 7 1 2 90064 22057
0 22059 7 1 2 90062 22058
0 22060 5 1 1 22059
0 22061 7 1 2 22054 22060
0 22062 5 1 1 22061
0 22063 7 1 2 66830 22062
0 22064 5 1 1 22063
0 22065 7 1 2 66694 22064
0 22066 7 1 2 22027 22065
0 22067 5 1 1 22066
0 22068 7 1 2 85633 89856
0 22069 5 1 1 22068
0 22070 7 1 2 85085 89868
0 22071 5 1 1 22070
0 22072 7 1 2 22069 22071
0 22073 5 1 1 22072
0 22074 7 1 2 63885 22073
0 22075 5 1 1 22074
0 22076 7 1 2 77006 89869
0 22077 5 1 1 22076
0 22078 7 1 2 22075 22077
0 22079 5 1 1 22078
0 22080 7 1 2 59802 22079
0 22081 5 1 1 22080
0 22082 7 1 2 71816 72804
0 22083 7 1 2 89256 22082
0 22084 7 1 2 85481 22083
0 22085 5 1 1 22084
0 22086 7 1 2 22081 22085
0 22087 5 1 1 22086
0 22088 7 1 2 61279 22087
0 22089 5 1 1 22088
0 22090 7 11 2 65900 66433
0 22091 7 1 2 81836 90068
0 22092 7 1 2 80990 22091
0 22093 5 1 1 22092
0 22094 7 1 2 22089 22093
0 22095 5 1 1 22094
0 22096 7 1 2 60914 22095
0 22097 5 1 1 22096
0 22098 7 1 2 85690 86207
0 22099 5 1 1 22098
0 22100 7 1 2 89550 22099
0 22101 5 1 1 22100
0 22102 7 1 2 64523 22101
0 22103 5 1 1 22102
0 22104 7 1 2 65038 85976
0 22105 5 1 1 22104
0 22106 7 1 2 22103 22105
0 22107 5 1 1 22106
0 22108 7 1 2 63252 22107
0 22109 5 1 1 22108
0 22110 7 1 2 85639 86208
0 22111 5 1 1 22110
0 22112 7 1 2 22109 22111
0 22113 5 1 1 22112
0 22114 7 1 2 66434 22113
0 22115 5 1 1 22114
0 22116 7 1 2 22097 22115
0 22117 5 1 1 22116
0 22118 7 1 2 66213 22117
0 22119 5 1 1 22118
0 22120 7 1 2 86212 18261
0 22121 5 1 1 22120
0 22122 7 1 2 76194 77864
0 22123 7 1 2 22121 22122
0 22124 5 1 1 22123
0 22125 7 2 2 77357 74127
0 22126 5 1 1 90079
0 22127 7 1 2 84983 90080
0 22128 5 2 1 22127
0 22129 7 5 2 59803 67188
0 22130 7 1 2 80805 90083
0 22131 5 3 1 22130
0 22132 7 1 2 90081 90088
0 22133 5 1 1 22132
0 22134 7 1 2 65901 22133
0 22135 5 1 1 22134
0 22136 7 1 2 64302 75573
0 22137 7 1 2 89535 22136
0 22138 7 1 2 89676 22137
0 22139 5 1 1 22138
0 22140 7 1 2 22135 22139
0 22141 7 1 2 22124 22140
0 22142 5 1 1 22141
0 22143 7 1 2 89641 22142
0 22144 5 1 1 22143
0 22145 7 1 2 22119 22144
0 22146 5 1 1 22145
0 22147 7 1 2 89038 22146
0 22148 5 1 1 22147
0 22149 7 1 2 80970 81310
0 22150 5 1 1 22149
0 22151 7 1 2 75517 78556
0 22152 5 1 1 22151
0 22153 7 1 2 22150 22152
0 22154 5 1 1 22153
0 22155 7 1 2 66435 22154
0 22156 5 1 1 22155
0 22157 7 1 2 89050 89485
0 22158 5 1 1 22157
0 22159 7 1 2 22156 22158
0 22160 5 1 1 22159
0 22161 7 1 2 84656 22160
0 22162 5 1 1 22161
0 22163 7 1 2 59804 84371
0 22164 5 2 1 22163
0 22165 7 1 2 79406 90091
0 22166 5 1 1 22165
0 22167 7 1 2 58507 22166
0 22168 5 1 1 22167
0 22169 7 1 2 73375 86956
0 22170 5 1 1 22169
0 22171 7 1 2 22168 22170
0 22172 5 1 1 22171
0 22173 7 1 2 89466 22172
0 22174 5 1 1 22173
0 22175 7 6 2 64303 79336
0 22176 5 1 1 90093
0 22177 7 1 2 63886 85623
0 22178 7 1 2 90094 22177
0 22179 5 1 1 22178
0 22180 7 1 2 22174 22179
0 22181 5 1 1 22180
0 22182 7 1 2 66214 22181
0 22183 5 1 1 22182
0 22184 7 3 2 58508 81499
0 22185 5 1 1 90099
0 22186 7 1 2 89493 90100
0 22187 5 1 1 22186
0 22188 7 1 2 61799 22187
0 22189 7 1 2 22183 22188
0 22190 5 1 1 22189
0 22191 7 1 2 75004 87445
0 22192 7 1 2 89540 22191
0 22193 5 1 1 22192
0 22194 7 1 2 66436 22193
0 22195 5 1 1 22194
0 22196 7 1 2 65902 22195
0 22197 7 1 2 22190 22196
0 22198 5 1 1 22197
0 22199 7 1 2 22162 22198
0 22200 5 1 1 22199
0 22201 7 1 2 79973 22200
0 22202 5 1 1 22201
0 22203 7 8 2 60003 82801
0 22204 7 2 2 64524 82681
0 22205 7 6 2 61800 67927
0 22206 7 1 2 90110 90112
0 22207 7 1 2 90102 22206
0 22208 7 1 2 89556 22207
0 22209 5 1 1 22208
0 22210 7 1 2 22202 22209
0 22211 5 1 1 22210
0 22212 7 1 2 66586 22211
0 22213 5 1 1 22212
0 22214 7 1 2 62078 22213
0 22215 7 1 2 22148 22214
0 22216 5 1 1 22215
0 22217 7 1 2 62402 22216
0 22218 7 1 2 22067 22217
0 22219 5 1 1 22218
0 22220 7 1 2 66215 89541
0 22221 5 1 1 22220
0 22222 7 1 2 87102 81354
0 22223 5 1 1 22222
0 22224 7 1 2 22221 22223
0 22225 5 1 1 22224
0 22226 7 1 2 65903 22225
0 22227 5 1 1 22226
0 22228 7 2 2 72086 84657
0 22229 7 1 2 89713 90118
0 22230 5 1 1 22229
0 22231 7 1 2 22227 22230
0 22232 5 2 1 22231
0 22233 7 1 2 76135 90120
0 22234 5 1 1 22233
0 22235 7 2 2 77343 87197
0 22236 7 1 2 82668 90122
0 22237 5 1 1 22236
0 22238 7 1 2 65584 86709
0 22239 7 1 2 89967 22238
0 22240 5 1 1 22239
0 22241 7 1 2 22237 22240
0 22242 5 2 1 22241
0 22243 7 1 2 69271 90124
0 22244 5 1 1 22243
0 22245 7 1 2 64043 83029
0 22246 7 1 2 85515 22245
0 22247 5 1 1 22246
0 22248 7 1 2 22244 22247
0 22249 5 1 1 22248
0 22250 7 1 2 62686 22249
0 22251 5 1 1 22250
0 22252 7 2 2 61599 71059
0 22253 7 1 2 73421 90126
0 22254 7 1 2 83581 22253
0 22255 5 1 1 22254
0 22256 7 1 2 84276 81395
0 22257 7 1 2 69676 22256
0 22258 5 1 1 22257
0 22259 7 1 2 22255 22258
0 22260 5 1 1 22259
0 22261 7 1 2 63887 22260
0 22262 5 1 1 22261
0 22263 7 1 2 84125 69352
0 22264 5 1 1 22263
0 22265 7 1 2 22262 22264
0 22266 5 1 1 22265
0 22267 7 1 2 65904 22266
0 22268 5 1 1 22267
0 22269 7 8 2 66216 71274
0 22270 5 1 1 90128
0 22271 7 1 2 73621 69677
0 22272 7 1 2 90129 22271
0 22273 5 1 1 22272
0 22274 7 1 2 22268 22273
0 22275 7 1 2 22251 22274
0 22276 5 1 1 22275
0 22277 7 1 2 60342 22276
0 22278 5 1 1 22277
0 22279 7 1 2 82248 89704
0 22280 5 1 1 22279
0 22281 7 6 2 65905 66695
0 22282 7 3 2 82711 90136
0 22283 7 1 2 62687 69938
0 22284 7 1 2 90142 22283
0 22285 7 1 2 84257 22284
0 22286 5 1 1 22285
0 22287 7 1 2 22280 22286
0 22288 7 1 2 22278 22287
0 22289 5 1 1 22288
0 22290 7 1 2 75656 22289
0 22291 5 1 1 22290
0 22292 7 1 2 22234 22291
0 22293 5 1 1 22292
0 22294 7 1 2 61801 22293
0 22295 5 1 1 22294
0 22296 7 1 2 81926 20094
0 22297 5 1 1 22296
0 22298 7 1 2 62956 22297
0 22299 5 1 1 22298
0 22300 7 1 2 74982 82051
0 22301 5 1 1 22300
0 22302 7 1 2 22299 22301
0 22303 5 1 1 22302
0 22304 7 1 2 71817 22303
0 22305 5 1 1 22304
0 22306 7 1 2 79997 83130
0 22307 5 1 1 22306
0 22308 7 1 2 22305 22307
0 22309 5 1 1 22308
0 22310 7 1 2 67189 22309
0 22311 5 1 1 22310
0 22312 7 1 2 77303 82035
0 22313 7 1 2 79476 22312
0 22314 5 1 1 22313
0 22315 7 1 2 22311 22314
0 22316 5 1 1 22315
0 22317 7 1 2 89663 22316
0 22318 5 1 1 22317
0 22319 7 1 2 22295 22318
0 22320 5 1 1 22319
0 22321 7 1 2 58509 22320
0 22322 5 1 1 22321
0 22323 7 4 2 60343 62079
0 22324 7 2 2 61935 77424
0 22325 7 1 2 90145 90149
0 22326 7 1 2 83564 22325
0 22327 7 1 2 89691 22326
0 22328 5 1 1 22327
0 22329 7 1 2 22322 22328
0 22330 5 1 1 22329
0 22331 7 1 2 59805 22330
0 22332 5 1 1 22331
0 22333 7 1 2 61802 90121
0 22334 5 1 1 22333
0 22335 7 7 2 77585 89642
0 22336 7 5 2 62688 60344
0 22337 5 4 1 90158
0 22338 7 1 2 75461 90159
0 22339 7 1 2 72087 22338
0 22340 7 1 2 90151 22339
0 22341 5 1 1 22340
0 22342 7 1 2 22334 22341
0 22343 5 1 1 22342
0 22344 7 1 2 74280 22343
0 22345 5 1 1 22344
0 22346 7 1 2 60345 90125
0 22347 5 1 1 22346
0 22348 7 2 2 71404 86557
0 22349 7 1 2 84255 90167
0 22350 5 1 1 22349
0 22351 7 1 2 22347 22350
0 22352 5 1 1 22351
0 22353 7 1 2 62689 22352
0 22354 5 1 1 22353
0 22355 7 1 2 69787 86694
0 22356 7 1 2 78729 22355
0 22357 5 1 1 22356
0 22358 7 1 2 22354 22357
0 22359 5 1 1 22358
0 22360 7 1 2 61803 22359
0 22361 5 1 1 22360
0 22362 7 2 2 70294 89686
0 22363 7 1 2 89983 90169
0 22364 5 1 1 22363
0 22365 7 1 2 22361 22364
0 22366 5 1 1 22365
0 22367 7 1 2 74411 22366
0 22368 5 1 1 22367
0 22369 7 1 2 22345 22368
0 22370 5 1 1 22369
0 22371 7 1 2 76636 22370
0 22372 5 1 1 22371
0 22373 7 1 2 78440 77904
0 22374 5 1 1 22373
0 22375 7 1 2 64044 22374
0 22376 5 1 1 22375
0 22377 7 1 2 78026 22376
0 22378 5 1 1 22377
0 22379 7 14 2 60346 66437
0 22380 7 1 2 84162 90171
0 22381 7 2 2 22378 22380
0 22382 7 1 2 66831 90185
0 22383 5 1 1 22382
0 22384 7 6 2 71176 89583
0 22385 5 1 1 90187
0 22386 7 1 2 75901 90188
0 22387 5 1 1 22386
0 22388 7 1 2 87288 89862
0 22389 5 1 1 22388
0 22390 7 1 2 22387 22389
0 22391 5 1 1 22390
0 22392 7 1 2 65585 22391
0 22393 5 1 1 22392
0 22394 7 3 2 60915 89584
0 22395 7 3 2 59562 70058
0 22396 7 1 2 90193 90196
0 22397 5 1 1 22396
0 22398 7 1 2 22393 22397
0 22399 5 1 1 22398
0 22400 7 2 2 67519 22399
0 22401 7 1 2 66774 90199
0 22402 5 1 1 22401
0 22403 7 1 2 22383 22402
0 22404 5 1 1 22403
0 22405 7 1 2 65906 22404
0 22406 5 1 1 22405
0 22407 7 2 2 82379 74281
0 22408 5 1 1 90201
0 22409 7 1 2 64045 74412
0 22410 7 1 2 87773 22409
0 22411 5 1 1 22410
0 22412 7 1 2 22408 22411
0 22413 5 1 1 22412
0 22414 7 1 2 62957 22413
0 22415 5 1 1 22414
0 22416 7 2 2 87755 84025
0 22417 7 1 2 83654 90203
0 22418 5 1 1 22417
0 22419 7 1 2 22415 22418
0 22420 5 1 1 22419
0 22421 7 1 2 60347 22420
0 22422 5 1 1 22421
0 22423 7 2 2 60565 74473
0 22424 7 2 2 79770 90205
0 22425 7 5 2 61600 67520
0 22426 7 1 2 77344 90209
0 22427 7 1 2 90207 22426
0 22428 5 1 1 22427
0 22429 7 1 2 22422 22428
0 22430 5 1 1 22429
0 22431 7 1 2 89501 22430
0 22432 5 1 1 22431
0 22433 7 1 2 22406 22432
0 22434 5 1 1 22433
0 22435 7 1 2 62690 22434
0 22436 5 1 1 22435
0 22437 7 1 2 84896 79786
0 22438 5 1 1 22437
0 22439 7 1 2 19120 22438
0 22440 5 1 1 22439
0 22441 7 5 2 65907 67469
0 22442 7 1 2 89585 90214
0 22443 7 2 2 22440 22442
0 22444 7 1 2 83655 90219
0 22445 5 1 1 22444
0 22446 7 1 2 86352 89529
0 22447 5 4 1 22446
0 22448 7 5 2 66438 67521
0 22449 7 8 2 62958 61601
0 22450 7 1 2 90225 90230
0 22451 7 2 2 90221 22450
0 22452 7 1 2 83013 90238
0 22453 5 1 1 22452
0 22454 7 1 2 22445 22453
0 22455 5 1 1 22454
0 22456 7 1 2 59360 22455
0 22457 5 1 1 22456
0 22458 7 3 2 78984 89586
0 22459 5 3 1 90240
0 22460 7 1 2 77345 90241
0 22461 5 1 1 22460
0 22462 7 6 2 65908 77981
0 22463 5 4 1 90246
0 22464 7 1 2 14144 90252
0 22465 5 1 1 22464
0 22466 7 1 2 66439 90231
0 22467 7 1 2 22465 22466
0 22468 5 1 1 22467
0 22469 7 1 2 22461 22468
0 22470 5 1 1 22469
0 22471 7 1 2 74248 81916
0 22472 7 1 2 22470 22471
0 22473 5 1 1 22472
0 22474 7 1 2 22457 22473
0 22475 7 1 2 22436 22474
0 22476 5 1 1 22475
0 22477 7 1 2 76734 22476
0 22478 5 1 1 22477
0 22479 7 1 2 62691 74888
0 22480 7 10 2 60004 66217
0 22481 7 1 2 88693 90256
0 22482 7 1 2 22479 22481
0 22483 7 1 2 85238 22482
0 22484 5 1 1 22483
0 22485 7 1 2 78159 77231
0 22486 7 1 2 81355 88907
0 22487 7 1 2 22485 22486
0 22488 7 1 2 74306 22487
0 22489 5 1 1 22488
0 22490 7 1 2 22484 22489
0 22491 5 1 1 22490
0 22492 7 1 2 90222 22491
0 22493 5 1 1 22492
0 22494 7 3 2 75518 90172
0 22495 7 2 2 74927 81500
0 22496 7 1 2 77709 90269
0 22497 5 1 1 22496
0 22498 7 1 2 72088 73171
0 22499 7 1 2 84126 22498
0 22500 5 1 1 22499
0 22501 7 1 2 22497 22500
0 22502 5 2 1 22501
0 22503 7 1 2 74413 90271
0 22504 5 1 1 22503
0 22505 7 2 2 67470 81501
0 22506 7 1 2 59563 74421
0 22507 7 1 2 90273 22506
0 22508 5 1 1 22507
0 22509 7 1 2 22504 22508
0 22510 5 1 1 22509
0 22511 7 1 2 62692 22510
0 22512 5 1 1 22511
0 22513 7 1 2 70713 70692
0 22514 5 2 1 22513
0 22515 7 1 2 90275 90202
0 22516 5 1 1 22515
0 22517 7 1 2 22512 22516
0 22518 5 1 1 22517
0 22519 7 1 2 65909 22518
0 22520 5 1 1 22519
0 22521 7 1 2 84658 67522
0 22522 7 2 2 86904 22521
0 22523 7 1 2 90277 90208
0 22524 5 1 1 22523
0 22525 7 1 2 22520 22524
0 22526 5 1 1 22525
0 22527 7 1 2 90266 22526
0 22528 5 1 1 22527
0 22529 7 1 2 22493 22528
0 22530 7 1 2 22478 22529
0 22531 7 1 2 22372 22530
0 22532 5 1 1 22531
0 22533 7 1 2 70503 22532
0 22534 5 1 1 22533
0 22535 7 1 2 79967 90186
0 22536 5 1 1 22535
0 22537 7 1 2 82065 90200
0 22538 5 1 1 22537
0 22539 7 1 2 22536 22538
0 22540 5 1 1 22539
0 22541 7 1 2 65910 22540
0 22542 5 1 1 22541
0 22543 7 3 2 86330 82617
0 22544 7 1 2 82249 90279
0 22545 5 1 1 22544
0 22546 7 1 2 64304 77000
0 22547 7 1 2 79149 22546
0 22548 7 3 2 64814 70295
0 22549 7 4 2 66696 82655
0 22550 7 1 2 90282 90285
0 22551 7 1 2 22547 22550
0 22552 5 1 1 22551
0 22553 7 1 2 22545 22552
0 22554 5 1 1 22553
0 22555 7 1 2 62959 22554
0 22556 5 1 1 22555
0 22557 7 3 2 71134 81889
0 22558 7 1 2 90289 90204
0 22559 5 1 1 22558
0 22560 7 1 2 22556 22559
0 22561 5 1 1 22560
0 22562 7 1 2 60348 22561
0 22563 5 1 1 22562
0 22564 7 1 2 69577 88238
0 22565 7 1 2 84227 81822
0 22566 7 1 2 22564 22565
0 22567 5 1 1 22566
0 22568 7 1 2 22563 22567
0 22569 5 1 1 22568
0 22570 7 1 2 89502 22569
0 22571 5 1 1 22570
0 22572 7 1 2 22542 22571
0 22573 5 1 1 22572
0 22574 7 1 2 62693 22573
0 22575 5 1 1 22574
0 22576 7 1 2 90290 90220
0 22577 5 1 1 22576
0 22578 7 2 2 80254 83518
0 22579 7 1 2 90239 90292
0 22580 5 1 1 22579
0 22581 7 1 2 22577 22580
0 22582 5 1 1 22581
0 22583 7 1 2 59361 22582
0 22584 5 1 1 22583
0 22585 7 1 2 70654 89626
0 22586 5 1 1 22585
0 22587 7 2 2 75462 89643
0 22588 5 1 1 90294
0 22589 7 1 2 71818 90295
0 22590 5 1 1 22589
0 22591 7 1 2 22586 22590
0 22592 5 1 1 22591
0 22593 7 1 2 77270 22592
0 22594 5 1 1 22593
0 22595 7 1 2 66832 89762
0 22596 5 1 1 22595
0 22597 7 1 2 22594 22596
0 22598 5 1 1 22597
0 22599 7 1 2 59564 22598
0 22600 5 1 1 22599
0 22601 7 1 2 66587 72089
0 22602 7 1 2 87685 89922
0 22603 7 1 2 22601 22602
0 22604 5 1 1 22603
0 22605 7 1 2 22600 22604
0 22606 5 1 1 22605
0 22607 7 1 2 69223 22606
0 22608 5 1 1 22607
0 22609 7 1 2 22584 22608
0 22610 7 1 2 22575 22609
0 22611 5 1 1 22610
0 22612 7 1 2 76735 22611
0 22613 5 1 1 22612
0 22614 7 1 2 81770 90272
0 22615 5 1 1 22614
0 22616 7 2 2 59362 77505
0 22617 7 2 2 63487 61602
0 22618 7 1 2 72436 90298
0 22619 7 1 2 76084 22618
0 22620 7 1 2 90296 22619
0 22621 5 1 1 22620
0 22622 7 1 2 22615 22621
0 22623 5 1 1 22622
0 22624 7 1 2 62694 22623
0 22625 5 1 1 22624
0 22626 7 1 2 84026 90291
0 22627 7 1 2 90276 22626
0 22628 5 1 1 22627
0 22629 7 1 2 22625 22628
0 22630 5 1 1 22629
0 22631 7 1 2 65911 22630
0 22632 5 1 1 22631
0 22633 7 1 2 70296 83114
0 22634 7 1 2 90278 22633
0 22635 5 1 1 22634
0 22636 7 1 2 22632 22635
0 22637 5 1 1 22636
0 22638 7 1 2 90267 22637
0 22639 5 1 1 22638
0 22640 7 5 2 63488 64305
0 22641 7 5 2 60124 66218
0 22642 7 1 2 62695 90305
0 22643 7 1 2 90300 22642
0 22644 7 4 2 58860 59806
0 22645 7 3 2 58510 90310
0 22646 7 1 2 88860 90314
0 22647 7 1 2 22643 22646
0 22648 5 1 1 22647
0 22649 7 2 2 90127 90226
0 22650 7 8 2 64525 82802
0 22651 5 1 1 90319
0 22652 7 1 2 73422 74415
0 22653 7 1 2 90320 22652
0 22654 7 1 2 90317 22653
0 22655 5 1 1 22654
0 22656 7 1 2 22648 22655
0 22657 5 1 1 22656
0 22658 7 1 2 90223 22657
0 22659 5 1 1 22658
0 22660 7 1 2 64876 22659
0 22661 7 1 2 22639 22660
0 22662 7 1 2 22613 22661
0 22663 7 1 2 22534 22662
0 22664 7 1 2 22332 22663
0 22665 7 1 2 22219 22664
0 22666 5 1 1 22665
0 22667 7 1 2 63682 22666
0 22668 7 1 2 21758 22667
0 22669 5 1 1 22668
0 22670 7 2 2 86119 82380
0 22671 5 1 1 90327
0 22672 7 1 2 59363 79787
0 22673 5 1 1 22672
0 22674 7 1 2 70714 22673
0 22675 5 1 1 22674
0 22676 7 1 2 90328 22675
0 22677 5 1 1 22676
0 22678 7 3 2 62403 66219
0 22679 7 1 2 89543 90329
0 22680 5 1 1 22679
0 22681 7 1 2 22677 22680
0 22682 5 1 1 22681
0 22683 7 1 2 64877 89310
0 22684 7 1 2 22682 22683
0 22685 5 1 1 22684
0 22686 7 4 2 67747 76195
0 22687 5 2 1 90332
0 22688 7 2 2 78480 88239
0 22689 7 2 2 64306 60183
0 22690 7 3 2 88718 90340
0 22691 7 1 2 90338 90342
0 22692 7 1 2 90333 22691
0 22693 5 1 1 22692
0 22694 7 1 2 22685 22693
0 22695 5 1 1 22694
0 22696 7 1 2 58511 22695
0 22697 5 1 1 22696
0 22698 7 10 2 65266 61603
0 22699 7 3 2 65039 90345
0 22700 5 2 1 90355
0 22701 7 2 2 63253 84174
0 22702 5 2 1 90360
0 22703 7 1 2 90358 90362
0 22704 5 1 1 22703
0 22705 7 1 2 68233 22704
0 22706 5 1 1 22705
0 22707 7 1 2 81191 87188
0 22708 7 1 2 75836 22707
0 22709 5 1 1 22708
0 22710 7 1 2 22706 22709
0 22711 5 1 1 22710
0 22712 7 1 2 61280 22711
0 22713 5 1 1 22712
0 22714 7 1 2 86468 77902
0 22715 5 1 1 22714
0 22716 7 1 2 22713 22715
0 22717 5 1 1 22716
0 22718 7 1 2 60916 22717
0 22719 5 1 1 22718
0 22720 7 2 2 13568 86736
0 22721 5 4 1 90364
0 22722 7 1 2 61604 90366
0 22723 5 1 1 22722
0 22724 7 1 2 22719 22723
0 22725 5 2 1 22724
0 22726 7 1 2 62960 90370
0 22727 5 1 1 22726
0 22728 7 4 2 62404 77896
0 22729 5 4 1 90372
0 22730 7 2 2 74337 84794
0 22731 7 1 2 90373 90380
0 22732 5 1 1 22731
0 22733 7 1 2 22727 22732
0 22734 5 1 1 22733
0 22735 7 1 2 67190 22734
0 22736 5 1 1 22735
0 22737 7 4 2 68234 71405
0 22738 7 1 2 90381 90382
0 22739 5 1 1 22738
0 22740 7 1 2 22736 22739
0 22741 5 1 1 22740
0 22742 7 1 2 60184 88719
0 22743 7 1 2 22741 22742
0 22744 5 1 1 22743
0 22745 7 1 2 22697 22744
0 22746 5 1 1 22745
0 22747 7 1 2 59807 22746
0 22748 5 1 1 22747
0 22749 7 5 2 60185 61936
0 22750 7 1 2 77013 3632
0 22751 5 1 1 22750
0 22752 7 1 2 89801 22751
0 22753 5 1 1 22752
0 22754 7 1 2 81837 82873
0 22755 5 1 1 22754
0 22756 7 1 2 22753 22755
0 22757 5 1 1 22756
0 22758 7 1 2 60917 22757
0 22759 5 1 1 22758
0 22760 7 2 2 72797 84175
0 22761 5 1 1 90391
0 22762 7 1 2 22759 22761
0 22763 5 1 1 22762
0 22764 7 1 2 65912 22763
0 22765 5 1 1 22764
0 22766 7 1 2 85108 87332
0 22767 5 1 1 22766
0 22768 7 1 2 22765 22767
0 22769 5 1 1 22768
0 22770 7 1 2 61804 22769
0 22771 5 1 1 22770
0 22772 7 2 2 79488 90025
0 22773 5 1 1 90393
0 22774 7 1 2 63254 77950
0 22775 7 1 2 90394 22774
0 22776 5 1 1 22775
0 22777 7 1 2 22771 22776
0 22778 5 1 1 22777
0 22779 7 1 2 76196 22778
0 22780 5 1 1 22779
0 22781 7 1 2 69788 85444
0 22782 5 1 1 22781
0 22783 7 1 2 21627 22782
0 22784 5 1 1 22783
0 22785 7 1 2 60918 22784
0 22786 5 1 1 22785
0 22787 7 1 2 60349 85396
0 22788 5 1 1 22787
0 22789 7 1 2 22786 22788
0 22790 5 1 1 22789
0 22791 7 1 2 66220 22790
0 22792 5 1 1 22791
0 22793 7 1 2 89795 22792
0 22794 5 1 1 22793
0 22795 7 1 2 84984 22794
0 22796 5 1 1 22795
0 22797 7 2 2 77425 82874
0 22798 7 1 2 86132 90395
0 22799 5 1 1 22798
0 22800 7 1 2 22796 22799
0 22801 5 1 1 22800
0 22802 7 1 2 61805 22801
0 22803 5 1 1 22802
0 22804 7 1 2 86539 70985
0 22805 5 1 1 22804
0 22806 7 1 2 84567 22805
0 22807 5 1 1 22806
0 22808 7 1 2 64307 22807
0 22809 5 1 1 22808
0 22810 7 1 2 70736 79360
0 22811 5 1 1 22810
0 22812 7 1 2 22809 22811
0 22813 5 1 1 22812
0 22814 7 1 2 61281 22813
0 22815 5 1 1 22814
0 22816 7 1 2 84032 84410
0 22817 5 2 1 22816
0 22818 7 1 2 22815 90397
0 22819 5 1 1 22818
0 22820 7 1 2 80806 89644
0 22821 7 1 2 22819 22820
0 22822 5 1 1 22821
0 22823 7 2 2 22803 22822
0 22824 5 1 1 90399
0 22825 7 1 2 22780 90400
0 22826 5 1 1 22825
0 22827 7 1 2 64526 22826
0 22828 5 1 1 22827
0 22829 7 3 2 67191 80760
0 22830 7 1 2 89799 90401
0 22831 5 1 1 22830
0 22832 7 1 2 22828 22831
0 22833 5 1 1 22832
0 22834 7 1 2 90386 22833
0 22835 5 1 1 22834
0 22836 7 1 2 22748 22835
0 22837 5 1 1 22836
0 22838 7 1 2 63683 22837
0 22839 5 1 1 22838
0 22840 7 1 2 77007 89721
0 22841 5 1 1 22840
0 22842 7 1 2 87314 73525
0 22843 5 7 1 22842
0 22844 7 1 2 75075 90404
0 22845 5 1 1 22844
0 22846 7 1 2 22841 22845
0 22847 5 1 1 22846
0 22848 7 1 2 62405 22847
0 22849 5 1 1 22848
0 22850 7 1 2 75440 78481
0 22851 7 1 2 86640 22850
0 22852 5 1 1 22851
0 22853 7 1 2 22849 22852
0 22854 5 1 1 22853
0 22855 7 1 2 61605 22854
0 22856 5 1 1 22855
0 22857 7 1 2 86120 81467
0 22858 7 1 2 89431 22857
0 22859 5 1 1 22858
0 22860 7 1 2 22856 22859
0 22861 5 1 1 22860
0 22862 7 1 2 60919 22861
0 22863 5 1 1 22862
0 22864 7 3 2 60350 85723
0 22865 7 1 2 88551 90411
0 22866 5 1 1 22865
0 22867 7 1 2 22863 22866
0 22868 5 1 1 22867
0 22869 7 1 2 61806 22868
0 22870 5 1 1 22869
0 22871 7 1 2 86600 89807
0 22872 7 1 2 90170 22871
0 22873 5 1 1 22872
0 22874 7 1 2 22870 22873
0 22875 5 1 1 22874
0 22876 7 1 2 76197 22875
0 22877 5 1 1 22876
0 22878 7 1 2 64527 22824
0 22879 5 1 1 22878
0 22880 7 1 2 59808 90371
0 22881 5 1 1 22880
0 22882 7 1 2 85513 90392
0 22883 5 1 1 22882
0 22884 7 1 2 22881 22883
0 22885 5 1 1 22884
0 22886 7 1 2 61807 80867
0 22887 7 1 2 22885 22886
0 22888 5 1 1 22887
0 22889 7 1 2 22879 22888
0 22890 7 1 2 22877 22889
0 22891 5 1 1 22890
0 22892 7 1 2 61937 88387
0 22893 7 1 2 22891 22892
0 22894 5 1 1 22893
0 22895 7 1 2 22839 22894
0 22896 5 1 1 22895
0 22897 7 1 2 62080 22896
0 22898 5 1 1 22897
0 22899 7 3 2 67523 88123
0 22900 7 1 2 71782 79414
0 22901 5 1 1 22900
0 22902 7 1 2 89945 22901
0 22903 5 1 1 22902
0 22904 7 1 2 60351 22903
0 22905 5 1 1 22904
0 22906 7 1 2 87419 74956
0 22907 5 1 1 22906
0 22908 7 1 2 22905 22907
0 22909 5 1 1 22908
0 22910 7 1 2 88552 22909
0 22911 5 1 1 22910
0 22912 7 2 2 78578 82553
0 22913 5 1 1 90417
0 22914 7 3 2 62961 85624
0 22915 7 1 2 90418 90419
0 22916 7 1 2 89615 22915
0 22917 5 1 1 22916
0 22918 7 1 2 22911 22917
0 22919 5 1 1 22918
0 22920 7 1 2 61282 22919
0 22921 5 1 1 22920
0 22922 7 6 2 65913 75519
0 22923 7 2 2 71177 82682
0 22924 5 2 1 90428
0 22925 7 1 2 60566 90429
0 22926 5 1 1 22925
0 22927 7 1 2 75902 84127
0 22928 5 1 1 22927
0 22929 7 1 2 22926 22928
0 22930 5 1 1 22929
0 22931 7 1 2 65586 22930
0 22932 5 1 1 22931
0 22933 7 2 2 86934 81517
0 22934 5 1 1 90432
0 22935 7 1 2 69924 89564
0 22936 5 1 1 22935
0 22937 7 1 2 22934 22936
0 22938 5 1 1 22937
0 22939 7 1 2 62406 22938
0 22940 5 1 1 22939
0 22941 7 1 2 63888 90433
0 22942 5 1 1 22941
0 22943 7 2 2 71406 81396
0 22944 5 2 1 90434
0 22945 7 1 2 22942 90436
0 22946 7 1 2 22940 22945
0 22947 5 1 1 22946
0 22948 7 1 2 65267 22947
0 22949 5 1 1 22948
0 22950 7 1 2 22932 22949
0 22951 5 1 1 22950
0 22952 7 1 2 90422 22951
0 22953 5 1 1 22952
0 22954 7 1 2 22921 22953
0 22955 5 1 1 22954
0 22956 7 1 2 62696 22955
0 22957 5 1 1 22956
0 22958 7 1 2 81333 81654
0 22959 5 2 1 22958
0 22960 7 1 2 90430 90438
0 22961 5 1 1 22960
0 22962 7 1 2 62407 22961
0 22963 5 1 1 22962
0 22964 7 1 2 69789 84056
0 22965 5 1 1 22964
0 22966 7 1 2 22963 22965
0 22967 5 1 1 22966
0 22968 7 1 2 83456 22967
0 22969 5 1 1 22968
0 22970 7 5 2 62408 58287
0 22971 7 2 2 69391 90440
0 22972 7 1 2 90270 90445
0 22973 5 1 1 22972
0 22974 7 1 2 22969 22973
0 22975 5 1 1 22974
0 22976 7 1 2 65914 22975
0 22977 5 1 1 22976
0 22978 7 1 2 63889 90446
0 22979 7 1 2 90123 22978
0 22980 5 1 1 22979
0 22981 7 1 2 22977 22980
0 22982 5 1 1 22981
0 22983 7 1 2 75520 22982
0 22984 5 1 1 22983
0 22985 7 1 2 22957 22984
0 22986 5 1 1 22985
0 22987 7 1 2 61808 22986
0 22988 5 1 1 22987
0 22989 7 1 2 79290 90026
0 22990 7 1 2 90049 22989
0 22991 5 1 1 22990
0 22992 7 1 2 22988 22991
0 22993 5 1 1 22992
0 22994 7 1 2 90414 22993
0 22995 5 1 1 22994
0 22996 7 1 2 22898 22995
0 22997 5 1 1 22996
0 22998 7 1 2 70504 22997
0 22999 5 1 1 22998
0 23000 7 4 2 60920 66440
0 23001 7 2 2 86646 90447
0 23002 7 1 2 74437 90451
0 23003 5 1 1 23002
0 23004 7 3 2 80832 88694
0 23005 5 1 1 90453
0 23006 7 1 2 23003 23005
0 23007 5 1 1 23006
0 23008 7 1 2 62409 23007
0 23009 5 1 1 23008
0 23010 7 1 2 86546 89001
0 23011 5 2 1 23010
0 23012 7 1 2 84446 90173
0 23013 5 1 1 23012
0 23014 7 1 2 90456 23013
0 23015 5 1 1 23014
0 23016 7 1 2 62962 23015
0 23017 5 1 1 23016
0 23018 7 1 2 23009 23017
0 23019 5 1 1 23018
0 23020 7 1 2 67192 23019
0 23021 5 1 1 23020
0 23022 7 7 2 59809 87016
0 23023 7 1 2 83930 89217
0 23024 7 1 2 90458 23023
0 23025 5 1 1 23024
0 23026 7 1 2 23021 23025
0 23027 5 1 1 23026
0 23028 7 1 2 60567 23027
0 23029 5 1 1 23028
0 23030 7 1 2 65587 83933
0 23031 5 1 1 23030
0 23032 7 1 2 67193 90454
0 23033 7 1 2 23031 23032
0 23034 5 1 1 23033
0 23035 7 1 2 23029 23034
0 23036 5 1 1 23035
0 23037 7 1 2 89114 23036
0 23038 5 1 1 23037
0 23039 7 1 2 70689 88908
0 23040 7 1 2 85263 23039
0 23041 5 1 1 23040
0 23042 7 1 2 89175 90457
0 23043 5 3 1 23042
0 23044 7 1 2 64046 89176
0 23045 5 1 1 23044
0 23046 7 1 2 60568 78801
0 23047 7 1 2 23045 23046
0 23048 7 1 2 90465 23047
0 23049 5 1 1 23048
0 23050 7 1 2 23041 23049
0 23051 5 1 1 23050
0 23052 7 1 2 88350 23051
0 23053 5 1 1 23052
0 23054 7 1 2 89115 90466
0 23055 5 1 1 23054
0 23056 7 1 2 23053 23055
0 23057 5 1 1 23056
0 23058 7 1 2 62963 23057
0 23059 5 1 1 23058
0 23060 7 1 2 67194 90467
0 23061 5 1 1 23060
0 23062 7 1 2 68706 90452
0 23063 5 1 1 23062
0 23064 7 1 2 23061 23063
0 23065 5 1 1 23064
0 23066 7 1 2 89116 23065
0 23067 5 1 1 23066
0 23068 7 1 2 23059 23067
0 23069 5 1 1 23068
0 23070 7 1 2 60352 23069
0 23071 5 1 1 23070
0 23072 7 3 2 61809 77210
0 23073 7 3 2 75521 90468
0 23074 5 1 1 90471
0 23075 7 2 2 89117 90472
0 23076 5 1 1 90474
0 23077 7 1 2 62964 90475
0 23078 5 1 1 23077
0 23079 7 2 2 87017 67524
0 23080 7 1 2 73376 89022
0 23081 7 1 2 90476 23080
0 23082 5 1 1 23081
0 23083 7 1 2 23076 23082
0 23084 5 1 1 23083
0 23085 7 1 2 62697 23084
0 23086 5 1 1 23085
0 23087 7 2 2 88994 89290
0 23088 7 1 2 77031 90478
0 23089 5 1 1 23088
0 23090 7 1 2 23086 23089
0 23091 5 1 1 23090
0 23092 7 1 2 64047 23091
0 23093 5 1 1 23092
0 23094 7 1 2 23078 23093
0 23095 7 1 2 23071 23094
0 23096 5 1 1 23095
0 23097 7 1 2 62410 23096
0 23098 5 1 1 23097
0 23099 7 1 2 59364 72769
0 23100 5 1 1 23099
0 23101 7 1 2 90479 23100
0 23102 5 1 1 23101
0 23103 7 1 2 73172 89159
0 23104 7 1 2 90174 23103
0 23105 7 1 2 90477 23104
0 23106 5 1 1 23105
0 23107 7 1 2 23102 23106
0 23108 5 1 1 23107
0 23109 7 1 2 62698 23108
0 23110 5 1 1 23109
0 23111 7 4 2 61810 88990
0 23112 7 1 2 80807 67471
0 23113 7 1 2 90480 23112
0 23114 5 1 1 23113
0 23115 7 1 2 23110 23114
0 23116 5 1 1 23115
0 23117 7 1 2 72090 23116
0 23118 5 1 1 23117
0 23119 7 1 2 23098 23118
0 23120 5 1 1 23119
0 23121 7 1 2 64308 23120
0 23122 5 1 1 23121
0 23123 7 1 2 23038 23122
0 23124 5 1 1 23123
0 23125 7 1 2 65915 23124
0 23126 5 1 1 23125
0 23127 7 1 2 89432 88832
0 23128 5 1 1 23127
0 23129 7 1 2 89177 23128
0 23130 5 1 1 23129
0 23131 7 1 2 85691 23130
0 23132 5 1 1 23131
0 23133 7 1 2 74096 88695
0 23134 7 1 2 87252 23133
0 23135 5 1 1 23134
0 23136 7 1 2 23132 23135
0 23137 5 1 1 23136
0 23138 7 1 2 62411 23137
0 23139 5 1 1 23138
0 23140 7 1 2 74017 77608
0 23141 7 1 2 89002 23140
0 23142 5 1 1 23141
0 23143 7 1 2 23139 23142
0 23144 5 1 1 23143
0 23145 7 1 2 86209 89118
0 23146 7 1 2 23144 23145
0 23147 5 1 1 23146
0 23148 7 1 2 23126 23147
0 23149 5 1 1 23148
0 23150 7 1 2 66221 23149
0 23151 5 1 1 23150
0 23152 7 2 2 84659 89928
0 23153 5 1 1 90484
0 23154 7 1 2 86469 74599
0 23155 7 1 2 83854 23154
0 23156 5 1 1 23155
0 23157 7 1 2 23153 23156
0 23158 5 1 1 23157
0 23159 7 1 2 67195 23158
0 23160 5 1 1 23159
0 23161 7 2 2 62965 84660
0 23162 5 3 1 90486
0 23163 7 1 2 70170 86470
0 23164 5 2 1 23163
0 23165 7 1 2 90488 90491
0 23166 5 1 1 23165
0 23167 7 1 2 60569 23166
0 23168 5 1 1 23167
0 23169 7 3 2 61606 73310
0 23170 7 1 2 75076 90493
0 23171 5 1 1 23170
0 23172 7 1 2 23168 23171
0 23173 5 1 1 23172
0 23174 7 1 2 63255 23173
0 23175 5 1 1 23174
0 23176 7 1 2 23160 23175
0 23177 5 1 1 23176
0 23178 7 1 2 89119 23177
0 23179 5 1 1 23178
0 23180 7 1 2 81838 87198
0 23181 5 1 1 23180
0 23182 7 1 2 89766 23181
0 23183 5 1 1 23182
0 23184 7 1 2 64048 23183
0 23185 5 1 1 23184
0 23186 7 1 2 73256 81356
0 23187 5 1 1 23186
0 23188 7 1 2 23185 23187
0 23189 5 1 1 23188
0 23190 7 1 2 62699 23189
0 23191 5 1 1 23190
0 23192 7 1 2 78550 71607
0 23193 7 1 2 86471 23192
0 23194 5 1 1 23193
0 23195 7 1 2 23191 23194
0 23196 5 1 1 23195
0 23197 7 1 2 77782 88351
0 23198 7 1 2 23196 23197
0 23199 5 1 1 23198
0 23200 7 1 2 23179 23199
0 23201 5 1 1 23200
0 23202 7 1 2 64528 23201
0 23203 5 1 1 23202
0 23204 7 2 2 59810 60186
0 23205 7 1 2 61283 82181
0 23206 7 1 2 90496 23205
0 23207 7 2 2 70297 75396
0 23208 7 1 2 81663 90498
0 23209 7 1 2 23206 23208
0 23210 5 1 1 23209
0 23211 7 1 2 23203 23210
0 23212 5 1 1 23211
0 23213 7 1 2 62412 23212
0 23214 5 1 1 23213
0 23215 7 1 2 76198 90119
0 23216 5 1 1 23215
0 23217 7 1 2 21457 23216
0 23218 5 1 1 23217
0 23219 7 2 2 75522 89120
0 23220 7 1 2 23218 90500
0 23221 5 1 1 23220
0 23222 7 1 2 23214 23221
0 23223 5 1 1 23222
0 23224 7 1 2 88696 23223
0 23225 5 1 1 23224
0 23226 7 6 2 64049 60187
0 23227 7 2 2 83022 90502
0 23228 7 1 2 79998 83202
0 23229 7 1 2 90508 23228
0 23230 5 1 1 23229
0 23231 7 2 2 60570 88352
0 23232 7 1 2 58512 72285
0 23233 7 1 2 81429 23232
0 23234 7 1 2 90510 23233
0 23235 5 1 1 23234
0 23236 7 1 2 23230 23235
0 23237 5 1 1 23236
0 23238 7 1 2 67748 23237
0 23239 5 1 1 23238
0 23240 7 2 2 87900 76869
0 23241 7 1 2 70655 90512
0 23242 5 1 1 23241
0 23243 7 3 2 65040 89121
0 23244 5 1 1 90514
0 23245 7 1 2 23242 23244
0 23246 5 1 1 23245
0 23247 7 1 2 62413 23246
0 23248 5 1 1 23247
0 23249 7 1 2 81676 90513
0 23250 5 1 1 23249
0 23251 7 1 2 23248 23250
0 23252 5 1 1 23251
0 23253 7 1 2 90101 23252
0 23254 5 1 1 23253
0 23255 7 1 2 23239 23254
0 23256 5 1 1 23255
0 23257 7 1 2 65916 23256
0 23258 5 1 1 23257
0 23259 7 2 2 58288 88353
0 23260 7 2 2 74983 81468
0 23261 7 1 2 70737 90519
0 23262 5 1 1 23261
0 23263 7 1 2 82001 81357
0 23264 5 1 1 23263
0 23265 7 1 2 23262 23264
0 23266 5 1 1 23265
0 23267 7 1 2 90517 23266
0 23268 5 1 1 23267
0 23269 7 4 2 62414 89122
0 23270 7 1 2 71819 81397
0 23271 7 1 2 90521 23270
0 23272 5 1 1 23271
0 23273 7 1 2 23268 23272
0 23274 5 1 1 23273
0 23275 7 1 2 80559 23274
0 23276 5 1 1 23275
0 23277 7 1 2 23258 23276
0 23278 5 1 1 23277
0 23279 7 1 2 59811 88909
0 23280 7 1 2 23278 23279
0 23281 5 1 1 23280
0 23282 7 1 2 23225 23281
0 23283 5 1 1 23282
0 23284 7 1 2 59565 23283
0 23285 5 1 1 23284
0 23286 7 4 2 60188 60353
0 23287 7 1 2 76591 90525
0 23288 5 1 1 23287
0 23289 7 3 2 60571 72311
0 23290 7 1 2 64878 86284
0 23291 7 1 2 90529 23290
0 23292 5 1 1 23291
0 23293 7 1 2 23288 23292
0 23294 5 1 1 23293
0 23295 7 1 2 62415 23294
0 23296 5 1 1 23295
0 23297 7 3 2 62081 90526
0 23298 5 1 1 90532
0 23299 7 1 2 87131 90533
0 23300 5 1 1 23299
0 23301 7 1 2 23296 23300
0 23302 5 1 1 23301
0 23303 7 1 2 89224 23302
0 23304 5 1 1 23303
0 23305 7 1 2 72091 89123
0 23306 5 1 1 23305
0 23307 7 3 2 62416 64879
0 23308 7 4 2 66697 90535
0 23309 7 1 2 72764 90538
0 23310 5 1 1 23309
0 23311 7 1 2 23306 23310
0 23312 5 1 1 23311
0 23313 7 1 2 90268 23312
0 23314 5 1 1 23313
0 23315 7 1 2 23304 23314
0 23316 5 1 1 23315
0 23317 7 1 2 61284 23316
0 23318 5 1 1 23317
0 23319 7 9 2 65917 62082
0 23320 7 2 2 60572 90542
0 23321 7 4 2 62417 77032
0 23322 5 6 1 90553
0 23323 7 1 2 89225 90527
0 23324 7 1 2 90554 23323
0 23325 7 1 2 90551 23324
0 23326 5 1 1 23325
0 23327 7 1 2 23318 23326
0 23328 5 1 1 23327
0 23329 7 1 2 64309 23328
0 23330 5 1 1 23329
0 23331 7 3 2 61811 84452
0 23332 7 2 2 62083 90563
0 23333 7 3 2 60189 65918
0 23334 7 1 2 86641 90568
0 23335 7 1 2 90566 23334
0 23336 5 1 1 23335
0 23337 7 1 2 23330 23336
0 23338 5 1 1 23337
0 23339 7 1 2 62966 23338
0 23340 5 1 1 23339
0 23341 7 1 2 79379 88475
0 23342 7 2 2 64310 88855
0 23343 7 5 2 61285 68235
0 23344 7 1 2 90571 90573
0 23345 7 1 2 23341 23344
0 23346 5 1 1 23345
0 23347 7 1 2 23340 23346
0 23348 5 1 1 23347
0 23349 7 1 2 67196 23348
0 23350 5 1 1 23349
0 23351 7 2 2 62418 87018
0 23352 7 3 2 63890 60190
0 23353 7 1 2 90572 90580
0 23354 7 1 2 90578 23353
0 23355 7 1 2 85598 23354
0 23356 5 1 1 23355
0 23357 7 1 2 23350 23356
0 23358 5 1 1 23357
0 23359 7 1 2 82097 23358
0 23360 5 1 1 23359
0 23361 7 1 2 23285 23360
0 23362 7 1 2 23151 23361
0 23363 5 1 1 23362
0 23364 7 1 2 63684 23363
0 23365 5 1 1 23364
0 23366 7 1 2 77358 80544
0 23367 5 2 1 23366
0 23368 7 1 2 85600 90583
0 23369 5 1 1 23368
0 23370 7 1 2 59566 23369
0 23371 5 1 1 23370
0 23372 7 6 2 70298 79489
0 23373 5 1 1 90585
0 23374 7 1 2 58513 23373
0 23375 5 1 1 23374
0 23376 7 1 2 87495 23375
0 23377 5 1 1 23376
0 23378 7 1 2 23371 23377
0 23379 5 1 1 23378
0 23380 7 1 2 61607 23379
0 23381 5 1 1 23380
0 23382 7 10 2 66222 76673
0 23383 7 1 2 82002 72861
0 23384 5 1 1 23383
0 23385 7 1 2 60354 90423
0 23386 5 1 1 23385
0 23387 7 1 2 23384 23386
0 23388 5 1 1 23387
0 23389 7 1 2 90591 23388
0 23390 5 1 1 23389
0 23391 7 1 2 23381 23390
0 23392 5 1 1 23391
0 23393 7 1 2 77426 23392
0 23394 5 1 1 23393
0 23395 7 3 2 63256 79162
0 23396 7 3 2 60921 86558
0 23397 7 1 2 90601 90604
0 23398 5 1 1 23397
0 23399 7 1 2 23394 23398
0 23400 5 1 1 23399
0 23401 7 1 2 64050 23400
0 23402 5 1 1 23401
0 23403 7 1 2 86968 79329
0 23404 5 1 1 23403
0 23405 7 1 2 86353 89792
0 23406 5 2 1 23405
0 23407 7 1 2 88553 90607
0 23408 5 1 1 23407
0 23409 7 1 2 23404 23408
0 23410 5 1 1 23409
0 23411 7 1 2 76199 23410
0 23412 5 1 1 23411
0 23413 7 1 2 75523 86236
0 23414 7 1 2 86710 23413
0 23415 5 1 1 23414
0 23416 7 1 2 23412 23415
0 23417 7 1 2 23402 23416
0 23418 5 1 1 23417
0 23419 7 1 2 88697 23418
0 23420 5 1 1 23419
0 23421 7 1 2 60355 85942
0 23422 5 1 1 23421
0 23423 7 1 2 73068 23422
0 23424 5 1 1 23423
0 23425 7 4 2 59812 70299
0 23426 5 1 1 90609
0 23427 7 1 2 58514 89605
0 23428 7 1 2 90610 23427
0 23429 7 1 2 23424 23428
0 23430 5 1 1 23429
0 23431 7 1 2 23420 23430
0 23432 5 1 1 23431
0 23433 7 1 2 63891 23432
0 23434 5 1 1 23433
0 23435 7 1 2 86213 89793
0 23436 5 2 1 23435
0 23437 7 1 2 76200 90613
0 23438 5 1 1 23437
0 23439 7 1 2 89513 23438
0 23440 5 1 1 23439
0 23441 7 1 2 66223 23440
0 23442 5 1 1 23441
0 23443 7 1 2 89520 23442
0 23444 5 1 1 23443
0 23445 7 1 2 89172 23444
0 23446 5 1 1 23445
0 23447 7 1 2 23434 23446
0 23448 5 1 1 23447
0 23449 7 1 2 62419 23448
0 23450 5 1 1 23449
0 23451 7 5 2 61608 88698
0 23452 7 1 2 72862 90615
0 23453 5 2 1 23452
0 23454 7 4 2 86559 88910
0 23455 5 1 1 90622
0 23456 7 1 2 90620 23455
0 23457 5 2 1 23456
0 23458 7 1 2 76637 90626
0 23459 5 1 1 23458
0 23460 7 5 2 64311 66441
0 23461 7 6 2 61286 82098
0 23462 7 2 2 90628 90633
0 23463 7 1 2 89433 90639
0 23464 5 1 1 23463
0 23465 7 1 2 23459 23464
0 23466 5 1 1 23465
0 23467 7 1 2 60573 23466
0 23468 5 1 1 23467
0 23469 7 1 2 78391 90640
0 23470 5 1 1 23469
0 23471 7 1 2 23468 23470
0 23472 5 1 1 23471
0 23473 7 1 2 60356 23472
0 23474 5 1 1 23473
0 23475 7 2 2 78392 88699
0 23476 7 1 2 86560 90641
0 23477 5 1 1 23476
0 23478 7 1 2 23474 23477
0 23479 5 1 1 23478
0 23480 7 1 2 62967 23479
0 23481 5 1 1 23480
0 23482 7 2 2 66588 73086
0 23483 7 1 2 81398 88970
0 23484 7 1 2 90643 23483
0 23485 5 1 1 23484
0 23486 7 1 2 23481 23485
0 23487 5 1 1 23486
0 23488 7 1 2 64051 23487
0 23489 5 1 1 23488
0 23490 7 1 2 80836 89601
0 23491 7 1 2 90224 23490
0 23492 5 1 1 23491
0 23493 7 1 2 23489 23492
0 23494 5 1 1 23493
0 23495 7 1 2 62700 23494
0 23496 5 1 1 23495
0 23497 7 1 2 70171 86695
0 23498 5 2 1 23497
0 23499 7 1 2 84405 90645
0 23500 5 1 1 23499
0 23501 7 1 2 90473 23500
0 23502 5 1 1 23501
0 23503 7 1 2 65588 86935
0 23504 7 1 2 69164 89424
0 23505 7 1 2 23503 23504
0 23506 5 1 1 23505
0 23507 7 1 2 23074 23506
0 23508 5 1 1 23507
0 23509 7 1 2 62968 23508
0 23510 5 1 1 23509
0 23511 7 1 2 80837 90469
0 23512 5 1 1 23511
0 23513 7 1 2 23510 23512
0 23514 5 1 1 23513
0 23515 7 1 2 65919 23514
0 23516 5 1 1 23515
0 23517 7 3 2 61287 73717
0 23518 5 2 1 90647
0 23519 7 1 2 63257 90470
0 23520 7 1 2 90648 23519
0 23521 5 1 1 23520
0 23522 7 1 2 23516 23521
0 23523 5 1 1 23522
0 23524 7 1 2 66224 23523
0 23525 5 1 1 23524
0 23526 7 3 2 72863 86577
0 23527 5 1 1 90652
0 23528 7 1 2 80468 90653
0 23529 7 1 2 90616 23528
0 23530 5 1 1 23529
0 23531 7 1 2 23525 23530
0 23532 5 1 1 23531
0 23533 7 1 2 67197 23532
0 23534 5 1 1 23533
0 23535 7 1 2 23502 23534
0 23536 5 1 1 23535
0 23537 7 1 2 67749 23536
0 23538 5 1 1 23537
0 23539 7 2 2 74154 83180
0 23540 5 1 1 90655
0 23541 7 1 2 84406 23540
0 23542 5 1 1 23541
0 23543 7 1 2 90642 23542
0 23544 5 1 1 23543
0 23545 7 1 2 23538 23544
0 23546 7 1 2 23496 23545
0 23547 7 1 2 23450 23546
0 23548 5 2 1 23547
0 23549 7 1 2 89097 90657
0 23550 5 1 1 23549
0 23551 7 1 2 23365 23550
0 23552 5 1 1 23551
0 23553 7 1 2 69537 23552
0 23554 5 1 1 23553
0 23555 7 4 2 61609 85692
0 23556 7 2 2 89843 90659
0 23557 7 3 2 60191 61288
0 23558 7 1 2 90663 90665
0 23559 5 1 1 23558
0 23560 7 8 2 61812 66698
0 23561 7 3 2 81113 90668
0 23562 7 2 2 90053 90676
0 23563 7 1 2 75397 90679
0 23564 5 1 1 23563
0 23565 7 2 2 67472 89895
0 23566 7 1 2 59365 85775
0 23567 7 1 2 90681 23566
0 23568 5 2 1 23567
0 23569 7 1 2 23564 90683
0 23570 5 1 1 23569
0 23571 7 1 2 71820 23570
0 23572 5 1 1 23571
0 23573 7 7 2 61813 67525
0 23574 7 2 2 62969 90685
0 23575 7 2 2 82683 90692
0 23576 7 1 2 61289 90694
0 23577 5 1 1 23576
0 23578 7 1 2 90684 23577
0 23579 5 1 1 23578
0 23580 7 1 2 62701 23579
0 23581 5 1 1 23580
0 23582 7 1 2 23572 23581
0 23583 5 1 1 23582
0 23584 7 1 2 59567 23583
0 23585 5 1 1 23584
0 23586 7 2 2 86472 81655
0 23587 7 1 2 68707 90669
0 23588 7 1 2 90696 23587
0 23589 7 1 2 84397 23588
0 23590 5 1 1 23589
0 23591 7 1 2 23585 23590
0 23592 5 1 1 23591
0 23593 7 1 2 62420 23592
0 23594 5 1 1 23593
0 23595 7 2 2 66442 67473
0 23596 7 4 2 86561 90698
0 23597 7 1 2 80892 90700
0 23598 5 1 1 23597
0 23599 7 5 2 88396 90210
0 23600 7 1 2 84190 90160
0 23601 7 1 2 90704 23600
0 23602 5 1 1 23601
0 23603 7 1 2 23598 23602
0 23604 5 1 1 23603
0 23605 7 1 2 58289 23604
0 23606 5 1 1 23605
0 23607 7 1 2 83911 90686
0 23608 7 1 2 90697 23607
0 23609 5 1 1 23608
0 23610 7 1 2 23606 23609
0 23611 7 1 2 23594 23610
0 23612 5 1 1 23611
0 23613 7 1 2 64880 23612
0 23614 5 1 1 23613
0 23615 7 1 2 23559 23614
0 23616 5 1 1 23615
0 23617 7 1 2 65589 23616
0 23618 5 1 1 23617
0 23619 7 1 2 82182 90569
0 23620 7 1 2 76201 23619
0 23621 5 1 1 23620
0 23622 7 2 2 78447 75481
0 23623 7 1 2 61290 75129
0 23624 7 3 2 64052 64881
0 23625 7 5 2 66225 66699
0 23626 7 1 2 90711 90714
0 23627 7 1 2 23623 23626
0 23628 7 1 2 90709 23627
0 23629 5 1 1 23628
0 23630 7 1 2 23621 23629
0 23631 5 1 1 23630
0 23632 7 1 2 61938 89671
0 23633 7 1 2 23631 23632
0 23634 5 1 1 23633
0 23635 7 1 2 23618 23634
0 23636 5 1 1 23635
0 23637 7 1 2 63685 23636
0 23638 5 1 1 23637
0 23639 7 1 2 76149 14140
0 23640 5 1 1 23639
0 23641 7 1 2 85724 89098
0 23642 7 1 2 89400 23641
0 23643 7 1 2 23640 23642
0 23644 5 1 1 23643
0 23645 7 1 2 23638 23644
0 23646 5 1 1 23645
0 23647 7 1 2 70505 23646
0 23648 5 1 1 23647
0 23649 7 4 2 66589 89878
0 23650 7 1 2 73594 89124
0 23651 5 1 1 23650
0 23652 7 8 2 62421 68085
0 23653 5 1 1 90723
0 23654 7 1 2 64312 88354
0 23655 7 1 2 72244 23654
0 23656 7 1 2 90724 23655
0 23657 5 1 1 23656
0 23658 7 1 2 23651 23657
0 23659 5 1 1 23658
0 23660 7 1 2 69538 23659
0 23661 5 1 1 23660
0 23662 7 1 2 68665 88746
0 23663 7 1 2 73595 23662
0 23664 5 1 1 23663
0 23665 7 1 2 23661 23664
0 23666 5 1 1 23665
0 23667 7 1 2 62970 23666
0 23668 5 1 1 23667
0 23669 7 2 2 62084 88754
0 23670 7 1 2 77910 90731
0 23671 5 1 1 23670
0 23672 7 1 2 23668 23671
0 23673 5 1 1 23672
0 23674 7 1 2 90719 23673
0 23675 5 1 1 23674
0 23676 7 1 2 73596 71783
0 23677 5 1 1 23676
0 23678 7 1 2 78525 84411
0 23679 5 1 1 23678
0 23680 7 1 2 23677 23679
0 23681 5 1 1 23680
0 23682 7 1 2 90695 23681
0 23683 5 1 1 23682
0 23684 7 1 2 62422 84953
0 23685 7 1 2 90682 23684
0 23686 5 1 1 23685
0 23687 7 1 2 23683 23686
0 23688 5 1 1 23687
0 23689 7 1 2 64882 23688
0 23690 5 1 1 23689
0 23691 7 1 2 60574 90581
0 23692 7 1 2 90664 23691
0 23693 5 1 1 23692
0 23694 7 1 2 23690 23693
0 23695 5 1 1 23694
0 23696 7 1 2 70506 23695
0 23697 5 1 1 23696
0 23698 7 1 2 87896 71060
0 23699 7 1 2 80645 23698
0 23700 7 1 2 90227 23699
0 23701 5 1 1 23700
0 23702 7 1 2 84277 84163
0 23703 7 1 2 88763 23702
0 23704 5 1 1 23703
0 23705 7 1 2 23701 23704
0 23706 5 1 1 23705
0 23707 7 1 2 77666 23706
0 23708 5 1 1 23707
0 23709 7 1 2 59568 83804
0 23710 5 1 1 23709
0 23711 7 1 2 63892 23710
0 23712 5 1 1 23711
0 23713 7 1 2 81162 23712
0 23714 5 1 1 23713
0 23715 7 2 2 82183 88700
0 23716 7 1 2 64053 90733
0 23717 7 1 2 88755 23716
0 23718 7 1 2 23714 23717
0 23719 5 1 1 23718
0 23720 7 1 2 23708 23719
0 23721 5 1 1 23720
0 23722 7 1 2 60357 23721
0 23723 5 1 1 23722
0 23724 7 1 2 23697 23723
0 23725 7 1 2 23675 23724
0 23726 5 1 1 23725
0 23727 7 1 2 65920 23726
0 23728 5 1 1 23727
0 23729 7 1 2 85004 88355
0 23730 5 1 1 23729
0 23731 7 1 2 60192 80006
0 23732 5 1 1 23731
0 23733 7 1 2 23730 23732
0 23734 5 1 1 23733
0 23735 7 1 2 59569 23734
0 23736 5 1 1 23735
0 23737 7 1 2 74454 90515
0 23738 5 1 1 23737
0 23739 7 1 2 23736 23738
0 23740 5 1 1 23739
0 23741 7 1 2 61610 23740
0 23742 5 1 1 23741
0 23743 7 1 2 66700 87901
0 23744 7 1 2 80868 23743
0 23745 5 1 1 23744
0 23746 7 1 2 76202 89125
0 23747 7 1 2 89467 23746
0 23748 5 1 1 23747
0 23749 7 1 2 23745 23748
0 23750 5 1 1 23749
0 23751 7 1 2 81334 23750
0 23752 5 1 1 23751
0 23753 7 1 2 23742 23752
0 23754 5 1 1 23753
0 23755 7 1 2 62423 23754
0 23756 5 1 1 23755
0 23757 7 1 2 66226 85475
0 23758 5 1 1 23757
0 23759 7 2 2 87189 23758
0 23760 7 1 2 80007 90582
0 23761 7 1 2 90735 23760
0 23762 5 1 1 23761
0 23763 7 1 2 23756 23762
0 23764 5 1 1 23763
0 23765 7 1 2 72744 23764
0 23766 5 1 1 23765
0 23767 7 4 2 59570 82684
0 23768 5 2 1 90737
0 23769 7 1 2 70948 90738
0 23770 5 1 1 23769
0 23771 7 1 2 76884 81335
0 23772 5 1 1 23771
0 23773 7 1 2 23770 23772
0 23774 5 2 1 23773
0 23775 7 1 2 90732 90743
0 23776 5 1 1 23775
0 23777 7 1 2 71407 84176
0 23778 5 2 1 23777
0 23779 7 1 2 82398 90745
0 23780 5 1 1 23779
0 23781 7 1 2 84602 90065
0 23782 7 1 2 90511 23781
0 23783 7 1 2 23780 23782
0 23784 5 1 1 23783
0 23785 7 1 2 23776 23784
0 23786 5 1 1 23785
0 23787 7 1 2 66590 23786
0 23788 5 1 1 23787
0 23789 7 1 2 23766 23788
0 23790 5 1 1 23789
0 23791 7 1 2 88397 23790
0 23792 5 1 1 23791
0 23793 7 1 2 23728 23792
0 23794 5 1 1 23793
0 23795 7 1 2 63686 23794
0 23796 5 1 1 23795
0 23797 7 1 2 86245 90736
0 23798 5 1 1 23797
0 23799 7 1 2 78553 90660
0 23800 5 1 1 23799
0 23801 7 1 2 23798 23800
0 23802 5 1 1 23801
0 23803 7 1 2 60575 23802
0 23804 5 1 1 23803
0 23805 7 1 2 87591 90359
0 23806 5 1 1 23805
0 23807 7 1 2 90574 23806
0 23808 5 1 1 23807
0 23809 7 1 2 23804 23808
0 23810 5 1 1 23809
0 23811 7 1 2 72745 23810
0 23812 5 1 1 23811
0 23813 7 1 2 61291 90744
0 23814 5 1 1 23813
0 23815 7 2 2 71275 77667
0 23816 5 1 1 90747
0 23817 7 4 2 70013 75130
0 23818 5 5 1 90749
0 23819 7 1 2 23816 90753
0 23820 5 1 1 23819
0 23821 7 1 2 60576 23820
0 23822 5 1 1 23821
0 23823 7 1 2 84833 67865
0 23824 5 1 1 23823
0 23825 7 1 2 23822 23824
0 23826 5 1 1 23825
0 23827 7 1 2 60358 23826
0 23828 5 1 1 23827
0 23829 7 1 2 84381 23828
0 23830 5 1 1 23829
0 23831 7 1 2 86473 23830
0 23832 5 1 1 23831
0 23833 7 1 2 23814 23832
0 23834 5 1 1 23833
0 23835 7 1 2 84223 23834
0 23836 5 1 1 23835
0 23837 7 1 2 23812 23836
0 23838 5 1 1 23837
0 23839 7 1 2 61814 89099
0 23840 7 1 2 23838 23839
0 23841 5 1 1 23840
0 23842 7 1 2 23796 23841
0 23843 5 1 1 23842
0 23844 7 1 2 60922 23843
0 23845 5 1 1 23844
0 23846 7 2 2 66591 88398
0 23847 7 1 2 80469 90661
0 23848 5 1 1 23847
0 23849 7 1 2 76885 82518
0 23850 5 1 1 23849
0 23851 7 1 2 23848 23850
0 23852 5 1 1 23851
0 23853 7 1 2 90758 23852
0 23854 5 1 1 23853
0 23855 7 1 2 73759 71995
0 23856 7 1 2 90623 23855
0 23857 5 1 1 23856
0 23858 7 1 2 23854 23857
0 23859 5 1 1 23858
0 23860 7 1 2 67750 23859
0 23861 5 1 1 23860
0 23862 7 1 2 65921 90374
0 23863 5 1 1 23862
0 23864 7 1 2 15467 23863
0 23865 5 1 1 23864
0 23866 7 1 2 67198 23865
0 23867 5 1 1 23866
0 23868 7 1 2 78448 86629
0 23869 5 1 1 23868
0 23870 7 1 2 23867 23869
0 23871 5 1 1 23870
0 23872 7 1 2 90720 23871
0 23873 5 1 1 23872
0 23874 7 2 2 73311 89606
0 23875 5 1 1 90760
0 23876 7 1 2 78526 69361
0 23877 7 1 2 90761 23876
0 23878 5 1 1 23877
0 23879 7 1 2 23873 23878
0 23880 7 1 2 23861 23879
0 23881 5 1 1 23880
0 23882 7 5 2 69337 89155
0 23883 5 1 1 90762
0 23884 7 1 2 69539 88592
0 23885 5 1 1 23884
0 23886 7 1 2 23883 23885
0 23887 5 1 1 23886
0 23888 7 1 2 23881 23887
0 23889 5 1 1 23888
0 23890 7 5 2 61939 89896
0 23891 7 2 2 71178 90767
0 23892 5 1 1 90772
0 23893 7 1 2 75102 90773
0 23894 5 1 1 23893
0 23895 7 1 2 81444 88701
0 23896 7 1 2 86015 23895
0 23897 5 1 1 23896
0 23898 7 1 2 23894 23897
0 23899 5 1 1 23898
0 23900 7 1 2 62424 23899
0 23901 5 1 1 23900
0 23902 7 2 2 84177 88911
0 23903 7 1 2 78527 79771
0 23904 7 1 2 90774 23903
0 23905 5 1 1 23904
0 23906 7 1 2 23901 23905
0 23907 5 1 1 23906
0 23908 7 1 2 65922 78802
0 23909 7 1 2 88513 23908
0 23910 7 1 2 23907 23909
0 23911 5 1 1 23910
0 23912 7 1 2 23889 23911
0 23913 7 1 2 23845 23912
0 23914 7 1 2 23648 23913
0 23915 5 1 1 23914
0 23916 7 1 2 76736 23915
0 23917 5 1 1 23916
0 23918 7 1 2 90658 90763
0 23919 5 1 1 23918
0 23920 7 1 2 23917 23919
0 23921 7 1 2 23554 23920
0 23922 7 1 2 22999 23921
0 23923 5 1 1 23922
0 23924 7 1 2 66902 23923
0 23925 5 1 1 23924
0 23926 7 1 2 22669 23925
0 23927 7 1 2 21756 23926
0 23928 5 1 1 23927
0 23929 7 1 2 68831 23928
0 23930 5 1 1 23929
0 23931 7 3 2 63258 89831
0 23932 5 1 1 90776
0 23933 7 1 2 88614 23932
0 23934 5 2 1 23933
0 23935 7 2 2 86896 90779
0 23936 5 1 1 90781
0 23937 7 1 2 84661 80971
0 23938 5 1 1 23937
0 23939 7 1 2 23936 23938
0 23940 5 1 1 23939
0 23941 7 1 2 60923 23940
0 23942 5 1 1 23941
0 23943 7 1 2 83683 85965
0 23944 5 1 1 23943
0 23945 7 3 2 65923 82919
0 23946 5 2 1 90783
0 23947 7 9 2 65590 85146
0 23948 5 1 1 90788
0 23949 7 1 2 65041 90789
0 23950 5 2 1 23949
0 23951 7 1 2 90786 90797
0 23952 5 1 1 23951
0 23953 7 1 2 64529 85782
0 23954 7 1 2 23952 23953
0 23955 5 1 1 23954
0 23956 7 1 2 23944 23955
0 23957 5 1 1 23956
0 23958 7 1 2 66227 23957
0 23959 5 1 1 23958
0 23960 7 1 2 65924 82947
0 23961 5 5 1 23960
0 23962 7 1 2 75452 78507
0 23963 5 7 1 23962
0 23964 7 4 2 60359 84240
0 23965 5 1 1 90811
0 23966 7 1 2 90804 90812
0 23967 5 1 1 23966
0 23968 7 1 2 61292 23967
0 23969 7 1 2 90798 23968
0 23970 5 1 1 23969
0 23971 7 1 2 90799 23970
0 23972 5 1 1 23971
0 23973 7 1 2 59813 23972
0 23974 5 1 1 23973
0 23975 7 1 2 73027 86214
0 23976 5 3 1 23975
0 23977 7 1 2 58515 90815
0 23978 5 1 1 23977
0 23979 7 3 2 65042 73312
0 23980 7 1 2 78499 90818
0 23981 5 1 1 23980
0 23982 7 1 2 64530 23981
0 23983 7 1 2 23978 23982
0 23984 5 1 1 23983
0 23985 7 1 2 61611 23984
0 23986 7 1 2 23974 23985
0 23987 5 1 1 23986
0 23988 7 1 2 23959 23987
0 23989 5 1 1 23988
0 23990 7 1 2 64054 23989
0 23991 5 1 1 23990
0 23992 7 1 2 23942 23991
0 23993 5 1 1 23992
0 23994 7 1 2 89100 23993
0 23995 5 1 1 23994
0 23996 7 1 2 77793 80968
0 23997 5 5 1 23996
0 23998 7 2 2 73116 84662
0 23999 5 4 1 90826
0 24000 7 1 2 89702 90828
0 24001 5 2 1 24000
0 24002 7 1 2 88356 90832
0 24003 7 1 2 90821 24002
0 24004 5 1 1 24003
0 24005 7 5 2 62085 90666
0 24006 7 3 2 85336 88240
0 24007 7 1 2 90805 90839
0 24008 7 1 2 90834 24007
0 24009 5 1 1 24008
0 24010 7 1 2 24004 24009
0 24011 5 2 1 24010
0 24012 7 1 2 62425 90842
0 24013 5 1 1 24012
0 24014 7 1 2 78183 78052
0 24015 5 4 1 24014
0 24016 7 5 2 62086 90570
0 24017 7 1 2 88554 90848
0 24018 7 1 2 90844 24017
0 24019 5 1 1 24018
0 24020 7 1 2 24013 24019
0 24021 5 1 1 24020
0 24022 7 1 2 60360 24021
0 24023 5 1 1 24022
0 24024 7 1 2 79840 69156
0 24025 7 1 2 90341 24024
0 24026 5 1 1 24025
0 24027 7 2 2 58516 86442
0 24028 5 4 1 90853
0 24029 7 2 2 63259 74146
0 24030 5 2 1 90859
0 24031 7 1 2 90539 90861
0 24032 7 1 2 90855 24031
0 24033 5 1 1 24032
0 24034 7 1 2 24026 24033
0 24035 5 1 1 24034
0 24036 7 1 2 61293 24035
0 24037 5 1 1 24036
0 24038 7 4 2 63260 60193
0 24039 7 1 2 65925 90863
0 24040 7 1 2 75118 24039
0 24041 5 1 1 24040
0 24042 7 1 2 59814 24041
0 24043 7 1 2 24037 24042
0 24044 5 1 1 24043
0 24045 7 1 2 73257 89126
0 24046 5 1 1 24045
0 24047 7 3 2 64883 61294
0 24048 7 1 2 78717 83392
0 24049 7 1 2 90867 24048
0 24050 5 1 1 24049
0 24051 7 1 2 24046 24050
0 24052 5 1 1 24051
0 24053 7 1 2 58517 24052
0 24054 5 1 1 24053
0 24055 7 2 2 69817 75022
0 24056 5 1 1 90870
0 24057 7 1 2 90849 90871
0 24058 5 1 1 24057
0 24059 7 1 2 64531 24058
0 24060 7 1 2 24054 24059
0 24061 5 1 1 24060
0 24062 7 1 2 62971 24061
0 24063 7 1 2 24044 24062
0 24064 5 1 1 24063
0 24065 7 1 2 64055 90816
0 24066 5 1 1 24065
0 24067 7 1 2 90253 24066
0 24068 5 1 1 24067
0 24069 7 2 2 62087 77865
0 24070 7 1 2 60194 90872
0 24071 7 1 2 24068 24070
0 24072 5 1 1 24071
0 24073 7 1 2 24064 24072
0 24074 5 1 1 24073
0 24075 7 1 2 61612 24074
0 24076 5 1 1 24075
0 24077 7 1 2 76674 90039
0 24078 5 1 1 24077
0 24079 7 1 2 13483 24078
0 24080 5 1 1 24079
0 24081 7 1 2 71408 24080
0 24082 5 1 1 24081
0 24083 7 1 2 74547 90042
0 24084 5 2 1 24083
0 24085 7 1 2 75524 90874
0 24086 5 1 1 24085
0 24087 7 1 2 24082 24086
0 24088 5 1 1 24087
0 24089 7 1 2 90835 24088
0 24090 5 1 1 24089
0 24091 7 1 2 85586 88357
0 24092 7 2 2 72810 24091
0 24093 5 1 1 90876
0 24094 7 1 2 24090 24093
0 24095 5 1 1 24094
0 24096 7 1 2 66228 24095
0 24097 5 1 1 24096
0 24098 7 1 2 24076 24097
0 24099 7 1 2 24023 24098
0 24100 5 1 1 24099
0 24101 7 1 2 63687 24100
0 24102 5 1 1 24101
0 24103 7 1 2 23995 24102
0 24104 5 1 1 24103
0 24105 7 1 2 62702 24104
0 24106 5 1 1 24105
0 24107 7 2 2 64056 82875
0 24108 5 1 1 90878
0 24109 7 4 2 62426 82685
0 24110 7 1 2 58518 90880
0 24111 5 1 1 24110
0 24112 7 1 2 24108 24111
0 24113 5 1 1 24112
0 24114 7 1 2 79781 24113
0 24115 5 1 1 24114
0 24116 7 3 2 64313 82201
0 24117 5 1 1 90884
0 24118 7 1 2 90420 90885
0 24119 5 1 1 24118
0 24120 7 3 2 63261 79325
0 24121 5 1 1 90887
0 24122 7 2 2 59571 89802
0 24123 5 1 1 90890
0 24124 7 1 2 90888 90891
0 24125 5 1 1 24124
0 24126 7 1 2 24119 24125
0 24127 7 1 2 24115 24126
0 24128 5 1 1 24127
0 24129 7 1 2 61295 24128
0 24130 5 1 1 24129
0 24131 7 1 2 64057 90782
0 24132 5 1 1 24131
0 24133 7 1 2 24130 24132
0 24134 5 1 1 24133
0 24135 7 1 2 60924 24134
0 24136 5 1 1 24135
0 24137 7 1 2 85372 85776
0 24138 5 1 1 24137
0 24139 7 1 2 62972 90817
0 24140 5 1 1 24139
0 24141 7 2 2 89514 24140
0 24142 5 1 1 90892
0 24143 7 1 2 76737 24142
0 24144 5 1 1 24143
0 24145 7 1 2 24138 24144
0 24146 5 1 1 24145
0 24147 7 1 2 61613 24146
0 24148 5 1 1 24147
0 24149 7 1 2 62973 90614
0 24150 5 1 1 24149
0 24151 7 1 2 89515 24150
0 24152 5 1 1 24151
0 24153 7 1 2 88555 24152
0 24154 5 1 1 24153
0 24155 7 1 2 24148 24154
0 24156 7 1 2 24136 24155
0 24157 5 1 1 24156
0 24158 7 1 2 88593 24157
0 24159 5 1 1 24158
0 24160 7 1 2 24106 24159
0 24161 5 1 1 24160
0 24162 7 1 2 66443 24161
0 24163 5 1 1 24162
0 24164 7 6 2 66229 89226
0 24165 7 3 2 71276 73258
0 24166 5 2 1 90900
0 24167 7 1 2 14571 90903
0 24168 5 1 1 24167
0 24169 7 2 2 62427 60195
0 24170 7 1 2 63688 90905
0 24171 7 1 2 24168 24170
0 24172 5 1 1 24171
0 24173 7 1 2 68086 85725
0 24174 5 2 1 24173
0 24175 7 1 2 60925 85943
0 24176 5 1 1 24175
0 24177 7 1 2 90907 24176
0 24178 5 1 1 24177
0 24179 7 1 2 58913 90536
0 24180 7 1 2 24178 24179
0 24181 5 1 1 24180
0 24182 7 1 2 24172 24181
0 24183 5 1 1 24182
0 24184 7 1 2 90146 24183
0 24185 5 1 1 24184
0 24186 7 2 2 62703 63689
0 24187 7 2 2 62974 64884
0 24188 7 6 2 66701 90911
0 24189 7 1 2 73007 90913
0 24190 5 2 1 24189
0 24191 7 1 2 60361 90836
0 24192 5 1 1 24191
0 24193 7 1 2 90919 24192
0 24194 5 1 1 24193
0 24195 7 1 2 62428 24194
0 24196 5 1 1 24195
0 24197 7 2 2 62975 86936
0 24198 7 1 2 66702 90868
0 24199 7 1 2 90921 24198
0 24200 5 1 1 24199
0 24201 7 1 2 24196 24200
0 24202 5 1 1 24201
0 24203 7 1 2 65591 24202
0 24204 5 1 1 24203
0 24205 7 1 2 75482 81134
0 24206 7 1 2 90850 24205
0 24207 5 1 1 24206
0 24208 7 1 2 24204 24207
0 24209 5 1 1 24208
0 24210 7 1 2 90909 24209
0 24211 5 1 1 24210
0 24212 7 1 2 24185 24211
0 24213 5 1 1 24212
0 24214 7 1 2 58519 24213
0 24215 5 1 1 24214
0 24216 7 1 2 78500 88323
0 24217 7 2 2 71996 90543
0 24218 7 1 2 90725 90923
0 24219 7 1 2 24216 24218
0 24220 5 1 1 24219
0 24221 7 1 2 24215 24220
0 24222 5 1 1 24221
0 24223 7 1 2 90894 24222
0 24224 5 1 1 24223
0 24225 7 1 2 24163 24224
0 24226 5 1 1 24225
0 24227 7 1 2 66775 24226
0 24228 5 1 1 24227
0 24229 7 2 2 77982 80669
0 24230 5 1 1 90925
0 24231 7 2 2 65926 73173
0 24232 5 8 1 90927
0 24233 7 1 2 85663 81135
0 24234 7 1 2 90929 24233
0 24235 5 1 1 24234
0 24236 7 1 2 24230 24235
0 24237 5 1 1 24236
0 24238 7 1 2 62704 24237
0 24239 5 2 1 24238
0 24240 7 1 2 71409 72927
0 24241 5 2 1 24240
0 24242 7 1 2 90937 90939
0 24243 5 1 1 24242
0 24244 7 2 2 90567 24243
0 24245 7 3 2 61614 88324
0 24246 7 1 2 79569 90943
0 24247 7 1 2 90941 24246
0 24248 5 1 1 24247
0 24249 7 1 2 24228 24248
0 24250 5 1 1 24249
0 24251 7 1 2 61940 24250
0 24252 5 1 1 24251
0 24253 7 2 2 85567 90734
0 24254 7 2 2 71410 83660
0 24255 7 4 2 86666 90948
0 24256 7 1 2 85796 88325
0 24257 7 1 2 90950 24256
0 24258 7 1 2 90946 24257
0 24259 5 1 1 24258
0 24260 7 1 2 24252 24259
0 24261 5 1 1 24260
0 24262 7 1 2 70507 24261
0 24263 5 1 1 24262
0 24264 7 1 2 72777 89681
0 24265 5 1 1 24264
0 24266 7 2 2 66444 86801
0 24267 7 1 2 80424 90954
0 24268 5 1 1 24267
0 24269 7 1 2 24265 24268
0 24270 5 1 1 24269
0 24271 7 1 2 59572 24270
0 24272 5 2 1 24271
0 24273 7 1 2 62976 89665
0 24274 5 1 1 24273
0 24275 7 1 2 64314 89627
0 24276 5 1 1 24275
0 24277 7 1 2 24274 24276
0 24278 5 1 1 24277
0 24279 7 1 2 60926 24278
0 24280 5 1 1 24279
0 24281 7 1 2 64058 89621
0 24282 5 1 1 24281
0 24283 7 1 2 24280 24282
0 24284 5 1 1 24283
0 24285 7 1 2 58520 24284
0 24286 5 1 1 24285
0 24287 7 1 2 90956 24286
0 24288 5 1 1 24287
0 24289 7 1 2 59815 24288
0 24290 5 1 1 24289
0 24291 7 2 2 73718 81254
0 24292 5 1 1 90958
0 24293 7 4 2 60927 89503
0 24294 7 1 2 90959 90960
0 24295 5 1 1 24294
0 24296 7 1 2 24290 24295
0 24297 5 1 1 24296
0 24298 7 1 2 63690 89127
0 24299 5 1 1 24298
0 24300 7 1 2 89112 24299
0 24301 5 1 1 24300
0 24302 7 1 2 24297 24301
0 24303 5 1 1 24302
0 24304 7 1 2 66445 90843
0 24305 5 1 1 24304
0 24306 7 2 2 65927 81136
0 24307 7 1 2 58521 90964
0 24308 5 1 1 24307
0 24309 7 1 2 18278 24308
0 24310 5 1 1 24309
0 24311 7 1 2 66230 88856
0 24312 7 1 2 90497 24311
0 24313 7 1 2 24310 24312
0 24314 5 1 1 24313
0 24315 7 1 2 24305 24314
0 24316 5 1 1 24315
0 24317 7 1 2 63691 24316
0 24318 5 1 1 24317
0 24319 7 1 2 89684 90035
0 24320 5 1 1 24319
0 24321 7 1 2 78501 24320
0 24322 5 1 1 24321
0 24323 7 1 2 64059 89669
0 24324 5 1 1 24323
0 24325 7 1 2 89623 24324
0 24326 5 1 1 24325
0 24327 7 1 2 58522 24326
0 24328 5 1 1 24327
0 24329 7 1 2 24322 24328
0 24330 5 1 1 24329
0 24331 7 1 2 59816 89101
0 24332 7 1 2 24330 24331
0 24333 5 1 1 24332
0 24334 7 1 2 24318 24333
0 24335 5 1 1 24334
0 24336 7 1 2 62705 24335
0 24337 5 1 1 24336
0 24338 7 1 2 24303 24337
0 24339 5 1 1 24338
0 24340 7 1 2 62429 24339
0 24341 5 1 1 24340
0 24342 7 2 2 64885 89016
0 24343 7 1 2 74128 75463
0 24344 7 6 2 62706 58523
0 24345 7 1 2 90670 90968
0 24346 7 1 2 24343 24345
0 24347 7 1 2 90966 24346
0 24348 5 1 1 24347
0 24349 7 2 2 86897 88594
0 24350 7 4 2 71493 73174
0 24351 5 4 1 90976
0 24352 7 2 2 84635 90977
0 24353 5 2 1 90984
0 24354 7 1 2 89080 90986
0 24355 7 1 2 90974 24354
0 24356 5 1 1 24355
0 24357 7 1 2 24348 24356
0 24358 5 1 1 24357
0 24359 7 1 2 66231 24358
0 24360 5 1 1 24359
0 24361 7 1 2 24341 24360
0 24362 5 1 1 24361
0 24363 7 1 2 69540 24362
0 24364 5 1 1 24363
0 24365 7 1 2 78042 89081
0 24366 5 1 1 24365
0 24367 7 1 2 75453 87421
0 24368 5 7 1 24367
0 24369 7 4 2 62430 61815
0 24370 7 1 2 59817 90995
0 24371 7 1 2 90988 24370
0 24372 5 1 1 24371
0 24373 7 1 2 24366 24372
0 24374 5 1 1 24373
0 24375 7 1 2 68087 24374
0 24376 5 1 1 24375
0 24377 7 5 2 63262 66446
0 24378 7 1 2 85439 90999
0 24379 5 1 1 24378
0 24380 7 1 2 85264 90996
0 24381 7 1 2 85693 24380
0 24382 5 1 1 24381
0 24383 7 1 2 24379 24382
0 24384 7 1 2 24376 24383
0 24385 5 1 1 24384
0 24386 7 1 2 65928 24385
0 24387 5 1 1 24386
0 24388 7 4 2 58524 73377
0 24389 5 1 1 91004
0 24390 7 1 2 85834 90997
0 24391 7 1 2 91005 24390
0 24392 5 1 1 24391
0 24393 7 1 2 24387 24392
0 24394 5 1 1 24393
0 24395 7 1 2 66232 24394
0 24396 5 1 1 24395
0 24397 7 1 2 77840 90092
0 24398 5 1 1 24397
0 24399 7 1 2 84241 90027
0 24400 7 1 2 80853 24399
0 24401 7 1 2 24398 24400
0 24402 5 1 1 24401
0 24403 7 1 2 24396 24402
0 24404 5 1 1 24403
0 24405 7 1 2 90764 24404
0 24406 5 1 1 24405
0 24407 7 1 2 24364 24406
0 24408 5 1 1 24407
0 24409 7 1 2 60362 24408
0 24410 5 1 1 24409
0 24411 7 3 2 59818 72778
0 24412 7 1 2 86725 88542
0 24413 5 1 1 24412
0 24414 7 2 2 64315 88144
0 24415 7 3 2 62431 80425
0 24416 7 1 2 86621 91013
0 24417 7 1 2 91011 24416
0 24418 5 1 1 24417
0 24419 7 1 2 24413 24418
0 24420 5 1 1 24419
0 24421 7 1 2 91008 24420
0 24422 5 1 1 24421
0 24423 7 2 2 77586 90544
0 24424 7 1 2 88515 91016
0 24425 5 1 1 24424
0 24426 7 1 2 88326 91017
0 24427 5 1 1 24426
0 24428 7 2 2 83393 88124
0 24429 7 1 2 79216 73622
0 24430 7 1 2 91018 24429
0 24431 5 1 1 24430
0 24432 7 1 2 24427 24431
0 24433 5 1 1 24432
0 24434 7 1 2 69541 24433
0 24435 5 1 1 24434
0 24436 7 1 2 24425 24435
0 24437 5 1 1 24436
0 24438 7 1 2 76738 24437
0 24439 5 1 1 24438
0 24440 7 1 2 24422 24439
0 24441 5 1 1 24440
0 24442 7 1 2 89645 24441
0 24443 5 1 1 24442
0 24444 7 1 2 87485 90579
0 24445 7 2 2 78078 87876
0 24446 7 3 2 63621 63692
0 24447 7 2 2 90671 91022
0 24448 7 1 2 91020 91025
0 24449 7 1 2 24444 24448
0 24450 5 1 1 24449
0 24451 7 1 2 24443 24450
0 24452 5 1 1 24451
0 24453 7 1 2 62707 24452
0 24454 5 1 1 24453
0 24455 7 1 2 24410 24454
0 24456 5 1 1 24455
0 24457 7 1 2 66833 24456
0 24458 5 1 1 24457
0 24459 7 1 2 67928 88327
0 24460 5 1 1 24459
0 24461 7 1 2 58914 87861
0 24462 5 1 1 24461
0 24463 7 1 2 24460 24462
0 24464 5 2 1 24463
0 24465 7 1 2 86331 87911
0 24466 7 1 2 91027 24465
0 24467 7 1 2 90942 24466
0 24468 5 1 1 24467
0 24469 7 1 2 24458 24468
0 24470 5 1 1 24469
0 24471 7 1 2 61941 24470
0 24472 5 1 1 24471
0 24473 7 4 2 80808 79451
0 24474 5 1 1 91029
0 24475 7 2 2 84003 85797
0 24476 5 1 1 91033
0 24477 7 1 2 91030 91034
0 24478 7 1 2 88523 24477
0 24479 7 1 2 90947 24478
0 24480 5 1 1 24479
0 24481 7 1 2 24472 24480
0 24482 7 1 2 24263 24481
0 24483 5 1 1 24482
0 24484 7 1 2 68832 24483
0 24485 5 1 1 24484
0 24486 7 2 2 82524 88912
0 24487 7 1 2 58290 77346
0 24488 7 1 2 91035 24487
0 24489 5 1 1 24488
0 24490 7 1 2 71411 90721
0 24491 7 1 2 90046 24490
0 24492 5 1 1 24491
0 24493 7 1 2 24489 24492
0 24494 5 1 1 24493
0 24495 7 1 2 83080 24494
0 24496 5 1 1 24495
0 24497 7 1 2 70656 86937
0 24498 7 1 2 91036 24497
0 24499 5 1 1 24498
0 24500 7 1 2 24496 24499
0 24501 5 1 1 24500
0 24502 7 1 2 88358 24501
0 24503 5 1 1 24502
0 24504 7 1 2 65592 71010
0 24505 5 3 1 24504
0 24506 7 1 2 78181 91037
0 24507 5 1 1 24506
0 24508 7 1 2 71494 24507
0 24509 5 2 1 24508
0 24510 7 1 2 84164 88768
0 24511 7 1 2 91040 24510
0 24512 5 1 1 24511
0 24513 7 1 2 24503 24512
0 24514 5 1 1 24513
0 24515 7 1 2 65929 24514
0 24516 5 1 1 24515
0 24517 7 1 2 82392 90746
0 24518 5 1 1 24517
0 24519 7 2 2 63766 24518
0 24520 5 1 1 91042
0 24521 7 1 2 90741 24520
0 24522 5 1 1 24521
0 24523 7 1 2 89128 24522
0 24524 5 1 1 24523
0 24525 7 1 2 81550 89129
0 24526 5 1 1 24525
0 24527 7 1 2 77618 90518
0 24528 7 1 2 90739 24527
0 24529 5 1 1 24528
0 24530 7 1 2 24526 24529
0 24531 5 1 1 24530
0 24532 7 1 2 62432 24531
0 24533 5 1 1 24532
0 24534 7 1 2 24524 24533
0 24535 5 1 1 24534
0 24536 7 1 2 60928 24535
0 24537 5 1 1 24536
0 24538 7 2 2 79490 81009
0 24539 5 1 1 91044
0 24540 7 1 2 90509 91045
0 24541 5 1 1 24540
0 24542 7 1 2 24537 24541
0 24543 5 1 1 24542
0 24544 7 1 2 62189 24543
0 24545 5 1 1 24544
0 24546 7 3 2 60929 78290
0 24547 5 1 1 91046
0 24548 7 1 2 82381 91047
0 24549 5 1 1 24548
0 24550 7 1 2 59366 72199
0 24551 5 2 1 24550
0 24552 7 1 2 60930 91049
0 24553 5 1 1 24552
0 24554 7 1 2 75413 24553
0 24555 5 1 1 24554
0 24556 7 1 2 84128 24555
0 24557 5 1 1 24556
0 24558 7 1 2 24549 24557
0 24559 5 1 1 24558
0 24560 7 1 2 89130 24559
0 24561 5 1 1 24560
0 24562 7 1 2 24545 24561
0 24563 5 1 1 24562
0 24564 7 1 2 90759 24563
0 24565 5 1 1 24564
0 24566 7 1 2 24516 24565
0 24567 5 1 1 24566
0 24568 7 1 2 63693 24567
0 24569 5 1 1 24568
0 24570 7 1 2 65930 91041
0 24571 5 1 1 24570
0 24572 7 2 2 73046 77729
0 24573 5 1 1 91051
0 24574 7 1 2 60931 91052
0 24575 5 1 1 24574
0 24576 7 1 2 24571 24575
0 24577 5 1 1 24576
0 24578 7 1 2 61615 24577
0 24579 5 1 1 24578
0 24580 7 2 2 72200 87949
0 24581 5 3 1 91053
0 24582 7 1 2 60932 91055
0 24583 5 1 1 24582
0 24584 7 1 2 59367 24583
0 24585 5 1 1 24584
0 24586 7 3 2 71412 84663
0 24587 5 1 1 91058
0 24588 7 1 2 91038 91059
0 24589 7 1 2 24585 24588
0 24590 5 1 1 24589
0 24591 7 1 2 24579 24590
0 24592 5 1 1 24591
0 24593 7 1 2 88388 89291
0 24594 7 1 2 24592 24593
0 24595 5 1 1 24594
0 24596 7 1 2 24569 24595
0 24597 5 1 1 24596
0 24598 7 1 2 62708 24597
0 24599 5 1 1 24598
0 24600 7 2 2 77347 86648
0 24601 5 2 1 91061
0 24602 7 1 2 86513 90829
0 24603 5 2 1 24602
0 24604 7 1 2 64316 77395
0 24605 7 1 2 91065 24604
0 24606 5 1 1 24605
0 24607 7 1 2 91063 24606
0 24608 5 1 1 24607
0 24609 7 1 2 78291 24608
0 24610 5 1 1 24609
0 24611 7 1 2 62433 71413
0 24612 7 1 2 91066 24611
0 24613 5 1 1 24612
0 24614 7 1 2 62190 91062
0 24615 5 1 1 24614
0 24616 7 1 2 24613 24615
0 24617 5 1 1 24616
0 24618 7 1 2 69029 24617
0 24619 5 1 1 24618
0 24620 7 2 2 64060 77092
0 24621 5 2 1 91067
0 24622 7 1 2 59573 91069
0 24623 5 1 1 24622
0 24624 7 1 2 73259 90232
0 24625 7 1 2 24623 24624
0 24626 5 1 1 24625
0 24627 7 1 2 24619 24626
0 24628 7 1 2 24610 24627
0 24629 5 1 1 24628
0 24630 7 1 2 88595 88702
0 24631 7 1 2 24629 24630
0 24632 5 1 1 24631
0 24633 7 1 2 24599 24632
0 24634 5 1 1 24633
0 24635 7 1 2 69542 24634
0 24636 5 1 1 24635
0 24637 7 3 2 60363 86474
0 24638 5 2 1 91071
0 24639 7 1 2 62434 86687
0 24640 5 1 1 24639
0 24641 7 1 2 91074 24640
0 24642 5 1 1 24641
0 24643 7 1 2 68833 24642
0 24644 5 1 1 24643
0 24645 7 2 2 66233 70638
0 24646 7 1 2 87697 91076
0 24647 5 1 1 24646
0 24648 7 1 2 86514 86691
0 24649 5 4 1 24648
0 24650 7 1 2 62709 91078
0 24651 5 1 1 24650
0 24652 7 1 2 24647 24651
0 24653 7 1 2 24644 24652
0 24654 5 1 1 24653
0 24655 7 1 2 62977 24654
0 24656 5 1 1 24655
0 24657 7 2 2 62710 73008
0 24658 5 1 1 91082
0 24659 7 1 2 24658 24573
0 24660 5 1 1 24659
0 24661 7 1 2 61616 24660
0 24662 5 1 1 24661
0 24663 7 1 2 24656 24662
0 24664 5 1 1 24663
0 24665 7 1 2 64061 24664
0 24666 5 1 1 24665
0 24667 7 1 2 62191 91043
0 24668 5 1 1 24667
0 24669 7 1 2 79217 81336
0 24670 5 2 1 24669
0 24671 7 1 2 90742 91084
0 24672 5 1 1 24671
0 24673 7 1 2 68834 24672
0 24674 5 1 1 24673
0 24675 7 1 2 24123 24674
0 24676 7 1 2 24668 24675
0 24677 5 1 1 24676
0 24678 7 1 2 90054 24677
0 24679 5 1 1 24678
0 24680 7 1 2 16493 24679
0 24681 7 1 2 24666 24680
0 24682 5 1 1 24681
0 24683 7 1 2 60933 24682
0 24684 5 1 1 24683
0 24685 7 1 2 58032 85926
0 24686 5 1 1 24685
0 24687 7 1 2 86963 24686
0 24688 5 1 1 24687
0 24689 7 1 2 58291 87190
0 24690 5 1 1 24689
0 24691 7 1 2 67199 24690
0 24692 7 1 2 71004 24691
0 24693 7 1 2 91079 24692
0 24694 5 1 1 24693
0 24695 7 1 2 24688 24694
0 24696 7 1 2 24684 24695
0 24697 5 1 1 24696
0 24698 7 1 2 88516 89292
0 24699 7 1 2 24697 24698
0 24700 5 1 1 24699
0 24701 7 1 2 24636 24700
0 24702 5 1 1 24701
0 24703 7 1 2 76739 24702
0 24704 5 1 1 24703
0 24705 7 1 2 62978 90627
0 24706 5 1 1 24705
0 24707 7 3 2 73009 90768
0 24708 5 1 1 91086
0 24709 7 1 2 24706 24708
0 24710 5 1 1 24709
0 24711 7 3 2 60934 24710
0 24712 5 1 1 91089
0 24713 7 1 2 62711 91087
0 24714 5 1 1 24713
0 24715 7 1 2 24712 24714
0 24716 5 1 1 24715
0 24717 7 1 2 64062 24716
0 24718 5 1 1 24717
0 24719 7 2 2 62979 73010
0 24720 5 1 1 91092
0 24721 7 1 2 89607 91093
0 24722 5 1 1 24721
0 24723 7 1 2 24718 24722
0 24724 5 1 1 24723
0 24725 7 1 2 88543 24724
0 24726 5 1 1 24725
0 24727 7 1 2 89897 90055
0 24728 7 1 2 91023 24727
0 24729 7 1 2 64886 69715
0 24730 7 1 2 80893 24729
0 24731 7 1 2 67550 24730
0 24732 7 1 2 24728 24731
0 24733 5 1 1 24732
0 24734 7 1 2 24726 24733
0 24735 5 1 1 24734
0 24736 7 1 2 68835 24735
0 24737 5 1 1 24736
0 24738 7 2 2 61942 89131
0 24739 7 2 2 66447 91094
0 24740 7 3 2 73047 81399
0 24741 5 1 1 91098
0 24742 7 1 2 91096 91099
0 24743 5 1 1 24742
0 24744 7 1 2 63767 75084
0 24745 7 1 2 89986 24744
0 24746 5 1 1 24745
0 24747 7 1 2 23875 24746
0 24748 5 1 1 24747
0 24749 7 1 2 77609 90914
0 24750 7 1 2 24748 24749
0 24751 5 1 1 24750
0 24752 7 1 2 24743 24751
0 24753 5 1 1 24752
0 24754 7 1 2 88509 24753
0 24755 5 1 1 24754
0 24756 7 1 2 88521 18911
0 24757 5 1 1 24756
0 24758 7 1 2 88996 91100
0 24759 7 1 2 24757 24758
0 24760 5 1 1 24759
0 24761 7 1 2 24755 24760
0 24762 5 1 1 24761
0 24763 7 1 2 64063 24762
0 24764 5 1 1 24763
0 24765 7 1 2 24737 24764
0 24766 5 1 1 24765
0 24767 7 1 2 60364 24766
0 24768 5 1 1 24767
0 24769 7 1 2 77621 90163
0 24770 5 1 1 24769
0 24771 7 1 2 62192 24770
0 24772 5 1 1 24771
0 24773 7 1 2 83278 24772
0 24774 5 1 1 24773
0 24775 7 1 2 88544 91090
0 24776 5 1 1 24775
0 24777 7 2 2 63694 90537
0 24778 7 2 2 74129 89475
0 24779 7 1 2 91101 91103
0 24780 7 1 2 90318 24779
0 24781 5 1 1 24780
0 24782 7 1 2 24776 24781
0 24783 5 1 1 24782
0 24784 7 1 2 24774 24783
0 24785 5 1 1 24784
0 24786 7 1 2 87585 91088
0 24787 5 1 1 24786
0 24788 7 1 2 83907 23653
0 24789 5 1 1 24788
0 24790 7 1 2 91091 24789
0 24791 5 1 1 24790
0 24792 7 1 2 24787 24791
0 24793 5 1 1 24792
0 24794 7 1 2 88545 24793
0 24795 5 1 1 24794
0 24796 7 1 2 24785 24795
0 24797 7 1 2 24768 24796
0 24798 5 1 1 24797
0 24799 7 1 2 76638 24798
0 24800 5 1 1 24799
0 24801 7 1 2 87199 88999
0 24802 5 1 1 24801
0 24803 7 5 2 66592 66703
0 24804 7 1 2 61816 91105
0 24805 7 2 2 90047 24804
0 24806 7 5 2 64532 64887
0 24807 7 1 2 78985 86802
0 24808 7 1 2 91112 24807
0 24809 7 1 2 91110 24808
0 24810 5 1 1 24809
0 24811 7 1 2 24802 24810
0 24812 5 1 1 24811
0 24813 7 1 2 59574 24812
0 24814 5 1 1 24813
0 24815 7 1 2 61296 90516
0 24816 5 1 1 24815
0 24817 7 1 2 90920 24816
0 24818 5 1 1 24817
0 24819 7 6 2 59819 82656
0 24820 7 2 2 65593 66448
0 24821 7 1 2 85625 91123
0 24822 7 1 2 91117 24821
0 24823 7 1 2 24818 24822
0 24824 5 1 1 24823
0 24825 7 1 2 24814 24824
0 24826 5 1 1 24825
0 24827 7 1 2 62712 24826
0 24828 5 1 1 24827
0 24829 7 1 2 89767 90830
0 24830 5 1 1 24829
0 24831 7 1 2 59575 24830
0 24832 5 1 1 24831
0 24833 7 1 2 89545 90130
0 24834 5 1 1 24833
0 24835 7 1 2 24832 24834
0 24836 5 2 1 24835
0 24837 7 1 2 89005 91095
0 24838 7 1 2 91125 24837
0 24839 5 1 1 24838
0 24840 7 1 2 24828 24839
0 24841 5 1 1 24840
0 24842 7 1 2 63695 24841
0 24843 5 1 1 24842
0 24844 7 1 2 62713 90875
0 24845 5 1 1 24844
0 24846 7 1 2 65043 82699
0 24847 5 1 1 24846
0 24848 7 1 2 79410 24847
0 24849 7 1 2 24845 24848
0 24850 5 1 1 24849
0 24851 7 1 2 84664 24850
0 24852 5 1 1 24851
0 24853 7 1 2 89521 24852
0 24854 5 1 1 24853
0 24855 7 2 2 89027 24854
0 24856 7 1 2 58915 76639
0 24857 7 1 2 91127 24856
0 24858 5 1 1 24857
0 24859 7 1 2 24843 24858
0 24860 5 1 1 24859
0 24861 7 1 2 69543 24860
0 24862 5 1 1 24861
0 24863 7 1 2 89020 91128
0 24864 5 1 1 24863
0 24865 7 1 2 24862 24864
0 24866 5 1 1 24865
0 24867 7 1 2 83081 24866
0 24868 5 1 1 24867
0 24869 7 1 2 89634 22773
0 24870 5 1 1 24869
0 24871 7 1 2 62980 24870
0 24872 5 1 1 24871
0 24873 7 6 2 61817 81870
0 24874 7 1 2 61297 91129
0 24875 5 1 1 24874
0 24876 7 1 2 24872 24875
0 24877 5 1 1 24876
0 24878 7 1 2 75772 24877
0 24879 5 1 1 24878
0 24880 7 1 2 79224 3536
0 24881 5 1 1 24880
0 24882 7 8 2 65931 61818
0 24883 7 1 2 84178 91135
0 24884 7 1 2 24881 24883
0 24885 5 1 1 24884
0 24886 7 1 2 24879 24885
0 24887 5 1 1 24886
0 24888 7 1 2 64064 24887
0 24889 5 1 1 24888
0 24890 7 1 2 61819 84404
0 24891 5 1 1 24890
0 24892 7 1 2 24889 24891
0 24893 5 1 1 24892
0 24894 7 1 2 60935 24893
0 24895 5 1 1 24894
0 24896 7 1 2 65594 75492
0 24897 5 3 1 24896
0 24898 7 1 2 64065 91143
0 24899 5 1 1 24898
0 24900 7 5 2 60936 68836
0 24901 5 4 1 91146
0 24902 7 1 2 62435 91147
0 24903 5 3 1 24902
0 24904 7 1 2 24899 91155
0 24905 5 1 1 24904
0 24906 7 1 2 91130 24905
0 24907 5 1 1 24906
0 24908 7 1 2 71681 91131
0 24909 5 1 1 24908
0 24910 7 2 2 66449 69030
0 24911 7 1 2 78579 90233
0 24912 7 1 2 91158 24911
0 24913 5 1 1 24912
0 24914 7 1 2 24909 24913
0 24915 5 1 1 24914
0 24916 7 1 2 62193 24915
0 24917 5 1 1 24916
0 24918 7 3 2 79491 89646
0 24919 7 1 2 62436 81010
0 24920 7 1 2 91160 24919
0 24921 5 1 1 24920
0 24922 7 1 2 24917 24921
0 24923 5 1 1 24922
0 24924 7 1 2 70204 24923
0 24925 5 1 1 24924
0 24926 7 1 2 24907 24925
0 24927 5 1 1 24926
0 24928 7 1 2 61298 24927
0 24929 5 1 1 24928
0 24930 7 2 2 61820 86562
0 24931 7 1 2 72786 91054
0 24932 5 1 1 24931
0 24933 7 1 2 78043 24932
0 24934 5 1 1 24933
0 24935 7 1 2 71495 24934
0 24936 5 1 1 24935
0 24937 7 1 2 91163 24936
0 24938 5 1 1 24937
0 24939 7 1 2 24929 24938
0 24940 5 1 1 24939
0 24941 7 1 2 62714 24940
0 24942 5 1 1 24941
0 24943 7 1 2 24895 24942
0 24944 5 1 1 24943
0 24945 7 1 2 88524 24944
0 24946 5 1 1 24945
0 24947 7 2 2 70639 88525
0 24948 7 1 2 90037 90922
0 24949 7 1 2 91165 24948
0 24950 5 1 1 24949
0 24951 7 1 2 24946 24950
0 24952 5 1 1 24951
0 24953 7 1 2 75525 67474
0 24954 7 1 2 24952 24953
0 24955 5 1 1 24954
0 24956 7 1 2 24868 24955
0 24957 7 1 2 24800 24956
0 24958 7 1 2 24704 24957
0 24959 5 1 1 24958
0 24960 7 1 2 66903 24959
0 24961 5 1 1 24960
0 24962 7 2 2 71179 66776
0 24963 7 1 2 89160 91167
0 24964 7 1 2 91111 24963
0 24965 5 1 1 24964
0 24966 7 1 2 71277 88991
0 24967 7 1 2 74249 24966
0 24968 7 1 2 89218 24967
0 24969 5 1 1 24968
0 24970 7 1 2 24965 24969
0 24971 5 1 1 24970
0 24972 7 1 2 58525 24971
0 24973 5 1 1 24972
0 24974 7 1 2 63263 79337
0 24975 5 2 1 24974
0 24976 7 1 2 73719 90040
0 24977 5 1 1 24976
0 24978 7 1 2 91169 24977
0 24979 5 1 1 24978
0 24980 7 1 2 62981 24979
0 24981 5 1 1 24980
0 24982 7 1 2 77983 77799
0 24983 5 1 1 24982
0 24984 7 1 2 24981 24983
0 24985 5 1 1 24984
0 24986 7 2 2 66834 91097
0 24987 7 1 2 24985 91171
0 24988 5 1 1 24987
0 24989 7 1 2 24973 24988
0 24990 5 1 1 24989
0 24991 7 1 2 62715 24990
0 24992 5 1 1 24991
0 24993 7 1 2 78160 87426
0 24994 5 1 1 24993
0 24995 7 3 2 71278 77866
0 24996 7 1 2 90980 91173
0 24997 5 1 1 24996
0 24998 7 1 2 24994 24997
0 24999 5 1 1 24998
0 25000 7 1 2 91172 24999
0 25001 5 1 1 25000
0 25002 7 1 2 24992 25001
0 25003 5 1 1 25002
0 25004 7 1 2 63696 25003
0 25005 5 1 1 25004
0 25006 7 1 2 77867 82294
0 25007 7 1 2 82861 25006
0 25008 5 1 1 25007
0 25009 7 1 2 90082 25008
0 25010 5 1 1 25009
0 25011 7 1 2 66450 75657
0 25012 7 1 2 89102 25011
0 25013 7 1 2 25010 25012
0 25014 5 1 1 25013
0 25015 7 1 2 25005 25014
0 25016 5 1 1 25015
0 25017 7 1 2 65932 25016
0 25018 5 1 1 25017
0 25019 7 1 2 67200 85147
0 25020 5 1 1 25019
0 25021 7 3 2 82948 25020
0 25022 5 7 1 91176
0 25023 7 1 2 59820 91179
0 25024 5 1 1 25023
0 25025 7 1 2 77818 85694
0 25026 5 1 1 25025
0 25027 7 1 2 25024 25026
0 25028 5 1 1 25027
0 25029 7 1 2 67956 89504
0 25030 7 1 2 82280 25029
0 25031 7 1 2 88328 25030
0 25032 7 1 2 25028 25031
0 25033 5 1 1 25032
0 25034 7 1 2 25018 25033
0 25035 5 1 1 25034
0 25036 7 1 2 61617 25035
0 25037 5 1 1 25036
0 25038 7 1 2 90877 90910
0 25039 5 1 1 25038
0 25040 7 1 2 73916 80972
0 25041 5 1 1 25040
0 25042 7 1 2 72027 80991
0 25043 5 1 1 25042
0 25044 7 1 2 25041 25043
0 25045 5 1 1 25044
0 25046 7 1 2 80030 88329
0 25047 7 1 2 25045 25046
0 25048 5 1 1 25047
0 25049 7 1 2 25039 25048
0 25050 5 1 1 25049
0 25051 7 2 2 66234 66835
0 25052 7 1 2 88913 91186
0 25053 7 1 2 25050 25052
0 25054 5 1 1 25053
0 25055 7 1 2 25037 25054
0 25056 5 1 1 25055
0 25057 7 1 2 69544 25056
0 25058 5 1 1 25057
0 25059 7 1 2 58033 79350
0 25060 5 1 1 25059
0 25061 7 1 2 79345 90043
0 25062 5 1 1 25061
0 25063 7 1 2 81337 25062
0 25064 7 1 2 25060 25063
0 25065 5 1 1 25064
0 25066 7 1 2 89779 25065
0 25067 5 1 1 25066
0 25068 7 1 2 61299 25067
0 25069 5 1 1 25068
0 25070 7 2 2 59821 86475
0 25071 7 1 2 59576 73922
0 25072 5 1 1 25071
0 25073 7 1 2 91188 25072
0 25074 5 1 1 25073
0 25075 7 1 2 25069 25074
0 25076 5 1 1 25075
0 25077 7 1 2 62982 25076
0 25078 5 1 1 25077
0 25079 7 1 2 73623 79841
0 25080 5 2 1 25079
0 25081 7 1 2 90254 91190
0 25082 5 1 1 25081
0 25083 7 1 2 62716 25082
0 25084 5 1 1 25083
0 25085 7 2 2 64066 73260
0 25086 5 2 1 91192
0 25087 7 2 2 86215 91194
0 25088 5 1 1 91196
0 25089 7 1 2 64317 25088
0 25090 5 1 1 25089
0 25091 7 1 2 25084 25090
0 25092 5 1 1 25091
0 25093 7 1 2 82554 25092
0 25094 5 1 1 25093
0 25095 7 1 2 25078 25094
0 25096 5 1 1 25095
0 25097 7 1 2 63264 25096
0 25098 5 1 1 25097
0 25099 7 1 2 85626 82514
0 25100 5 1 1 25099
0 25101 7 1 2 60937 72805
0 25102 5 1 1 25101
0 25103 7 1 2 90044 25102
0 25104 5 1 1 25103
0 25105 7 1 2 66235 85148
0 25106 7 1 2 25104 25105
0 25107 5 1 1 25106
0 25108 7 1 2 25100 25107
0 25109 5 1 1 25108
0 25110 7 1 2 61300 25109
0 25111 5 1 1 25110
0 25112 7 2 2 58526 77984
0 25113 5 1 1 91198
0 25114 7 1 2 76983 24056
0 25115 5 1 1 25114
0 25116 7 1 2 62983 25115
0 25117 5 1 1 25116
0 25118 7 1 2 25113 25117
0 25119 5 1 1 25118
0 25120 7 1 2 86476 25119
0 25121 5 1 1 25120
0 25122 7 1 2 25111 25121
0 25123 5 1 1 25122
0 25124 7 1 2 62717 25123
0 25125 5 1 1 25124
0 25126 7 1 2 63265 91126
0 25127 5 1 1 25126
0 25128 7 1 2 74732 91197
0 25129 5 1 1 25128
0 25130 7 1 2 89777 25129
0 25131 5 1 1 25130
0 25132 7 1 2 87026 81551
0 25133 5 1 1 25132
0 25134 7 1 2 25131 25133
0 25135 5 1 1 25134
0 25136 7 1 2 58527 25135
0 25137 5 1 1 25136
0 25138 7 1 2 25127 25137
0 25139 7 1 2 25125 25138
0 25140 5 1 1 25139
0 25141 7 1 2 64533 25140
0 25142 5 1 1 25141
0 25143 7 2 2 65595 84778
0 25144 7 1 2 85005 79658
0 25145 7 1 2 91200 25144
0 25146 5 1 1 25145
0 25147 7 1 2 25142 25146
0 25148 7 1 2 25098 25147
0 25149 5 1 1 25148
0 25150 7 2 2 60125 83552
0 25151 7 3 2 60005 64888
0 25152 7 3 2 63697 91204
0 25153 7 2 2 91202 91207
0 25154 5 1 1 91210
0 25155 7 1 2 88997 91211
0 25156 7 1 2 25149 25155
0 25157 5 1 1 25156
0 25158 7 1 2 25058 25157
0 25159 5 1 1 25158
0 25160 7 1 2 83082 25159
0 25161 5 1 1 25160
0 25162 7 2 2 63698 88158
0 25163 5 1 1 91212
0 25164 7 1 2 18913 25163
0 25165 5 5 1 25164
0 25166 7 1 2 89707 91144
0 25167 5 1 1 25166
0 25168 7 1 2 57421 80601
0 25169 5 2 1 25168
0 25170 7 3 2 81588 91219
0 25171 5 1 1 91221
0 25172 7 1 2 71414 89257
0 25173 7 1 2 91222 25172
0 25174 5 1 1 25173
0 25175 7 1 2 25167 25174
0 25176 5 1 1 25175
0 25177 7 1 2 58528 25176
0 25178 5 1 1 25177
0 25179 7 1 2 79659 91148
0 25180 5 1 1 25179
0 25181 7 1 2 75005 86011
0 25182 5 1 1 25181
0 25183 7 1 2 79782 25182
0 25184 5 1 1 25183
0 25185 7 1 2 25180 25184
0 25186 5 1 1 25185
0 25187 7 1 2 91000 25186
0 25188 5 1 1 25187
0 25189 7 1 2 25178 25188
0 25190 5 1 1 25189
0 25191 7 1 2 64067 25190
0 25192 5 1 1 25191
0 25193 7 1 2 61821 68837
0 25194 7 1 2 85265 25193
0 25195 5 1 1 25194
0 25196 7 2 2 66451 80833
0 25197 5 1 1 91224
0 25198 7 1 2 25195 25197
0 25199 5 1 1 25198
0 25200 7 1 2 59577 25199
0 25201 5 1 1 25200
0 25202 7 2 2 74191 89258
0 25203 5 1 1 91226
0 25204 7 1 2 69313 91227
0 25205 5 1 1 25204
0 25206 7 1 2 25201 25205
0 25207 5 1 1 25206
0 25208 7 1 2 62437 25207
0 25209 5 1 1 25208
0 25210 7 1 2 25192 25209
0 25211 5 1 1 25210
0 25212 7 1 2 66236 25211
0 25213 5 1 1 25212
0 25214 7 1 2 71496 77841
0 25215 5 1 1 25214
0 25216 7 5 2 85212 25215
0 25217 7 4 2 61618 78851
0 25218 7 2 2 62438 66452
0 25219 7 2 2 91233 91237
0 25220 7 1 2 91228 91239
0 25221 5 1 1 25220
0 25222 7 1 2 63768 79326
0 25223 7 1 2 89455 25222
0 25224 7 1 2 91132 25223
0 25225 5 1 1 25224
0 25226 7 1 2 25221 25225
0 25227 5 1 1 25226
0 25228 7 1 2 70205 25227
0 25229 5 1 1 25228
0 25230 7 1 2 61301 25229
0 25231 7 1 2 25213 25230
0 25232 5 1 1 25231
0 25233 7 1 2 89051 91056
0 25234 5 1 1 25233
0 25235 7 2 2 65044 89259
0 25236 7 1 2 64068 84453
0 25237 7 1 2 91241 25236
0 25238 5 1 1 25237
0 25239 7 1 2 25234 25238
0 25240 5 1 1 25239
0 25241 7 1 2 71279 25240
0 25242 5 1 1 25241
0 25243 7 1 2 72779 89052
0 25244 5 1 1 25243
0 25245 7 1 2 25242 25244
0 25246 5 1 1 25245
0 25247 7 1 2 60938 25246
0 25248 5 1 1 25247
0 25249 7 1 2 75441 89227
0 25250 5 1 1 25249
0 25251 7 1 2 78718 89082
0 25252 7 1 2 86788 25251
0 25253 5 1 1 25252
0 25254 7 1 2 25250 25253
0 25255 5 1 1 25254
0 25256 7 1 2 62984 25255
0 25257 5 1 1 25256
0 25258 7 1 2 25248 25257
0 25259 5 1 1 25258
0 25260 7 1 2 66237 25259
0 25261 5 1 1 25260
0 25262 7 1 2 90845 91240
0 25263 5 1 1 25262
0 25264 7 9 2 65596 89587
0 25265 5 2 1 91243
0 25266 7 1 2 72987 91244
0 25267 5 1 1 25266
0 25268 7 1 2 25263 25267
0 25269 5 1 1 25268
0 25270 7 1 2 76740 25269
0 25271 5 1 1 25270
0 25272 7 1 2 65933 25271
0 25273 7 1 2 25261 25272
0 25274 5 1 1 25273
0 25275 7 1 2 62718 25274
0 25276 7 1 2 25232 25275
0 25277 5 1 1 25276
0 25278 7 4 2 82407 89445
0 25279 7 1 2 74480 75773
0 25280 5 1 1 25279
0 25281 7 1 2 73075 25280
0 25282 5 1 1 25281
0 25283 7 1 2 60939 25282
0 25284 5 1 1 25283
0 25285 7 1 2 72898 90930
0 25286 7 1 2 71005 25285
0 25287 5 1 1 25286
0 25288 7 1 2 25284 25287
0 25289 5 1 1 25288
0 25290 7 1 2 91254 25289
0 25291 5 1 1 25290
0 25292 7 2 2 68838 75483
0 25293 5 2 1 91258
0 25294 7 1 2 70172 91260
0 25295 5 2 1 25294
0 25296 7 1 2 89964 91262
0 25297 5 1 1 25296
0 25298 7 2 2 76640 86440
0 25299 7 1 2 91264 91259
0 25300 5 1 1 25299
0 25301 7 1 2 25297 25300
0 25302 5 1 1 25301
0 25303 7 1 2 61619 25302
0 25304 5 1 1 25303
0 25305 7 1 2 89813 90879
0 25306 5 1 1 25305
0 25307 7 1 2 61302 25306
0 25308 7 1 2 25304 25307
0 25309 5 1 1 25308
0 25310 7 1 2 88007 91263
0 25311 5 1 1 25310
0 25312 7 1 2 72724 78788
0 25313 7 1 2 88556 25312
0 25314 5 1 1 25313
0 25315 7 1 2 25311 25314
0 25316 5 1 1 25315
0 25317 7 1 2 64318 25316
0 25318 5 1 1 25317
0 25319 7 3 2 68839 77868
0 25320 7 1 2 73117 90881
0 25321 7 1 2 91266 25320
0 25322 5 1 1 25321
0 25323 7 1 2 65934 25322
0 25324 7 1 2 25318 25323
0 25325 5 1 1 25324
0 25326 7 1 2 66453 25325
0 25327 7 1 2 25309 25326
0 25328 5 1 1 25327
0 25329 7 1 2 25291 25328
0 25330 5 1 1 25329
0 25331 7 1 2 62985 25330
0 25332 5 1 1 25331
0 25333 7 3 2 89647 89808
0 25334 5 1 1 91269
0 25335 7 1 2 89744 25334
0 25336 5 4 1 25335
0 25337 7 1 2 58529 91272
0 25338 5 1 1 25337
0 25339 7 3 2 61620 77800
0 25340 5 1 1 91276
0 25341 7 1 2 90175 91277
0 25342 5 1 1 25341
0 25343 7 1 2 25338 25342
0 25344 5 3 1 25343
0 25345 7 3 2 61303 68840
0 25346 5 1 1 91282
0 25347 7 1 2 73118 83327
0 25348 7 1 2 91283 25347
0 25349 7 1 2 91279 25348
0 25350 5 1 1 25349
0 25351 7 1 2 25332 25350
0 25352 7 1 2 25277 25351
0 25353 5 1 1 25352
0 25354 7 1 2 67475 25353
0 25355 5 1 1 25354
0 25356 7 1 2 77427 86976
0 25357 7 2 2 78580 25356
0 25358 7 4 2 86604 72312
0 25359 7 1 2 88720 91287
0 25360 7 1 2 91285 25359
0 25361 5 1 1 25360
0 25362 7 1 2 25355 25361
0 25363 5 1 1 25362
0 25364 7 1 2 91214 25363
0 25365 5 1 1 25364
0 25366 7 1 2 90492 90831
0 25367 5 1 1 25366
0 25368 7 2 2 67526 88892
0 25369 7 2 2 91113 91291
0 25370 7 4 2 58034 63699
0 25371 7 1 2 80809 91295
0 25372 7 1 2 91293 25371
0 25373 5 1 1 25372
0 25374 7 3 2 62088 91215
0 25375 7 3 2 66593 91299
0 25376 7 1 2 71006 89053
0 25377 7 1 2 91302 25376
0 25378 5 1 1 25377
0 25379 7 1 2 25373 25378
0 25380 5 1 1 25379
0 25381 7 1 2 59578 25380
0 25382 5 1 1 25381
0 25383 7 2 2 70640 88330
0 25384 7 2 2 75526 88703
0 25385 7 1 2 90147 91307
0 25386 7 1 2 91305 25385
0 25387 5 1 1 25386
0 25388 7 3 2 67527 89023
0 25389 7 3 2 58035 62986
0 25390 7 2 2 58530 63700
0 25391 7 1 2 59822 91315
0 25392 7 1 2 91312 25391
0 25393 7 1 2 91309 25392
0 25394 5 1 1 25393
0 25395 7 1 2 25387 25394
0 25396 5 1 1 25395
0 25397 7 1 2 59579 25396
0 25398 5 1 1 25397
0 25399 7 1 2 75442 73964
0 25400 7 1 2 91296 25399
0 25401 7 1 2 91310 25400
0 25402 5 1 1 25401
0 25403 7 1 2 25398 25402
0 25404 5 1 1 25403
0 25405 7 1 2 69545 25404
0 25406 5 1 1 25405
0 25407 7 6 2 60126 61822
0 25408 7 1 2 81917 91317
0 25409 7 1 2 80898 25408
0 25410 7 1 2 89156 25409
0 25411 7 1 2 77050 25410
0 25412 5 1 1 25411
0 25413 7 1 2 25406 25412
0 25414 5 1 1 25413
0 25415 7 1 2 79888 25414
0 25416 5 1 1 25415
0 25417 7 1 2 63266 78930
0 25418 7 1 2 91297 25417
0 25419 7 1 2 91294 25418
0 25420 5 1 1 25419
0 25421 7 1 2 25416 25420
0 25422 7 1 2 25382 25421
0 25423 5 1 1 25422
0 25424 7 1 2 25367 25423
0 25425 5 1 1 25424
0 25426 7 2 2 62089 81303
0 25427 7 1 2 91323 91166
0 25428 5 1 1 25427
0 25429 7 1 2 64889 74941
0 25430 7 1 2 80170 25429
0 25431 7 2 2 63769 91024
0 25432 7 1 2 75411 91325
0 25433 7 1 2 25430 25432
0 25434 5 1 1 25433
0 25435 7 1 2 25428 25434
0 25436 5 1 1 25435
0 25437 7 4 2 79850 79552
0 25438 7 1 2 90063 91327
0 25439 7 1 2 25436 25438
0 25440 5 1 1 25439
0 25441 7 1 2 86446 90705
0 25442 5 1 1 25441
0 25443 7 1 2 62439 72988
0 25444 7 1 2 91072 25443
0 25445 5 1 1 25444
0 25446 7 1 2 1633 87735
0 25447 5 2 1 25446
0 25448 7 1 2 66238 72509
0 25449 7 1 2 91331 25448
0 25450 5 1 1 25449
0 25451 7 1 2 25445 25450
0 25452 5 1 1 25451
0 25453 7 1 2 65597 25452
0 25454 5 1 1 25453
0 25455 7 1 2 73069 79845
0 25456 5 1 1 25455
0 25457 7 1 2 62987 25456
0 25458 5 1 1 25457
0 25459 7 1 2 73119 85789
0 25460 5 1 1 25459
0 25461 7 1 2 25458 25460
0 25462 5 1 1 25461
0 25463 7 1 2 62719 25462
0 25464 5 1 1 25463
0 25465 7 1 2 74725 78683
0 25466 5 1 1 25465
0 25467 7 1 2 25464 25466
0 25468 5 1 1 25467
0 25469 7 1 2 66239 25468
0 25470 5 1 1 25469
0 25471 7 1 2 25454 25470
0 25472 5 1 1 25471
0 25473 7 1 2 89315 25472
0 25474 5 1 1 25473
0 25475 7 1 2 25442 25474
0 25476 5 1 1 25475
0 25477 7 1 2 20891 88052
0 25478 5 1 1 25477
0 25479 7 1 2 64890 25478
0 25480 5 1 1 25479
0 25481 7 1 2 19075 25480
0 25482 5 1 1 25481
0 25483 7 1 2 63701 25482
0 25484 5 1 1 25483
0 25485 7 1 2 19086 25484
0 25486 5 2 1 25485
0 25487 7 1 2 68841 91333
0 25488 7 1 2 25476 25487
0 25489 5 1 1 25488
0 25490 7 1 2 25440 25489
0 25491 7 1 2 25425 25490
0 25492 7 1 2 25365 25491
0 25493 7 1 2 25161 25492
0 25494 7 1 2 24961 25493
0 25495 7 1 2 24485 25494
0 25496 7 2 2 87182 86578
0 25497 7 1 2 76488 91335
0 25498 5 1 1 25497
0 25499 7 3 2 62440 85149
0 25500 5 2 1 91337
0 25501 7 1 2 75272 82876
0 25502 5 1 1 25501
0 25503 7 1 2 89827 25502
0 25504 5 1 1 25503
0 25505 7 1 2 71415 25504
0 25506 5 1 1 25505
0 25507 7 1 2 68842 89832
0 25508 5 1 1 25507
0 25509 7 1 2 87302 25508
0 25510 7 1 2 25506 25509
0 25511 5 1 1 25510
0 25512 7 1 2 91338 25511
0 25513 5 1 1 25512
0 25514 7 1 2 25498 25513
0 25515 5 1 1 25514
0 25516 7 1 2 62720 25515
0 25517 5 1 1 25516
0 25518 7 1 2 75527 90131
0 25519 5 1 1 25518
0 25520 7 1 2 25517 25519
0 25521 5 1 1 25520
0 25522 7 1 2 64069 25521
0 25523 5 1 1 25522
0 25524 7 1 2 62988 89833
0 25525 5 1 1 25524
0 25526 7 2 2 79163 84179
0 25527 5 1 1 91342
0 25528 7 1 2 25525 25527
0 25529 5 1 1 25528
0 25530 7 2 2 63267 68843
0 25531 7 1 2 25529 91344
0 25532 5 2 1 25531
0 25533 7 1 2 86862 79447
0 25534 5 1 1 25533
0 25535 7 1 2 91346 25534
0 25536 5 1 1 25535
0 25537 7 1 2 62441 25536
0 25538 5 1 1 25537
0 25539 7 1 2 25523 25538
0 25540 5 1 1 25539
0 25541 7 1 2 60940 25540
0 25542 5 1 1 25541
0 25543 7 1 2 80931 85327
0 25544 5 1 1 25543
0 25545 7 1 2 91170 25544
0 25546 5 1 1 25545
0 25547 7 1 2 90234 25546
0 25548 5 1 1 25547
0 25549 7 1 2 85328 82686
0 25550 5 1 1 25549
0 25551 7 1 2 65598 68844
0 25552 7 1 2 87351 25551
0 25553 5 1 1 25552
0 25554 7 1 2 25550 25553
0 25555 5 1 1 25554
0 25556 7 1 2 62989 25555
0 25557 5 1 1 25556
0 25558 7 1 2 25557 91347
0 25559 5 1 1 25558
0 25560 7 1 2 62442 25559
0 25561 5 1 1 25560
0 25562 7 1 2 25548 25561
0 25563 5 1 1 25562
0 25564 7 1 2 68088 25563
0 25565 5 1 1 25564
0 25566 7 1 2 66240 82920
0 25567 7 1 2 74838 25566
0 25568 5 1 1 25567
0 25569 7 2 2 59580 81502
0 25570 5 1 1 91348
0 25571 7 1 2 72780 91349
0 25572 5 1 1 25571
0 25573 7 1 2 25568 25572
0 25574 5 1 1 25573
0 25575 7 1 2 62721 25574
0 25576 5 1 1 25575
0 25577 7 1 2 87806 25576
0 25578 5 1 1 25577
0 25579 7 1 2 64534 25578
0 25580 5 1 1 25579
0 25581 7 1 2 25565 25580
0 25582 7 1 2 25542 25581
0 25583 5 1 1 25582
0 25584 7 1 2 89844 25583
0 25585 5 1 1 25584
0 25586 7 1 2 60196 25585
0 25587 5 1 1 25586
0 25588 7 1 2 90602 90687
0 25589 5 1 1 25588
0 25590 7 4 2 63770 66454
0 25591 7 1 2 62090 75398
0 25592 7 1 2 91350 25591
0 25593 7 1 2 89284 25592
0 25594 5 1 1 25593
0 25595 7 1 2 25589 25594
0 25596 5 1 1 25595
0 25597 7 1 2 62194 25596
0 25598 5 1 1 25597
0 25599 7 2 2 66704 75528
0 25600 7 1 2 69031 88721
0 25601 7 1 2 91354 25600
0 25602 5 1 1 25601
0 25603 7 1 2 76641 90699
0 25604 5 1 1 25603
0 25605 7 1 2 25602 25604
0 25606 5 1 1 25605
0 25607 7 1 2 64319 25606
0 25608 5 1 1 25607
0 25609 7 1 2 25598 25608
0 25610 5 1 1 25609
0 25611 7 1 2 65599 25610
0 25612 5 1 1 25611
0 25613 7 3 2 65045 67476
0 25614 7 1 2 73120 89006
0 25615 7 1 2 91356 25614
0 25616 5 1 1 25615
0 25617 7 1 2 25612 25616
0 25618 5 1 1 25617
0 25619 7 1 2 62990 25618
0 25620 5 1 1 25619
0 25621 7 1 2 87810 71360
0 25622 7 1 2 91265 25621
0 25623 5 1 1 25622
0 25624 7 1 2 25620 25623
0 25625 5 1 1 25624
0 25626 7 1 2 62443 25625
0 25627 5 1 1 25626
0 25628 7 1 2 68500 79703
0 25629 7 4 2 63268 89809
0 25630 5 1 1 91359
0 25631 7 1 2 90688 91360
0 25632 7 1 2 25628 25631
0 25633 5 1 1 25632
0 25634 7 1 2 25627 25633
0 25635 5 1 1 25634
0 25636 7 1 2 62722 25635
0 25637 5 1 1 25636
0 25638 7 1 2 80213 89316
0 25639 7 1 2 90019 25638
0 25640 5 1 1 25639
0 25641 7 1 2 25637 25640
0 25642 5 1 1 25641
0 25643 7 1 2 66241 25642
0 25644 5 1 1 25643
0 25645 7 3 2 59823 79218
0 25646 7 1 2 82864 89317
0 25647 7 1 2 91363 25646
0 25648 5 1 1 25647
0 25649 7 2 2 63269 90689
0 25650 7 5 2 63771 64535
0 25651 5 1 1 91368
0 25652 7 6 2 62195 91369
0 25653 5 1 1 91373
0 25654 7 1 2 84057 91374
0 25655 7 1 2 91366 25654
0 25656 5 1 1 25655
0 25657 7 1 2 25648 25656
0 25658 5 1 1 25657
0 25659 7 1 2 78789 25658
0 25660 5 1 1 25659
0 25661 7 1 2 64891 25660
0 25662 7 1 2 25644 25661
0 25663 5 1 1 25662
0 25664 7 1 2 65935 25663
0 25665 7 1 2 25587 25664
0 25666 5 1 1 25665
0 25667 7 2 2 81871 89024
0 25668 7 3 2 66594 91379
0 25669 5 1 1 91381
0 25670 7 1 2 64070 91382
0 25671 5 1 1 25670
0 25672 7 1 2 68501 88241
0 25673 7 1 2 90343 25672
0 25674 5 1 1 25673
0 25675 7 1 2 25671 25674
0 25676 5 1 1 25675
0 25677 7 1 2 60365 25676
0 25678 5 1 1 25677
0 25679 7 2 2 60366 88242
0 25680 7 1 2 90344 91384
0 25681 5 1 1 25680
0 25682 7 1 2 62723 91383
0 25683 5 1 1 25682
0 25684 7 1 2 25681 25683
0 25685 5 1 1 25684
0 25686 7 1 2 62444 25685
0 25687 5 1 1 25686
0 25688 7 1 2 25678 25687
0 25689 5 1 1 25688
0 25690 7 1 2 58531 25689
0 25691 5 1 1 25690
0 25692 7 2 2 81114 88769
0 25693 7 2 2 68845 77464
0 25694 5 1 1 91388
0 25695 7 1 2 59368 25694
0 25696 5 1 1 25695
0 25697 7 3 2 88628 25696
0 25698 5 1 1 91390
0 25699 7 1 2 69742 91391
0 25700 5 1 1 25699
0 25701 7 1 2 58036 3666
0 25702 5 1 1 25701
0 25703 7 1 2 71007 25702
0 25704 7 1 2 89943 25703
0 25705 5 1 1 25704
0 25706 7 1 2 25700 25705
0 25707 5 1 1 25706
0 25708 7 1 2 91386 25707
0 25709 5 1 1 25708
0 25710 7 1 2 25691 25709
0 25711 5 1 1 25710
0 25712 7 1 2 59824 25711
0 25713 5 1 1 25712
0 25714 7 1 2 75529 90152
0 25715 5 1 1 25714
0 25716 7 2 2 63270 85099
0 25717 7 2 2 89648 91393
0 25718 7 1 2 60941 91395
0 25719 5 1 1 25718
0 25720 7 1 2 64320 91245
0 25721 5 1 1 25720
0 25722 7 1 2 25719 25721
0 25723 5 1 1 25722
0 25724 7 3 2 68846 76675
0 25725 7 1 2 78646 91397
0 25726 7 1 2 25723 25725
0 25727 5 1 1 25726
0 25728 7 1 2 25715 25727
0 25729 5 1 1 25728
0 25730 7 1 2 62724 25729
0 25731 5 1 1 25730
0 25732 7 3 2 61823 82525
0 25733 7 1 2 83912 91400
0 25734 7 1 2 91398 25733
0 25735 5 1 1 25734
0 25736 7 1 2 25731 25735
0 25737 5 1 1 25736
0 25738 7 1 2 62445 25737
0 25739 5 1 1 25738
0 25740 7 1 2 65600 90164
0 25741 5 1 1 25740
0 25742 7 1 2 90153 25741
0 25743 5 1 1 25742
0 25744 7 1 2 91252 25743
0 25745 5 1 1 25744
0 25746 7 1 2 75530 25745
0 25747 5 1 1 25746
0 25748 7 1 2 25739 25747
0 25749 5 1 1 25748
0 25750 7 1 2 90387 25749
0 25751 5 1 1 25750
0 25752 7 1 2 25713 25751
0 25753 5 1 1 25752
0 25754 7 1 2 62991 25753
0 25755 5 1 1 25754
0 25756 7 1 2 87897 89969
0 25757 7 1 2 81829 25756
0 25758 5 1 1 25757
0 25759 7 2 2 75531 90388
0 25760 7 1 2 77985 91403
0 25761 7 1 2 91234 25760
0 25762 5 1 1 25761
0 25763 7 1 2 25758 25762
0 25764 5 1 1 25763
0 25765 7 1 2 66455 25764
0 25766 5 1 1 25765
0 25767 7 2 2 61621 75443
0 25768 5 2 1 91405
0 25769 7 6 2 59825 61943
0 25770 7 1 2 74984 88770
0 25771 7 1 2 91409 25770
0 25772 7 1 2 91406 25771
0 25773 5 1 1 25772
0 25774 7 1 2 25766 25773
0 25775 5 1 1 25774
0 25776 7 1 2 64071 25775
0 25777 5 1 1 25776
0 25778 7 1 2 88214 90629
0 25779 7 1 2 89285 25778
0 25780 5 1 1 25779
0 25781 7 5 2 61944 78852
0 25782 7 3 2 64536 61824
0 25783 7 1 2 90864 91420
0 25784 7 1 2 91415 25783
0 25785 5 1 1 25784
0 25786 7 1 2 25780 25785
0 25787 5 1 1 25786
0 25788 7 1 2 82526 25787
0 25789 5 1 1 25788
0 25790 7 1 2 25777 25789
0 25791 5 1 1 25790
0 25792 7 1 2 62446 25791
0 25793 5 1 1 25792
0 25794 7 3 2 61945 89588
0 25795 7 1 2 73720 90865
0 25796 7 1 2 91423 25795
0 25797 5 1 1 25796
0 25798 7 1 2 86083 91387
0 25799 5 1 1 25798
0 25800 7 1 2 25669 25799
0 25801 5 1 1 25800
0 25802 7 1 2 76642 75399
0 25803 7 1 2 25801 25802
0 25804 5 1 1 25803
0 25805 7 1 2 25797 25804
0 25806 5 1 1 25805
0 25807 7 1 2 60942 25806
0 25808 5 1 1 25807
0 25809 7 1 2 25793 25808
0 25810 5 1 1 25809
0 25811 7 1 2 62725 25810
0 25812 5 1 1 25811
0 25813 7 1 2 74130 91261
0 25814 5 1 1 25813
0 25815 7 1 2 78006 1243
0 25816 7 1 2 82202 25815
0 25817 7 1 2 25814 25816
0 25818 5 1 1 25817
0 25819 7 3 2 59826 81503
0 25820 7 1 2 64321 91426
0 25821 5 1 1 25820
0 25822 7 1 2 25818 25821
0 25823 5 1 1 25822
0 25824 7 1 2 88722 90866
0 25825 7 1 2 25823 25824
0 25826 5 1 1 25825
0 25827 7 1 2 25812 25826
0 25828 7 1 2 25755 25827
0 25829 5 1 1 25828
0 25830 7 1 2 62091 25829
0 25831 5 1 1 25830
0 25832 7 1 2 84242 90154
0 25833 5 1 1 25832
0 25834 7 1 2 86938 91246
0 25835 5 1 1 25834
0 25836 7 1 2 25833 25835
0 25837 5 1 1 25836
0 25838 7 1 2 68847 25837
0 25839 5 1 1 25838
0 25840 7 3 2 60943 70641
0 25841 5 2 1 91429
0 25842 7 1 2 60367 90155
0 25843 7 1 2 91430 25842
0 25844 5 1 1 25843
0 25845 7 1 2 25839 25844
0 25846 5 1 1 25845
0 25847 7 1 2 75532 25846
0 25848 5 1 1 25847
0 25849 7 2 2 77986 85337
0 25850 5 1 1 91434
0 25851 7 1 2 78116 89879
0 25852 7 1 2 91435 25851
0 25853 5 1 1 25852
0 25854 7 1 2 25848 25853
0 25855 5 1 1 25854
0 25856 7 1 2 88359 90150
0 25857 7 1 2 25855 25856
0 25858 5 1 1 25857
0 25859 7 1 2 25831 25858
0 25860 5 1 1 25859
0 25861 7 1 2 61304 25860
0 25862 5 1 1 25861
0 25863 7 1 2 67957 88992
0 25864 7 1 2 79226 25863
0 25865 7 2 2 85109 81668
0 25866 7 1 2 90156 91436
0 25867 7 1 2 25864 25866
0 25868 5 1 1 25867
0 25869 7 1 2 25862 25868
0 25870 7 1 2 25666 25869
0 25871 5 1 1 25870
0 25872 7 1 2 63702 25871
0 25873 5 1 1 25872
0 25874 7 2 2 61305 71682
0 25875 5 2 1 91438
0 25876 7 1 2 88070 24539
0 25877 5 2 1 25876
0 25878 7 1 2 62196 91442
0 25879 5 1 1 25878
0 25880 7 1 2 91440 25879
0 25881 5 1 1 25880
0 25882 7 1 2 78044 25881
0 25883 5 1 1 25882
0 25884 7 1 2 86266 25883
0 25885 5 1 1 25884
0 25886 7 1 2 62447 25885
0 25887 5 1 1 25886
0 25888 7 1 2 72864 79999
0 25889 5 2 1 25888
0 25890 7 1 2 25887 91444
0 25891 5 1 1 25890
0 25892 7 1 2 62726 25891
0 25893 5 1 1 25892
0 25894 7 1 2 18631 25893
0 25895 5 1 1 25894
0 25896 7 1 2 91396 25895
0 25897 5 1 1 25896
0 25898 7 1 2 82221 89525
0 25899 5 1 1 25898
0 25900 7 1 2 82921 25899
0 25901 5 1 1 25900
0 25902 7 2 2 68502 90330
0 25903 7 1 2 80785 91446
0 25904 5 1 1 25903
0 25905 7 1 2 87183 91009
0 25906 5 1 1 25905
0 25907 7 1 2 25904 25906
0 25908 5 1 1 25907
0 25909 7 1 2 62727 25908
0 25910 5 1 1 25909
0 25911 7 1 2 25901 25910
0 25912 5 1 1 25911
0 25913 7 1 2 61306 25912
0 25914 5 1 1 25913
0 25915 7 4 2 64537 86477
0 25916 7 1 2 62992 86905
0 25917 7 1 2 91448 25916
0 25918 5 1 1 25917
0 25919 7 1 2 65601 25918
0 25920 7 1 2 25914 25919
0 25921 5 1 1 25920
0 25922 7 1 2 85996 87310
0 25923 5 1 1 25922
0 25924 7 4 2 58532 73510
0 25925 5 1 1 91452
0 25926 7 1 2 79219 91453
0 25927 5 1 1 25926
0 25928 7 1 2 25923 25927
0 25929 5 1 1 25928
0 25930 7 1 2 61622 25929
0 25931 5 1 1 25930
0 25932 7 4 2 62448 65936
0 25933 7 3 2 66242 68848
0 25934 7 1 2 91456 91460
0 25935 7 1 2 80992 25934
0 25936 5 1 1 25935
0 25937 7 1 2 25931 25936
0 25938 5 1 1 25937
0 25939 7 1 2 60368 25938
0 25940 5 1 1 25939
0 25941 7 1 2 59581 87453
0 25942 5 1 1 25941
0 25943 7 1 2 15912 25942
0 25944 5 1 1 25943
0 25945 7 1 2 68089 25944
0 25946 5 1 1 25945
0 25947 7 3 2 64072 66243
0 25948 7 1 2 85424 77555
0 25949 5 1 1 25948
0 25950 7 1 2 85434 25949
0 25951 5 1 1 25950
0 25952 7 1 2 91463 25951
0 25953 5 1 1 25952
0 25954 7 3 2 62449 76203
0 25955 7 1 2 68849 82555
0 25956 7 1 2 91466 25955
0 25957 5 1 1 25956
0 25958 7 1 2 25953 25957
0 25959 5 1 1 25958
0 25960 7 1 2 65937 25959
0 25961 5 1 1 25960
0 25962 7 1 2 25946 25961
0 25963 5 1 1 25962
0 25964 7 1 2 63271 25963
0 25965 5 1 1 25964
0 25966 7 1 2 62197 82203
0 25967 5 1 1 25966
0 25968 7 1 2 82592 25967
0 25969 5 2 1 25968
0 25970 7 5 2 62198 61623
0 25971 5 1 1 91471
0 25972 7 1 2 58977 25971
0 25973 5 1 1 25972
0 25974 7 1 2 79295 91083
0 25975 7 1 2 25973 25974
0 25976 7 1 2 91469 25975
0 25977 5 1 1 25976
0 25978 7 1 2 60944 25977
0 25979 7 1 2 25965 25978
0 25980 7 1 2 25940 25979
0 25981 5 1 1 25980
0 25982 7 1 2 25921 25981
0 25983 5 1 1 25982
0 25984 7 1 2 71029 82838
0 25985 5 1 1 25984
0 25986 7 1 2 71497 25985
0 25987 5 1 1 25986
0 25988 7 2 2 66244 25987
0 25989 7 1 2 90424 91476
0 25990 5 1 1 25989
0 25991 7 1 2 59827 85988
0 25992 5 1 1 25991
0 25993 7 2 2 90367 25992
0 25994 7 2 2 75774 84180
0 25995 7 1 2 91478 91480
0 25996 5 1 1 25995
0 25997 7 1 2 59828 90365
0 25998 5 1 1 25997
0 25999 7 1 2 64538 73690
0 26000 5 6 1 25999
0 26001 7 1 2 61624 79990
0 26002 7 1 2 91482 26001
0 26003 7 1 2 78347 26002
0 26004 7 1 2 25998 26003
0 26005 5 1 1 26004
0 26006 7 1 2 25996 26005
0 26007 5 1 1 26006
0 26008 7 1 2 62993 26007
0 26009 5 1 1 26008
0 26010 7 2 2 75775 88557
0 26011 5 1 1 91488
0 26012 7 1 2 90412 91489
0 26013 5 1 1 26012
0 26014 7 1 2 26009 26013
0 26015 5 1 1 26014
0 26016 7 1 2 68090 26015
0 26017 5 1 1 26016
0 26018 7 1 2 25990 26017
0 26019 7 1 2 25983 26018
0 26020 5 1 1 26019
0 26021 7 1 2 61825 26020
0 26022 5 1 1 26021
0 26023 7 1 2 25897 26022
0 26024 5 1 1 26023
0 26025 7 1 2 89011 26024
0 26026 5 1 1 26025
0 26027 7 3 2 68503 86478
0 26028 7 1 2 78790 91490
0 26029 5 1 1 26028
0 26030 7 3 2 62728 77730
0 26031 5 1 1 91493
0 26032 7 1 2 90833 91494
0 26033 5 1 1 26032
0 26034 7 1 2 26029 26033
0 26035 5 1 1 26034
0 26036 7 1 2 64322 26035
0 26037 5 1 1 26036
0 26038 7 3 2 60945 86479
0 26039 7 1 2 65046 79677
0 26040 7 1 2 91496 26039
0 26041 5 1 1 26040
0 26042 7 1 2 26037 26041
0 26043 5 1 1 26042
0 26044 7 1 2 90693 26043
0 26045 5 1 1 26044
0 26046 7 1 2 75153 81994
0 26047 5 1 1 26046
0 26048 7 1 2 62450 26047
0 26049 5 1 1 26048
0 26050 7 1 2 7004 81995
0 26051 5 1 1 26050
0 26052 7 1 2 68850 26051
0 26053 5 1 1 26052
0 26054 7 1 2 26049 26053
0 26055 5 1 1 26054
0 26056 7 1 2 90680 26055
0 26057 5 1 1 26056
0 26058 7 1 2 58292 78791
0 26059 5 1 1 26058
0 26060 7 1 2 65047 71091
0 26061 5 1 1 26060
0 26062 7 1 2 26059 26061
0 26063 5 1 1 26062
0 26064 7 1 2 75722 90701
0 26065 7 1 2 26063 26064
0 26066 5 1 1 26065
0 26067 7 1 2 77428 83490
0 26068 7 1 2 90706 26067
0 26069 5 1 1 26068
0 26070 7 1 2 26066 26069
0 26071 7 1 2 26057 26070
0 26072 5 1 1 26071
0 26073 7 1 2 59582 26072
0 26074 5 1 1 26073
0 26075 7 1 2 26045 26074
0 26076 5 1 1 26075
0 26077 7 1 2 88125 26076
0 26078 5 1 1 26077
0 26079 7 1 2 85408 86589
0 26080 5 1 1 26079
0 26081 7 1 2 90908 26080
0 26082 5 1 1 26081
0 26083 7 1 2 70642 26082
0 26084 5 1 1 26083
0 26085 7 1 2 68504 90901
0 26086 5 1 1 26085
0 26087 7 1 2 26084 26086
0 26088 5 1 1 26087
0 26089 7 1 2 60369 26088
0 26090 5 1 1 26089
0 26091 7 1 2 68851 90726
0 26092 5 1 1 26091
0 26093 7 1 2 58293 26092
0 26094 5 1 1 26093
0 26095 7 1 2 85726 26094
0 26096 5 1 1 26095
0 26097 7 1 2 68005 75784
0 26098 5 1 1 26097
0 26099 7 1 2 90247 26098
0 26100 5 1 1 26099
0 26101 7 1 2 61625 85415
0 26102 7 1 2 26100 26101
0 26103 7 1 2 26096 26102
0 26104 7 1 2 26090 26103
0 26105 5 1 1 26104
0 26106 7 2 2 68091 80426
0 26107 5 1 1 91499
0 26108 7 1 2 71416 91500
0 26109 5 2 1 26108
0 26110 7 1 2 66245 91501
0 26111 5 1 1 26110
0 26112 7 2 2 62092 88140
0 26113 7 1 2 88723 91503
0 26114 7 1 2 26111 26113
0 26115 7 1 2 26105 26114
0 26116 5 1 1 26115
0 26117 7 1 2 26078 26116
0 26118 5 1 1 26117
0 26119 7 1 2 77869 88317
0 26120 7 1 2 26118 26119
0 26121 5 1 1 26120
0 26122 7 1 2 26026 26121
0 26123 7 1 2 25873 26122
0 26124 5 1 1 26123
0 26125 7 1 2 79889 26124
0 26126 5 1 1 26125
0 26127 7 1 2 91306 91324
0 26128 5 1 1 26127
0 26129 7 2 2 64073 74942
0 26130 5 1 1 91505
0 26131 7 1 2 74950 91506
0 26132 7 1 2 88585 26131
0 26133 5 1 1 26132
0 26134 7 1 2 26128 26133
0 26135 5 1 1 26134
0 26136 7 1 2 89987 90951
0 26137 7 1 2 26135 26136
0 26138 5 1 1 26137
0 26139 7 1 2 26126 26138
0 26140 5 1 1 26139
0 26141 7 1 2 70508 26140
0 26142 5 1 1 26141
0 26143 7 1 2 68777 84248
0 26144 5 2 1 26143
0 26145 7 1 2 66246 70206
0 26146 7 1 2 67477 26145
0 26147 7 4 2 91507 26146
0 26148 7 2 2 88662 91509
0 26149 7 1 2 88209 91513
0 26150 5 1 1 26149
0 26151 7 2 2 87856 87922
0 26152 5 1 1 91515
0 26153 7 1 2 91514 91516
0 26154 5 1 1 26153
0 26155 7 3 2 60127 74293
0 26156 5 1 1 91517
0 26157 7 1 2 60946 88960
0 26158 5 1 1 26157
0 26159 7 1 2 26156 26158
0 26160 5 1 1 26159
0 26161 7 1 2 64074 26160
0 26162 5 1 1 26161
0 26163 7 2 2 71997 66971
0 26164 5 1 1 91520
0 26165 7 1 2 83903 91521
0 26166 5 1 1 26165
0 26167 7 1 2 65048 68940
0 26168 5 1 1 26167
0 26169 7 1 2 26166 26168
0 26170 7 1 2 26162 26169
0 26171 5 1 1 26170
0 26172 7 1 2 62451 26171
0 26173 5 1 1 26172
0 26174 7 1 2 64075 83491
0 26175 5 1 1 26174
0 26176 7 2 2 88634 26175
0 26177 5 1 1 91522
0 26178 7 1 2 67049 26177
0 26179 5 1 1 26178
0 26180 7 1 2 26173 26179
0 26181 5 1 1 26180
0 26182 7 1 2 63622 26181
0 26183 5 1 1 26182
0 26184 7 3 2 61946 70454
0 26185 7 1 2 62452 78792
0 26186 5 1 1 26185
0 26187 7 1 2 91523 26186
0 26188 5 1 1 26187
0 26189 7 1 2 91524 26188
0 26190 5 1 1 26189
0 26191 7 1 2 26183 26190
0 26192 5 1 1 26191
0 26193 7 1 2 88008 26192
0 26194 5 1 1 26193
0 26195 7 3 2 66247 70509
0 26196 7 2 2 84873 85100
0 26197 7 1 2 74294 91530
0 26198 7 1 2 91527 26197
0 26199 5 1 1 26198
0 26200 7 1 2 26194 26199
0 26201 5 1 1 26200
0 26202 7 1 2 61826 26201
0 26203 5 1 1 26202
0 26204 7 2 2 77465 91416
0 26205 7 1 2 88984 89994
0 26206 7 1 2 91532 26205
0 26207 5 1 1 26206
0 26208 7 1 2 26203 26207
0 26209 5 1 1 26208
0 26210 7 1 2 66705 26209
0 26211 5 1 1 26210
0 26212 7 1 2 70510 89007
0 26213 7 1 2 91510 26212
0 26214 5 1 1 26213
0 26215 7 1 2 26211 26214
0 26216 5 1 1 26215
0 26217 7 1 2 66904 26216
0 26218 5 1 1 26217
0 26219 7 1 2 85380 91511
0 26220 5 1 1 26219
0 26221 7 2 2 70643 88009
0 26222 5 1 1 91534
0 26223 7 1 2 26011 26222
0 26224 5 1 1 26223
0 26225 7 1 2 60370 26224
0 26226 5 1 1 26225
0 26227 7 1 2 84454 87300
0 26228 5 1 1 26227
0 26229 7 1 2 26226 26228
0 26230 5 1 1 26229
0 26231 7 1 2 65602 67528
0 26232 7 2 2 26230 26231
0 26233 7 1 2 79922 91536
0 26234 5 1 1 26233
0 26235 7 1 2 26220 26234
0 26236 5 1 1 26235
0 26237 7 1 2 66456 26236
0 26238 5 1 1 26237
0 26239 7 1 2 79920 90690
0 26240 7 2 2 58533 85338
0 26241 7 3 2 64707 82527
0 26242 7 1 2 91538 91540
0 26243 7 1 2 26239 26242
0 26244 5 1 1 26243
0 26245 7 1 2 26238 26244
0 26246 5 1 1 26245
0 26247 7 1 2 70511 26246
0 26248 5 1 1 26247
0 26249 7 1 2 88060 91512
0 26250 5 1 1 26249
0 26251 7 1 2 62729 82066
0 26252 7 1 2 91537 26251
0 26253 5 1 1 26252
0 26254 7 1 2 26250 26253
0 26255 5 1 1 26254
0 26256 7 1 2 66457 26255
0 26257 5 1 1 26256
0 26258 7 1 2 80459 90084
0 26259 7 1 2 91247 26258
0 26260 7 1 2 83153 26259
0 26261 5 1 1 26260
0 26262 7 1 2 26257 26261
0 26263 7 1 2 26248 26262
0 26264 7 1 2 26218 26263
0 26265 5 1 1 26264
0 26266 7 1 2 64892 26265
0 26267 5 1 1 26266
0 26268 7 1 2 26154 26267
0 26269 5 1 1 26268
0 26270 7 1 2 63703 26269
0 26271 5 1 1 26270
0 26272 7 1 2 26150 26271
0 26273 5 1 1 26272
0 26274 7 1 2 61307 26273
0 26275 5 1 1 26274
0 26276 7 1 2 68505 69546
0 26277 7 1 2 89976 26276
0 26278 7 1 2 87871 26277
0 26279 5 1 1 26278
0 26280 7 1 2 89898 91417
0 26281 7 1 2 88110 26280
0 26282 5 1 1 26281
0 26283 7 1 2 26279 26282
0 26284 5 1 1 26283
0 26285 7 1 2 82123 26284
0 26286 5 1 1 26285
0 26287 7 2 2 82408 88914
0 26288 5 1 1 91543
0 26289 7 1 2 77359 90617
0 26290 5 1 1 26289
0 26291 7 1 2 26288 26290
0 26292 5 1 1 26291
0 26293 7 1 2 63272 26292
0 26294 5 1 1 26293
0 26295 7 1 2 77819 89608
0 26296 5 1 1 26295
0 26297 7 1 2 26294 26296
0 26298 5 1 1 26297
0 26299 7 1 2 79890 26298
0 26300 5 1 1 26299
0 26301 7 3 2 65049 79823
0 26302 7 1 2 76921 90722
0 26303 7 1 2 91545 26302
0 26304 5 1 1 26303
0 26305 7 1 2 26300 26304
0 26306 5 1 1 26305
0 26307 7 1 2 81069 69547
0 26308 7 1 2 26306 26307
0 26309 5 1 1 26308
0 26310 7 1 2 26286 26309
0 26311 5 1 1 26310
0 26312 7 1 2 90137 91102
0 26313 7 1 2 26311 26312
0 26314 5 1 1 26313
0 26315 7 1 2 26275 26314
0 26316 5 1 1 26315
0 26317 7 1 2 87933 26316
0 26318 5 1 1 26317
0 26319 7 1 2 26142 26318
0 26320 7 1 2 25495 26319
0 26321 7 1 2 67201 79053
0 26322 5 1 1 26321
0 26323 7 1 2 70409 26322
0 26324 5 1 1 26323
0 26325 7 1 2 62453 26324
0 26326 5 1 1 26325
0 26327 7 1 2 15763 26326
0 26328 5 1 1 26327
0 26329 7 1 2 88596 26328
0 26330 5 1 1 26329
0 26331 7 3 2 70014 83461
0 26332 7 1 2 63704 90915
0 26333 7 1 2 91548 26332
0 26334 5 1 1 26333
0 26335 7 1 2 26330 26334
0 26336 5 1 1 26335
0 26337 7 2 2 77987 84665
0 26338 5 1 1 91551
0 26339 7 1 2 26336 91552
0 26340 5 1 1 26339
0 26341 7 1 2 84500 90522
0 26342 5 1 1 26341
0 26343 7 1 2 70644 88360
0 26344 7 1 2 74674 26343
0 26345 5 1 1 26344
0 26346 7 1 2 26342 26345
0 26347 5 1 1 26346
0 26348 7 1 2 62730 26347
0 26349 5 1 1 26348
0 26350 7 1 2 71280 90851
0 26351 5 1 1 26350
0 26352 7 1 2 26349 26351
0 26353 5 1 1 26352
0 26354 7 1 2 60371 26353
0 26355 5 1 1 26354
0 26356 7 1 2 65938 81163
0 26357 5 1 1 26356
0 26358 7 1 2 72899 89132
0 26359 7 1 2 26357 26358
0 26360 5 1 1 26359
0 26361 7 1 2 26355 26360
0 26362 5 1 1 26361
0 26363 7 1 2 63705 26362
0 26364 5 1 1 26363
0 26365 7 2 2 70924 83276
0 26366 5 1 1 91553
0 26367 7 2 2 65939 16186
0 26368 5 1 1 91555
0 26369 7 1 2 81164 91556
0 26370 7 1 2 26366 26369
0 26371 5 1 1 26370
0 26372 7 1 2 72900 89103
0 26373 7 1 2 26371 26372
0 26374 5 1 1 26373
0 26375 7 1 2 26364 26374
0 26376 5 1 1 26375
0 26377 7 1 2 64076 26376
0 26378 5 1 1 26377
0 26379 7 3 2 68506 79492
0 26380 5 1 1 91557
0 26381 7 1 2 82841 26380
0 26382 5 1 1 26381
0 26383 7 1 2 88597 91457
0 26384 7 1 2 26382 26383
0 26385 5 1 1 26384
0 26386 7 1 2 26378 26385
0 26387 5 1 1 26386
0 26388 7 1 2 60947 26387
0 26389 5 1 1 26388
0 26390 7 1 2 80932 73011
0 26391 5 1 1 26390
0 26392 7 1 2 91191 26391
0 26393 5 1 1 26392
0 26394 7 1 2 62731 26393
0 26395 5 1 1 26394
0 26396 7 1 2 90893 26395
0 26397 5 1 1 26396
0 26398 7 1 2 88598 26397
0 26399 5 1 1 26398
0 26400 7 3 2 73012 75144
0 26401 5 1 1 91560
0 26402 7 2 2 68092 68507
0 26403 7 1 2 88371 91563
0 26404 7 1 2 91561 26403
0 26405 5 1 1 26404
0 26406 7 1 2 26399 26405
0 26407 5 1 1 26406
0 26408 7 1 2 62454 26407
0 26409 5 1 1 26408
0 26410 7 1 2 71417 86121
0 26411 7 1 2 88599 26410
0 26412 5 1 1 26411
0 26413 7 1 2 26409 26412
0 26414 7 1 2 26389 26413
0 26415 5 1 1 26414
0 26416 7 1 2 61626 26415
0 26417 5 1 1 26416
0 26418 7 1 2 26340 26417
0 26419 5 1 1 26418
0 26420 7 1 2 76741 26419
0 26421 5 1 1 26420
0 26422 7 1 2 88941 89693
0 26423 5 1 1 26422
0 26424 7 1 2 60372 90827
0 26425 5 1 1 26424
0 26426 7 1 2 26423 26425
0 26427 5 1 1 26426
0 26428 7 1 2 59583 26427
0 26429 5 1 1 26428
0 26430 7 1 2 68508 91193
0 26431 5 1 1 26430
0 26432 7 1 2 62455 86210
0 26433 5 1 1 26432
0 26434 7 1 2 26431 26433
0 26435 5 1 1 26434
0 26436 7 1 2 71281 26435
0 26437 5 1 1 26436
0 26438 7 1 2 71418 84501
0 26439 5 1 1 26438
0 26440 7 1 2 26437 26439
0 26441 5 1 1 26440
0 26442 7 1 2 66248 26441
0 26443 5 1 1 26442
0 26444 7 1 2 26429 26443
0 26445 5 1 1 26444
0 26446 7 1 2 64539 26445
0 26447 5 1 1 26446
0 26448 7 1 2 76489 91364
0 26449 7 1 2 91497 26448
0 26450 5 1 1 26449
0 26451 7 1 2 26447 26450
0 26452 5 1 1 26451
0 26453 7 1 2 63273 26452
0 26454 5 1 1 26453
0 26455 7 1 2 77587 84795
0 26456 7 1 2 90459 26455
0 26457 5 1 1 26456
0 26458 7 1 2 26454 26457
0 26459 5 1 1 26458
0 26460 7 1 2 88600 26459
0 26461 5 1 1 26460
0 26462 7 1 2 81669 84740
0 26463 5 2 1 26462
0 26464 7 1 2 79584 91565
0 26465 5 1 1 26464
0 26466 7 1 2 82556 26465
0 26467 5 1 1 26466
0 26468 7 2 2 79173 74985
0 26469 7 1 2 68509 91567
0 26470 5 1 1 26469
0 26471 7 1 2 79585 26470
0 26472 5 1 1 26471
0 26473 7 1 2 90592 26472
0 26474 5 1 1 26473
0 26475 7 1 2 26467 26474
0 26476 5 1 1 26475
0 26477 7 1 2 61308 26476
0 26478 5 1 1 26477
0 26479 7 1 2 76490 90095
0 26480 5 1 1 26479
0 26481 7 1 2 22126 26480
0 26482 5 1 1 26481
0 26483 7 1 2 86480 26482
0 26484 5 1 1 26483
0 26485 7 1 2 26478 26484
0 26486 5 1 1 26485
0 26487 7 1 2 62994 26486
0 26488 5 1 1 26487
0 26489 7 2 2 59829 68510
0 26490 7 1 2 87776 91569
0 26491 5 1 1 26490
0 26492 7 1 2 82877 87427
0 26493 5 1 1 26492
0 26494 7 1 2 26491 26493
0 26495 5 1 1 26494
0 26496 7 1 2 61309 26495
0 26497 5 1 1 26496
0 26498 7 1 2 26488 26497
0 26499 5 1 1 26498
0 26500 7 1 2 64077 26499
0 26501 5 1 1 26500
0 26502 7 3 2 81011 89408
0 26503 7 2 2 86122 82557
0 26504 7 1 2 91571 91574
0 26505 5 1 1 26504
0 26506 7 1 2 26501 26505
0 26507 5 1 1 26506
0 26508 7 1 2 62456 88601
0 26509 7 1 2 26507 26508
0 26510 5 1 1 26509
0 26511 7 2 2 70207 87446
0 26512 5 1 1 91576
0 26513 7 1 2 90975 91577
0 26514 5 1 1 26513
0 26515 7 1 2 62995 74986
0 26516 7 1 2 87043 26515
0 26517 7 2 2 61310 88921
0 26518 7 1 2 89166 91578
0 26519 7 1 2 26516 26518
0 26520 5 1 1 26519
0 26521 7 1 2 26514 26520
0 26522 5 1 1 26521
0 26523 7 1 2 70645 26522
0 26524 5 1 1 26523
0 26525 7 2 2 85636 88126
0 26526 7 1 2 72725 73313
0 26527 7 1 2 80810 90715
0 26528 7 1 2 26526 26527
0 26529 7 1 2 91580 26528
0 26530 5 1 1 26529
0 26531 7 1 2 26524 26530
0 26532 7 1 2 26510 26531
0 26533 5 1 1 26532
0 26534 7 1 2 62732 26533
0 26535 5 1 1 26534
0 26536 7 1 2 26461 26535
0 26537 7 1 2 26421 26536
0 26538 5 1 1 26537
0 26539 7 1 2 66458 26538
0 26540 5 1 1 26539
0 26541 7 3 2 89805 91001
0 26542 5 1 1 91582
0 26543 7 1 2 89245 26542
0 26544 5 2 1 26543
0 26545 7 1 2 74539 85835
0 26546 5 1 1 26545
0 26547 7 5 2 71282 90981
0 26548 7 1 2 65940 91587
0 26549 5 1 1 26548
0 26550 7 1 2 26546 26549
0 26551 5 1 1 26550
0 26552 7 1 2 88346 26551
0 26553 5 1 1 26552
0 26554 7 5 2 65941 88922
0 26555 7 1 2 74131 88127
0 26556 7 1 2 84395 26555
0 26557 7 1 2 91592 26556
0 26558 5 1 1 26557
0 26559 7 1 2 26553 26558
0 26560 5 1 1 26559
0 26561 7 1 2 91585 26560
0 26562 5 1 1 26561
0 26563 7 1 2 87030 77557
0 26564 5 1 1 26563
0 26565 7 1 2 87725 26564
0 26566 5 1 1 26565
0 26567 7 1 2 74839 90969
0 26568 7 1 2 90965 26567
0 26569 5 1 1 26568
0 26570 7 1 2 26566 26569
0 26571 5 1 1 26570
0 26572 7 1 2 88602 26571
0 26573 5 1 1 26572
0 26574 7 2 2 62733 87727
0 26575 5 2 1 91597
0 26576 7 1 2 87416 88372
0 26577 7 1 2 91598 26576
0 26578 7 1 2 71008 26577
0 26579 5 1 1 26578
0 26580 7 1 2 26573 26579
0 26581 5 1 1 26580
0 26582 7 1 2 66249 26581
0 26583 5 1 1 26582
0 26584 7 2 2 68511 78684
0 26585 5 3 1 91601
0 26586 7 1 2 88128 91602
0 26587 7 1 2 86289 91593
0 26588 7 1 2 26586 26587
0 26589 5 1 1 26588
0 26590 7 1 2 26583 26589
0 26591 5 1 1 26590
0 26592 7 1 2 89228 26591
0 26593 5 1 1 26592
0 26594 7 1 2 26562 26593
0 26595 7 1 2 26540 26594
0 26596 5 1 1 26595
0 26597 7 1 2 66777 26596
0 26598 5 1 1 26597
0 26599 7 2 2 71419 80670
0 26600 5 1 1 91606
0 26601 7 1 2 90938 26600
0 26602 5 1 1 26601
0 26603 7 1 2 70646 26602
0 26604 5 1 1 26603
0 26605 7 1 2 86051 77405
0 26606 5 1 1 26605
0 26607 7 1 2 26604 26606
0 26608 5 1 1 26607
0 26609 7 1 2 60373 26608
0 26610 5 1 1 26609
0 26611 7 1 2 26610 91502
0 26612 5 1 1 26611
0 26613 7 1 2 61627 88857
0 26614 7 2 2 26612 26613
0 26615 7 1 2 85381 88331
0 26616 7 1 2 91608 26615
0 26617 5 1 1 26616
0 26618 7 1 2 26598 26617
0 26619 5 1 1 26618
0 26620 7 1 2 70512 26619
0 26621 5 1 1 26620
0 26622 7 1 2 82558 75484
0 26623 7 1 2 90856 26622
0 26624 5 1 1 26623
0 26625 7 1 2 26512 26624
0 26626 5 1 1 26625
0 26627 7 1 2 62996 26626
0 26628 5 1 1 26627
0 26629 7 1 2 72941 88558
0 26630 5 1 1 26629
0 26631 7 1 2 26628 26630
0 26632 5 1 1 26631
0 26633 7 1 2 62734 26632
0 26634 5 1 1 26633
0 26635 7 1 2 87825 90882
0 26636 5 1 1 26635
0 26637 7 1 2 80838 91464
0 26638 5 1 1 26637
0 26639 7 1 2 26636 26638
0 26640 5 1 1 26639
0 26641 7 1 2 60948 26640
0 26642 5 1 1 26641
0 26643 7 1 2 26634 26642
0 26644 5 1 1 26643
0 26645 7 1 2 66459 26644
0 26646 5 1 1 26645
0 26647 7 1 2 77466 91280
0 26648 5 1 1 26647
0 26649 7 3 2 64540 89899
0 26650 7 1 2 80811 91610
0 26651 5 1 1 26650
0 26652 7 1 2 26648 26651
0 26653 5 1 1 26652
0 26654 7 1 2 81137 26653
0 26655 5 1 1 26654
0 26656 7 2 2 77467 89589
0 26657 7 1 2 73378 78502
0 26658 7 1 2 91613 26657
0 26659 5 1 1 26658
0 26660 7 1 2 26655 26659
0 26661 7 1 2 26646 26660
0 26662 5 1 1 26661
0 26663 7 1 2 89104 26662
0 26664 5 1 1 26663
0 26665 7 2 2 65603 90916
0 26666 5 1 1 91615
0 26667 7 1 2 23298 26666
0 26668 5 1 1 26667
0 26669 7 1 2 62735 26668
0 26670 5 1 1 26669
0 26671 7 1 2 64078 91616
0 26672 5 1 1 26671
0 26673 7 1 2 26670 26672
0 26674 5 1 1 26673
0 26675 7 1 2 64323 26674
0 26676 5 1 1 26675
0 26677 7 1 2 60949 73597
0 26678 7 1 2 90534 26677
0 26679 5 1 1 26678
0 26680 7 1 2 26676 26679
0 26681 5 1 1 26680
0 26682 7 1 2 58534 26681
0 26683 5 1 1 26682
0 26684 7 1 2 75023 88361
0 26685 7 1 2 82903 26684
0 26686 5 1 1 26685
0 26687 7 1 2 26683 26686
0 26688 5 1 1 26687
0 26689 7 1 2 62457 89260
0 26690 7 1 2 26688 26689
0 26691 5 1 1 26690
0 26692 7 2 2 63274 81138
0 26693 5 1 1 91617
0 26694 7 1 2 58294 26693
0 26695 5 1 1 26694
0 26696 7 2 2 90857 26695
0 26697 7 1 2 62736 91619
0 26698 5 2 1 26697
0 26699 7 1 2 87765 91621
0 26700 5 1 1 26699
0 26701 7 1 2 90176 90523
0 26702 7 1 2 26700 26701
0 26703 5 1 1 26702
0 26704 7 1 2 64079 89874
0 26705 5 1 1 26704
0 26706 7 2 2 63275 79220
0 26707 7 1 2 68093 90630
0 26708 7 1 2 91623 26707
0 26709 5 1 1 26708
0 26710 7 1 2 26705 26709
0 26711 5 1 1 26710
0 26712 7 1 2 65604 26711
0 26713 5 1 1 26712
0 26714 7 1 2 78685 89875
0 26715 5 1 1 26714
0 26716 7 1 2 26713 26715
0 26717 5 1 1 26716
0 26718 7 1 2 88362 26717
0 26719 5 1 1 26718
0 26720 7 1 2 26703 26719
0 26721 5 1 1 26720
0 26722 7 1 2 59830 26721
0 26723 5 1 1 26722
0 26724 7 1 2 61628 26723
0 26725 7 1 2 26691 26724
0 26726 5 1 1 26725
0 26727 7 2 2 70208 89083
0 26728 5 1 1 91625
0 26729 7 3 2 61827 83328
0 26730 7 1 2 73379 91627
0 26731 5 1 1 26730
0 26732 7 1 2 26728 26731
0 26733 5 1 1 26732
0 26734 7 1 2 89133 26733
0 26735 5 1 1 26734
0 26736 7 1 2 75444 71998
0 26737 7 1 2 89161 90672
0 26738 7 1 2 26736 26737
0 26739 5 1 1 26738
0 26740 7 1 2 26735 26739
0 26741 5 1 1 26740
0 26742 7 1 2 62997 26741
0 26743 5 1 1 26742
0 26744 7 1 2 81139 89461
0 26745 5 1 1 26744
0 26746 7 1 2 64324 91626
0 26747 5 1 1 26746
0 26748 7 1 2 26745 26747
0 26749 5 1 1 26748
0 26750 7 1 2 89134 26749
0 26751 5 1 1 26750
0 26752 7 1 2 26743 26751
0 26753 5 1 1 26752
0 26754 7 1 2 62737 26753
0 26755 5 1 1 26754
0 26756 7 1 2 89084 89135
0 26757 7 1 2 91588 26756
0 26758 5 1 1 26757
0 26759 7 1 2 66250 26758
0 26760 7 1 2 26755 26759
0 26761 5 1 1 26760
0 26762 7 1 2 63706 26761
0 26763 7 1 2 26726 26762
0 26764 5 1 1 26763
0 26765 7 1 2 26664 26764
0 26766 5 1 1 26765
0 26767 7 1 2 68512 26766
0 26768 5 1 1 26767
0 26769 7 1 2 75119 90906
0 26770 5 1 1 26769
0 26771 7 1 2 64893 77588
0 26772 7 1 2 76413 26771
0 26773 5 1 1 26772
0 26774 7 1 2 26770 26773
0 26775 5 1 1 26774
0 26776 7 1 2 89085 26775
0 26777 5 1 1 26776
0 26778 7 1 2 65605 78079
0 26779 7 1 2 78117 87902
0 26780 7 1 2 90673 26779
0 26781 7 1 2 26778 26780
0 26782 5 1 1 26781
0 26783 7 1 2 26777 26782
0 26784 5 1 1 26783
0 26785 7 1 2 62738 26784
0 26786 5 1 1 26785
0 26787 7 1 2 81140 89136
0 26788 7 1 2 91586 26787
0 26789 5 1 1 26788
0 26790 7 1 2 26786 26789
0 26791 5 1 1 26790
0 26792 7 1 2 63707 26791
0 26793 5 1 1 26792
0 26794 7 1 2 81141 89054
0 26795 5 1 1 26794
0 26796 7 1 2 84636 81132
0 26797 5 1 1 26796
0 26798 7 1 2 91583 26797
0 26799 5 1 1 26798
0 26800 7 1 2 26795 26799
0 26801 5 1 1 26800
0 26802 7 1 2 89105 26801
0 26803 5 1 1 26802
0 26804 7 1 2 26793 26803
0 26805 5 1 1 26804
0 26806 7 1 2 66251 26805
0 26807 5 1 1 26806
0 26808 7 2 2 77870 82687
0 26809 5 1 1 91630
0 26810 7 1 2 87811 81142
0 26811 7 1 2 88332 26810
0 26812 7 1 2 91631 26811
0 26813 5 1 1 26812
0 26814 7 1 2 26807 26813
0 26815 5 1 1 26814
0 26816 7 1 2 62998 26815
0 26817 5 1 1 26816
0 26818 7 1 2 90194 91539
0 26819 5 1 1 26818
0 26820 7 1 2 85568 87308
0 26821 5 1 1 26820
0 26822 7 1 2 60374 90840
0 26823 5 1 1 26822
0 26824 7 1 2 26821 26823
0 26825 5 1 1 26824
0 26826 7 1 2 63276 26825
0 26827 5 1 1 26826
0 26828 7 1 2 73121 85086
0 26829 7 1 2 87258 26828
0 26830 5 1 1 26829
0 26831 7 1 2 26827 26830
0 26832 5 1 1 26831
0 26833 7 1 2 66460 26832
0 26834 5 1 1 26833
0 26835 7 1 2 26819 26834
0 26836 5 1 1 26835
0 26837 7 1 2 64325 88603
0 26838 7 1 2 26836 26837
0 26839 5 1 1 26838
0 26840 7 1 2 26817 26839
0 26841 7 1 2 26768 26840
0 26842 5 1 1 26841
0 26843 7 1 2 69548 26842
0 26844 5 1 1 26843
0 26845 7 1 2 76340 77801
0 26846 5 1 1 26845
0 26847 7 1 2 67202 91199
0 26848 5 1 1 26847
0 26849 7 1 2 26846 26848
0 26850 5 1 1 26849
0 26851 7 1 2 62999 26850
0 26852 5 1 1 26851
0 26853 7 1 2 77988 76742
0 26854 5 1 1 26853
0 26855 7 1 2 26852 26854
0 26856 5 1 1 26855
0 26857 7 1 2 74840 26856
0 26858 5 1 1 26857
0 26859 7 1 2 77871 78123
0 26860 5 1 1 26859
0 26861 7 1 2 26858 26860
0 26862 5 1 1 26861
0 26863 7 1 2 89727 26862
0 26864 5 1 1 26863
0 26865 7 1 2 58295 77558
0 26866 5 3 1 26865
0 26867 7 1 2 91632 91281
0 26868 5 1 1 26867
0 26869 7 2 2 66461 70647
0 26870 7 2 2 80812 82204
0 26871 5 1 1 91637
0 26872 7 1 2 91635 91638
0 26873 5 1 1 26872
0 26874 7 1 2 26868 26873
0 26875 5 1 1 26874
0 26876 7 1 2 81143 26875
0 26877 5 1 1 26876
0 26878 7 1 2 87420 77556
0 26879 5 1 1 26878
0 26880 7 1 2 73122 75445
0 26881 5 1 1 26880
0 26882 7 1 2 26879 26881
0 26883 5 1 1 26882
0 26884 7 1 2 89229 26883
0 26885 5 1 1 26884
0 26886 7 1 2 71283 84631
0 26887 5 1 1 26886
0 26888 7 1 2 3954 26887
0 26889 5 1 1 26888
0 26890 7 1 2 75533 91636
0 26891 7 1 2 26889 26890
0 26892 5 1 1 26891
0 26893 7 1 2 26885 26892
0 26894 5 1 1 26893
0 26895 7 1 2 66252 26894
0 26896 5 1 1 26895
0 26897 7 1 2 26877 26896
0 26898 7 1 2 26864 26897
0 26899 5 1 1 26898
0 26900 7 1 2 90765 26899
0 26901 5 1 1 26900
0 26902 7 1 2 65942 26901
0 26903 7 1 2 26844 26902
0 26904 5 1 1 26903
0 26905 7 4 2 78171 89850
0 26906 5 3 1 91639
0 26907 7 2 2 63772 90806
0 26908 7 1 2 81020 91646
0 26909 5 1 1 26908
0 26910 7 1 2 91640 26909
0 26911 5 1 1 26910
0 26912 7 1 2 89834 26911
0 26913 5 1 1 26912
0 26914 7 1 2 90889 91477
0 26915 5 1 1 26914
0 26916 7 1 2 26915 24292
0 26917 7 1 2 26913 26916
0 26918 5 1 1 26917
0 26919 7 1 2 88546 26918
0 26920 5 1 1 26919
0 26921 7 1 2 90431 91085
0 26922 5 2 1 26921
0 26923 7 1 2 68513 91648
0 26924 5 1 1 26923
0 26925 7 1 2 90740 90441
0 26926 5 1 1 26925
0 26927 7 1 2 26924 26926
0 26928 5 1 1 26927
0 26929 7 1 2 77872 26928
0 26930 5 1 1 26929
0 26931 7 1 2 87184 90460
0 26932 7 1 2 71009 26931
0 26933 5 1 1 26932
0 26934 7 1 2 26930 26933
0 26935 5 1 1 26934
0 26936 7 2 2 88145 90066
0 26937 7 1 2 26935 91650
0 26938 5 1 1 26937
0 26939 7 1 2 26920 26938
0 26940 5 1 1 26939
0 26941 7 1 2 66462 26940
0 26942 5 1 1 26941
0 26943 7 1 2 72653 89741
0 26944 7 1 2 88547 26943
0 26945 5 1 1 26944
0 26946 7 1 2 26942 26945
0 26947 5 1 1 26946
0 26948 7 1 2 64080 26947
0 26949 5 1 1 26948
0 26950 7 1 2 89935 90970
0 26951 7 1 2 88548 26950
0 26952 5 1 1 26951
0 26953 7 1 2 26949 26952
0 26954 5 1 1 26953
0 26955 7 1 2 60950 26954
0 26956 5 1 1 26955
0 26957 7 1 2 76643 91401
0 26958 7 1 2 91633 26957
0 26959 7 1 2 88549 26958
0 26960 5 1 1 26959
0 26961 7 1 2 61311 26960
0 26962 7 1 2 26956 26961
0 26963 5 1 1 26962
0 26964 7 1 2 66836 26963
0 26965 7 1 2 26904 26964
0 26966 5 1 1 26965
0 26967 7 9 2 66778 75534
0 26968 7 1 2 91652 91028
0 26969 7 1 2 91609 26968
0 26970 5 1 1 26969
0 26971 7 1 2 26966 26970
0 26972 7 1 2 26621 26971
0 26973 5 1 1 26972
0 26974 7 1 2 61947 26973
0 26975 5 1 1 26974
0 26976 7 5 2 87136 88243
0 26977 5 1 1 91661
0 26978 7 1 2 80681 91662
0 26979 5 1 1 26978
0 26980 7 2 2 77820 91080
0 26981 5 1 1 91666
0 26982 7 4 2 63277 72865
0 26983 5 1 1 91668
0 26984 7 1 2 82409 91669
0 26985 5 1 1 26984
0 26986 7 1 2 26981 26985
0 26987 5 1 1 26986
0 26988 7 1 2 60951 26987
0 26989 5 1 1 26988
0 26990 7 1 2 74481 91278
0 26991 5 1 1 26990
0 26992 7 1 2 26989 26991
0 26993 5 1 1 26992
0 26994 7 1 2 63000 26993
0 26995 5 1 1 26994
0 26996 7 1 2 81400 90649
0 26997 5 1 1 26996
0 26998 7 2 2 64081 78080
0 26999 7 1 2 86481 91672
0 27000 5 1 1 26999
0 27001 7 1 2 26997 27000
0 27002 5 1 1 27001
0 27003 7 1 2 63278 27002
0 27004 5 1 1 27003
0 27005 7 3 2 86482 87821
0 27006 5 1 1 91674
0 27007 7 1 2 64082 91675
0 27008 5 1 1 27007
0 27009 7 1 2 27004 27008
0 27010 7 1 2 26995 27009
0 27011 5 1 1 27010
0 27012 7 1 2 60375 27011
0 27013 5 1 1 27012
0 27014 7 1 2 86649 91229
0 27015 5 1 1 27014
0 27016 7 1 2 27013 27015
0 27017 5 1 1 27016
0 27018 7 1 2 64708 27017
0 27019 5 1 1 27018
0 27020 7 1 2 26979 27019
0 27021 5 1 1 27020
0 27022 7 1 2 63489 27021
0 27023 5 1 1 27022
0 27024 7 4 2 86667 84796
0 27025 7 1 2 91031 91677
0 27026 5 1 1 27025
0 27027 7 1 2 27023 27026
0 27028 5 1 1 27027
0 27029 7 1 2 67050 27028
0 27030 5 1 1 27029
0 27031 7 1 2 73070 73340
0 27032 5 1 1 27031
0 27033 7 1 2 63001 27032
0 27034 5 1 1 27033
0 27035 7 1 2 59369 85397
0 27036 5 1 1 27035
0 27037 7 1 2 27034 27036
0 27038 5 2 1 27037
0 27039 7 1 2 84181 91681
0 27040 5 1 1 27039
0 27041 7 1 2 90646 27040
0 27042 5 1 1 27041
0 27043 7 1 2 64541 27042
0 27044 5 1 1 27043
0 27045 7 1 2 63002 73087
0 27046 5 3 1 27045
0 27047 7 1 2 64083 86592
0 27048 5 1 1 27047
0 27049 7 1 2 91683 27048
0 27050 5 1 1 27049
0 27051 7 1 2 82559 27050
0 27052 5 1 1 27051
0 27053 7 1 2 27044 27052
0 27054 5 1 1 27053
0 27055 7 1 2 64709 27054
0 27056 5 1 1 27055
0 27057 7 2 2 64542 86016
0 27058 7 1 2 91663 91686
0 27059 5 1 1 27058
0 27060 7 1 2 27056 27059
0 27061 5 1 1 27060
0 27062 7 1 2 63490 27061
0 27063 5 1 1 27062
0 27064 7 1 2 71420 79145
0 27065 7 1 2 91678 27064
0 27066 5 1 1 27065
0 27067 7 1 2 27063 27066
0 27068 5 1 1 27067
0 27069 7 1 2 66595 27068
0 27070 5 1 1 27069
0 27071 7 2 2 64084 86483
0 27072 5 1 1 91688
0 27073 7 1 2 26338 27072
0 27074 5 1 1 27073
0 27075 7 1 2 63003 27074
0 27076 5 1 1 27075
0 27077 7 1 2 77589 86484
0 27078 5 2 1 27077
0 27079 7 1 2 27076 91690
0 27080 5 1 1 27079
0 27081 7 1 2 60376 27080
0 27082 5 1 1 27081
0 27083 7 1 2 73048 88244
0 27084 5 2 1 27083
0 27085 7 1 2 27082 91692
0 27086 5 1 1 27085
0 27087 7 1 2 59831 27086
0 27088 5 1 1 27087
0 27089 7 1 2 86368 86597
0 27090 5 1 1 27089
0 27091 7 1 2 27088 27090
0 27092 5 1 1 27091
0 27093 7 1 2 75658 27092
0 27094 5 1 1 27093
0 27095 7 1 2 63279 27094
0 27096 7 1 2 27070 27095
0 27097 5 1 1 27096
0 27098 7 1 2 77332 83676
0 27099 5 1 1 27098
0 27100 7 1 2 63004 73511
0 27101 7 1 2 27099 27100
0 27102 5 1 1 27101
0 27103 7 1 2 76003 83677
0 27104 5 1 1 27103
0 27105 7 1 2 61312 79783
0 27106 7 1 2 27104 27105
0 27107 5 1 1 27106
0 27108 7 1 2 27102 27107
0 27109 5 1 1 27108
0 27110 7 1 2 61629 27109
0 27111 5 1 1 27110
0 27112 7 2 2 58745 86680
0 27113 5 1 1 91694
0 27114 7 1 2 3596 18584
0 27115 5 1 1 27114
0 27116 7 1 2 91695 27115
0 27117 5 1 1 27116
0 27118 7 1 2 79258 74664
0 27119 5 1 1 27118
0 27120 7 1 2 27117 27119
0 27121 5 1 1 27120
0 27122 7 1 2 84666 74438
0 27123 7 1 2 27121 27122
0 27124 5 1 1 27123
0 27125 7 1 2 27111 27124
0 27126 5 1 1 27125
0 27127 7 1 2 60952 27126
0 27128 5 1 1 27127
0 27129 7 1 2 81826 90644
0 27130 5 1 1 27129
0 27131 7 2 2 86123 75958
0 27132 7 1 2 85857 91696
0 27133 5 1 1 27132
0 27134 7 1 2 27130 27133
0 27135 5 1 1 27134
0 27136 7 1 2 87259 27135
0 27137 5 1 1 27136
0 27138 7 1 2 58535 27137
0 27139 7 1 2 27128 27138
0 27140 5 1 1 27139
0 27141 7 1 2 64815 27140
0 27142 7 1 2 27097 27141
0 27143 5 1 1 27142
0 27144 7 1 2 27030 27143
0 27145 5 1 1 27144
0 27146 7 1 2 66463 27145
0 27147 5 1 1 27146
0 27148 7 3 2 59832 85458
0 27149 7 3 2 71284 73417
0 27150 5 1 1 91701
0 27151 7 1 2 90862 91702
0 27152 5 1 1 27151
0 27153 7 2 2 64085 73624
0 27154 5 1 1 91704
0 27155 7 1 2 58536 91705
0 27156 5 1 1 27155
0 27157 7 1 2 27152 27156
0 27158 5 1 1 27157
0 27159 7 1 2 91698 27158
0 27160 5 1 1 27159
0 27161 7 1 2 27150 27154
0 27162 5 1 1 27161
0 27163 7 1 2 64543 27162
0 27164 5 1 1 27163
0 27165 7 1 2 79704 80671
0 27166 5 1 1 27165
0 27167 7 1 2 27164 27166
0 27168 5 2 1 27167
0 27169 7 1 2 63280 91706
0 27170 5 1 1 27169
0 27171 7 2 2 73625 91687
0 27172 5 1 1 91708
0 27173 7 1 2 27170 27172
0 27174 5 1 1 27173
0 27175 7 1 2 85311 27174
0 27176 5 1 1 27175
0 27177 7 1 2 27160 27176
0 27178 5 1 1 27177
0 27179 7 1 2 91424 27178
0 27180 5 1 1 27179
0 27181 7 1 2 27147 27180
0 27182 5 1 1 27181
0 27183 7 1 2 63623 27182
0 27184 5 1 1 27183
0 27185 7 1 2 58537 89666
0 27186 5 1 1 27185
0 27187 7 2 2 61313 90177
0 27188 7 1 2 86859 91710
0 27189 5 1 1 27188
0 27190 7 1 2 27186 27189
0 27191 5 1 1 27190
0 27192 7 1 2 60953 27191
0 27193 5 2 1 27192
0 27194 7 1 2 86133 90955
0 27195 5 1 1 27194
0 27196 7 1 2 91712 27195
0 27197 5 1 1 27196
0 27198 7 1 2 63005 27197
0 27199 5 1 1 27198
0 27200 7 5 2 61828 81187
0 27201 7 2 2 70209 85727
0 27202 7 1 2 91714 91719
0 27203 5 1 1 27202
0 27204 7 3 2 63281 86124
0 27205 5 1 1 91721
0 27206 7 1 2 90157 91722
0 27207 5 1 1 27206
0 27208 7 1 2 27203 27207
0 27209 7 1 2 90957 27208
0 27210 7 1 2 27199 27209
0 27211 5 1 1 27210
0 27212 7 1 2 59833 27211
0 27213 5 1 1 27212
0 27214 7 1 2 70906 91081
0 27215 5 1 1 27214
0 27216 7 1 2 91691 27215
0 27217 5 1 1 27216
0 27218 7 1 2 60377 27217
0 27219 5 1 1 27218
0 27220 7 1 2 91693 27219
0 27221 5 1 1 27220
0 27222 7 1 2 58538 27221
0 27223 5 1 1 27222
0 27224 7 1 2 63282 86939
0 27225 7 1 2 87200 27224
0 27226 5 1 1 27225
0 27227 7 1 2 27223 27226
0 27228 5 1 1 27227
0 27229 7 1 2 89261 27228
0 27230 5 1 1 27229
0 27231 7 1 2 27213 27230
0 27232 5 2 1 27231
0 27233 7 1 2 63491 91724
0 27234 5 1 1 27233
0 27235 7 1 2 66952 27234
0 27236 5 1 1 27235
0 27237 7 1 2 89590 91707
0 27238 5 1 1 27237
0 27239 7 3 2 61630 71421
0 27240 7 2 2 90961 91726
0 27241 5 1 1 91729
0 27242 7 1 2 64544 91730
0 27243 5 1 1 27242
0 27244 7 1 2 27238 27243
0 27245 5 1 1 27244
0 27246 7 1 2 63283 27245
0 27247 5 1 1 27246
0 27248 7 1 2 89591 91709
0 27249 5 1 1 27248
0 27250 7 1 2 66801 27249
0 27251 7 1 2 27247 27250
0 27252 5 1 1 27251
0 27253 7 1 2 91525 27252
0 27254 7 1 2 27236 27253
0 27255 5 1 1 27254
0 27256 7 1 2 27184 27255
0 27257 5 1 1 27256
0 27258 7 1 2 62093 27257
0 27259 5 1 1 27258
0 27260 7 1 2 69939 83661
0 27261 7 1 2 86684 27260
0 27262 7 1 2 90677 90926
0 27263 7 1 2 27261 27262
0 27264 5 1 1 27263
0 27265 7 1 2 27259 27264
0 27266 5 1 1 27265
0 27267 7 1 2 88389 27266
0 27268 5 1 1 27267
0 27269 7 2 2 88399 90389
0 27270 7 1 2 85370 91731
0 27271 5 1 1 27270
0 27272 7 1 2 85087 89162
0 27273 7 1 2 89311 27272
0 27274 7 1 2 91332 27273
0 27275 5 1 1 27274
0 27276 7 1 2 27271 27275
0 27277 5 1 1 27276
0 27278 7 1 2 64326 27277
0 27279 5 1 1 27278
0 27280 7 1 2 91732 91394
0 27281 5 1 1 27280
0 27282 7 1 2 27279 27281
0 27283 5 1 1 27282
0 27284 7 1 2 66253 27283
0 27285 5 1 1 27284
0 27286 7 2 2 82099 90069
0 27287 7 1 2 88215 89970
0 27288 7 1 2 91733 27287
0 27289 5 1 1 27288
0 27290 7 1 2 27285 27289
0 27291 5 1 1 27290
0 27292 7 1 2 65606 27291
0 27293 5 1 1 27292
0 27294 7 1 2 89592 91703
0 27295 5 1 1 27294
0 27296 7 1 2 27241 27295
0 27297 5 1 1 27296
0 27298 7 1 2 27297 91404
0 27299 5 1 1 27298
0 27300 7 2 2 85798 89163
0 27301 7 3 2 66254 89312
0 27302 7 1 2 63006 72654
0 27303 7 1 2 91737 27302
0 27304 7 1 2 91735 27303
0 27305 5 1 1 27304
0 27306 7 1 2 27299 27305
0 27307 7 1 2 27293 27306
0 27308 5 1 1 27307
0 27309 7 1 2 64816 27308
0 27310 5 1 1 27309
0 27311 7 3 2 60378 82657
0 27312 7 4 2 58539 73831
0 27313 7 1 2 91740 91743
0 27314 5 1 1 27313
0 27315 7 1 2 86977 82100
0 27316 7 1 2 87851 27315
0 27317 5 1 1 27316
0 27318 7 1 2 27314 27317
0 27319 5 1 1 27318
0 27320 7 1 2 88747 90962
0 27321 7 1 2 27319 27320
0 27322 5 1 1 27321
0 27323 7 1 2 27310 27322
0 27324 5 1 1 27323
0 27325 7 1 2 62094 27324
0 27326 5 1 1 27325
0 27327 7 1 2 90678 90421
0 27328 7 3 2 61314 74987
0 27329 7 1 2 91747 91021
0 27330 7 1 2 27327 27329
0 27331 5 1 1 27330
0 27332 7 1 2 27326 27331
0 27333 5 1 1 27332
0 27334 7 1 2 79891 27333
0 27335 5 1 1 27334
0 27336 7 3 2 64545 73088
0 27337 5 1 1 91750
0 27338 7 1 2 73123 89722
0 27339 5 1 1 27338
0 27340 7 1 2 27337 27339
0 27341 5 1 1 27340
0 27342 7 1 2 81255 27341
0 27343 5 1 1 27342
0 27344 7 1 2 73261 82593
0 27345 5 1 1 27344
0 27346 7 1 2 84435 72901
0 27347 7 1 2 27345 27346
0 27348 7 1 2 90777 27347
0 27349 5 1 1 27348
0 27350 7 1 2 27343 27349
0 27351 5 1 1 27350
0 27352 7 1 2 89318 27351
0 27353 5 1 1 27352
0 27354 7 1 2 64327 86978
0 27355 7 1 2 89810 27354
0 27356 7 1 2 84797 90691
0 27357 7 1 2 27355 27356
0 27358 5 1 1 27357
0 27359 7 1 2 27353 27358
0 27360 5 1 1 27359
0 27361 7 1 2 85459 27360
0 27362 5 1 1 27361
0 27363 7 1 2 80021 90248
0 27364 7 7 2 63492 86668
0 27365 7 3 2 63284 89900
0 27366 7 1 2 91753 91760
0 27367 7 1 2 27363 27366
0 27368 5 1 1 27367
0 27369 7 1 2 85110 89649
0 27370 5 2 1 27369
0 27371 7 1 2 65607 91133
0 27372 5 1 1 27371
0 27373 7 1 2 91763 27372
0 27374 5 1 1 27373
0 27375 7 1 2 74482 27374
0 27376 5 1 1 27375
0 27377 7 1 2 91713 27376
0 27378 5 1 1 27377
0 27379 7 1 2 59834 27378
0 27380 5 1 1 27379
0 27381 7 1 2 60954 90178
0 27382 7 1 2 91667 27381
0 27383 5 1 1 27382
0 27384 7 1 2 27380 27383
0 27385 5 1 1 27384
0 27386 7 1 2 76606 74889
0 27387 7 1 2 27385 27386
0 27388 5 1 1 27387
0 27389 7 1 2 27368 27388
0 27390 5 1 1 27389
0 27391 7 1 2 61948 27390
0 27392 5 1 1 27391
0 27393 7 1 2 27362 27392
0 27394 5 1 1 27393
0 27395 7 1 2 63007 27394
0 27396 5 1 1 27395
0 27397 7 1 2 86698 86965
0 27398 5 3 1 27397
0 27399 7 2 2 70173 91765
0 27400 5 1 1 91768
0 27401 7 1 2 66972 91769
0 27402 5 1 1 27401
0 27403 7 1 2 84182 67051
0 27404 7 1 2 86369 27403
0 27405 5 1 1 27404
0 27406 7 1 2 27402 27405
0 27407 5 1 1 27406
0 27408 7 1 2 75535 27407
0 27409 5 1 1 27408
0 27410 7 1 2 67052 89789
0 27411 5 1 1 27410
0 27412 7 4 2 61315 66596
0 27413 7 7 2 64817 91770
0 27414 5 1 1 91774
0 27415 7 1 2 74540 91775
0 27416 5 1 1 27415
0 27417 7 1 2 27411 27416
0 27418 5 1 1 27417
0 27419 7 1 2 64086 27418
0 27420 5 1 1 27419
0 27421 7 1 2 89473 27420
0 27422 5 1 1 27421
0 27423 7 8 2 61631 75574
0 27424 5 2 1 91781
0 27425 7 1 2 27422 91782
0 27426 5 1 1 27425
0 27427 7 1 2 27409 27426
0 27428 5 1 1 27427
0 27429 7 1 2 89990 27428
0 27430 5 1 1 27429
0 27431 7 1 2 67053 91255
0 27432 7 1 2 91720 27431
0 27433 5 1 1 27432
0 27434 7 1 2 27430 27433
0 27435 5 1 1 27434
0 27436 7 1 2 66837 27435
0 27437 5 1 1 27436
0 27438 7 1 2 64546 27400
0 27439 5 1 1 27438
0 27440 7 1 2 59835 91064
0 27441 5 1 1 27440
0 27442 7 1 2 63285 27441
0 27443 7 1 2 27439 27442
0 27444 5 1 1 27443
0 27445 7 2 2 58540 79981
0 27446 5 1 1 91791
0 27447 7 1 2 77348 84779
0 27448 7 1 2 91792 27447
0 27449 5 1 1 27448
0 27450 7 1 2 27444 27449
0 27451 5 1 1 27450
0 27452 7 8 2 66464 66779
0 27453 7 1 2 67435 91793
0 27454 7 1 2 27451 27453
0 27455 5 1 1 27454
0 27456 7 1 2 27437 27455
0 27457 5 1 1 27456
0 27458 7 1 2 62095 27457
0 27459 5 1 1 27458
0 27460 7 1 2 27396 27459
0 27461 5 1 1 27460
0 27462 7 1 2 64894 27461
0 27463 5 1 1 27462
0 27464 7 3 2 66780 87857
0 27465 5 1 1 91801
0 27466 7 1 2 67958 91802
0 27467 7 1 2 91725 27466
0 27468 5 1 1 27467
0 27469 7 1 2 58861 27468
0 27470 7 1 2 27463 27469
0 27471 7 1 2 27335 27470
0 27472 5 1 1 27471
0 27473 7 1 2 58541 89835
0 27474 5 1 1 27473
0 27475 7 1 2 77802 84183
0 27476 5 1 1 27475
0 27477 7 1 2 27474 27476
0 27478 5 2 1 27477
0 27479 7 1 2 90837 91804
0 27480 5 1 1 27479
0 27481 7 1 2 63286 79399
0 27482 7 1 2 87898 90138
0 27483 7 1 2 27481 27482
0 27484 5 1 1 27483
0 27485 7 1 2 27480 27484
0 27486 5 1 1 27485
0 27487 7 1 2 91794 27486
0 27488 5 1 1 27487
0 27489 7 2 2 61632 90674
0 27490 7 1 2 85799 90712
0 27491 7 1 2 85382 27490
0 27492 7 1 2 91806 27491
0 27493 5 1 1 27492
0 27494 7 1 2 27488 27493
0 27495 5 1 1 27494
0 27496 7 1 2 64328 27495
0 27497 5 1 1 27496
0 27498 7 1 2 85678 90852
0 27499 7 1 2 91273 27498
0 27500 5 1 1 27499
0 27501 7 1 2 27497 27500
0 27502 5 1 1 27501
0 27503 7 1 2 63008 27502
0 27504 5 1 1 27503
0 27505 7 1 2 78081 89628
0 27506 5 1 1 27505
0 27507 7 1 2 73721 90028
0 27508 5 1 1 27507
0 27509 7 1 2 27506 27508
0 27510 5 1 1 27509
0 27511 7 1 2 58542 27510
0 27512 5 1 1 27511
0 27513 7 1 2 59584 89505
0 27514 7 1 2 90778 27513
0 27515 5 1 1 27514
0 27516 7 1 2 27512 27515
0 27517 5 1 1 27516
0 27518 7 1 2 66781 89137
0 27519 7 1 2 27517 27518
0 27520 5 1 1 27519
0 27521 7 1 2 89667 90501
0 27522 5 1 1 27521
0 27523 7 1 2 87044 91736
0 27524 7 1 2 91807 27523
0 27525 5 1 1 27524
0 27526 7 1 2 27522 27525
0 27527 5 1 1 27526
0 27528 7 1 2 63009 27527
0 27529 5 1 1 27528
0 27530 7 1 2 62096 73013
0 27531 7 1 2 82878 27530
0 27532 7 1 2 90481 27531
0 27533 5 1 1 27532
0 27534 7 1 2 27529 27533
0 27535 5 1 1 27534
0 27536 7 1 2 66905 27535
0 27537 5 1 1 27536
0 27538 7 1 2 27520 27537
0 27539 7 1 2 27504 27538
0 27540 5 1 1 27539
0 27541 7 1 2 61949 27540
0 27542 5 1 1 27541
0 27543 7 1 2 76644 86264
0 27544 5 1 1 27543
0 27545 7 1 2 76743 87738
0 27546 5 1 1 27545
0 27547 7 1 2 27544 27546
0 27548 5 1 1 27547
0 27549 7 1 2 79150 89025
0 27550 7 1 2 84165 27549
0 27551 7 1 2 27548 27550
0 27552 5 1 1 27551
0 27553 7 1 2 60128 27552
0 27554 7 1 2 27542 27553
0 27555 5 1 1 27554
0 27556 7 1 2 71422 89836
0 27557 5 1 1 27556
0 27558 7 1 2 58543 87354
0 27559 7 1 2 27557 27558
0 27560 5 1 1 27559
0 27561 7 1 2 61633 73832
0 27562 5 2 1 27561
0 27563 7 1 2 63287 91808
0 27564 5 1 1 27563
0 27565 7 1 2 75659 27564
0 27566 7 1 2 27560 27565
0 27567 5 1 1 27566
0 27568 7 1 2 79259 91741
0 27569 5 1 1 27568
0 27570 7 1 2 85101 82116
0 27571 5 1 1 27570
0 27572 7 1 2 27569 27571
0 27573 5 1 1 27572
0 27574 7 1 2 58544 74665
0 27575 5 1 1 27574
0 27576 7 1 2 24474 27575
0 27577 5 1 1 27576
0 27578 7 1 2 27573 27577
0 27579 5 1 1 27578
0 27580 7 1 2 83634 91742
0 27581 5 1 1 27580
0 27582 7 2 2 61634 82618
0 27583 7 1 2 86017 91810
0 27584 5 1 1 27583
0 27585 7 1 2 27581 27584
0 27586 5 1 1 27585
0 27587 7 1 2 87173 27586
0 27588 5 1 1 27587
0 27589 7 2 2 82101 83662
0 27590 7 1 2 85339 77506
0 27591 7 1 2 91812 27590
0 27592 5 1 1 27591
0 27593 7 1 2 27588 27592
0 27594 7 1 2 27579 27593
0 27595 7 1 2 27567 27594
0 27596 5 1 1 27595
0 27597 7 1 2 87812 27596
0 27598 5 1 1 27597
0 27599 7 2 2 77590 90111
0 27600 7 1 2 81827 91814
0 27601 7 1 2 91367 27600
0 27602 5 1 1 27601
0 27603 7 1 2 27598 27602
0 27604 5 1 1 27603
0 27605 7 1 2 90667 27604
0 27606 5 1 1 27605
0 27607 7 1 2 63010 87813
0 27608 7 1 2 90503 27607
0 27609 7 1 2 90280 27608
0 27610 5 1 1 27609
0 27611 7 2 2 71423 89880
0 27612 7 1 2 81918 91816
0 27613 5 1 1 27612
0 27614 7 1 2 23892 27613
0 27615 5 1 1 27614
0 27616 7 2 2 66706 88216
0 27617 7 1 2 79892 91818
0 27618 7 1 2 27615 27617
0 27619 5 1 1 27618
0 27620 7 1 2 27610 27619
0 27621 5 1 1 27620
0 27622 7 1 2 76744 27621
0 27623 5 1 1 27622
0 27624 7 1 2 89846 91544
0 27625 5 1 1 27624
0 27626 7 1 2 77791 89558
0 27627 5 1 1 27626
0 27628 7 1 2 27625 27627
0 27629 5 1 1 27628
0 27630 7 1 2 66906 27629
0 27631 5 1 1 27630
0 27632 7 2 2 66255 84004
0 27633 7 1 2 88915 91032
0 27634 7 1 2 91820 27633
0 27635 5 1 1 27634
0 27636 7 1 2 74905 90618
0 27637 7 1 2 81053 27636
0 27638 5 1 1 27637
0 27639 7 1 2 27635 27638
0 27640 7 1 2 27631 27639
0 27641 5 1 1 27640
0 27642 7 1 2 91819 27641
0 27643 5 1 1 27642
0 27644 7 1 2 63011 91274
0 27645 5 1 1 27644
0 27646 7 1 2 64329 89742
0 27647 5 1 1 27646
0 27648 7 1 2 27645 27647
0 27649 5 1 1 27648
0 27650 7 12 2 58545 58746
0 27651 5 1 1 91822
0 27652 7 1 2 74796 90390
0 27653 7 1 2 91823 27652
0 27654 7 1 2 27649 27653
0 27655 5 1 1 27654
0 27656 7 1 2 27643 27655
0 27657 7 1 2 27623 27656
0 27658 5 1 1 27657
0 27659 7 1 2 65943 27658
0 27660 5 1 1 27659
0 27661 7 1 2 64818 27660
0 27662 7 1 2 27606 27661
0 27663 5 1 1 27662
0 27664 7 1 2 60955 27663
0 27665 7 1 2 27555 27664
0 27666 5 1 1 27665
0 27667 7 1 2 88748 88043
0 27668 5 1 1 27667
0 27669 7 1 2 75536 91803
0 27670 5 1 1 27669
0 27671 7 1 2 27668 27670
0 27672 5 1 1 27671
0 27673 7 1 2 86611 91682
0 27674 7 1 2 27672 27673
0 27675 5 1 1 27674
0 27676 7 3 2 61950 86485
0 27677 7 1 2 90504 91834
0 27678 7 1 2 85460 27677
0 27679 7 1 2 87826 27678
0 27680 5 1 1 27679
0 27681 7 1 2 27675 27680
0 27682 5 1 1 27681
0 27683 7 1 2 60379 27682
0 27684 5 1 1 27683
0 27685 7 1 2 66838 88749
0 27686 5 1 1 27685
0 27687 7 1 2 27465 27686
0 27688 5 1 1 27687
0 27689 7 2 2 77873 75464
0 27690 5 1 1 91837
0 27691 7 1 2 80633 85587
0 27692 5 1 1 27691
0 27693 7 1 2 27690 27692
0 27694 5 1 1 27693
0 27695 7 1 2 59585 27694
0 27696 5 1 1 27695
0 27697 7 1 2 65944 80965
0 27698 5 1 1 27697
0 27699 7 1 2 27696 27698
0 27700 5 1 1 27699
0 27701 7 1 2 27688 27700
0 27702 5 1 1 27701
0 27703 7 5 2 58546 79893
0 27704 7 1 2 59836 74132
0 27705 7 1 2 74155 88750
0 27706 7 1 2 27704 27705
0 27707 7 1 2 91839 27706
0 27708 5 1 1 27707
0 27709 7 1 2 27702 27708
0 27710 5 1 1 27709
0 27711 7 1 2 82102 27710
0 27712 5 1 1 27711
0 27713 7 1 2 27684 27712
0 27714 5 1 1 27713
0 27715 7 1 2 66465 27714
0 27716 5 1 1 27715
0 27717 7 2 2 75537 85728
0 27718 5 1 1 91844
0 27719 7 1 2 63012 91479
0 27720 5 1 1 27719
0 27721 7 1 2 27718 27720
0 27722 5 1 1 27721
0 27723 7 1 2 85312 27722
0 27724 5 1 1 27723
0 27725 7 2 2 74133 87728
0 27726 5 1 1 91846
0 27727 7 5 2 58547 73691
0 27728 5 1 1 91848
0 27729 7 1 2 80446 91849
0 27730 5 1 1 27729
0 27731 7 1 2 27726 27730
0 27732 5 1 1 27731
0 27733 7 1 2 91699 27732
0 27734 5 1 1 27733
0 27735 7 1 2 27724 27734
0 27736 5 1 1 27735
0 27737 7 1 2 90505 91425
0 27738 7 1 2 27736 27737
0 27739 5 1 1 27738
0 27740 7 1 2 27716 27739
0 27741 5 1 1 27740
0 27742 7 1 2 62097 27741
0 27743 5 1 1 27742
0 27744 7 1 2 63624 27743
0 27745 7 1 2 27666 27744
0 27746 5 1 1 27745
0 27747 7 1 2 63708 27746
0 27748 7 1 2 27472 27747
0 27749 5 1 1 27748
0 27750 7 1 2 27268 27749
0 27751 5 1 1 27750
0 27752 7 1 2 82725 27751
0 27753 5 1 1 27752
0 27754 7 1 2 26975 27753
0 27755 7 1 2 26320 27754
0 27756 5 1 1 27755
0 27757 7 1 2 70815 27756
0 27758 5 1 1 27757
0 27759 7 1 2 80361 20030
0 27760 5 1 1 27759
0 27761 7 1 2 62739 27760
0 27762 5 1 1 27761
0 27763 7 1 2 81934 80259
0 27764 5 1 1 27763
0 27765 7 1 2 27762 27764
0 27766 5 1 1 27765
0 27767 7 1 2 60577 27766
0 27768 5 1 1 27767
0 27769 7 1 2 68236 75359
0 27770 5 2 1 27769
0 27771 7 1 2 27768 91853
0 27772 5 1 1 27771
0 27773 7 1 2 58296 27772
0 27774 5 1 1 27773
0 27775 7 1 2 84923 78371
0 27776 5 3 1 27775
0 27777 7 1 2 91313 91855
0 27778 5 1 1 27777
0 27779 7 1 2 27774 27778
0 27780 5 1 1 27779
0 27781 7 1 2 82205 27780
0 27782 5 1 1 27781
0 27783 7 2 2 71739 70048
0 27784 5 1 1 91858
0 27785 7 1 2 72726 27784
0 27786 5 1 1 27785
0 27787 7 1 2 57422 27786
0 27788 5 1 1 27787
0 27789 7 2 2 71891 78316
0 27790 5 1 1 91860
0 27791 7 1 2 88261 27790
0 27792 7 1 2 27788 27791
0 27793 5 1 1 27792
0 27794 7 1 2 58037 27793
0 27795 5 1 1 27794
0 27796 7 1 2 86889 27795
0 27797 5 2 1 27796
0 27798 7 2 2 61635 91862
0 27799 7 1 2 86579 91864
0 27800 5 1 1 27799
0 27801 7 1 2 27782 27800
0 27802 5 1 1 27801
0 27803 7 1 2 64330 27802
0 27804 5 1 1 27803
0 27805 7 1 2 79418 91865
0 27806 5 1 1 27805
0 27807 7 1 2 27804 27806
0 27808 5 1 1 27807
0 27809 7 1 2 63288 27808
0 27810 5 1 1 27809
0 27811 7 2 2 71424 88611
0 27812 7 1 2 91866 91863
0 27813 5 1 1 27812
0 27814 7 1 2 27810 27813
0 27815 5 1 1 27814
0 27816 7 1 2 88704 27815
0 27817 5 1 1 27816
0 27818 7 1 2 62740 81469
0 27819 7 1 2 89173 27818
0 27820 5 1 1 27819
0 27821 7 1 2 72552 90161
0 27822 5 1 1 27821
0 27823 7 1 2 79683 80702
0 27824 5 1 1 27823
0 27825 7 1 2 27822 27824
0 27826 5 1 1 27825
0 27827 7 1 2 88010 88705
0 27828 7 1 2 27826 27827
0 27829 5 1 1 27828
0 27830 7 1 2 27820 27829
0 27831 5 1 1 27830
0 27832 7 1 2 87934 27831
0 27833 5 1 1 27832
0 27834 7 1 2 59128 90021
0 27835 5 1 1 27834
0 27836 7 1 2 85239 73348
0 27837 5 1 1 27836
0 27838 7 1 2 27835 27837
0 27839 5 1 1 27838
0 27840 7 1 2 73404 90769
0 27841 7 1 2 27839 27840
0 27842 5 1 1 27841
0 27843 7 1 2 27833 27842
0 27844 7 1 2 27817 27843
0 27845 5 1 1 27844
0 27846 7 1 2 61316 27845
0 27847 5 1 1 27846
0 27848 7 2 2 61951 90070
0 27849 7 2 2 65268 87935
0 27850 7 1 2 66256 79655
0 27851 5 1 1 27850
0 27852 7 2 2 59837 81445
0 27853 5 5 1 91872
0 27854 7 1 2 59129 91873
0 27855 5 1 1 27854
0 27856 7 1 2 27851 27855
0 27857 5 1 1 27856
0 27858 7 1 2 57704 27857
0 27859 5 1 1 27858
0 27860 7 1 2 70721 82560
0 27861 5 1 1 27860
0 27862 7 1 2 27859 27861
0 27863 5 1 1 27862
0 27864 7 1 2 58548 27863
0 27865 5 1 1 27864
0 27866 7 4 2 63289 82410
0 27867 5 1 1 91879
0 27868 7 1 2 69191 91880
0 27869 5 1 1 27868
0 27870 7 1 2 27865 27869
0 27871 5 1 1 27870
0 27872 7 1 2 78503 27871
0 27873 5 1 1 27872
0 27874 7 1 2 58549 82606
0 27875 5 3 1 27874
0 27876 7 1 2 72845 82879
0 27877 5 2 1 27876
0 27878 7 1 2 91883 91886
0 27879 5 2 1 27878
0 27880 7 1 2 58038 91888
0 27881 5 1 1 27880
0 27882 7 1 2 67663 89353
0 27883 5 2 1 27882
0 27884 7 1 2 27881 91890
0 27885 5 1 1 27884
0 27886 7 1 2 68619 27885
0 27887 5 1 1 27886
0 27888 7 1 2 86844 89373
0 27889 5 1 1 27888
0 27890 7 1 2 27887 27889
0 27891 7 1 2 27873 27890
0 27892 5 1 1 27891
0 27893 7 1 2 91870 27892
0 27894 5 1 1 27893
0 27895 7 2 2 58039 87936
0 27896 7 1 2 67664 89328
0 27897 5 1 1 27896
0 27898 7 1 2 68620 89381
0 27899 5 1 1 27898
0 27900 7 2 2 58550 89294
0 27901 5 1 1 91894
0 27902 7 1 2 61636 91895
0 27903 5 1 1 27902
0 27904 7 1 2 27899 27903
0 27905 5 1 1 27904
0 27906 7 1 2 68374 27905
0 27907 5 1 1 27906
0 27908 7 1 2 27897 27907
0 27909 5 1 1 27908
0 27910 7 1 2 91892 27909
0 27911 5 1 1 27910
0 27912 7 3 2 62741 81038
0 27913 7 1 2 78528 82561
0 27914 7 1 2 91896 27913
0 27915 5 1 1 27914
0 27916 7 3 2 59838 90346
0 27917 7 2 2 70871 77545
0 27918 5 1 1 91902
0 27919 7 1 2 68375 72655
0 27920 7 1 2 91903 27919
0 27921 7 1 2 91899 27920
0 27922 5 1 1 27921
0 27923 7 1 2 27915 27922
0 27924 7 1 2 27911 27923
0 27925 7 1 2 27894 27924
0 27926 5 1 1 27925
0 27927 7 1 2 91868 27926
0 27928 5 1 1 27927
0 27929 7 1 2 79327 89609
0 27930 5 1 1 27929
0 27931 7 1 2 79856 90619
0 27932 5 1 1 27931
0 27933 7 1 2 27930 27932
0 27934 5 1 1 27933
0 27935 7 1 2 62742 27934
0 27936 5 1 1 27935
0 27937 7 4 2 62458 86642
0 27938 7 1 2 90775 91904
0 27939 5 1 1 27938
0 27940 7 1 2 27936 27939
0 27941 5 1 1 27940
0 27942 7 1 2 87937 27941
0 27943 5 1 1 27942
0 27944 7 2 2 69392 78082
0 27945 5 1 1 91908
0 27946 7 1 2 89610 90442
0 27947 7 1 2 91909 27946
0 27948 5 1 1 27947
0 27949 7 1 2 27943 27948
0 27950 5 1 1 27949
0 27951 7 1 2 61317 27950
0 27952 5 1 1 27951
0 27953 7 1 2 62743 82562
0 27954 5 1 1 27953
0 27955 7 2 2 64547 81470
0 27956 5 2 1 91910
0 27957 7 1 2 87298 91912
0 27958 5 1 1 27957
0 27959 7 1 2 62459 27958
0 27960 5 1 1 27959
0 27961 7 1 2 27954 27960
0 27962 5 1 1 27961
0 27963 7 2 2 60380 71180
0 27964 7 1 2 91914 91869
0 27965 7 1 2 27962 27964
0 27966 5 1 1 27965
0 27967 7 1 2 27952 27966
0 27968 5 1 1 27967
0 27969 7 1 2 58551 27968
0 27970 5 1 1 27969
0 27971 7 1 2 86940 90443
0 27972 7 1 2 90624 27971
0 27973 5 1 1 27972
0 27974 7 2 2 61829 84780
0 27975 7 1 2 77290 87938
0 27976 7 1 2 91916 27975
0 27977 5 1 1 27976
0 27978 7 1 2 27973 27977
0 27979 5 1 1 27978
0 27980 7 1 2 59839 27979
0 27981 5 1 1 27980
0 27982 7 2 2 59130 79164
0 27983 7 1 2 85800 80889
0 27984 7 1 2 89602 27983
0 27985 7 1 2 91918 27984
0 27986 5 1 1 27985
0 27987 7 1 2 27981 27986
0 27988 5 1 1 27987
0 27989 7 1 2 89929 27988
0 27990 5 1 1 27989
0 27991 7 1 2 27970 27990
0 27992 5 1 1 27991
0 27993 7 1 2 68852 27992
0 27994 5 1 1 27993
0 27995 7 1 2 78449 91481
0 27996 5 1 1 27995
0 27997 7 1 2 72678 90347
0 27998 7 1 2 89378 27997
0 27999 5 1 1 27998
0 28000 7 1 2 27996 27999
0 28001 5 1 1 28000
0 28002 7 1 2 76645 28001
0 28003 5 1 1 28002
0 28004 7 2 2 57705 71586
0 28005 7 1 2 77874 87234
0 28006 7 1 2 91920 28005
0 28007 5 1 1 28006
0 28008 7 1 2 28003 28007
0 28009 5 1 1 28008
0 28010 7 1 2 88916 28009
0 28011 5 1 1 28010
0 28012 7 1 2 60578 88975
0 28013 5 1 1 28012
0 28014 7 1 2 80187 28013
0 28015 5 1 1 28014
0 28016 7 2 2 70925 69790
0 28017 5 1 1 91922
0 28018 7 1 2 83510 91923
0 28019 5 1 1 28018
0 28020 7 1 2 28015 28019
0 28021 5 1 1 28020
0 28022 7 1 2 66257 90455
0 28023 7 1 2 28021 28022
0 28024 5 1 1 28023
0 28025 7 1 2 28011 28024
0 28026 5 1 1 28025
0 28027 7 1 2 73089 28026
0 28028 5 1 1 28027
0 28029 7 1 2 27994 28028
0 28030 7 1 2 27928 28029
0 28031 7 1 2 27847 28030
0 28032 5 1 1 28031
0 28033 7 1 2 88373 28032
0 28034 5 1 1 28033
0 28035 7 2 2 65945 83472
0 28036 5 3 1 91924
0 28037 7 2 2 59586 84310
0 28038 7 1 2 91925 91929
0 28039 5 1 1 28038
0 28040 7 2 2 60579 72276
0 28041 5 1 1 91931
0 28042 7 1 2 65269 6106
0 28043 5 1 1 28042
0 28044 7 1 2 28041 28043
0 28045 5 1 1 28044
0 28046 7 1 2 65050 28045
0 28047 5 1 1 28046
0 28048 7 1 2 75249 83893
0 28049 7 1 2 28047 28048
0 28050 5 2 1 28049
0 28051 7 1 2 84754 91933
0 28052 5 1 1 28051
0 28053 7 1 2 28039 28052
0 28054 5 1 1 28053
0 28055 7 1 2 91308 28054
0 28056 5 1 1 28055
0 28057 7 1 2 73662 90770
0 28058 5 1 1 28057
0 28059 7 1 2 90621 28058
0 28060 5 1 1 28059
0 28061 7 1 2 68237 88932
0 28062 5 1 1 28061
0 28063 7 1 2 77875 28062
0 28064 7 1 2 28060 28063
0 28065 5 1 1 28064
0 28066 7 1 2 69420 89174
0 28067 7 1 2 86711 28066
0 28068 5 1 1 28067
0 28069 7 1 2 28065 28068
0 28070 7 1 2 28056 28069
0 28071 5 1 1 28070
0 28072 7 2 2 62098 28071
0 28073 7 1 2 88333 91935
0 28074 5 1 1 28073
0 28075 7 1 2 28034 28074
0 28076 5 1 1 28075
0 28077 7 1 2 69549 28076
0 28078 5 1 1 28077
0 28079 7 1 2 88517 91936
0 28080 5 1 1 28079
0 28081 7 1 2 63290 87356
0 28082 5 1 1 28081
0 28083 7 1 2 64548 86969
0 28084 5 1 1 28083
0 28085 7 1 2 28082 28084
0 28086 5 1 1 28085
0 28087 7 1 2 88604 28086
0 28088 5 1 1 28087
0 28089 7 1 2 59587 81949
0 28090 5 1 1 28089
0 28091 7 1 2 83765 28090
0 28092 5 2 1 28091
0 28093 7 1 2 63013 91937
0 28094 5 1 1 28093
0 28095 7 2 2 74928 77468
0 28096 5 1 1 91939
0 28097 7 1 2 78939 28096
0 28098 5 1 1 28097
0 28099 7 1 2 81950 28098
0 28100 5 1 1 28099
0 28101 7 1 2 28094 28100
0 28102 5 1 1 28101
0 28103 7 1 2 61318 28102
0 28104 5 1 1 28103
0 28105 7 4 2 60580 73014
0 28106 7 2 2 63014 77668
0 28107 5 1 1 91945
0 28108 7 1 2 79054 83777
0 28109 5 1 1 28108
0 28110 7 1 2 28107 28109
0 28111 5 2 1 28110
0 28112 7 1 2 91941 91947
0 28113 5 1 1 28112
0 28114 7 1 2 28104 28113
0 28115 5 1 1 28114
0 28116 7 1 2 66258 28115
0 28117 5 1 1 28116
0 28118 7 1 2 68853 69393
0 28119 5 2 1 28118
0 28120 7 1 2 58040 91949
0 28121 5 1 1 28120
0 28122 7 3 2 73663 81430
0 28123 5 1 1 91951
0 28124 7 1 2 28121 91952
0 28125 5 1 1 28124
0 28126 7 1 2 28117 28125
0 28127 5 1 1 28126
0 28128 7 1 2 64549 28127
0 28129 5 1 1 28128
0 28130 7 2 2 60581 83778
0 28131 5 1 1 91954
0 28132 7 1 2 77093 91955
0 28133 5 1 1 28132
0 28134 7 1 2 77433 28133
0 28135 5 2 1 28134
0 28136 7 1 2 87185 87496
0 28137 7 1 2 91956 28136
0 28138 5 1 1 28137
0 28139 7 1 2 28129 28138
0 28140 5 1 1 28139
0 28141 7 1 2 63291 28140
0 28142 5 1 1 28141
0 28143 7 1 2 91676 91957
0 28144 5 1 1 28143
0 28145 7 1 2 28142 28144
0 28146 5 1 1 28145
0 28147 7 1 2 88374 28146
0 28148 5 1 1 28147
0 28149 7 1 2 28088 28148
0 28150 5 1 1 28149
0 28151 7 1 2 88724 28150
0 28152 5 1 1 28151
0 28153 7 2 2 59840 77149
0 28154 5 1 1 91958
0 28155 7 1 2 61637 91959
0 28156 5 2 1 28155
0 28157 7 1 2 81935 82206
0 28158 5 1 1 28157
0 28159 7 1 2 91960 28158
0 28160 5 1 1 28159
0 28161 7 1 2 58552 28160
0 28162 5 1 1 28161
0 28163 7 1 2 81936 91881
0 28164 5 1 1 28163
0 28165 7 1 2 28162 28164
0 28166 5 1 1 28165
0 28167 7 1 2 68376 28166
0 28168 5 1 1 28167
0 28169 7 1 2 60381 78588
0 28170 7 1 2 89329 28169
0 28171 5 1 1 28170
0 28172 7 1 2 91891 28171
0 28173 7 1 2 28168 28172
0 28174 5 1 1 28173
0 28175 7 1 2 59588 28174
0 28176 5 1 1 28175
0 28177 7 1 2 79493 86643
0 28178 7 1 2 90331 90971
0 28179 7 1 2 28177 28178
0 28180 5 1 1 28179
0 28181 7 1 2 28176 28180
0 28182 5 1 1 28181
0 28183 7 1 2 65946 28182
0 28184 5 1 1 28183
0 28185 7 5 2 66259 73498
0 28186 7 1 2 85088 69775
0 28187 7 1 2 71647 28186
0 28188 7 1 2 91962 28187
0 28189 5 1 1 28188
0 28190 7 1 2 28184 28189
0 28191 5 1 1 28190
0 28192 7 6 2 66466 88129
0 28193 7 3 2 60582 67478
0 28194 7 1 2 91967 91973
0 28195 7 1 2 28191 28194
0 28196 5 1 1 28195
0 28197 7 1 2 28152 28196
0 28198 5 1 1 28197
0 28199 7 1 2 70513 28198
0 28200 5 1 1 28199
0 28201 7 1 2 28080 28200
0 28202 7 1 2 28078 28201
0 28203 5 1 1 28202
0 28204 7 1 2 66907 28203
0 28205 5 1 1 28204
0 28206 7 3 2 61319 77876
0 28207 5 1 1 91976
0 28208 7 1 2 69986 91977
0 28209 5 1 1 28208
0 28210 7 2 2 75538 73664
0 28211 7 1 2 19515 91979
0 28212 5 1 1 28211
0 28213 7 1 2 28209 28212
0 28214 5 1 1 28213
0 28215 7 1 2 57706 28214
0 28216 5 1 1 28215
0 28217 7 1 2 84108 91980
0 28218 5 1 1 28217
0 28219 7 1 2 28216 28218
0 28220 5 1 1 28219
0 28221 7 1 2 66467 28220
0 28222 5 1 1 28221
0 28223 7 1 2 83473 91136
0 28224 7 1 2 89971 28223
0 28225 5 1 1 28224
0 28226 7 1 2 28222 28225
0 28227 5 1 1 28226
0 28228 7 1 2 84311 28227
0 28229 5 1 1 28228
0 28230 7 1 2 75446 73499
0 28231 7 1 2 91934 28230
0 28232 5 1 1 28231
0 28233 7 1 2 85777 89965
0 28234 7 1 2 91932 28233
0 28235 5 1 1 28234
0 28236 7 1 2 28232 28235
0 28237 5 1 1 28236
0 28238 7 1 2 61830 28237
0 28239 5 1 1 28238
0 28240 7 1 2 61320 86340
0 28241 5 1 1 28240
0 28242 7 1 2 72798 79857
0 28243 7 1 2 90179 28242
0 28244 7 1 2 91926 28243
0 28245 7 1 2 28241 28244
0 28246 5 1 1 28245
0 28247 7 1 2 28239 28246
0 28248 5 1 1 28247
0 28249 7 1 2 66260 28248
0 28250 5 1 1 28249
0 28251 7 1 2 28229 28250
0 28252 5 1 1 28251
0 28253 7 1 2 91300 28252
0 28254 5 1 1 28253
0 28255 7 1 2 78292 84667
0 28256 7 1 2 87939 28255
0 28257 5 1 1 28256
0 28258 7 1 2 59589 83482
0 28259 7 1 2 91073 28258
0 28260 5 1 1 28259
0 28261 7 1 2 28257 28260
0 28262 5 1 1 28261
0 28263 7 1 2 64550 28262
0 28264 5 1 1 28263
0 28265 7 2 2 63015 84264
0 28266 5 1 1 91981
0 28267 7 1 2 91575 91982
0 28268 5 1 1 28267
0 28269 7 1 2 28264 28268
0 28270 5 1 1 28269
0 28271 7 1 2 62199 28270
0 28272 5 1 1 28271
0 28273 7 1 2 78303 87454
0 28274 7 1 2 87940 28273
0 28275 5 1 1 28274
0 28276 7 1 2 28272 28275
0 28277 5 1 1 28276
0 28278 7 1 2 66468 28277
0 28279 5 1 1 28278
0 28280 7 2 2 73965 81872
0 28281 7 1 2 77094 91137
0 28282 7 1 2 91983 28281
0 28283 5 1 1 28282
0 28284 7 1 2 28279 28283
0 28285 5 1 1 28284
0 28286 7 1 2 59131 28285
0 28287 5 1 1 28286
0 28288 7 2 2 73833 80156
0 28289 7 1 2 90242 91985
0 28290 5 1 1 28289
0 28291 7 1 2 28287 28290
0 28292 5 1 1 28291
0 28293 7 1 2 60583 28292
0 28294 5 1 1 28293
0 28295 7 2 2 75183 91871
0 28296 7 1 2 89687 91905
0 28297 7 1 2 91987 28296
0 28298 5 1 1 28297
0 28299 7 1 2 28294 28298
0 28300 5 1 1 28299
0 28301 7 1 2 63292 28300
0 28302 5 1 1 28301
0 28303 7 1 2 90575 91988
0 28304 5 1 1 28303
0 28305 7 1 2 74580 87729
0 28306 7 1 2 91558 28305
0 28307 5 1 1 28306
0 28308 7 1 2 28304 28307
0 28309 5 1 1 28308
0 28310 7 1 2 81256 89262
0 28311 7 1 2 28309 28310
0 28312 5 1 1 28311
0 28313 7 1 2 62744 28312
0 28314 7 1 2 28302 28313
0 28315 5 1 1 28314
0 28316 7 1 2 74726 82563
0 28317 5 1 1 28316
0 28318 7 1 2 86515 87930
0 28319 5 1 1 28318
0 28320 7 1 2 64551 86901
0 28321 7 1 2 21574 28320
0 28322 7 1 2 28319 28321
0 28323 5 1 1 28322
0 28324 7 1 2 28317 28323
0 28325 5 1 1 28324
0 28326 7 1 2 91351 28325
0 28327 5 1 1 28326
0 28328 7 2 2 83826 89629
0 28329 5 1 1 91989
0 28330 7 1 2 28327 28329
0 28331 5 1 1 28330
0 28332 7 5 2 62200 68238
0 28333 7 2 2 69394 91991
0 28334 7 1 2 28331 91996
0 28335 5 1 1 28334
0 28336 7 1 2 81873 86580
0 28337 7 1 2 91138 28336
0 28338 7 1 2 91856 28337
0 28339 5 1 1 28338
0 28340 7 1 2 28335 28339
0 28341 5 1 1 28340
0 28342 7 1 2 63293 28341
0 28343 5 1 1 28342
0 28344 7 4 2 57707 79165
0 28345 7 1 2 77546 90180
0 28346 7 1 2 79105 28345
0 28347 7 1 2 91998 28346
0 28348 5 1 1 28347
0 28349 7 1 2 65051 70976
0 28350 5 1 1 28349
0 28351 7 1 2 73293 76549
0 28352 7 1 2 28350 28351
0 28353 5 1 1 28352
0 28354 7 1 2 61831 83827
0 28355 7 1 2 28353 28354
0 28356 5 1 1 28355
0 28357 7 1 2 28348 28356
0 28358 5 1 1 28357
0 28359 7 1 2 61321 28358
0 28360 5 1 1 28359
0 28361 7 2 2 71110 81012
0 28362 5 1 1 92002
0 28363 7 1 2 66469 89811
0 28364 7 1 2 91942 28363
0 28365 7 1 2 92003 28364
0 28366 5 1 1 28365
0 28367 7 1 2 28360 28366
0 28368 5 1 1 28367
0 28369 7 1 2 81257 28368
0 28370 5 1 1 28369
0 28371 7 1 2 58041 28370
0 28372 7 1 2 28343 28371
0 28373 5 1 1 28372
0 28374 7 1 2 28315 28373
0 28375 5 1 1 28374
0 28376 7 1 2 87975 91893
0 28377 5 1 1 28376
0 28378 7 2 2 75184 77469
0 28379 7 1 2 71181 92004
0 28380 5 1 1 28379
0 28381 7 1 2 28377 28380
0 28382 5 1 1 28381
0 28383 7 1 2 61638 28382
0 28384 5 1 1 28383
0 28385 7 1 2 77470 81552
0 28386 7 1 2 79287 28385
0 28387 5 1 1 28386
0 28388 7 1 2 28384 28387
0 28389 5 1 1 28388
0 28390 7 1 2 64552 28389
0 28391 5 1 1 28390
0 28392 7 1 2 91336 92005
0 28393 5 1 1 28392
0 28394 7 1 2 28391 28393
0 28395 5 1 1 28394
0 28396 7 1 2 65947 28395
0 28397 5 1 1 28396
0 28398 7 1 2 58042 86104
0 28399 7 2 2 70591 28398
0 28400 5 1 1 92006
0 28401 7 1 2 61639 79666
0 28402 7 1 2 92007 28401
0 28403 5 1 1 28402
0 28404 7 1 2 28397 28403
0 28405 5 1 1 28404
0 28406 7 1 2 63294 28405
0 28407 5 1 1 28406
0 28408 7 1 2 87094 91458
0 28409 5 1 1 28408
0 28410 7 1 2 28400 28409
0 28411 5 1 1 28410
0 28412 7 1 2 28411 91867
0 28413 5 1 1 28412
0 28414 7 1 2 28407 28413
0 28415 5 1 1 28414
0 28416 7 1 2 66470 28415
0 28417 5 1 1 28416
0 28418 7 1 2 58297 90405
0 28419 5 2 1 28418
0 28420 7 1 2 73090 86581
0 28421 5 1 1 28420
0 28422 7 1 2 92008 28421
0 28423 5 1 1 28422
0 28424 7 1 2 58553 28423
0 28425 5 1 1 28424
0 28426 7 1 2 82904 87497
0 28427 5 1 1 28426
0 28428 7 1 2 28425 28427
0 28429 5 1 1 28428
0 28430 7 1 2 91614 28429
0 28431 5 1 1 28430
0 28432 7 1 2 28417 28431
0 28433 5 1 1 28432
0 28434 7 1 2 74590 28433
0 28435 5 1 1 28434
0 28436 7 1 2 78365 89915
0 28437 5 1 1 28436
0 28438 7 1 2 74000 89650
0 28439 7 1 2 81690 28438
0 28440 5 1 1 28439
0 28441 7 1 2 28437 28440
0 28442 5 1 1 28441
0 28443 7 1 2 71892 28442
0 28444 5 1 1 28443
0 28445 7 1 2 84916 89916
0 28446 5 1 1 28445
0 28447 7 1 2 28444 28446
0 28448 5 1 1 28447
0 28449 7 1 2 63016 28448
0 28450 5 1 1 28449
0 28451 7 1 2 58298 91715
0 28452 7 1 2 91997 28451
0 28453 5 1 1 28452
0 28454 7 1 2 28450 28453
0 28455 5 1 1 28454
0 28456 7 1 2 58043 28455
0 28457 5 1 1 28456
0 28458 7 2 2 69794 78853
0 28459 5 1 1 92010
0 28460 7 1 2 62745 77710
0 28461 7 1 2 89917 28460
0 28462 7 1 2 92011 28461
0 28463 5 1 1 28462
0 28464 7 1 2 28457 28463
0 28465 5 1 1 28464
0 28466 7 1 2 90406 28465
0 28467 5 1 1 28466
0 28468 7 1 2 71587 77877
0 28469 7 1 2 91857 28468
0 28470 5 1 1 28469
0 28471 7 1 2 18777 28459
0 28472 5 1 1 28471
0 28473 7 1 2 60584 84732
0 28474 7 1 2 90461 28473
0 28475 7 1 2 28472 28474
0 28476 5 1 1 28475
0 28477 7 1 2 28470 28476
0 28478 5 1 1 28477
0 28479 7 1 2 89593 28478
0 28480 5 1 1 28479
0 28481 7 1 2 71893 89185
0 28482 7 1 2 72835 28481
0 28483 7 1 2 91270 28482
0 28484 5 1 1 28483
0 28485 7 1 2 28480 28484
0 28486 5 1 1 28485
0 28487 7 1 2 73091 28486
0 28488 5 1 1 28487
0 28489 7 4 2 57708 58554
0 28490 7 3 2 84150 92012
0 28491 7 2 2 58978 92016
0 28492 7 2 2 59590 89295
0 28493 7 1 2 84298 88400
0 28494 7 1 2 92021 28493
0 28495 7 1 2 92019 28494
0 28496 5 1 1 28495
0 28497 7 1 2 28488 28496
0 28498 7 1 2 28467 28497
0 28499 7 1 2 28435 28498
0 28500 7 1 2 28375 28499
0 28501 5 1 1 28500
0 28502 7 1 2 88375 88835
0 28503 7 1 2 28501 28502
0 28504 5 1 1 28503
0 28505 7 1 2 28254 28504
0 28506 5 1 1 28505
0 28507 7 1 2 66597 28506
0 28508 5 1 1 28507
0 28509 7 1 2 87968 91824
0 28510 5 1 1 28509
0 28511 7 2 2 63493 71373
0 28512 7 1 2 80957 92023
0 28513 5 1 1 28512
0 28514 7 1 2 28510 28513
0 28515 5 1 1 28514
0 28516 7 1 2 64895 28515
0 28517 5 1 1 28516
0 28518 7 1 2 26152 28517
0 28519 5 1 1 28518
0 28520 7 1 2 63709 28519
0 28521 5 1 1 28520
0 28522 7 1 2 19084 28521
0 28523 5 1 1 28522
0 28524 7 1 2 86105 88736
0 28525 5 1 1 28524
0 28526 7 2 2 65948 74906
0 28527 7 1 2 83462 89857
0 28528 7 1 2 92025 28527
0 28529 5 1 1 28528
0 28530 7 1 2 28525 28529
0 28531 5 1 1 28530
0 28532 7 1 2 28523 28531
0 28533 5 1 1 28532
0 28534 7 2 2 58555 79025
0 28535 5 3 1 92027
0 28536 7 1 2 20695 92029
0 28537 5 5 1 28536
0 28538 7 2 2 86106 88732
0 28539 7 1 2 89333 92037
0 28540 5 1 1 28539
0 28541 7 4 2 60006 70514
0 28542 7 1 2 90162 90071
0 28543 7 1 2 76897 28542
0 28544 7 1 2 92039 28543
0 28545 5 1 1 28544
0 28546 7 1 2 28540 28545
0 28547 5 1 1 28546
0 28548 7 1 2 64896 28547
0 28549 5 1 1 28548
0 28550 7 1 2 63625 88199
0 28551 7 1 2 92038 28550
0 28552 5 1 1 28551
0 28553 7 1 2 28549 28552
0 28554 5 1 1 28553
0 28555 7 1 2 63710 28554
0 28556 5 1 1 28555
0 28557 7 3 2 65052 79301
0 28558 7 1 2 67429 88401
0 28559 7 1 2 88390 28558
0 28560 7 1 2 92043 28559
0 28561 5 1 1 28560
0 28562 7 1 2 28556 28561
0 28563 5 1 1 28562
0 28564 7 1 2 92032 28563
0 28565 5 1 1 28564
0 28566 7 1 2 28533 28565
0 28567 5 1 1 28566
0 28568 7 1 2 62099 28567
0 28569 5 1 1 28568
0 28570 7 5 2 69421 78854
0 28571 7 1 2 74696 87736
0 28572 5 4 1 28571
0 28573 7 2 2 61832 92051
0 28574 7 1 2 91651 92055
0 28575 7 1 2 87889 28574
0 28576 7 1 2 92046 28575
0 28577 5 1 1 28576
0 28578 7 1 2 28569 28577
0 28579 5 1 1 28578
0 28580 7 1 2 66598 28579
0 28581 5 1 1 28580
0 28582 7 1 2 90462 91139
0 28583 5 1 1 28582
0 28584 7 4 2 64553 89506
0 28585 7 1 2 63295 83483
0 28586 7 1 2 92057 28585
0 28587 5 1 1 28586
0 28588 7 1 2 28583 28587
0 28589 5 1 1 28588
0 28590 7 1 2 62201 28589
0 28591 5 1 1 28590
0 28592 7 1 2 58979 78699
0 28593 5 2 1 28592
0 28594 7 2 2 92052 92061
0 28595 7 1 2 89055 92063
0 28596 5 1 1 28595
0 28597 7 1 2 28591 28596
0 28598 5 1 1 28597
0 28599 7 1 2 60585 28598
0 28600 5 1 1 28599
0 28601 7 1 2 63296 80890
0 28602 7 1 2 92058 28601
0 28603 5 1 1 28602
0 28604 7 1 2 28600 28603
0 28605 5 1 1 28604
0 28606 7 1 2 86064 28605
0 28607 5 1 1 28606
0 28608 7 4 2 60129 88971
0 28609 5 1 1 92065
0 28610 7 1 2 87730 92066
0 28611 5 1 1 28610
0 28612 7 2 2 79180 89507
0 28613 7 1 2 58299 84519
0 28614 7 1 2 92069 28613
0 28615 5 1 1 28614
0 28616 7 1 2 28611 28615
0 28617 5 1 1 28616
0 28618 7 1 2 62202 28617
0 28619 5 1 1 28618
0 28620 7 1 2 92067 92064
0 28621 5 1 1 28620
0 28622 7 1 2 28619 28621
0 28623 5 1 1 28622
0 28624 7 1 2 60586 28623
0 28625 5 1 1 28624
0 28626 7 1 2 92070 91897
0 28627 5 1 1 28626
0 28628 7 1 2 28625 28627
0 28629 5 1 1 28628
0 28630 7 1 2 63626 28629
0 28631 5 1 1 28630
0 28632 7 4 2 63297 79858
0 28633 5 1 1 92071
0 28634 7 1 2 70455 92072
0 28635 7 1 2 27918 28634
0 28636 7 1 2 92056 28635
0 28637 5 1 1 28636
0 28638 7 1 2 28631 28637
0 28639 5 1 1 28638
0 28640 7 1 2 66908 28639
0 28641 5 1 1 28640
0 28642 7 1 2 28607 28641
0 28643 5 1 1 28642
0 28644 7 1 2 90415 28643
0 28645 5 1 1 28644
0 28646 7 1 2 28581 28645
0 28647 5 1 1 28646
0 28648 7 1 2 66261 28647
0 28649 5 1 1 28648
0 28650 7 2 2 75185 74687
0 28651 7 1 2 85901 92075
0 28652 5 1 1 28651
0 28653 7 1 2 91599 28652
0 28654 5 1 1 28653
0 28655 7 1 2 88893 28654
0 28656 5 1 1 28655
0 28657 7 1 2 87731 88829
0 28658 7 1 2 89369 28657
0 28659 5 1 1 28658
0 28660 7 1 2 28656 28659
0 28661 5 1 1 28660
0 28662 7 1 2 61952 28661
0 28663 5 1 1 28662
0 28664 7 1 2 88869 92076
0 28665 5 1 1 28664
0 28666 7 1 2 77640 87964
0 28667 7 1 2 91352 28666
0 28668 7 1 2 92026 28667
0 28669 5 1 1 28668
0 28670 7 1 2 28665 28669
0 28671 5 1 1 28670
0 28672 7 1 2 84540 28671
0 28673 5 1 1 28672
0 28674 7 1 2 28663 28673
0 28675 5 1 1 28674
0 28676 7 1 2 88011 88376
0 28677 7 1 2 28675 28676
0 28678 5 1 1 28677
0 28679 7 1 2 28649 28678
0 28680 5 1 1 28679
0 28681 7 1 2 64331 28680
0 28682 5 1 1 28681
0 28683 7 2 2 58300 86486
0 28684 5 2 1 92077
0 28685 7 1 2 90489 92079
0 28686 5 3 1 28685
0 28687 7 1 2 67054 92081
0 28688 5 1 1 28687
0 28689 7 1 2 80933 67114
0 28690 7 1 2 92078 28689
0 28691 5 1 1 28690
0 28692 7 1 2 28688 28691
0 28693 5 1 1 28692
0 28694 7 1 2 89086 28693
0 28695 5 1 1 28694
0 28696 7 1 2 86522 89437
0 28697 7 2 2 92047 28696
0 28698 7 1 2 90463 92084
0 28699 5 1 1 28698
0 28700 7 1 2 28695 28699
0 28701 5 1 1 28700
0 28702 7 1 2 62746 28701
0 28703 5 1 1 28702
0 28704 7 1 2 91002 91375
0 28705 5 1 1 28704
0 28706 7 1 2 89064 28705
0 28707 5 1 1 28706
0 28708 7 1 2 90487 28707
0 28709 5 1 1 28708
0 28710 7 1 2 78986 90003
0 28711 5 1 1 28710
0 28712 7 1 2 28709 28711
0 28713 5 1 1 28712
0 28714 7 3 2 60130 68708
0 28715 7 1 2 28713 92086
0 28716 5 1 1 28715
0 28717 7 1 2 28703 28716
0 28718 5 1 1 28717
0 28719 7 1 2 63627 28718
0 28720 5 1 1 28719
0 28721 7 1 2 77008 89230
0 28722 5 2 1 28721
0 28723 7 2 2 84874 89263
0 28724 5 1 1 92091
0 28725 7 1 2 92089 28724
0 28726 5 1 1 28725
0 28727 7 1 2 92082 28726
0 28728 5 1 1 28727
0 28729 7 1 2 78482 91572
0 28730 7 1 2 91611 28729
0 28731 5 1 1 28730
0 28732 7 1 2 28728 28731
0 28733 5 2 1 28732
0 28734 7 1 2 84768 92093
0 28735 5 1 1 28734
0 28736 7 1 2 28720 28735
0 28737 5 1 1 28736
0 28738 7 1 2 66782 28737
0 28739 5 1 1 28738
0 28740 7 2 2 72553 88917
0 28741 7 1 2 85461 92095
0 28742 5 1 1 28741
0 28743 7 1 2 87683 89439
0 28744 5 1 1 28743
0 28745 7 1 2 28742 28744
0 28746 5 1 1 28745
0 28747 7 1 2 63628 28746
0 28748 5 1 1 28747
0 28749 7 1 2 88285 92096
0 28750 5 1 1 28749
0 28751 7 1 2 28748 28750
0 28752 5 1 1 28751
0 28753 7 1 2 61640 75465
0 28754 7 1 2 28752 28753
0 28755 5 1 1 28754
0 28756 7 3 2 61833 88405
0 28757 7 1 2 78987 81471
0 28758 7 1 2 92097 28757
0 28759 5 1 1 28758
0 28760 7 1 2 28755 28759
0 28761 5 1 1 28760
0 28762 7 1 2 60382 28761
0 28763 5 1 1 28762
0 28764 7 1 2 90243 22588
0 28765 5 1 1 28764
0 28766 7 1 2 60587 28765
0 28767 7 1 2 88406 28766
0 28768 5 1 1 28767
0 28769 7 6 2 61641 79894
0 28770 7 1 2 75466 92100
0 28771 5 1 1 28770
0 28772 7 1 2 86125 87235
0 28773 7 1 2 75387 28772
0 28774 5 1 1 28773
0 28775 7 1 2 28771 28774
0 28776 5 1 1 28775
0 28777 7 1 2 61834 84541
0 28778 7 1 2 28776 28777
0 28779 5 1 1 28778
0 28780 7 1 2 28768 28779
0 28781 5 1 1 28780
0 28782 7 1 2 68854 28781
0 28783 5 1 1 28782
0 28784 7 1 2 63773 65949
0 28785 7 1 2 79237 28784
0 28786 7 1 2 80994 28785
0 28787 7 1 2 89603 92044
0 28788 7 1 2 28786 28787
0 28789 5 1 1 28788
0 28790 7 1 2 28783 28789
0 28791 7 1 2 28763 28790
0 28792 5 1 1 28791
0 28793 7 1 2 77878 28792
0 28794 5 1 1 28793
0 28795 7 1 2 89067 92094
0 28796 5 1 1 28795
0 28797 7 1 2 89403 92073
0 28798 5 1 1 28797
0 28799 7 1 2 63629 90972
0 28800 7 1 2 89952 28799
0 28801 5 1 1 28800
0 28802 7 1 2 28798 28801
0 28803 5 1 1 28802
0 28804 7 1 2 92083 28803
0 28805 5 1 1 28804
0 28806 7 2 2 61322 89901
0 28807 7 1 2 69550 86582
0 28808 7 1 2 84523 28807
0 28809 7 1 2 92106 28808
0 28810 5 1 1 28809
0 28811 7 1 2 28805 28810
0 28812 5 1 1 28811
0 28813 7 1 2 61953 28812
0 28814 5 1 1 28813
0 28815 7 1 2 80834 88197
0 28816 7 1 2 92085 28815
0 28817 5 1 1 28816
0 28818 7 1 2 28814 28817
0 28819 5 1 1 28818
0 28820 7 1 2 66909 28819
0 28821 5 1 1 28820
0 28822 7 1 2 28796 28821
0 28823 7 1 2 28794 28822
0 28824 7 1 2 28739 28823
0 28825 5 1 1 28824
0 28826 7 1 2 91019 28825
0 28827 5 1 1 28826
0 28828 7 1 2 28682 28827
0 28829 5 1 1 28828
0 28830 7 1 2 67751 28829
0 28831 5 1 1 28830
0 28832 7 1 2 58044 78416
0 28833 5 1 1 28832
0 28834 7 1 2 60588 78988
0 28835 7 1 2 28833 28834
0 28836 5 1 1 28835
0 28837 7 1 2 65270 92053
0 28838 7 1 2 83763 28837
0 28839 5 1 1 28838
0 28840 7 1 2 28836 28839
0 28841 5 1 1 28840
0 28842 7 1 2 89594 28841
0 28843 5 1 1 28842
0 28844 7 1 2 74372 91946
0 28845 5 1 1 28844
0 28846 7 1 2 80484 83779
0 28847 5 1 1 28846
0 28848 7 1 2 28845 28847
0 28849 5 1 1 28848
0 28850 7 1 2 89688 28849
0 28851 5 1 1 28850
0 28852 7 1 2 28843 28851
0 28853 5 1 1 28852
0 28854 7 1 2 88363 28853
0 28855 5 1 1 28854
0 28856 7 1 2 89138 89630
0 28857 5 1 1 28856
0 28858 7 1 2 28855 28857
0 28859 5 1 1 28858
0 28860 7 1 2 63711 28859
0 28861 5 1 1 28860
0 28862 7 1 2 89106 91164
0 28863 5 1 1 28862
0 28864 7 1 2 28861 28863
0 28865 5 1 1 28864
0 28866 7 1 2 59591 28865
0 28867 5 1 1 28866
0 28868 7 1 2 78700 90029
0 28869 5 1 1 28868
0 28870 7 1 2 90244 28869
0 28871 5 1 1 28870
0 28872 7 1 2 67860 28871
0 28873 5 1 1 28872
0 28874 7 1 2 77547 90030
0 28875 5 1 1 28874
0 28876 7 1 2 90245 28875
0 28877 5 1 1 28876
0 28878 7 1 2 57423 28877
0 28879 5 1 1 28878
0 28880 7 1 2 83923 89631
0 28881 5 1 1 28880
0 28882 7 1 2 28879 28881
0 28883 5 1 1 28882
0 28884 7 1 2 76074 28883
0 28885 5 1 1 28884
0 28886 7 1 2 28873 28885
0 28887 5 1 1 28886
0 28888 7 1 2 65271 28887
0 28889 5 1 1 28888
0 28890 7 1 2 76491 74688
0 28891 5 1 1 28890
0 28892 7 1 2 91600 28891
0 28893 5 1 1 28892
0 28894 7 1 2 60589 28893
0 28895 5 1 1 28894
0 28896 7 2 2 63017 68855
0 28897 5 1 1 92108
0 28898 7 1 2 86126 92109
0 28899 5 1 1 28898
0 28900 7 1 2 61323 83263
0 28901 5 1 1 28900
0 28902 7 1 2 28899 28901
0 28903 5 1 1 28902
0 28904 7 1 2 77669 28903
0 28905 5 1 1 28904
0 28906 7 1 2 28895 28905
0 28907 5 1 1 28906
0 28908 7 1 2 89651 28907
0 28909 5 1 1 28908
0 28910 7 1 2 28889 28909
0 28911 5 1 1 28910
0 28912 7 1 2 91012 28911
0 28913 5 1 1 28912
0 28914 7 1 2 28867 28913
0 28915 5 1 1 28914
0 28916 7 1 2 86065 28915
0 28917 5 1 1 28916
0 28918 7 1 2 68666 87607
0 28919 7 1 2 83635 91318
0 28920 7 1 2 28918 28919
0 28921 7 1 2 89376 28920
0 28922 5 1 1 28921
0 28923 7 1 2 28917 28922
0 28924 5 1 1 28923
0 28925 7 1 2 76745 28924
0 28926 5 1 1 28925
0 28927 7 2 2 83559 88130
0 28928 5 1 1 92110
0 28929 7 1 2 69422 89087
0 28930 5 1 1 28929
0 28931 7 1 2 89246 28930
0 28932 5 1 1 28931
0 28933 7 2 2 62100 28932
0 28934 7 1 2 92111 92112
0 28935 5 1 1 28934
0 28936 7 1 2 77670 89088
0 28937 5 1 1 28936
0 28938 7 1 2 92090 28937
0 28939 5 1 1 28938
0 28940 7 1 2 77095 28939
0 28941 5 1 1 28940
0 28942 7 1 2 60590 92092
0 28943 5 1 1 28942
0 28944 7 1 2 28941 28943
0 28945 5 1 1 28944
0 28946 7 1 2 58301 28945
0 28947 5 1 1 28946
0 28948 7 1 2 89264 91314
0 28949 7 1 2 84817 28948
0 28950 5 1 1 28949
0 28951 7 1 2 28947 28950
0 28952 5 1 1 28951
0 28953 7 1 2 88377 28952
0 28954 5 1 1 28953
0 28955 7 1 2 88334 92113
0 28956 5 1 1 28955
0 28957 7 1 2 28954 28956
0 28958 5 1 1 28957
0 28959 7 1 2 86066 28958
0 28960 5 1 1 28959
0 28961 7 1 2 28935 28960
0 28962 5 1 1 28961
0 28963 7 1 2 86712 28962
0 28964 5 1 1 28963
0 28965 7 1 2 89056 91938
0 28966 5 1 1 28965
0 28967 7 1 2 62747 78592
0 28968 5 1 1 28967
0 28969 7 2 2 70816 77096
0 28970 5 1 1 92114
0 28971 7 1 2 62460 92115
0 28972 5 1 1 28971
0 28973 7 1 2 28968 28972
0 28974 5 1 1 28973
0 28975 7 1 2 73722 91003
0 28976 7 1 2 28974 28975
0 28977 5 1 1 28976
0 28978 7 1 2 28966 28977
0 28979 5 1 1 28978
0 28980 7 1 2 63018 28979
0 28981 5 1 1 28980
0 28982 7 1 2 77783 77097
0 28983 7 1 2 89491 28982
0 28984 5 1 1 28983
0 28985 7 1 2 77453 89453
0 28986 7 1 2 77166 28985
0 28987 5 1 1 28986
0 28988 7 1 2 28984 28987
0 28989 5 1 1 28988
0 28990 7 1 2 62461 28989
0 28991 5 1 1 28990
0 28992 7 1 2 81039 89231
0 28993 7 1 2 86084 28992
0 28994 5 1 1 28993
0 28995 7 1 2 28991 28994
0 28996 5 1 1 28995
0 28997 7 1 2 60591 28996
0 28998 5 1 1 28997
0 28999 7 1 2 28981 28998
0 29000 5 1 1 28999
0 29001 7 1 2 61324 29000
0 29002 5 1 1 29001
0 29003 7 1 2 89057 91948
0 29004 5 1 1 29003
0 29005 7 1 2 62462 77098
0 29006 7 1 2 91225 29005
0 29007 5 1 1 29006
0 29008 7 1 2 29004 29007
0 29009 5 1 1 29008
0 29010 7 1 2 91943 29009
0 29011 5 1 1 29010
0 29012 7 1 2 66262 29011
0 29013 7 1 2 29002 29012
0 29014 5 1 1 29013
0 29015 7 2 2 86067 88146
0 29016 7 1 2 85737 74709
0 29017 5 1 1 29016
0 29018 7 1 2 70084 29017
0 29019 5 1 1 29018
0 29020 7 1 2 71588 73015
0 29021 5 1 1 29020
0 29022 7 1 2 29019 29021
0 29023 5 1 1 29022
0 29024 7 1 2 68377 29023
0 29025 5 1 1 29024
0 29026 7 2 2 69818 74689
0 29027 5 1 1 92118
0 29028 7 1 2 65950 76507
0 29029 7 1 2 87941 29028
0 29030 5 1 1 29029
0 29031 7 1 2 29027 29030
0 29032 5 1 1 29031
0 29033 7 1 2 67861 29032
0 29034 5 1 1 29033
0 29035 7 1 2 29025 29034
0 29036 5 1 1 29035
0 29037 7 1 2 89280 29036
0 29038 5 1 1 29037
0 29039 7 2 2 87498 89870
0 29040 7 1 2 91898 92120
0 29041 5 1 1 29040
0 29042 7 1 2 61642 29041
0 29043 7 1 2 29038 29042
0 29044 5 1 1 29043
0 29045 7 1 2 92116 29044
0 29046 7 1 2 29014 29045
0 29047 5 1 1 29046
0 29048 7 1 2 28964 29047
0 29049 7 1 2 28926 29048
0 29050 5 1 1 29049
0 29051 7 1 2 61954 29050
0 29052 5 1 1 29051
0 29053 7 1 2 28831 29052
0 29054 7 1 2 28508 29053
0 29055 7 1 2 28205 29054
0 29056 5 1 1 29055
0 29057 7 1 2 80136 29056
0 29058 5 1 1 29057
0 29059 7 1 2 79533 82306
0 29060 5 1 1 29059
0 29061 7 2 2 75959 82411
0 29062 5 1 1 92122
0 29063 7 1 2 85089 92123
0 29064 5 1 1 29063
0 29065 7 1 2 62748 77879
0 29066 7 2 2 87665 29065
0 29067 7 1 2 57709 92124
0 29068 5 1 1 29067
0 29069 7 1 2 29064 29068
0 29070 5 1 1 29069
0 29071 7 1 2 68856 29070
0 29072 5 1 1 29071
0 29073 7 1 2 88185 92125
0 29074 5 1 1 29073
0 29075 7 1 2 29072 29074
0 29076 5 1 1 29075
0 29077 7 1 2 73092 29076
0 29078 5 1 1 29077
0 29079 7 2 2 62463 79260
0 29080 7 1 2 72656 72969
0 29081 7 1 2 92126 29080
0 29082 5 1 1 29081
0 29083 7 1 2 62203 88564
0 29084 5 1 1 29083
0 29085 7 1 2 88568 29084
0 29086 5 2 1 29085
0 29087 7 1 2 73016 92128
0 29088 5 1 1 29087
0 29089 7 1 2 68857 74058
0 29090 5 1 1 29089
0 29091 7 1 2 29088 29090
0 29092 5 1 1 29091
0 29093 7 1 2 87675 77291
0 29094 7 1 2 29092 29093
0 29095 5 1 1 29094
0 29096 7 1 2 29082 29095
0 29097 5 1 1 29096
0 29098 7 1 2 66263 29097
0 29099 5 1 1 29098
0 29100 7 1 2 29078 29099
0 29101 5 1 1 29100
0 29102 7 1 2 63494 29101
0 29103 5 1 1 29102
0 29104 7 1 2 73049 87637
0 29105 5 2 1 29104
0 29106 7 1 2 79851 91449
0 29107 5 1 1 29106
0 29108 7 1 2 92130 29107
0 29109 5 1 1 29108
0 29110 7 1 2 58556 29109
0 29111 5 1 1 29110
0 29112 7 1 2 89526 90650
0 29113 5 1 1 29112
0 29114 7 2 2 12707 29113
0 29115 7 1 2 85094 92132
0 29116 5 1 1 29115
0 29117 7 1 2 29111 29116
0 29118 5 1 1 29117
0 29119 7 1 2 88022 29118
0 29120 5 1 1 29119
0 29121 7 2 2 68858 89790
0 29122 7 1 2 87656 92134
0 29123 5 1 1 29122
0 29124 7 1 2 29120 29123
0 29125 5 1 1 29124
0 29126 7 1 2 75682 29125
0 29127 5 1 1 29126
0 29128 7 1 2 29103 29127
0 29129 5 1 1 29128
0 29130 7 1 2 69551 29129
0 29131 5 1 1 29130
0 29132 7 1 2 63298 92133
0 29133 5 1 1 29132
0 29134 7 1 2 27006 29133
0 29135 5 1 1 29134
0 29136 7 1 2 88023 29135
0 29137 5 1 1 29136
0 29138 7 1 2 88559 92135
0 29139 5 1 1 29138
0 29140 7 1 2 29137 29139
0 29141 5 1 1 29140
0 29142 7 1 2 61955 86055
0 29143 7 1 2 29141 29142
0 29144 5 1 1 29143
0 29145 7 1 2 29131 29144
0 29146 5 1 1 29145
0 29147 7 1 2 64087 29146
0 29148 5 1 1 29147
0 29149 7 1 2 88571 90301
0 29150 7 1 2 87615 29149
0 29151 5 1 1 29150
0 29152 7 1 2 73665 83047
0 29153 7 1 2 88844 29152
0 29154 5 1 1 29153
0 29155 7 1 2 29151 29154
0 29156 5 1 1 29155
0 29157 7 1 2 78637 29156
0 29158 5 1 1 29157
0 29159 7 2 2 82274 87658
0 29160 5 1 1 92136
0 29161 7 3 2 61325 75186
0 29162 5 1 1 92138
0 29163 7 1 2 64332 75785
0 29164 7 1 2 87666 29163
0 29165 7 1 2 92139 29164
0 29166 5 1 1 29165
0 29167 7 1 2 29160 29166
0 29168 5 1 1 29167
0 29169 7 1 2 63495 29168
0 29170 5 1 1 29169
0 29171 7 4 2 58747 77507
0 29172 7 1 2 87659 92141
0 29173 5 1 1 29172
0 29174 7 1 2 29170 29173
0 29175 5 1 1 29174
0 29176 7 1 2 58045 29175
0 29177 5 1 1 29176
0 29178 7 1 2 29158 29177
0 29179 5 1 1 29178
0 29180 7 1 2 77880 29179
0 29181 5 1 1 29180
0 29182 7 1 2 63299 79656
0 29183 7 1 2 87679 29182
0 29184 7 1 2 82997 29183
0 29185 7 1 2 88186 29184
0 29186 5 1 1 29185
0 29187 7 1 2 29181 29186
0 29188 5 1 1 29187
0 29189 7 1 2 76411 29188
0 29190 5 1 1 29189
0 29191 7 1 2 29148 29190
0 29192 5 1 1 29191
0 29193 7 1 2 63019 29192
0 29194 5 1 1 29193
0 29195 7 1 2 72866 90085
0 29196 5 1 1 29195
0 29197 7 1 2 68006 91751
0 29198 5 1 1 29197
0 29199 7 1 2 29196 29198
0 29200 5 1 1 29199
0 29201 7 1 2 63300 29200
0 29202 5 1 1 29201
0 29203 7 1 2 85630 87321
0 29204 5 1 1 29203
0 29205 7 1 2 29202 29204
0 29206 5 1 1 29205
0 29207 7 1 2 88194 29206
0 29208 5 1 1 29207
0 29209 7 1 2 80899 84611
0 29210 7 1 2 88187 29209
0 29211 5 1 1 29210
0 29212 7 1 2 29208 29211
0 29213 5 1 1 29212
0 29214 7 1 2 90281 29213
0 29215 5 1 1 29214
0 29216 7 1 2 69314 88502
0 29217 5 2 1 29216
0 29218 7 1 2 59592 91068
0 29219 5 1 1 29218
0 29220 7 1 2 92145 29219
0 29221 5 1 1 29220
0 29222 7 5 2 61956 86563
0 29223 7 1 2 87868 92147
0 29224 7 1 2 29221 29223
0 29225 5 1 1 29224
0 29226 7 1 2 29215 29225
0 29227 5 1 1 29226
0 29228 7 1 2 82342 29227
0 29229 5 1 1 29228
0 29230 7 1 2 29194 29229
0 29231 5 1 1 29230
0 29232 7 1 2 88147 29231
0 29233 5 1 1 29232
0 29234 7 1 2 75400 83069
0 29235 5 1 1 29234
0 29236 7 1 2 76204 77271
0 29237 7 1 2 82827 29236
0 29238 5 1 1 29237
0 29239 7 1 2 29235 29238
0 29240 5 1 1 29239
0 29241 7 1 2 75539 29240
0 29242 5 1 1 29241
0 29243 7 9 2 59841 79895
0 29244 5 3 1 92152
0 29245 7 3 2 58557 92153
0 29246 5 3 1 92164
0 29247 7 1 2 70657 74439
0 29248 7 1 2 92165 29247
0 29249 5 1 1 29248
0 29250 7 1 2 29242 29249
0 29251 5 1 1 29250
0 29252 7 1 2 64819 29251
0 29253 5 1 1 29252
0 29254 7 2 2 60131 74440
0 29255 5 2 1 92170
0 29256 7 1 2 63496 70658
0 29257 7 1 2 87676 29256
0 29258 7 1 2 92171 29257
0 29259 5 1 1 29258
0 29260 7 1 2 29253 29259
0 29261 5 1 1 29260
0 29262 7 1 2 63630 29261
0 29263 5 1 1 29262
0 29264 7 1 2 77784 74441
0 29265 7 1 2 83118 29264
0 29266 7 1 2 89344 29265
0 29267 5 1 1 29266
0 29268 7 1 2 29263 29267
0 29269 5 1 1 29268
0 29270 7 1 2 68859 29269
0 29271 5 1 1 29270
0 29272 7 1 2 84213 90444
0 29273 7 1 2 88111 29272
0 29274 5 1 1 29273
0 29275 7 1 2 29271 29274
0 29276 5 1 1 29275
0 29277 7 1 2 66707 29276
0 29278 5 1 1 29277
0 29279 7 2 2 69678 72450
0 29280 7 1 2 88044 92174
0 29281 5 1 1 29280
0 29282 7 1 2 29278 29281
0 29283 5 1 1 29282
0 29284 7 1 2 88131 29283
0 29285 5 1 1 29284
0 29286 7 1 2 72451 91504
0 29287 7 1 2 88112 29286
0 29288 5 1 1 29287
0 29289 7 1 2 29285 29288
0 29290 5 1 1 29289
0 29291 7 1 2 86713 88318
0 29292 7 1 2 29290 29291
0 29293 5 1 1 29292
0 29294 7 1 2 29233 29293
0 29295 5 1 1 29294
0 29296 7 1 2 66471 29295
0 29297 5 1 1 29296
0 29298 7 5 2 64554 79896
0 29299 5 1 1 92176
0 29300 7 4 2 62101 69362
0 29301 7 2 2 88391 92181
0 29302 5 1 1 92185
0 29303 7 1 2 70659 88429
0 29304 5 1 1 29303
0 29305 7 1 2 78231 76847
0 29306 5 1 1 29305
0 29307 7 1 2 29304 29306
0 29308 5 2 1 29307
0 29309 7 1 2 88364 92187
0 29310 5 1 1 29309
0 29311 7 1 2 60197 92182
0 29312 5 1 1 29311
0 29313 7 1 2 29310 29312
0 29314 5 1 1 29313
0 29315 7 1 2 63712 29314
0 29316 5 1 1 29315
0 29317 7 1 2 29302 29316
0 29318 5 1 1 29317
0 29319 7 1 2 61326 29318
0 29320 5 1 1 29319
0 29321 7 1 2 63713 66708
0 29322 7 2 2 88430 29321
0 29323 7 1 2 87732 90713
0 29324 7 1 2 92189 29323
0 29325 5 1 1 29324
0 29326 7 1 2 29320 29325
0 29327 5 1 1 29326
0 29328 7 1 2 64333 29327
0 29329 5 1 1 29328
0 29330 7 2 2 59593 72781
0 29331 7 1 2 90869 92191
0 29332 7 1 2 92190 29331
0 29333 5 1 1 29332
0 29334 7 1 2 29329 29333
0 29335 5 1 1 29334
0 29336 7 1 2 69552 29335
0 29337 5 1 1 29336
0 29338 7 1 2 72867 69363
0 29339 7 1 2 90766 29338
0 29340 5 1 1 29339
0 29341 7 1 2 29337 29340
0 29342 5 1 1 29341
0 29343 7 1 2 92177 29342
0 29344 5 1 1 29343
0 29345 7 1 2 83617 79188
0 29346 7 1 2 88148 29345
0 29347 7 1 2 74707 29346
0 29348 7 1 2 78232 29347
0 29349 5 1 1 29348
0 29350 7 1 2 29344 29349
0 29351 5 1 1 29350
0 29352 7 1 2 63301 29351
0 29353 5 1 1 29352
0 29354 7 1 2 69578 92188
0 29355 5 1 1 29354
0 29356 7 1 2 69367 29355
0 29357 5 1 1 29356
0 29358 7 1 2 66783 29357
0 29359 5 1 1 29358
0 29360 7 1 2 79951 92183
0 29361 5 1 1 29360
0 29362 7 1 2 29359 29361
0 29363 5 1 1 29362
0 29364 7 1 2 64897 29363
0 29365 5 1 1 29364
0 29366 7 1 2 88085 92184
0 29367 5 1 1 29366
0 29368 7 1 2 29365 29367
0 29369 5 1 1 29368
0 29370 7 1 2 63714 29369
0 29371 5 1 1 29370
0 29372 7 1 2 88836 92186
0 29373 5 1 1 29372
0 29374 7 1 2 29371 29373
0 29375 5 1 1 29374
0 29376 7 1 2 77842 72902
0 29377 5 1 1 29376
0 29378 7 4 2 85537 91483
0 29379 7 1 2 29377 92193
0 29380 7 1 2 29375 29379
0 29381 5 1 1 29380
0 29382 7 1 2 88431 91010
0 29383 5 1 1 29382
0 29384 7 2 2 58302 79400
0 29385 7 1 2 78233 92197
0 29386 5 1 1 29385
0 29387 7 1 2 29383 29386
0 29388 5 1 1 29387
0 29389 7 1 2 73093 88980
0 29390 7 1 2 88450 88378
0 29391 7 1 2 29389 29390
0 29392 7 1 2 29388 29391
0 29393 5 1 1 29392
0 29394 7 1 2 29381 29393
0 29395 7 1 2 29353 29394
0 29396 5 1 1 29395
0 29397 7 1 2 66264 29396
0 29398 5 1 1 29397
0 29399 7 1 2 77349 88486
0 29400 5 1 1 29399
0 29401 7 1 2 92146 29400
0 29402 5 1 1 29401
0 29403 7 1 2 63020 29402
0 29404 5 1 1 29403
0 29405 7 1 2 58303 77591
0 29406 7 1 2 88487 29405
0 29407 5 1 1 29406
0 29408 7 1 2 29404 29407
0 29409 5 1 1 29408
0 29410 7 1 2 77881 29409
0 29411 5 1 1 29410
0 29412 7 1 2 78161 92198
0 29413 7 1 2 88503 29412
0 29414 5 1 1 29413
0 29415 7 1 2 29411 29414
0 29416 5 1 1 29415
0 29417 7 1 2 79897 29416
0 29418 5 1 1 29417
0 29419 7 2 2 79824 81040
0 29420 7 6 2 59594 92199
0 29421 5 2 1 92201
0 29422 7 1 2 75808 92202
0 29423 7 1 2 88504 29422
0 29424 5 1 1 29423
0 29425 7 1 2 29418 29424
0 29426 5 1 1 29425
0 29427 7 1 2 64898 88510
0 29428 7 1 2 91579 29427
0 29429 7 1 2 29426 29428
0 29430 5 1 1 29429
0 29431 7 1 2 29398 29430
0 29432 5 1 1 29431
0 29433 7 1 2 88706 29432
0 29434 5 1 1 29433
0 29435 7 1 2 29297 29434
0 29436 5 1 1 29435
0 29437 7 1 2 29060 29436
0 29438 5 1 1 29437
0 29439 7 1 2 78253 75006
0 29440 5 2 1 29439
0 29441 7 1 2 87853 88518
0 29442 5 1 1 29441
0 29443 7 1 2 63497 80813
0 29444 7 1 2 88335 29443
0 29445 7 1 2 79937 29444
0 29446 5 1 1 29445
0 29447 7 1 2 29442 29446
0 29448 5 1 1 29447
0 29449 7 1 2 77481 90707
0 29450 7 1 2 29448 29449
0 29451 5 1 1 29450
0 29452 7 3 2 75540 79452
0 29453 7 1 2 91208 92211
0 29454 7 1 2 90708 29453
0 29455 5 1 1 29454
0 29456 7 5 2 76646 88132
0 29457 7 1 2 72868 81125
0 29458 7 1 2 92214 29457
0 29459 7 1 2 88870 29458
0 29460 5 1 1 29459
0 29461 7 1 2 29455 29460
0 29462 5 1 1 29461
0 29463 7 1 2 70515 79227
0 29464 7 1 2 29462 29463
0 29465 5 1 1 29464
0 29466 7 1 2 29451 29465
0 29467 5 1 1 29466
0 29468 7 1 2 77491 29467
0 29469 5 1 1 29468
0 29470 7 2 2 83141 84469
0 29471 7 2 2 76028 82719
0 29472 7 1 2 92219 92221
0 29473 5 1 1 29472
0 29474 7 4 2 74654 67617
0 29475 5 1 1 92223
0 29476 7 1 2 79166 92224
0 29477 5 1 1 29476
0 29478 7 1 2 29473 29477
0 29479 5 1 1 29478
0 29480 7 1 2 62749 29479
0 29481 5 1 1 29480
0 29482 7 2 2 64820 84470
0 29483 7 3 2 63631 79261
0 29484 7 1 2 92227 92229
0 29485 5 1 1 29484
0 29486 7 2 2 60132 79199
0 29487 7 1 2 74768 90576
0 29488 7 1 2 92232 29487
0 29489 5 1 1 29488
0 29490 7 1 2 29485 29489
0 29491 5 1 1 29490
0 29492 7 1 2 64334 29491
0 29493 5 1 1 29492
0 29494 7 1 2 29481 29493
0 29495 5 1 1 29494
0 29496 7 1 2 63498 29495
0 29497 5 1 1 29496
0 29498 7 1 2 59595 89379
0 29499 5 2 1 29498
0 29500 7 3 2 84471 92234
0 29501 7 1 2 76109 89303
0 29502 7 1 2 92236 29501
0 29503 5 1 1 29502
0 29504 7 1 2 29497 29503
0 29505 5 1 1 29504
0 29506 7 1 2 63302 29505
0 29507 5 1 1 29506
0 29508 7 2 2 79898 92237
0 29509 7 1 2 77821 69553
0 29510 7 1 2 92239 29509
0 29511 5 1 1 29510
0 29512 7 1 2 29507 29511
0 29513 5 1 1 29512
0 29514 7 1 2 63021 29513
0 29515 5 1 1 29514
0 29516 7 2 2 87869 92220
0 29517 7 1 2 64335 90067
0 29518 7 1 2 92241 29517
0 29519 5 1 1 29518
0 29520 7 1 2 29515 29519
0 29521 5 1 1 29520
0 29522 7 1 2 88336 29521
0 29523 5 1 1 29522
0 29524 7 3 2 58862 77369
0 29525 7 1 2 84472 91209
0 29526 7 1 2 92243 29525
0 29527 7 1 2 92235 29526
0 29528 5 1 1 29527
0 29529 7 1 2 79167 72970
0 29530 7 1 2 88088 29529
0 29531 7 1 2 77671 88200
0 29532 7 1 2 29530 29531
0 29533 5 1 1 29532
0 29534 7 1 2 29528 29533
0 29535 5 1 1 29534
0 29536 7 1 2 63499 29535
0 29537 5 1 1 29536
0 29538 7 1 2 76059 83553
0 29539 7 1 2 89167 29538
0 29540 7 1 2 92238 29539
0 29541 5 1 1 29540
0 29542 7 1 2 29537 29541
0 29543 5 1 1 29542
0 29544 7 1 2 63303 29543
0 29545 5 1 1 29544
0 29546 7 1 2 67929 91114
0 29547 7 1 2 91316 29546
0 29548 7 1 2 92240 29547
0 29549 5 1 1 29548
0 29550 7 1 2 29545 29549
0 29551 5 1 1 29550
0 29552 7 1 2 63022 29551
0 29553 5 1 1 29552
0 29554 7 1 2 85374 89157
0 29555 7 1 2 92242 29554
0 29556 5 1 1 29555
0 29557 7 1 2 29553 29556
0 29558 7 1 2 29523 29557
0 29559 5 1 1 29558
0 29560 7 1 2 61643 29559
0 29561 5 1 1 29560
0 29562 7 1 2 80479 91684
0 29563 7 1 2 73094 84412
0 29564 5 2 1 29563
0 29565 7 1 2 65951 80541
0 29566 5 1 1 29565
0 29567 7 1 2 92246 29566
0 29568 7 1 2 29562 29567
0 29569 5 1 1 29568
0 29570 7 1 2 87890 29569
0 29571 5 1 1 29570
0 29572 7 1 2 87019 73363
0 29573 7 1 2 77628 29572
0 29574 5 1 1 29573
0 29575 7 2 2 62464 77429
0 29576 7 1 2 73500 86601
0 29577 7 1 2 92248 29576
0 29578 5 1 1 29577
0 29579 7 1 2 29574 29578
0 29580 5 1 1 29579
0 29581 7 1 2 66910 29580
0 29582 5 1 1 29581
0 29583 7 1 2 29571 29582
0 29584 5 1 1 29583
0 29585 7 1 2 86612 88526
0 29586 7 1 2 29584 29585
0 29587 5 1 1 29586
0 29588 7 1 2 29561 29587
0 29589 5 1 1 29588
0 29590 7 1 2 61835 29589
0 29591 5 1 1 29590
0 29592 7 1 2 87942 89168
0 29593 7 2 2 67752 80560
0 29594 5 1 1 92250
0 29595 7 1 2 91738 92251
0 29596 7 1 2 29592 29595
0 29597 5 1 1 29596
0 29598 7 1 2 86898 89232
0 29599 5 1 1 29598
0 29600 7 2 2 66472 68860
0 29601 7 1 2 64555 85645
0 29602 7 1 2 92252 29601
0 29603 5 1 1 29602
0 29604 7 1 2 29599 29603
0 29605 5 1 1 29604
0 29606 7 1 2 63304 29605
0 29607 5 1 1 29606
0 29608 7 1 2 87822 91140
0 29609 5 1 1 29608
0 29610 7 1 2 29607 29609
0 29611 5 1 1 29610
0 29612 7 2 2 61957 77672
0 29613 7 1 2 90944 92254
0 29614 7 1 2 29611 29613
0 29615 5 1 1 29614
0 29616 7 1 2 29597 29615
0 29617 5 1 1 29616
0 29618 7 1 2 66911 29617
0 29619 5 1 1 29618
0 29620 7 4 2 66473 67753
0 29621 5 1 1 92256
0 29622 7 2 2 86523 87943
0 29623 7 1 2 85383 88133
0 29624 7 1 2 92260 29623
0 29625 5 1 1 29624
0 29626 7 1 2 84574 79923
0 29627 7 1 2 87827 29626
0 29628 7 1 2 90945 29627
0 29629 5 1 1 29628
0 29630 7 1 2 29625 29629
0 29631 5 1 1 29630
0 29632 7 1 2 92257 29631
0 29633 5 1 1 29632
0 29634 7 9 2 61836 66839
0 29635 5 1 1 92262
0 29636 7 5 2 61644 75541
0 29637 7 1 2 86265 88337
0 29638 7 1 2 92271 29637
0 29639 7 1 2 92255 29638
0 29640 5 1 1 29639
0 29641 7 1 2 63023 72903
0 29642 7 1 2 91927 29641
0 29643 5 1 1 29642
0 29644 7 1 2 64336 92054
0 29645 5 1 1 29644
0 29646 7 1 2 92247 29645
0 29647 7 1 2 29643 29646
0 29648 5 1 1 29647
0 29649 7 1 2 86613 92215
0 29650 7 1 2 29648 29649
0 29651 5 1 1 29650
0 29652 7 1 2 29640 29651
0 29653 5 1 1 29652
0 29654 7 1 2 92263 29653
0 29655 5 1 1 29654
0 29656 7 1 2 29633 29655
0 29657 7 1 2 29619 29656
0 29658 5 1 1 29657
0 29659 7 1 2 70516 29658
0 29660 5 1 1 29659
0 29661 7 1 2 91754 92261
0 29662 5 1 1 29661
0 29663 7 1 2 71285 77241
0 29664 7 1 2 87621 29663
0 29665 5 1 1 29664
0 29666 7 1 2 29662 29665
0 29667 5 1 1 29666
0 29668 7 1 2 63305 29667
0 29669 5 1 1 29668
0 29670 7 1 2 90973 91835
0 29671 7 1 2 91328 29670
0 29672 5 1 1 29671
0 29673 7 1 2 29669 29672
0 29674 5 1 1 29673
0 29675 7 1 2 88527 92258
0 29676 7 1 2 29674 29675
0 29677 5 1 1 29676
0 29678 7 1 2 29660 29677
0 29679 7 1 2 29591 29678
0 29680 5 1 1 29679
0 29681 7 1 2 62102 29680
0 29682 5 1 1 29681
0 29683 7 1 2 29469 29682
0 29684 5 1 1 29683
0 29685 7 1 2 92209 29684
0 29686 5 1 1 29685
0 29687 7 1 2 70780 73626
0 29688 5 3 1 29687
0 29689 7 1 2 89530 92276
0 29690 5 1 1 29689
0 29691 7 1 2 64088 78234
0 29692 5 1 1 29691
0 29693 7 1 2 88434 29692
0 29694 5 1 1 29693
0 29695 7 1 2 90917 29694
0 29696 5 1 1 29695
0 29697 7 1 2 90148 90506
0 29698 5 1 1 29697
0 29699 7 1 2 29696 29698
0 29700 5 1 1 29699
0 29701 7 1 2 63715 29700
0 29702 5 1 1 29701
0 29703 7 1 2 75401 89107
0 29704 5 1 1 29703
0 29705 7 1 2 29702 29704
0 29706 5 1 1 29705
0 29707 7 1 2 82207 29706
0 29708 5 1 1 29707
0 29709 7 2 2 61645 88507
0 29710 7 1 2 89017 90918
0 29711 7 1 2 92279 29710
0 29712 5 1 1 29711
0 29713 7 1 2 29708 29712
0 29714 5 1 1 29713
0 29715 7 1 2 64337 29714
0 29716 5 1 1 29715
0 29717 7 1 2 64556 88379
0 29718 7 2 2 92280 29717
0 29719 7 1 2 71182 92281
0 29720 5 1 1 29719
0 29721 7 1 2 29716 29720
0 29722 5 1 1 29721
0 29723 7 1 2 63306 29722
0 29724 5 1 1 29723
0 29725 7 1 2 89847 92282
0 29726 5 1 1 29725
0 29727 7 1 2 29724 29726
0 29728 5 1 1 29727
0 29729 7 1 2 88707 29728
0 29730 5 1 1 29729
0 29731 7 3 2 66265 90022
0 29732 7 1 2 88024 92283
0 29733 5 1 1 29732
0 29734 7 1 2 86290 89822
0 29735 5 1 1 29734
0 29736 7 1 2 29733 29735
0 29737 5 1 1 29736
0 29738 7 2 2 63716 59370
0 29739 7 1 2 91311 92286
0 29740 7 1 2 29737 29739
0 29741 5 1 1 29740
0 29742 7 1 2 29730 29741
0 29743 5 1 1 29742
0 29744 7 1 2 69554 29743
0 29745 5 1 1 29744
0 29746 7 3 2 67479 89595
0 29747 7 1 2 69217 80958
0 29748 7 1 2 92288 29747
0 29749 7 1 2 91581 29748
0 29750 5 1 1 29749
0 29751 7 1 2 29745 29750
0 29752 5 1 1 29751
0 29753 7 1 2 66912 29752
0 29754 5 1 1 29753
0 29755 7 1 2 79288 89089
0 29756 5 1 1 29755
0 29757 7 1 2 89247 29756
0 29758 5 1 1 29757
0 29759 7 1 2 57710 29758
0 29760 5 1 1 29759
0 29761 7 2 2 61837 71740
0 29762 7 1 2 76647 92291
0 29763 5 1 1 29762
0 29764 7 1 2 62465 89186
0 29765 7 1 2 91242 29764
0 29766 5 1 1 29765
0 29767 7 1 2 89248 29766
0 29768 5 1 1 29767
0 29769 7 1 2 57424 29768
0 29770 5 1 1 29769
0 29771 7 1 2 29763 29770
0 29772 7 1 2 29760 29771
0 29773 5 1 1 29772
0 29774 7 1 2 81553 29773
0 29775 5 1 1 29774
0 29776 7 1 2 88188 89090
0 29777 5 1 1 29776
0 29778 7 1 2 89249 29777
0 29779 5 1 1 29778
0 29780 7 1 2 84058 29779
0 29781 5 1 1 29780
0 29782 7 1 2 29775 29781
0 29783 5 1 1 29782
0 29784 7 1 2 58046 29783
0 29785 5 1 1 29784
0 29786 7 1 2 68621 84059
0 29787 5 1 1 29786
0 29788 7 1 2 68778 81554
0 29789 5 1 1 29788
0 29790 7 1 2 29787 29789
0 29791 5 1 1 29790
0 29792 7 1 2 61838 85761
0 29793 7 1 2 74055 29792
0 29794 7 1 2 29791 29793
0 29795 5 1 1 29794
0 29796 7 1 2 29785 29795
0 29797 5 1 1 29796
0 29798 7 1 2 83675 29797
0 29799 5 1 1 29798
0 29800 7 1 2 88195 89923
0 29801 5 1 1 29800
0 29802 7 1 2 88445 90189
0 29803 5 1 1 29802
0 29804 7 1 2 29801 29803
0 29805 5 1 1 29804
0 29806 7 1 2 88957 29805
0 29807 5 1 1 29806
0 29808 7 1 2 74814 79842
0 29809 5 1 1 29808
0 29810 7 1 2 59371 78188
0 29811 5 1 1 29810
0 29812 7 1 2 29809 29811
0 29813 5 1 1 29812
0 29814 7 1 2 57425 29813
0 29815 5 1 1 29814
0 29816 7 1 2 58980 81484
0 29817 5 1 1 29816
0 29818 7 1 2 59372 88426
0 29819 5 1 1 29818
0 29820 7 1 2 29817 29819
0 29821 7 1 2 29815 29820
0 29822 5 1 1 29821
0 29823 7 1 2 90190 29822
0 29824 5 1 1 29823
0 29825 7 1 2 29807 29824
0 29826 5 1 1 29825
0 29827 7 1 2 77272 29826
0 29828 5 1 1 29827
0 29829 7 2 2 61646 88918
0 29830 7 1 2 85979 74422
0 29831 7 1 2 92293 29830
0 29832 5 1 1 29831
0 29833 7 1 2 29828 29832
0 29834 5 1 1 29833
0 29835 7 1 2 76746 29834
0 29836 5 1 1 29835
0 29837 7 1 2 85076 76051
0 29838 7 2 2 60007 60383
0 29839 7 3 2 64557 92295
0 29840 7 1 2 89611 92297
0 29841 7 1 2 29837 29840
0 29842 5 1 1 29841
0 29843 7 1 2 88958 89273
0 29844 5 1 1 29843
0 29845 7 1 2 74613 89241
0 29846 5 1 1 29845
0 29847 7 1 2 29844 29846
0 29848 5 1 1 29847
0 29849 7 1 2 75766 82396
0 29850 7 1 2 29848 29849
0 29851 5 1 1 29850
0 29852 7 1 2 29842 29851
0 29853 5 1 1 29852
0 29854 7 1 2 68861 29853
0 29855 5 1 1 29854
0 29856 7 1 2 81555 92129
0 29857 5 1 1 29856
0 29858 7 1 2 84060 88189
0 29859 5 1 1 29858
0 29860 7 1 2 29857 29859
0 29861 5 1 1 29860
0 29862 7 1 2 77295 29861
0 29863 5 1 1 29862
0 29864 7 1 2 75660 91649
0 29865 5 1 1 29864
0 29866 7 1 2 29863 29865
0 29867 5 1 1 29866
0 29868 7 1 2 89091 29867
0 29869 5 1 1 29868
0 29870 7 1 2 81556 88432
0 29871 5 1 1 29870
0 29872 7 1 2 58047 71011
0 29873 5 2 1 29872
0 29874 7 1 2 84061 92300
0 29875 5 1 1 29874
0 29876 7 1 2 29871 29875
0 29877 5 1 1 29876
0 29878 7 1 2 89192 29877
0 29879 5 1 1 29878
0 29880 7 1 2 29869 29879
0 29881 5 1 1 29880
0 29882 7 1 2 59373 29881
0 29883 5 1 1 29882
0 29884 7 1 2 29855 29883
0 29885 7 1 2 29836 29884
0 29886 7 1 2 29799 29885
0 29887 5 1 1 29886
0 29888 7 1 2 69272 29887
0 29889 5 1 1 29888
0 29890 7 1 2 79146 79262
0 29891 7 1 2 92289 29890
0 29892 5 1 1 29891
0 29893 7 1 2 64558 86332
0 29894 7 1 2 81979 29893
0 29895 7 1 2 90228 29894
0 29896 5 1 1 29895
0 29897 7 1 2 29892 29896
0 29898 5 1 1 29897
0 29899 7 1 2 58558 29898
0 29900 5 1 1 29899
0 29901 7 1 2 66474 74772
0 29902 7 8 2 58981 64559
0 29903 5 1 1 92302
0 29904 7 2 2 57426 92303
0 29905 5 1 1 92310
0 29906 7 1 2 81980 29905
0 29907 7 1 2 29901 29906
0 29908 7 1 2 88618 29907
0 29909 5 1 1 29908
0 29910 7 1 2 29900 29909
0 29911 5 1 1 29910
0 29912 7 1 2 60384 29911
0 29913 5 1 1 29912
0 29914 7 2 2 87531 79448
0 29915 7 1 2 84455 75809
0 29916 7 1 2 90229 29915
0 29917 7 1 2 92312 29916
0 29918 5 1 1 29917
0 29919 7 1 2 29913 29918
0 29920 5 1 1 29919
0 29921 7 1 2 64338 29920
0 29922 5 1 1 29921
0 29923 7 1 2 74773 81529
0 29924 7 2 2 73723 83663
0 29925 7 1 2 89728 92314
0 29926 7 1 2 29923 29925
0 29927 5 1 1 29926
0 29928 7 1 2 29922 29927
0 29929 5 1 1 29928
0 29930 7 1 2 70517 29929
0 29931 5 1 1 29930
0 29932 7 1 2 66784 69218
0 29933 7 1 2 76085 29932
0 29934 7 1 2 89918 91673
0 29935 7 1 2 29933 29934
0 29936 5 1 1 29935
0 29937 7 1 2 29931 29936
0 29938 7 1 2 29889 29937
0 29939 5 1 1 29938
0 29940 7 1 2 64899 29939
0 29941 5 1 1 29940
0 29942 7 2 2 89300 92290
0 29943 7 1 2 79494 90507
0 29944 7 1 2 89304 29943
0 29945 7 1 2 92316 29944
0 29946 5 1 1 29945
0 29947 7 1 2 29941 29946
0 29948 5 1 1 29947
0 29949 7 1 2 63717 29948
0 29950 5 1 1 29949
0 29951 7 2 2 58916 64339
0 29952 7 1 2 85340 92318
0 29953 7 1 2 87906 29952
0 29954 7 1 2 92317 29953
0 29955 5 1 1 29954
0 29956 7 1 2 29950 29955
0 29957 7 1 2 29754 29956
0 29958 5 1 1 29957
0 29959 7 1 2 29690 29958
0 29960 5 1 1 29959
0 29961 7 1 2 29686 29960
0 29962 7 1 2 29438 29961
0 29963 7 1 2 29058 29962
0 29964 7 1 2 66840 88756
0 29965 5 1 1 29964
0 29966 7 2 2 60198 86056
0 29967 5 1 1 92320
0 29968 7 1 2 29965 29967
0 29969 5 3 1 29968
0 29970 7 3 2 58559 91141
0 29971 5 1 1 92325
0 29972 7 1 2 69032 92326
0 29973 5 1 1 29972
0 29974 7 3 2 63024 86830
0 29975 7 1 2 91711 92328
0 29976 5 1 1 29975
0 29977 7 1 2 29973 29976
0 29978 5 1 1 29977
0 29979 7 1 2 62204 29978
0 29980 5 1 1 29979
0 29981 7 1 2 71683 92327
0 29982 5 1 1 29981
0 29983 7 1 2 29980 29982
0 29984 5 1 1 29983
0 29985 7 1 2 72092 29984
0 29986 5 1 1 29985
0 29987 7 1 2 63307 89508
0 29988 7 1 2 72765 29987
0 29989 5 1 1 29988
0 29990 7 1 2 29971 29989
0 29991 5 1 1 29990
0 29992 7 1 2 63025 29991
0 29993 5 1 1 29992
0 29994 7 1 2 29986 29993
0 29995 5 1 1 29994
0 29996 7 1 2 64340 29995
0 29997 5 1 1 29996
0 29998 7 1 2 84861 80561
0 29999 5 2 1 29998
0 30000 7 1 2 85751 87733
0 30001 5 1 1 30000
0 30002 7 1 2 92331 30001
0 30003 5 1 1 30002
0 30004 7 1 2 78855 30003
0 30005 5 1 1 30004
0 30006 7 1 2 63026 87050
0 30007 5 1 1 30006
0 30008 7 1 2 30005 30007
0 30009 5 1 1 30008
0 30010 7 1 2 61839 30009
0 30011 5 1 1 30010
0 30012 7 1 2 29997 30011
0 30013 5 1 1 30012
0 30014 7 1 2 59842 30013
0 30015 5 1 1 30014
0 30016 7 2 2 85061 87066
0 30017 5 1 1 92333
0 30018 7 1 2 59596 85062
0 30019 5 1 1 30018
0 30020 7 1 2 65608 80381
0 30021 5 1 1 30020
0 30022 7 1 2 30019 30021
0 30023 5 1 1 30022
0 30024 7 1 2 61327 30023
0 30025 5 1 1 30024
0 30026 7 1 2 65952 78032
0 30027 5 1 1 30026
0 30028 7 1 2 30025 30027
0 30029 5 3 1 30028
0 30030 7 1 2 63308 92335
0 30031 5 1 1 30030
0 30032 7 1 2 30017 30031
0 30033 5 1 1 30032
0 30034 7 1 2 89265 30033
0 30035 5 1 1 30034
0 30036 7 1 2 30015 30035
0 30037 5 1 1 30036
0 30038 7 1 2 92322 30037
0 30039 5 1 1 30038
0 30040 7 1 2 89425 88757
0 30041 7 1 2 92336 30040
0 30042 5 1 1 30041
0 30043 7 2 2 78856 70518
0 30044 7 1 2 87894 90482
0 30045 7 1 2 92338 30044
0 30046 5 1 1 30045
0 30047 7 1 2 30042 30046
0 30048 5 1 1 30047
0 30049 7 1 2 58560 30048
0 30050 5 1 1 30049
0 30051 7 2 2 63309 72093
0 30052 7 1 2 89723 92340
0 30053 5 1 1 30052
0 30054 7 1 2 79531 87322
0 30055 5 1 1 30054
0 30056 7 1 2 30053 30055
0 30057 5 1 1 30056
0 30058 7 1 2 63027 30057
0 30059 5 1 1 30058
0 30060 7 1 2 73071 85719
0 30061 5 2 1 30060
0 30062 7 1 2 64560 92341
0 30063 7 1 2 92342 30062
0 30064 5 1 1 30063
0 30065 7 1 2 30059 30064
0 30066 5 1 1 30065
0 30067 7 1 2 92339 30066
0 30068 5 1 1 30067
0 30069 7 1 2 84585 91845
0 30070 5 1 1 30069
0 30071 7 1 2 30068 30070
0 30072 5 1 1 30071
0 30073 7 1 2 88771 30072
0 30074 5 1 1 30073
0 30075 7 1 2 30050 30074
0 30076 5 1 1 30075
0 30077 7 1 2 66913 30076
0 30078 5 1 1 30077
0 30079 7 1 2 30039 30078
0 30080 5 1 1 30079
0 30081 7 1 2 62103 30080
0 30082 5 1 1 30081
0 30083 7 2 2 62104 87835
0 30084 7 2 2 88946 92344
0 30085 7 1 2 88045 92346
0 30086 5 1 1 30085
0 30087 7 1 2 66841 92347
0 30088 5 1 1 30087
0 30089 7 1 2 86669 79941
0 30090 7 2 2 89476 30089
0 30091 7 1 2 63310 80516
0 30092 7 1 2 92348 30091
0 30093 5 1 1 30092
0 30094 7 1 2 30088 30093
0 30095 5 1 1 30094
0 30096 7 1 2 63028 85208
0 30097 7 1 2 30095 30096
0 30098 5 1 1 30097
0 30099 7 1 2 30086 30098
0 30100 5 1 1 30099
0 30101 7 1 2 62205 30100
0 30102 5 1 1 30101
0 30103 7 1 2 60008 80786
0 30104 5 1 1 30103
0 30105 7 1 2 87167 30104
0 30106 5 1 1 30105
0 30107 7 1 2 58748 30106
0 30108 5 1 1 30107
0 30109 7 5 2 63500 79263
0 30110 5 3 1 92350
0 30111 7 1 2 58561 92351
0 30112 5 1 1 30111
0 30113 7 1 2 30108 30112
0 30114 5 2 1 30113
0 30115 7 1 2 79278 92345
0 30116 7 1 2 92358 30115
0 30117 5 1 1 30116
0 30118 7 3 2 64821 90139
0 30119 7 1 2 69033 92360
0 30120 7 1 2 90952 30119
0 30121 5 1 1 30120
0 30122 7 1 2 30117 30121
0 30123 5 1 1 30122
0 30124 7 1 2 60592 30123
0 30125 5 1 1 30124
0 30126 7 1 2 30102 30125
0 30127 5 1 1 30126
0 30128 7 1 2 58863 30127
0 30129 5 1 1 30128
0 30130 7 1 2 66914 90023
0 30131 5 1 1 30130
0 30132 7 1 2 18565 30131
0 30133 5 1 1 30132
0 30134 7 1 2 64822 30133
0 30135 5 1 1 30134
0 30136 7 3 2 60133 86670
0 30137 7 1 2 90949 92363
0 30138 5 1 1 30137
0 30139 7 1 2 30135 30138
0 30140 5 1 1 30139
0 30141 7 1 2 63632 90140
0 30142 7 1 2 79082 30141
0 30143 7 1 2 30140 30142
0 30144 5 1 1 30143
0 30145 7 1 2 30129 30144
0 30146 5 1 1 30145
0 30147 7 1 2 64900 30146
0 30148 5 1 1 30147
0 30149 7 1 2 64823 92359
0 30150 5 1 1 30149
0 30151 7 1 2 85201 80787
0 30152 5 1 1 30151
0 30153 7 1 2 30150 30152
0 30154 5 1 1 30153
0 30155 7 1 2 63633 30154
0 30156 5 1 1 30155
0 30157 7 1 2 80788 88286
0 30158 5 1 1 30157
0 30159 7 1 2 30156 30158
0 30160 5 1 1 30159
0 30161 7 1 2 88948 90838
0 30162 7 1 2 30160 30161
0 30163 5 1 1 30162
0 30164 7 1 2 30148 30163
0 30165 5 1 1 30164
0 30166 7 1 2 65609 30165
0 30167 5 1 1 30166
0 30168 7 1 2 73512 91345
0 30169 5 1 1 30168
0 30170 7 1 2 76747 72869
0 30171 5 1 1 30170
0 30172 7 1 2 30169 30171
0 30173 5 1 1 30172
0 30174 7 1 2 86057 30173
0 30175 5 1 1 30174
0 30176 7 1 2 90293 91978
0 30177 5 1 1 30176
0 30178 7 1 2 30175 30177
0 30179 5 1 1 30178
0 30180 7 1 2 63029 30179
0 30181 5 1 1 30180
0 30182 7 1 2 70519 87845
0 30183 7 1 2 5007 30182
0 30184 7 1 2 91752 30183
0 30185 5 1 1 30184
0 30186 7 1 2 30181 30185
0 30187 5 1 1 30186
0 30188 7 1 2 60385 30187
0 30189 5 1 1 30188
0 30190 7 4 2 62206 71286
0 30191 5 1 1 92366
0 30192 7 3 2 63774 92367
0 30193 5 1 1 92370
0 30194 7 1 2 86058 90425
0 30195 7 1 2 92371 30194
0 30196 5 1 1 30195
0 30197 7 1 2 30189 30196
0 30198 5 1 1 30197
0 30199 7 1 2 60199 30198
0 30200 5 1 1 30199
0 30201 7 2 2 88758 88046
0 30202 5 1 1 92373
0 30203 7 1 2 78857 86899
0 30204 5 1 1 30203
0 30205 7 1 2 86626 30204
0 30206 5 1 1 30205
0 30207 7 1 2 92374 30206
0 30208 5 1 1 30207
0 30209 7 1 2 64341 87903
0 30210 7 1 2 83560 30209
0 30211 7 1 2 91838 30210
0 30212 5 1 1 30211
0 30213 7 1 2 30208 30212
0 30214 7 1 2 30200 30213
0 30215 5 1 1 30214
0 30216 7 1 2 80008 30215
0 30217 5 1 1 30216
0 30218 7 1 2 30167 30217
0 30219 5 1 1 30218
0 30220 7 1 2 63893 30219
0 30221 5 1 1 30220
0 30222 7 1 2 75542 92321
0 30223 5 1 1 30222
0 30224 7 1 2 30202 30223
0 30225 5 1 1 30224
0 30226 7 1 2 80267 90902
0 30227 7 1 2 30225 30226
0 30228 5 1 1 30227
0 30229 7 1 2 80973 92323
0 30230 5 1 1 30229
0 30231 7 1 2 73834 88759
0 30232 7 1 2 91840 30231
0 30233 5 1 1 30232
0 30234 7 1 2 30230 30233
0 30235 5 1 1 30234
0 30236 7 1 2 62207 76393
0 30237 5 2 1 30236
0 30238 7 1 2 80079 92375
0 30239 5 2 1 30238
0 30240 7 1 2 61328 92377
0 30241 7 1 2 30235 30240
0 30242 5 1 1 30241
0 30243 7 1 2 30228 30242
0 30244 5 1 1 30243
0 30245 7 1 2 62105 30244
0 30246 5 1 1 30245
0 30247 7 1 2 66475 30246
0 30248 7 1 2 30221 30247
0 30249 5 1 1 30248
0 30250 7 1 2 63030 85752
0 30251 5 1 1 30250
0 30252 7 1 2 58562 80997
0 30253 5 1 1 30252
0 30254 7 1 2 30251 30253
0 30255 5 1 1 30254
0 30256 7 1 2 65953 30255
0 30257 5 1 1 30256
0 30258 7 1 2 92332 30257
0 30259 5 2 1 30258
0 30260 7 1 2 92324 92379
0 30261 5 1 1 30260
0 30262 7 4 2 63775 86791
0 30263 5 1 1 92381
0 30264 7 1 2 71938 92382
0 30265 5 1 1 30264
0 30266 7 1 2 71498 30265
0 30267 5 1 1 30266
0 30268 7 2 2 60200 89370
0 30269 7 1 2 63311 80427
0 30270 7 1 2 92385 30269
0 30271 7 1 2 30267 30270
0 30272 5 1 1 30271
0 30273 7 1 2 30261 30272
0 30274 5 1 1 30273
0 30275 7 1 2 59843 30274
0 30276 5 1 1 30275
0 30277 7 1 2 63312 73095
0 30278 5 1 1 30277
0 30279 7 2 2 85769 86737
0 30280 5 4 1 92387
0 30281 7 1 2 63031 92389
0 30282 5 1 1 30281
0 30283 7 2 2 30278 30282
0 30284 5 1 1 92393
0 30285 7 1 2 60956 30284
0 30286 5 1 1 30285
0 30287 7 1 2 68514 74988
0 30288 7 1 2 90807 30287
0 30289 5 1 1 30288
0 30290 7 1 2 61329 23948
0 30291 7 1 2 30289 30290
0 30292 5 1 1 30291
0 30293 7 1 2 71821 90800
0 30294 7 1 2 30292 30293
0 30295 5 1 1 30294
0 30296 7 1 2 30286 30295
0 30297 5 1 1 30296
0 30298 7 1 2 64561 30297
0 30299 5 1 1 30298
0 30300 7 1 2 84191 73627
0 30301 7 1 2 87785 30300
0 30302 5 1 1 30301
0 30303 7 1 2 30299 30302
0 30304 5 1 1 30303
0 30305 7 1 2 92386 30304
0 30306 5 1 1 30305
0 30307 7 1 2 30276 30306
0 30308 5 1 1 30307
0 30309 7 1 2 62106 30308
0 30310 5 1 1 30309
0 30311 7 2 2 78647 91267
0 30312 7 1 2 89820 92395
0 30313 5 1 1 30312
0 30314 7 2 2 62208 86831
0 30315 7 1 2 80653 92397
0 30316 5 1 1 30315
0 30317 7 1 2 30313 30316
0 30318 5 1 1 30317
0 30319 7 1 2 79899 30318
0 30320 5 1 1 30319
0 30321 7 3 2 62209 75080
0 30322 7 2 2 73380 87576
0 30323 7 1 2 85090 92402
0 30324 7 1 2 92399 30323
0 30325 5 1 1 30324
0 30326 7 1 2 30320 30325
0 30327 5 1 1 30326
0 30328 7 1 2 70520 30327
0 30329 5 1 1 30328
0 30330 7 1 2 85546 71999
0 30331 7 1 2 82067 30330
0 30332 7 1 2 91570 30331
0 30333 5 1 1 30332
0 30334 7 1 2 30329 30333
0 30335 5 1 1 30334
0 30336 7 1 2 71425 88365
0 30337 7 1 2 30335 30336
0 30338 5 1 1 30337
0 30339 7 1 2 61840 30338
0 30340 7 1 2 30310 30339
0 30341 5 1 1 30340
0 30342 7 1 2 62466 30341
0 30343 7 1 2 30249 30342
0 30344 5 1 1 30343
0 30345 7 1 2 30082 30344
0 30346 5 1 1 30345
0 30347 7 1 2 63718 30346
0 30348 5 1 1 30347
0 30349 7 1 2 77731 87603
0 30350 5 1 1 30349
0 30351 7 1 2 71499 30350
0 30352 5 1 1 30351
0 30353 7 1 2 90426 30352
0 30354 5 1 1 30353
0 30355 7 1 2 79221 76676
0 30356 7 1 2 91568 30355
0 30357 5 1 1 30356
0 30358 7 1 2 78398 30357
0 30359 5 1 1 30358
0 30360 7 1 2 71822 30359
0 30361 5 1 1 30360
0 30362 7 2 2 60957 78162
0 30363 5 1 1 92404
0 30364 7 1 2 64562 92405
0 30365 5 1 1 30364
0 30366 7 1 2 30361 30365
0 30367 5 1 1 30366
0 30368 7 1 2 63776 30367
0 30369 5 1 1 30368
0 30370 7 1 2 84862 91361
0 30371 5 1 1 30370
0 30372 7 1 2 30369 30371
0 30373 5 1 1 30372
0 30374 7 1 2 62210 30373
0 30375 5 1 1 30374
0 30376 7 5 2 63032 77732
0 30377 5 1 1 92406
0 30378 7 1 2 85958 30377
0 30379 5 1 1 30378
0 30380 7 1 2 85331 30379
0 30381 5 1 1 30380
0 30382 7 4 2 60593 76677
0 30383 7 1 2 76992 92411
0 30384 7 1 2 92407 30383
0 30385 5 1 1 30384
0 30386 7 1 2 30381 30385
0 30387 5 1 1 30386
0 30388 7 1 2 64342 30387
0 30389 5 1 1 30388
0 30390 7 1 2 84863 78293
0 30391 5 1 1 30390
0 30392 7 1 2 75154 30391
0 30393 5 1 1 30392
0 30394 7 1 2 75543 30393
0 30395 5 1 1 30394
0 30396 7 1 2 30389 30395
0 30397 7 1 2 30375 30396
0 30398 5 1 1 30397
0 30399 7 1 2 61330 30398
0 30400 5 1 1 30399
0 30401 7 1 2 30354 30400
0 30402 5 1 1 30401
0 30403 7 1 2 61841 70456
0 30404 7 1 2 30402 30403
0 30405 5 1 1 30404
0 30406 7 2 2 68239 88949
0 30407 5 2 1 92415
0 30408 7 1 2 80385 92417
0 30409 5 1 1 30408
0 30410 7 1 2 65610 30409
0 30411 5 1 1 30410
0 30412 7 2 2 60958 75799
0 30413 5 1 1 92419
0 30414 7 1 2 9346 30413
0 30415 5 1 1 30414
0 30416 7 1 2 59597 30415
0 30417 5 1 1 30416
0 30418 7 1 2 30411 30417
0 30419 5 1 1 30418
0 30420 7 1 2 58563 88851
0 30421 7 1 2 30419 30420
0 30422 5 1 1 30421
0 30423 7 1 2 84278 84043
0 30424 5 1 1 30423
0 30425 7 1 2 71500 30424
0 30426 5 1 1 30425
0 30427 7 1 2 63777 30426
0 30428 5 1 1 30427
0 30429 7 1 2 85980 30428
0 30430 5 1 1 30429
0 30431 7 1 2 62211 30430
0 30432 5 1 1 30431
0 30433 7 1 2 71426 78294
0 30434 5 1 1 30433
0 30435 7 1 2 30432 30434
0 30436 5 1 1 30435
0 30437 7 1 2 85496 91319
0 30438 7 1 2 30436 30437
0 30439 5 1 1 30438
0 30440 7 1 2 30422 30439
0 30441 5 1 1 30440
0 30442 7 1 2 59844 30441
0 30443 5 1 1 30442
0 30444 7 2 2 63894 85150
0 30445 7 1 2 60594 77733
0 30446 7 1 2 92421 30445
0 30447 5 1 1 30446
0 30448 7 1 2 80823 30447
0 30449 5 1 1 30448
0 30450 7 1 2 65611 30449
0 30451 5 1 1 30450
0 30452 7 1 2 91643 91048
0 30453 5 2 1 30452
0 30454 7 2 2 71823 75485
0 30455 5 1 1 92425
0 30456 7 1 2 91647 92426
0 30457 5 1 1 30456
0 30458 7 1 2 91641 30457
0 30459 5 1 1 30458
0 30460 7 1 2 60959 78839
0 30461 7 1 2 30459 30460
0 30462 5 1 1 30461
0 30463 7 1 2 92423 30462
0 30464 7 1 2 30451 30463
0 30465 5 1 1 30464
0 30466 7 1 2 64563 30465
0 30467 5 1 1 30466
0 30468 7 1 2 72799 78126
0 30469 7 1 2 92408 30468
0 30470 5 1 1 30469
0 30471 7 1 2 30467 30470
0 30472 5 1 1 30471
0 30473 7 1 2 91320 30472
0 30474 5 1 1 30473
0 30475 7 1 2 61331 30474
0 30476 7 1 2 30443 30475
0 30477 5 1 1 30476
0 30478 7 1 2 78118 89953
0 30479 5 1 1 30478
0 30480 7 1 2 28609 30479
0 30481 5 1 1 30480
0 30482 7 1 2 80268 30481
0 30483 5 1 1 30482
0 30484 7 1 2 71374 90564
0 30485 5 1 1 30484
0 30486 7 1 2 30483 30485
0 30487 5 1 1 30486
0 30488 7 1 2 87604 30487
0 30489 5 1 1 30488
0 30490 7 1 2 78033 89422
0 30491 5 1 1 30490
0 30492 7 1 2 71427 92068
0 30493 5 1 1 30492
0 30494 7 1 2 65954 30493
0 30495 7 1 2 30491 30494
0 30496 7 1 2 30489 30495
0 30497 5 1 1 30496
0 30498 7 1 2 63634 30497
0 30499 7 1 2 30477 30498
0 30500 5 1 1 30499
0 30501 7 1 2 30405 30500
0 30502 5 1 1 30501
0 30503 7 1 2 66915 30502
0 30504 5 1 1 30503
0 30505 7 2 2 86068 89233
0 30506 7 1 2 77734 92380
0 30507 5 1 1 30506
0 30508 7 1 2 85729 87020
0 30509 5 1 1 30508
0 30510 7 1 2 30507 30509
0 30511 5 1 1 30510
0 30512 7 1 2 92427 30511
0 30513 5 1 1 30512
0 30514 7 2 2 65612 88950
0 30515 5 2 1 92429
0 30516 7 1 2 80789 92430
0 30517 5 1 1 30516
0 30518 7 1 2 6479 30517
0 30519 5 1 1 30518
0 30520 7 1 2 63895 30519
0 30521 5 1 1 30520
0 30522 7 1 2 80974 92378
0 30523 5 1 1 30522
0 30524 7 1 2 30521 30523
0 30525 5 1 1 30524
0 30526 7 1 2 61332 30525
0 30527 5 1 1 30526
0 30528 7 1 2 80269 90427
0 30529 7 1 2 87605 30528
0 30530 5 1 1 30529
0 30531 7 1 2 30527 30530
0 30532 5 1 1 30531
0 30533 7 1 2 62467 30532
0 30534 5 1 1 30533
0 30535 7 1 2 64564 92334
0 30536 5 1 1 30535
0 30537 7 1 2 64565 92337
0 30538 5 1 1 30537
0 30539 7 1 2 85063 90654
0 30540 5 1 1 30539
0 30541 7 1 2 30538 30540
0 30542 5 1 1 30541
0 30543 7 1 2 63313 30542
0 30544 5 1 1 30543
0 30545 7 1 2 30536 30544
0 30546 7 1 2 30534 30545
0 30547 5 1 1 30546
0 30548 7 1 2 88894 30547
0 30549 5 1 1 30548
0 30550 7 1 2 30513 30549
0 30551 7 1 2 30504 30550
0 30552 5 1 1 30551
0 30553 7 1 2 89108 30552
0 30554 5 1 1 30553
0 30555 7 1 2 66266 30554
0 30556 7 1 2 30348 30555
0 30557 5 1 1 30556
0 30558 7 1 2 13185 88589
0 30559 5 1 1 30558
0 30560 7 1 2 79660 30559
0 30561 5 1 1 30560
0 30562 7 1 2 86942 88590
0 30563 5 1 1 30562
0 30564 7 1 2 76748 30563
0 30565 5 1 1 30564
0 30566 7 1 2 30561 30565
0 30567 5 1 1 30566
0 30568 7 1 2 91795 30567
0 30569 5 1 1 30568
0 30570 7 2 2 71684 88647
0 30571 5 1 1 92433
0 30572 7 2 2 60960 92434
0 30573 7 1 2 90321 92435
0 30574 5 1 1 30573
0 30575 7 1 2 73381 90631
0 30576 7 1 2 82134 30575
0 30577 5 1 1 30576
0 30578 7 1 2 30574 30577
0 30579 5 1 1 30578
0 30580 7 1 2 63033 30579
0 30581 5 1 1 30580
0 30582 7 2 2 64566 79453
0 30583 7 1 2 92436 92437
0 30584 5 1 1 30583
0 30585 7 4 2 63501 79825
0 30586 7 1 2 66476 72028
0 30587 7 1 2 92439 30586
0 30588 5 1 1 30587
0 30589 7 1 2 30584 30588
0 30590 5 1 1 30589
0 30591 7 1 2 63314 30590
0 30592 5 1 1 30591
0 30593 7 2 2 58564 83417
0 30594 5 1 1 92443
0 30595 7 2 2 73545 88663
0 30596 7 1 2 92444 92445
0 30597 5 1 1 30596
0 30598 7 1 2 30592 30597
0 30599 7 1 2 30581 30598
0 30600 5 1 1 30599
0 30601 7 1 2 62212 30600
0 30602 5 1 1 30601
0 30603 7 1 2 30569 30602
0 30604 5 1 1 30603
0 30605 7 1 2 62468 30604
0 30606 5 1 1 30605
0 30607 7 4 2 90103 91421
0 30608 5 1 1 92447
0 30609 7 1 2 70091 92448
0 30610 5 1 1 30609
0 30611 7 5 2 66477 76922
0 30612 7 1 2 79826 77099
0 30613 7 1 2 92451 30612
0 30614 5 1 1 30613
0 30615 7 1 2 30610 30614
0 30616 5 1 1 30615
0 30617 7 1 2 71428 30616
0 30618 5 1 1 30617
0 30619 7 1 2 77511 90181
0 30620 7 1 2 91268 30619
0 30621 5 1 1 30620
0 30622 7 1 2 30618 30621
0 30623 7 1 2 30606 30622
0 30624 5 1 1 30623
0 30625 7 1 2 89139 30624
0 30626 5 1 1 30625
0 30627 7 1 2 58749 88366
0 30628 7 1 2 88648 30627
0 30629 7 1 2 86634 91376
0 30630 7 1 2 30628 30629
0 30631 5 1 1 30630
0 30632 7 1 2 87163 90182
0 30633 7 1 2 92400 30632
0 30634 5 1 1 30633
0 30635 7 1 2 30608 30634
0 30636 5 1 1 30635
0 30637 7 1 2 85923 88581
0 30638 7 1 2 30636 30637
0 30639 5 1 1 30638
0 30640 7 1 2 30631 30639
0 30641 5 1 1 30640
0 30642 7 1 2 71429 30641
0 30643 5 1 1 30642
0 30644 7 1 2 30626 30643
0 30645 5 1 1 30644
0 30646 7 1 2 63896 30645
0 30647 5 1 1 30646
0 30648 7 2 2 77100 91796
0 30649 5 1 1 92456
0 30650 7 1 2 90524 92457
0 30651 7 1 2 91230 30650
0 30652 5 1 1 30651
0 30653 7 1 2 30647 30652
0 30654 5 1 1 30653
0 30655 7 1 2 60595 30654
0 30656 5 1 1 30655
0 30657 7 2 2 60961 75273
0 30658 5 2 1 92458
0 30659 7 1 2 59598 92459
0 30660 5 1 1 30659
0 30661 7 2 2 71287 77055
0 30662 5 1 1 92462
0 30663 7 1 2 76492 87126
0 30664 5 1 1 30663
0 30665 7 1 2 74548 30664
0 30666 5 1 1 30665
0 30667 7 1 2 62469 30666
0 30668 5 1 1 30667
0 30669 7 1 2 30662 30668
0 30670 7 1 2 30660 30669
0 30671 5 1 1 30670
0 30672 7 1 2 77822 30671
0 30673 5 1 1 30672
0 30674 7 2 2 85151 84629
0 30675 7 1 2 88943 92464
0 30676 5 1 1 30675
0 30677 7 2 2 60962 91644
0 30678 5 1 1 92466
0 30679 7 1 2 69034 92467
0 30680 5 1 1 30679
0 30681 7 1 2 30676 30680
0 30682 5 1 1 30681
0 30683 7 1 2 62213 30682
0 30684 5 1 1 30683
0 30685 7 1 2 63315 92463
0 30686 5 2 1 30685
0 30687 7 1 2 92424 92468
0 30688 7 1 2 30684 30687
0 30689 5 1 1 30688
0 30690 7 1 2 59845 30689
0 30691 5 1 1 30690
0 30692 7 1 2 30673 30691
0 30693 5 1 1 30692
0 30694 7 1 2 91797 30693
0 30695 5 1 1 30694
0 30696 7 1 2 71430 81589
0 30697 7 2 2 60963 74816
0 30698 5 2 1 92470
0 30699 7 1 2 57427 92472
0 30700 5 2 1 30699
0 30701 7 1 2 92449 92474
0 30702 7 1 2 30696 30701
0 30703 5 1 1 30702
0 30704 7 1 2 30695 30703
0 30705 5 1 1 30704
0 30706 7 1 2 89140 30705
0 30707 5 1 1 30706
0 30708 7 1 2 30656 30707
0 30709 5 1 1 30708
0 30710 7 1 2 63719 30709
0 30711 5 1 1 30710
0 30712 7 1 2 86356 92431
0 30713 5 1 1 30712
0 30714 7 1 2 79661 30713
0 30715 5 1 1 30714
0 30716 7 1 2 77578 92432
0 30717 5 1 1 30716
0 30718 7 1 2 76749 30717
0 30719 5 1 1 30718
0 30720 7 1 2 30715 30719
0 30721 5 1 1 30720
0 30722 7 1 2 63897 30721
0 30723 5 1 1 30722
0 30724 7 1 2 65613 91950
0 30725 5 4 1 30724
0 30726 7 1 2 91231 92476
0 30727 5 1 1 30726
0 30728 7 1 2 30723 30727
0 30729 5 1 1 30728
0 30730 7 1 2 62470 30729
0 30731 5 1 1 30730
0 30732 7 1 2 77056 91174
0 30733 5 1 1 30732
0 30734 7 1 2 72094 77101
0 30735 5 1 1 30734
0 30736 7 1 2 83573 30735
0 30737 5 1 1 30736
0 30738 7 1 2 91232 30737
0 30739 5 1 1 30738
0 30740 7 1 2 30733 30739
0 30741 7 1 2 30731 30740
0 30742 5 1 1 30741
0 30743 7 1 2 91798 30742
0 30744 5 1 1 30743
0 30745 7 1 2 72095 91508
0 30746 5 1 1 30745
0 30747 7 1 2 81847 30746
0 30748 5 1 1 30747
0 30749 7 1 2 64343 30748
0 30750 5 1 1 30749
0 30751 7 1 2 60386 81000
0 30752 5 1 1 30751
0 30753 7 1 2 30750 30752
0 30754 5 1 1 30753
0 30755 7 1 2 63034 30754
0 30756 5 1 1 30755
0 30757 7 2 2 76800 90586
0 30758 5 1 1 92480
0 30759 7 1 2 30756 30758
0 30760 5 1 1 30759
0 30761 7 1 2 92450 30760
0 30762 5 1 1 30761
0 30763 7 1 2 30744 30762
0 30764 5 1 1 30763
0 30765 7 1 2 89109 30764
0 30766 5 1 1 30765
0 30767 7 1 2 30711 30766
0 30768 5 1 1 30767
0 30769 7 1 2 61333 30768
0 30770 5 1 1 30769
0 30771 7 1 2 72096 87828
0 30772 5 1 1 30771
0 30773 7 1 2 79449 78129
0 30774 5 1 1 30773
0 30775 7 1 2 30772 30774
0 30776 5 1 1 30775
0 30777 7 1 2 68862 30776
0 30778 5 1 1 30777
0 30779 7 1 2 71824 77803
0 30780 5 2 1 30779
0 30781 7 1 2 68515 78113
0 30782 5 1 1 30781
0 30783 7 1 2 58565 72097
0 30784 5 1 1 30783
0 30785 7 1 2 30782 30784
0 30786 5 1 1 30785
0 30787 7 1 2 64567 30786
0 30788 5 1 1 30787
0 30789 7 1 2 92482 30788
0 30790 5 1 1 30789
0 30791 7 1 2 63035 30790
0 30792 5 1 1 30791
0 30793 7 1 2 3829 30792
0 30794 5 1 1 30793
0 30795 7 1 2 60387 30794
0 30796 5 1 1 30795
0 30797 7 1 2 30778 30796
0 30798 5 1 1 30797
0 30799 7 1 2 62471 30798
0 30800 5 1 1 30799
0 30801 7 1 2 71501 85058
0 30802 5 1 1 30801
0 30803 7 1 2 91175 30802
0 30804 5 1 1 30803
0 30805 7 1 2 30800 30804
0 30806 5 1 1 30805
0 30807 7 1 2 86040 88664
0 30808 7 1 2 30806 30807
0 30809 5 1 1 30808
0 30810 7 1 2 68516 77033
0 30811 7 1 2 89672 30810
0 30812 7 1 2 85384 90710
0 30813 7 1 2 30811 30812
0 30814 5 1 1 30813
0 30815 7 1 2 30809 30814
0 30816 5 1 1 30815
0 30817 7 1 2 88605 30816
0 30818 5 1 1 30817
0 30819 7 2 2 71771 73778
0 30820 5 1 1 92484
0 30821 7 1 2 12427 30820
0 30822 5 1 1 30821
0 30823 7 1 2 89141 30822
0 30824 5 1 1 30823
0 30825 7 1 2 69845 73050
0 30826 5 1 1 30825
0 30827 7 1 2 73779 78701
0 30828 5 1 1 30827
0 30829 7 1 2 30826 30828
0 30830 5 1 1 30829
0 30831 7 1 2 68517 30830
0 30832 5 1 1 30831
0 30833 7 1 2 69819 78483
0 30834 5 1 1 30833
0 30835 7 1 2 30832 30834
0 30836 5 1 1 30835
0 30837 7 1 2 68863 90540
0 30838 7 1 2 30836 30837
0 30839 5 1 1 30838
0 30840 7 1 2 30824 30839
0 30841 5 1 1 30840
0 30842 7 1 2 63898 30841
0 30843 5 1 1 30842
0 30844 7 1 2 74373 73051
0 30845 5 1 1 30844
0 30846 7 2 2 64344 75723
0 30847 5 1 1 92486
0 30848 7 1 2 65955 92487
0 30849 5 1 1 30848
0 30850 7 1 2 30845 30849
0 30851 5 1 1 30850
0 30852 7 1 2 89142 30851
0 30853 5 1 1 30852
0 30854 7 1 2 30843 30853
0 30855 5 1 1 30854
0 30856 7 1 2 60964 30855
0 30857 5 1 1 30856
0 30858 7 1 2 71894 78193
0 30859 5 1 1 30858
0 30860 7 2 2 81608 30859
0 30861 5 1 1 92488
0 30862 7 1 2 58304 30861
0 30863 5 1 1 30862
0 30864 7 1 2 73017 30863
0 30865 5 1 1 30864
0 30866 7 1 2 58305 83240
0 30867 5 2 1 30866
0 30868 7 1 2 73628 92490
0 30869 5 1 1 30868
0 30870 7 1 2 30865 30869
0 30871 5 1 1 30870
0 30872 7 1 2 89143 30871
0 30873 5 1 1 30872
0 30874 7 1 2 90541 91562
0 30875 7 1 2 78858 30874
0 30876 5 1 1 30875
0 30877 7 1 2 30873 30876
0 30878 7 1 2 30857 30877
0 30879 5 1 1 30878
0 30880 7 1 2 63720 30879
0 30881 5 1 1 30880
0 30882 7 2 2 65956 85959
0 30883 5 1 1 92492
0 30884 7 1 2 30847 92493
0 30885 5 1 1 30884
0 30886 7 1 2 85318 77539
0 30887 5 1 1 30886
0 30888 7 1 2 61334 30887
0 30889 5 1 1 30888
0 30890 7 1 2 60965 30889
0 30891 7 1 2 30885 30890
0 30892 5 1 1 30891
0 30893 7 1 2 85730 92491
0 30894 5 1 1 30893
0 30895 7 1 2 71614 86624
0 30896 5 1 1 30895
0 30897 7 1 2 30894 30896
0 30898 7 1 2 30892 30897
0 30899 5 1 1 30898
0 30900 7 1 2 89110 30899
0 30901 5 1 1 30900
0 30902 7 1 2 30881 30901
0 30903 5 1 1 30902
0 30904 7 1 2 76750 30903
0 30905 5 1 1 30904
0 30906 7 1 2 74374 80562
0 30907 5 1 1 30906
0 30908 7 1 2 63899 92485
0 30909 5 1 1 30908
0 30910 7 1 2 30907 30909
0 30911 5 1 1 30910
0 30912 7 1 2 64345 30911
0 30913 5 1 1 30912
0 30914 7 1 2 71030 86366
0 30915 5 1 1 30914
0 30916 7 1 2 86738 30915
0 30917 5 1 1 30916
0 30918 7 1 2 83083 30917
0 30919 5 1 1 30918
0 30920 7 1 2 30913 30919
0 30921 5 1 1 30920
0 30922 7 1 2 59846 30921
0 30923 5 1 1 30922
0 30924 7 1 2 74375 91454
0 30925 5 1 1 30924
0 30926 7 1 2 30923 30925
0 30927 5 1 1 30926
0 30928 7 1 2 60966 30927
0 30929 5 1 1 30928
0 30930 7 1 2 85605 92489
0 30931 5 1 1 30930
0 30932 7 1 2 71031 72000
0 30933 5 1 1 30932
0 30934 7 1 2 88229 30933
0 30935 5 1 1 30934
0 30936 7 1 2 90407 30935
0 30937 5 1 1 30936
0 30938 7 1 2 30931 30937
0 30939 7 1 2 30929 30938
0 30940 5 1 1 30939
0 30941 7 1 2 88606 30940
0 30942 5 1 1 30941
0 30943 7 1 2 72870 86285
0 30944 7 1 2 89169 30943
0 30945 7 1 2 90530 30944
0 30946 7 1 2 78348 30945
0 30947 5 1 1 30946
0 30948 7 1 2 30942 30947
0 30949 5 1 1 30948
0 30950 7 1 2 63036 30949
0 30951 5 1 1 30950
0 30952 7 1 2 80656 91559
0 30953 7 1 2 91906 30952
0 30954 7 1 2 88607 30953
0 30955 5 1 1 30954
0 30956 7 1 2 30951 30955
0 30957 7 1 2 30905 30956
0 30958 5 1 1 30957
0 30959 7 1 2 61842 30958
0 30960 5 1 1 30959
0 30961 7 1 2 75837 86341
0 30962 5 1 1 30961
0 30963 7 1 2 76814 30962
0 30964 5 1 1 30963
0 30965 7 1 2 60388 30964
0 30966 5 1 1 30965
0 30967 7 1 2 91432 30966
0 30968 5 1 1 30967
0 30969 7 1 2 88608 30968
0 30970 5 1 1 30969
0 30971 7 2 2 70926 87904
0 30972 7 1 2 63721 77492
0 30973 7 1 2 90531 30972
0 30974 7 1 2 92494 30973
0 30975 5 1 1 30974
0 30976 7 1 2 30970 30975
0 30977 5 1 1 30976
0 30978 7 1 2 80761 92059
0 30979 7 1 2 30977 30978
0 30980 5 1 1 30979
0 30981 7 1 2 30960 30980
0 30982 5 1 1 30981
0 30983 7 1 2 66916 30982
0 30984 5 1 1 30983
0 30985 7 1 2 30818 30984
0 30986 7 1 2 30770 30985
0 30987 5 1 1 30986
0 30988 7 1 2 70521 30987
0 30989 5 1 1 30988
0 30990 7 1 2 86080 74951
0 30991 5 1 1 30990
0 30992 7 1 2 86077 30991
0 30993 5 1 1 30992
0 30994 7 1 2 62214 30993
0 30995 5 1 1 30994
0 30996 7 1 2 72871 92471
0 30997 5 1 1 30996
0 30998 7 1 2 30995 30997
0 30999 5 1 1 30998
0 31000 7 1 2 63037 30999
0 31001 5 1 1 31000
0 31002 7 1 2 61335 92481
0 31003 5 1 1 31002
0 31004 7 1 2 31001 31003
0 31005 5 1 1 31004
0 31006 7 2 2 83664 88089
0 31007 7 1 2 88201 92496
0 31008 5 1 1 31007
0 31009 7 1 2 88338 89337
0 31010 5 1 1 31009
0 31011 7 1 2 31008 31010
0 31012 5 1 1 31011
0 31013 7 1 2 61843 31012
0 31014 7 1 2 31005 31013
0 31015 5 1 1 31014
0 31016 7 1 2 82068 88339
0 31017 5 1 1 31016
0 31018 7 1 2 25154 31017
0 31019 5 1 1 31018
0 31020 7 2 2 66478 31019
0 31021 7 1 2 91847 92416
0 31022 5 1 1 31021
0 31023 7 2 2 71655 83723
0 31024 5 1 1 92500
0 31025 7 1 2 77040 31024
0 31026 5 1 1 31025
0 31027 7 1 2 60596 31026
0 31028 5 1 1 31027
0 31029 7 1 2 59599 31028
0 31030 5 1 1 31029
0 31031 7 1 2 63038 31030
0 31032 5 1 1 31031
0 31033 7 1 2 77989 88174
0 31034 5 1 1 31033
0 31035 7 1 2 65957 31034
0 31036 7 1 2 31032 31035
0 31037 5 1 1 31036
0 31038 7 1 2 71288 69423
0 31039 5 1 1 31038
0 31040 7 1 2 92418 31039
0 31041 5 1 1 31040
0 31042 7 1 2 65614 31041
0 31043 5 1 1 31042
0 31044 7 1 2 83142 77574
0 31045 5 1 1 31044
0 31046 7 1 2 61336 31045
0 31047 7 1 2 31043 31046
0 31048 5 1 1 31047
0 31049 7 1 2 58566 31048
0 31050 7 1 2 31037 31049
0 31051 5 1 1 31050
0 31052 7 1 2 31022 31051
0 31053 5 1 1 31052
0 31054 7 1 2 92498 31053
0 31055 5 1 1 31054
0 31056 7 1 2 31015 31055
0 31057 5 1 1 31056
0 31058 7 1 2 64568 31057
0 31059 5 1 1 31058
0 31060 7 1 2 78045 88175
0 31061 5 1 1 31060
0 31062 7 1 2 71502 31061
0 31063 5 1 1 31062
0 31064 7 1 2 86726 31063
0 31065 5 1 1 31064
0 31066 7 1 2 69395 91645
0 31067 7 1 2 83143 31066
0 31068 5 1 1 31067
0 31069 7 1 2 88951 92465
0 31070 5 1 1 31069
0 31071 7 1 2 92469 31070
0 31072 7 1 2 31068 31071
0 31073 5 1 1 31072
0 31074 7 1 2 61337 31073
0 31075 5 1 1 31074
0 31076 7 1 2 31065 31075
0 31077 5 1 1 31076
0 31078 7 1 2 66842 89426
0 31079 7 1 2 88528 31078
0 31080 7 1 2 31077 31079
0 31081 5 1 1 31080
0 31082 7 1 2 31059 31081
0 31083 5 1 1 31082
0 31084 7 1 2 62107 31083
0 31085 5 1 1 31084
0 31086 7 1 2 27446 92483
0 31087 5 1 1 31086
0 31088 7 1 2 91459 31087
0 31089 5 1 1 31088
0 31090 7 1 2 79338 72872
0 31091 7 1 2 89456 31090
0 31092 5 1 1 31091
0 31093 7 1 2 31089 31092
0 31094 5 1 1 31093
0 31095 7 2 2 66843 87814
0 31096 7 1 2 31094 92502
0 31097 5 1 1 31096
0 31098 7 2 2 63900 79168
0 31099 7 1 2 79243 90565
0 31100 7 1 2 92504 31099
0 31101 7 1 2 90206 31100
0 31102 5 1 1 31101
0 31103 7 1 2 31097 31102
0 31104 5 1 1 31103
0 31105 7 1 2 88529 31104
0 31106 5 1 1 31105
0 31107 7 1 2 78484 79968
0 31108 7 1 2 88340 92505
0 31109 7 1 2 31107 31108
0 31110 5 1 1 31109
0 31111 7 1 2 58917 63901
0 31112 7 1 2 79859 31111
0 31113 7 1 2 83014 31112
0 31114 7 1 2 87866 31113
0 31115 5 1 1 31114
0 31116 7 1 2 31110 31115
0 31117 5 1 1 31116
0 31118 7 1 2 63316 88858
0 31119 7 1 2 31117 31118
0 31120 5 1 1 31119
0 31121 7 1 2 31106 31120
0 31122 5 1 1 31121
0 31123 7 1 2 63039 31122
0 31124 5 1 1 31123
0 31125 7 1 2 80428 84741
0 31126 5 1 1 31125
0 31127 7 1 2 68240 91944
0 31128 5 1 1 31127
0 31129 7 1 2 31126 31128
0 31130 5 1 1 31129
0 31131 7 1 2 90873 31130
0 31132 7 1 2 92499 31131
0 31133 5 1 1 31132
0 31134 7 1 2 31124 31133
0 31135 5 1 1 31134
0 31136 7 1 2 69035 31135
0 31137 5 1 1 31136
0 31138 7 2 2 63317 73780
0 31139 5 1 1 92506
0 31140 7 1 2 68199 92507
0 31141 5 1 1 31140
0 31142 7 1 2 16725 31141
0 31143 5 1 1 31142
0 31144 7 1 2 86583 31143
0 31145 5 1 1 31144
0 31146 7 1 2 72098 85446
0 31147 7 1 2 79776 31146
0 31148 5 1 1 31147
0 31149 7 1 2 86372 31148
0 31150 5 1 1 31149
0 31151 7 1 2 76751 31150
0 31152 5 1 1 31151
0 31153 7 1 2 31145 31152
0 31154 5 1 1 31153
0 31155 7 1 2 92503 31154
0 31156 5 1 1 31155
0 31157 7 3 2 64710 61844
0 31158 7 1 2 77396 76870
0 31159 7 1 2 92508 31158
0 31160 7 2 2 80429 87912
0 31161 7 1 2 86602 92511
0 31162 7 1 2 31159 31161
0 31163 5 1 1 31162
0 31164 7 1 2 31156 31163
0 31165 5 1 1 31164
0 31166 7 1 2 78295 88530
0 31167 7 1 2 31165 31166
0 31168 5 1 1 31167
0 31169 7 1 2 62215 88367
0 31170 7 1 2 90072 31169
0 31171 7 1 2 91326 31170
0 31172 7 1 2 84491 31171
0 31173 5 1 1 31172
0 31174 7 1 2 63040 90408
0 31175 5 1 1 31174
0 31176 7 1 2 28207 31175
0 31177 5 1 1 31176
0 31178 7 1 2 83084 88609
0 31179 7 1 2 89404 31178
0 31180 7 1 2 31177 31179
0 31181 5 1 1 31180
0 31182 7 1 2 31173 31181
0 31183 5 1 1 31182
0 31184 7 1 2 79900 31183
0 31185 5 1 1 31184
0 31186 7 1 2 68518 90073
0 31187 7 1 2 90822 31186
0 31188 7 1 2 92117 31187
0 31189 5 1 1 31188
0 31190 7 1 2 31185 31189
0 31191 5 1 1 31190
0 31192 7 1 2 88227 31191
0 31193 5 1 1 31192
0 31194 7 2 2 63722 66479
0 31195 7 1 2 69940 79244
0 31196 7 1 2 92513 31195
0 31197 7 1 2 90283 92495
0 31198 7 6 2 76648 66844
0 31199 7 2 2 63778 77897
0 31200 7 1 2 92515 92521
0 31201 7 1 2 31197 31200
0 31202 7 1 2 31196 31201
0 31203 5 1 1 31202
0 31204 7 1 2 61647 31203
0 31205 7 1 2 31193 31204
0 31206 7 1 2 31168 31205
0 31207 7 1 2 31137 31206
0 31208 7 1 2 31085 31207
0 31209 7 1 2 30989 31208
0 31210 5 1 1 31209
0 31211 7 1 2 30557 31210
0 31212 5 1 1 31211
0 31213 7 1 2 61958 31212
0 31214 5 1 1 31213
0 31215 7 2 2 79370 91039
0 31216 7 1 2 87969 89902
0 31217 7 1 2 92523 31216
0 31218 5 1 1 31217
0 31219 7 1 2 72727 87260
0 31220 7 1 2 90113 31219
0 31221 5 1 1 31220
0 31222 7 1 2 31218 31221
0 31223 5 1 1 31222
0 31224 7 1 2 58567 31223
0 31225 5 1 1 31224
0 31226 7 2 2 62472 87337
0 31227 5 1 1 92525
0 31228 7 1 2 87303 89828
0 31229 7 1 2 31227 31228
0 31230 5 1 1 31229
0 31231 7 1 2 63318 90114
0 31232 7 1 2 31230 31231
0 31233 5 1 1 31232
0 31234 7 1 2 31225 31233
0 31235 5 1 1 31234
0 31236 7 1 2 64901 31235
0 31237 5 1 1 31236
0 31238 7 1 2 72728 88012
0 31239 5 1 1 31238
0 31240 7 1 2 75544 91077
0 31241 5 1 1 31240
0 31242 7 1 2 31239 31241
0 31243 5 1 1 31242
0 31244 7 1 2 61845 87862
0 31245 7 1 2 31243 31244
0 31246 5 1 1 31245
0 31247 7 1 2 31237 31246
0 31248 5 1 1 31247
0 31249 7 1 2 64346 31248
0 31250 5 1 1 31249
0 31251 7 1 2 60597 91535
0 31252 5 1 1 31251
0 31253 7 2 2 62216 84456
0 31254 7 2 2 84184 91370
0 31255 5 1 1 92529
0 31256 7 1 2 92527 92530
0 31257 5 1 1 31256
0 31258 7 1 2 31252 31257
0 31259 5 1 1 31258
0 31260 7 1 2 60967 88764
0 31261 7 1 2 31259 31260
0 31262 5 1 1 31261
0 31263 7 1 2 31250 31262
0 31264 5 1 1 31263
0 31265 7 1 2 63723 31264
0 31266 5 1 1 31265
0 31267 7 3 2 61846 88093
0 31268 7 1 2 79982 91447
0 31269 5 1 1 31268
0 31270 7 1 2 89527 31269
0 31271 5 1 1 31270
0 31272 7 1 2 60389 31271
0 31273 5 1 1 31272
0 31274 7 2 2 79339 84312
0 31275 5 1 1 92534
0 31276 7 1 2 24117 31275
0 31277 5 1 1 31276
0 31278 7 1 2 70648 31277
0 31279 5 1 1 31278
0 31280 7 1 2 22913 31279
0 31281 7 1 2 31273 31280
0 31282 5 1 1 31281
0 31283 7 1 2 63319 31282
0 31284 5 1 1 31283
0 31285 7 1 2 59600 70322
0 31286 5 1 1 31285
0 31287 7 1 2 62473 31286
0 31288 5 1 1 31287
0 31289 7 2 2 72334 81670
0 31290 5 1 1 92536
0 31291 7 1 2 79503 31290
0 31292 7 1 2 31288 31291
0 31293 5 1 1 31292
0 31294 7 1 2 88612 31293
0 31295 5 1 1 31294
0 31296 7 1 2 31284 31295
0 31297 5 1 1 31296
0 31298 7 1 2 92531 31297
0 31299 5 1 1 31298
0 31300 7 1 2 31266 31299
0 31301 5 1 1 31300
0 31302 7 1 2 65958 31301
0 31303 5 1 1 31302
0 31304 7 1 2 87329 82539
0 31305 5 1 1 31304
0 31306 7 1 2 68519 77990
0 31307 7 1 2 91805 31306
0 31308 5 1 1 31307
0 31309 7 1 2 31305 31308
0 31310 5 1 1 31309
0 31311 7 1 2 61338 90998
0 31312 7 1 2 88531 31311
0 31313 7 1 2 31310 31312
0 31314 5 1 1 31313
0 31315 7 1 2 31303 31314
0 31316 5 1 1 31315
0 31317 7 1 2 63041 31316
0 31318 5 1 1 31317
0 31319 7 4 2 74338 89694
0 31320 5 1 1 92538
0 31321 7 1 2 75545 92539
0 31322 5 1 1 31321
0 31323 7 5 2 62217 61339
0 31324 5 1 1 92542
0 31325 7 1 2 81671 92543
0 31326 7 1 2 90780 31325
0 31327 5 1 1 31326
0 31328 7 1 2 31322 31327
0 31329 5 1 1 31328
0 31330 7 1 2 88532 91628
0 31331 7 1 2 31329 31330
0 31332 5 1 1 31331
0 31333 7 1 2 31318 31332
0 31334 5 1 1 31333
0 31335 7 1 2 66917 31334
0 31336 5 1 1 31335
0 31337 7 1 2 87891 88533
0 31338 5 1 1 31337
0 31339 7 1 2 79952 92216
0 31340 5 1 1 31339
0 31341 7 1 2 31338 31340
0 31342 5 2 1 31341
0 31343 7 1 2 78405 86593
0 31344 5 1 1 31343
0 31345 7 1 2 86256 31344
0 31346 5 1 1 31345
0 31347 7 1 2 66267 31346
0 31348 5 1 1 31347
0 31349 7 2 2 61648 72475
0 31350 7 1 2 85828 92549
0 31351 5 1 1 31350
0 31352 7 1 2 31348 31351
0 31353 5 1 1 31352
0 31354 7 1 2 61847 31353
0 31355 5 1 1 31354
0 31356 7 3 2 75264 91159
0 31357 7 1 2 78571 86650
0 31358 7 1 2 92551 31357
0 31359 5 1 1 31358
0 31360 7 1 2 31355 31359
0 31361 5 1 1 31360
0 31362 7 1 2 92547 31361
0 31363 5 1 1 31362
0 31364 7 1 2 88047 91817
0 31365 5 1 1 31364
0 31366 7 3 2 66268 74907
0 31367 5 1 1 92554
0 31368 7 1 2 92253 92315
0 31369 7 1 2 92555 31368
0 31370 5 1 1 31369
0 31371 7 1 2 31365 31370
0 31372 5 1 1 31371
0 31373 7 1 2 61340 31372
0 31374 5 1 1 31373
0 31375 7 1 2 70092 88871
0 31376 5 1 1 31375
0 31377 7 1 2 30649 31376
0 31378 5 1 1 31377
0 31379 7 1 2 91060 31378
0 31380 5 1 1 31379
0 31381 7 1 2 75274 91799
0 31382 5 1 1 31381
0 31383 7 1 2 20155 31382
0 31384 5 1 1 31383
0 31385 7 1 2 61649 87739
0 31386 7 1 2 31384 31385
0 31387 5 1 1 31386
0 31388 7 1 2 31380 31387
0 31389 5 1 1 31388
0 31390 7 1 2 76752 31389
0 31391 5 1 1 31390
0 31392 7 1 2 31374 31391
0 31393 5 1 1 31392
0 31394 7 1 2 60968 31393
0 31395 5 1 1 31394
0 31396 7 3 2 82528 90074
0 31397 7 1 2 90953 92557
0 31398 5 1 1 31397
0 31399 7 1 2 31395 31398
0 31400 5 1 1 31399
0 31401 7 1 2 88534 31400
0 31402 5 1 1 31401
0 31403 7 1 2 83656 89164
0 31404 7 1 2 92552 31403
0 31405 5 1 1 31404
0 31406 7 2 2 63042 90302
0 31407 7 1 2 64711 90483
0 31408 7 1 2 92560 31407
0 31409 5 1 1 31408
0 31410 7 1 2 31405 31409
0 31411 5 1 1 31410
0 31412 7 1 2 63724 31411
0 31413 5 1 1 31412
0 31414 7 1 2 88392 91422
0 31415 7 1 2 77643 31414
0 31416 5 1 1 31415
0 31417 7 1 2 31413 31416
0 31418 5 1 1 31417
0 31419 7 1 2 61650 31418
0 31420 5 1 1 31419
0 31421 7 1 2 77102 91187
0 31422 7 1 2 91968 31421
0 31423 7 1 2 79784 31422
0 31424 5 1 1 31423
0 31425 7 1 2 31420 31424
0 31426 5 1 1 31425
0 31427 7 1 2 63320 31426
0 31428 5 1 1 31427
0 31429 7 1 2 58750 87646
0 31430 5 1 1 31429
0 31431 7 2 2 79026 90257
0 31432 5 1 1 92562
0 31433 7 1 2 31430 31432
0 31434 5 1 1 31433
0 31435 7 1 2 59601 31434
0 31436 5 1 1 31435
0 31437 7 2 2 63043 79454
0 31438 7 1 2 91821 92564
0 31439 5 1 1 31438
0 31440 7 1 2 31436 31439
0 31441 5 1 1 31440
0 31442 7 1 2 77103 31441
0 31443 5 1 1 31442
0 31444 7 4 2 58751 63779
0 31445 7 2 2 62218 92566
0 31446 7 1 2 73724 87549
0 31447 7 1 2 92570 31446
0 31448 5 1 1 31447
0 31449 7 1 2 31443 31448
0 31450 5 1 1 31449
0 31451 7 1 2 58568 91969
0 31452 7 1 2 31450 31451
0 31453 5 1 1 31452
0 31454 7 1 2 31428 31453
0 31455 5 1 1 31454
0 31456 7 1 2 61341 31455
0 31457 5 1 1 31456
0 31458 7 2 2 65959 66845
0 31459 7 1 2 90235 91970
0 31460 7 1 2 92572 31459
0 31461 7 1 2 92396 31460
0 31462 5 1 1 31461
0 31463 7 1 2 31457 31462
0 31464 5 1 1 31463
0 31465 7 1 2 60969 31464
0 31466 5 1 1 31465
0 31467 7 2 2 71431 88134
0 31468 7 1 2 92558 92574
0 31469 7 1 2 88048 31468
0 31470 5 1 1 31469
0 31471 7 1 2 31466 31470
0 31472 5 1 1 31471
0 31473 7 1 2 70522 31472
0 31474 5 1 1 31473
0 31475 7 1 2 31402 31474
0 31476 5 1 1 31475
0 31477 7 1 2 60598 31476
0 31478 5 1 1 31477
0 31479 7 1 2 31363 31478
0 31480 5 1 1 31479
0 31481 7 1 2 63902 31480
0 31482 5 1 1 31481
0 31483 7 1 2 86941 87710
0 31484 5 1 1 31483
0 31485 7 1 2 26401 31484
0 31486 5 1 1 31485
0 31487 7 1 2 88049 91238
0 31488 7 1 2 31486 31487
0 31489 5 1 1 31488
0 31490 7 1 2 90464 92264
0 31491 7 1 2 90608 31490
0 31492 5 1 1 31491
0 31493 7 1 2 31489 31492
0 31494 5 1 1 31493
0 31495 7 1 2 66269 31494
0 31496 5 1 1 31495
0 31497 7 4 2 58569 79264
0 31498 7 3 2 83636 92576
0 31499 7 2 2 79020 89881
0 31500 7 1 2 92580 92583
0 31501 5 1 1 31500
0 31502 7 1 2 31496 31501
0 31503 5 1 1 31502
0 31504 7 1 2 64902 31503
0 31505 5 1 1 31504
0 31506 7 2 2 90051 91624
0 31507 7 1 2 79478 90528
0 31508 7 1 2 92585 31507
0 31509 5 1 1 31508
0 31510 7 1 2 31505 31509
0 31511 5 1 1 31510
0 31512 7 1 2 63725 31511
0 31513 5 1 1 31512
0 31514 7 1 2 91115 92319
0 31515 7 1 2 74914 31514
0 31516 7 1 2 92586 31515
0 31517 5 1 1 31516
0 31518 7 1 2 31513 31517
0 31519 5 1 1 31518
0 31520 7 1 2 70523 31519
0 31521 5 1 1 31520
0 31522 7 3 2 64712 86564
0 31523 7 2 2 66480 77641
0 31524 7 1 2 78581 92590
0 31525 7 1 2 92587 31524
0 31526 5 1 1 31525
0 31527 7 1 2 86699 90490
0 31528 5 1 1 31527
0 31529 7 1 2 74339 88872
0 31530 7 1 2 31528 31529
0 31531 5 1 1 31530
0 31532 7 1 2 31526 31531
0 31533 5 1 1 31532
0 31534 7 1 2 65615 31533
0 31535 5 1 1 31534
0 31536 7 1 2 88873 90168
0 31537 5 1 1 31536
0 31538 7 3 2 60009 89882
0 31539 5 1 1 92592
0 31540 7 1 2 92565 92593
0 31541 5 1 1 31540
0 31542 7 1 2 66270 89858
0 31543 7 1 2 77512 31542
0 31544 5 1 1 31543
0 31545 7 1 2 31541 31544
0 31546 5 1 1 31545
0 31547 7 1 2 91014 31546
0 31548 5 1 1 31547
0 31549 7 1 2 31537 31548
0 31550 5 1 1 31549
0 31551 7 1 2 60390 31550
0 31552 5 1 1 31551
0 31553 7 1 2 31535 31552
0 31554 5 1 1 31553
0 31555 7 1 2 75546 31554
0 31556 5 1 1 31555
0 31557 7 1 2 91015 92101
0 31558 5 1 1 31557
0 31559 7 1 2 86041 87532
0 31560 5 1 1 31559
0 31561 7 1 2 31558 31560
0 31562 5 1 1 31561
0 31563 7 1 2 79495 31562
0 31564 5 1 1 31563
0 31565 7 1 2 65272 87333
0 31566 7 1 2 82135 31565
0 31567 5 1 1 31566
0 31568 7 1 2 31564 31567
0 31569 5 1 1 31568
0 31570 7 1 2 63044 31569
0 31571 5 1 1 31570
0 31572 7 1 2 77513 92540
0 31573 5 1 1 31572
0 31574 7 1 2 31571 31573
0 31575 5 1 1 31574
0 31576 7 1 2 89058 31575
0 31577 5 1 1 31576
0 31578 7 1 2 31556 31577
0 31579 5 1 1 31578
0 31580 7 1 2 88535 31579
0 31581 5 1 1 31580
0 31582 7 1 2 67562 87201
0 31583 5 1 1 31582
0 31584 7 1 2 86516 31583
0 31585 5 1 1 31584
0 31586 7 1 2 90183 31585
0 31587 7 1 2 91216 31586
0 31588 5 1 1 31587
0 31589 7 3 2 88536 88874
0 31590 7 2 2 61651 92595
0 31591 7 1 2 65960 92598
0 31592 5 1 1 31591
0 31593 7 1 2 31588 31592
0 31594 5 1 1 31593
0 31595 7 1 2 71432 31594
0 31596 5 1 1 31595
0 31597 7 1 2 73052 90813
0 31598 7 1 2 92599 31597
0 31599 5 1 1 31598
0 31600 7 1 2 31596 31599
0 31601 5 1 1 31600
0 31602 7 1 2 76753 31601
0 31603 5 1 1 31602
0 31604 7 1 2 31581 31603
0 31605 7 1 2 31521 31604
0 31606 5 1 1 31605
0 31607 7 1 2 68864 31606
0 31608 5 1 1 31607
0 31609 7 1 2 86594 75486
0 31610 5 1 1 31609
0 31611 7 1 2 24720 31610
0 31612 5 1 1 31611
0 31613 7 1 2 59847 31612
0 31614 5 1 1 31613
0 31615 7 2 2 59602 77360
0 31616 7 1 2 73736 92600
0 31617 5 1 1 31616
0 31618 7 1 2 31614 31617
0 31619 5 1 1 31618
0 31620 7 1 2 68520 31619
0 31621 5 1 1 31620
0 31622 7 1 2 73028 86354
0 31623 5 1 1 31622
0 31624 7 1 2 91365 31623
0 31625 5 1 1 31624
0 31626 7 1 2 31621 31625
0 31627 5 1 1 31626
0 31628 7 1 2 58570 31627
0 31629 5 1 1 31628
0 31630 7 1 2 72476 86727
0 31631 7 1 2 91986 31630
0 31632 5 1 1 31631
0 31633 7 1 2 31629 31632
0 31634 5 1 1 31633
0 31635 7 1 2 61848 31634
0 31636 5 1 1 31635
0 31637 7 1 2 74727 89092
0 31638 7 1 2 92524 31637
0 31639 5 1 1 31638
0 31640 7 1 2 31636 31639
0 31641 5 1 1 31640
0 31642 7 1 2 66271 31641
0 31643 5 1 1 31642
0 31644 7 2 2 66481 80966
0 31645 7 1 2 68622 70351
0 31646 5 1 1 31645
0 31647 7 1 2 92602 31646
0 31648 5 1 1 31647
0 31649 7 2 2 74340 89495
0 31650 7 1 2 78119 73835
0 31651 7 1 2 92604 31650
0 31652 5 1 1 31651
0 31653 7 1 2 31648 31652
0 31654 5 1 1 31653
0 31655 7 1 2 86487 31654
0 31656 5 1 1 31655
0 31657 7 1 2 31643 31656
0 31658 5 1 1 31657
0 31659 7 1 2 91217 31658
0 31660 5 1 1 31659
0 31661 7 1 2 86069 88341
0 31662 5 1 1 31661
0 31663 7 1 2 31662 28928
0 31664 5 1 1 31663
0 31665 7 2 2 77397 84457
0 31666 7 1 2 84265 79983
0 31667 7 1 2 91917 31666
0 31668 7 1 2 92606 31667
0 31669 7 1 2 31664 31668
0 31670 5 1 1 31669
0 31671 7 1 2 31660 31670
0 31672 7 1 2 31608 31671
0 31673 7 1 2 31482 31672
0 31674 7 1 2 31336 31673
0 31675 5 1 1 31674
0 31676 7 1 2 62108 31675
0 31677 5 1 1 31676
0 31678 7 1 2 66918 90823
0 31679 5 1 1 31678
0 31680 7 1 2 6549 31679
0 31681 5 1 1 31680
0 31682 7 1 2 81504 87877
0 31683 7 1 2 91026 31682
0 31684 7 1 2 31681 31683
0 31685 5 1 1 31684
0 31686 7 1 2 62109 89903
0 31687 7 1 2 78046 31686
0 31688 7 1 2 91334 31687
0 31689 5 1 1 31688
0 31690 7 1 2 31685 31689
0 31691 5 1 1 31690
0 31692 7 1 2 88952 31691
0 31693 5 1 1 31692
0 31694 7 1 2 75374 92591
0 31695 5 1 1 31694
0 31696 7 1 2 87278 88875
0 31697 5 1 1 31696
0 31698 7 1 2 31695 31697
0 31699 5 1 1 31698
0 31700 7 1 2 88094 31699
0 31701 5 1 1 31700
0 31702 7 1 2 58752 89859
0 31703 7 1 2 90912 31702
0 31704 7 1 2 92040 31703
0 31705 5 1 1 31704
0 31706 7 1 2 78450 91800
0 31707 5 1 1 31706
0 31708 7 1 2 68865 88876
0 31709 5 1 1 31708
0 31710 7 1 2 31707 31709
0 31711 5 1 1 31710
0 31712 7 1 2 71289 88760
0 31713 7 1 2 31711 31712
0 31714 5 1 1 31713
0 31715 7 1 2 31705 31714
0 31716 5 1 1 31715
0 31717 7 1 2 63726 31716
0 31718 5 1 1 31717
0 31719 7 1 2 31701 31718
0 31720 5 1 1 31719
0 31721 7 1 2 60970 31720
0 31722 5 1 1 31721
0 31723 7 1 2 76898 86792
0 31724 7 1 2 92596 31723
0 31725 5 1 1 31724
0 31726 7 1 2 31722 31725
0 31727 5 1 1 31726
0 31728 7 1 2 88013 31727
0 31729 5 1 1 31728
0 31730 7 1 2 70911 86797
0 31731 5 1 1 31730
0 31732 7 1 2 61849 81472
0 31733 7 1 2 31731 31732
0 31734 7 1 2 92548 31733
0 31735 5 1 1 31734
0 31736 7 1 2 31729 31735
0 31737 5 1 1 31736
0 31738 7 1 2 62110 31737
0 31739 5 1 1 31738
0 31740 7 1 2 31693 31739
0 31741 5 1 1 31740
0 31742 7 1 2 65961 31741
0 31743 5 1 1 31742
0 31744 7 4 2 64569 87149
0 31745 7 1 2 83665 92608
0 31746 5 1 1 31745
0 31747 7 1 2 64713 76524
0 31748 7 1 2 92033 31747
0 31749 5 1 1 31748
0 31750 7 1 2 31746 31749
0 31751 5 2 1 31750
0 31752 7 1 2 88761 92612
0 31753 5 1 1 31752
0 31754 7 3 2 70524 88576
0 31755 7 1 2 92516 92614
0 31756 5 1 1 31755
0 31757 7 1 2 31753 31756
0 31758 5 1 1 31757
0 31759 7 1 2 61850 31758
0 31760 5 1 1 31759
0 31761 7 2 2 62219 66482
0 31762 7 1 2 60010 92617
0 31763 7 1 2 92034 31762
0 31764 7 1 2 92615 31763
0 31765 5 1 1 31764
0 31766 7 1 2 31760 31765
0 31767 5 1 1 31766
0 31768 7 1 2 63727 31767
0 31769 5 1 1 31768
0 31770 7 1 2 92532 92613
0 31771 5 1 1 31770
0 31772 7 1 2 31769 31771
0 31773 5 1 1 31772
0 31774 7 1 2 81874 31773
0 31775 5 1 1 31774
0 31776 7 1 2 62220 82382
0 31777 7 1 2 88877 31776
0 31778 5 1 1 31777
0 31779 7 1 2 81401 88665
0 31780 7 1 2 92561 31779
0 31781 5 1 1 31780
0 31782 7 1 2 31778 31781
0 31783 5 1 1 31782
0 31784 7 1 2 88537 31783
0 31785 5 1 1 31784
0 31786 7 2 2 89904 92616
0 31787 7 2 2 63728 64347
0 31788 7 3 2 63045 92621
0 31789 7 1 2 66846 92623
0 31790 7 1 2 92619 31789
0 31791 5 1 1 31790
0 31792 7 1 2 31785 31791
0 31793 5 1 1 31792
0 31794 7 1 2 69036 31793
0 31795 5 1 1 31794
0 31796 7 1 2 90435 92597
0 31797 5 1 1 31796
0 31798 7 1 2 62221 81557
0 31799 5 1 1 31798
0 31800 7 1 2 82393 31799
0 31801 5 1 1 31800
0 31802 7 1 2 66483 74466
0 31803 5 1 1 31802
0 31804 7 2 2 30571 31803
0 31805 5 1 1 92626
0 31806 7 1 2 63502 92627
0 31807 5 1 1 31806
0 31808 7 4 2 71685 92509
0 31809 5 1 1 92628
0 31810 7 1 2 58753 31809
0 31811 5 1 1 31810
0 31812 7 1 2 88538 31811
0 31813 7 1 2 31807 31812
0 31814 5 1 1 31813
0 31815 7 1 2 88577 92514
0 31816 7 1 2 79953 31815
0 31817 5 1 1 31816
0 31818 7 1 2 31814 31817
0 31819 5 1 1 31818
0 31820 7 1 2 31801 31819
0 31821 5 1 1 31820
0 31822 7 1 2 31797 31821
0 31823 7 1 2 31795 31822
0 31824 5 1 1 31823
0 31825 7 1 2 76754 31824
0 31826 5 1 1 31825
0 31827 7 1 2 59603 92620
0 31828 5 1 1 31827
0 31829 7 3 2 77398 87186
0 31830 7 1 2 88765 92632
0 31831 5 1 1 31830
0 31832 7 1 2 31828 31831
0 31833 5 1 1 31832
0 31834 7 1 2 63729 31833
0 31835 5 1 1 31834
0 31836 7 1 2 92633 92533
0 31837 5 1 1 31836
0 31838 7 1 2 31835 31837
0 31839 5 1 1 31838
0 31840 7 1 2 88050 31839
0 31841 5 1 1 31840
0 31842 7 1 2 89405 92634
0 31843 5 1 1 31842
0 31844 7 1 2 71960 82288
0 31845 7 1 2 89905 31844
0 31846 5 1 1 31845
0 31847 7 1 2 31843 31846
0 31848 5 1 1 31847
0 31849 7 1 2 88342 31848
0 31850 5 1 1 31849
0 31851 7 1 2 81025 89149
0 31852 7 1 2 91380 31851
0 31853 5 1 1 31852
0 31854 7 1 2 31850 31853
0 31855 5 1 1 31854
0 31856 7 1 2 91653 31855
0 31857 5 1 1 31856
0 31858 7 1 2 31841 31857
0 31859 5 1 1 31858
0 31860 7 1 2 69037 31859
0 31861 5 1 1 31860
0 31862 7 1 2 91727 92035
0 31863 5 1 1 31862
0 31864 7 2 2 82208 89409
0 31865 5 1 1 92635
0 31866 7 1 2 74666 92636
0 31867 5 1 1 31866
0 31868 7 1 2 31863 31867
0 31869 5 1 1 31868
0 31870 7 1 2 88539 31869
0 31871 5 1 1 31870
0 31872 7 1 2 84742 91825
0 31873 7 1 2 90967 31872
0 31874 7 1 2 91528 31873
0 31875 5 1 1 31874
0 31876 7 1 2 31871 31875
0 31877 5 1 1 31876
0 31878 7 1 2 31805 31877
0 31879 5 1 1 31878
0 31880 7 1 2 60134 92629
0 31881 5 1 1 31880
0 31882 7 1 2 76029 90448
0 31883 5 1 1 31882
0 31884 7 1 2 31881 31883
0 31885 5 1 1 31884
0 31886 7 1 2 87923 88343
0 31887 5 1 1 31886
0 31888 7 1 2 83554 92217
0 31889 5 1 1 31888
0 31890 7 1 2 31887 31889
0 31891 5 1 1 31890
0 31892 7 1 2 31885 31891
0 31893 5 1 1 31892
0 31894 7 1 2 87858 92630
0 31895 5 1 1 31894
0 31896 7 1 2 66484 76607
0 31897 7 1 2 88578 31896
0 31898 5 1 1 31897
0 31899 7 1 2 31895 31898
0 31900 5 1 1 31899
0 31901 7 1 2 63730 31900
0 31902 5 1 1 31901
0 31903 7 1 2 88205 92631
0 31904 5 1 1 31903
0 31905 7 1 2 31902 31904
0 31906 5 1 1 31905
0 31907 7 2 2 77810 79562
0 31908 5 1 1 92637
0 31909 7 1 2 79239 3356
0 31910 7 1 2 92638 31909
0 31911 7 1 2 31906 31910
0 31912 5 1 1 31911
0 31913 7 1 2 31893 31912
0 31914 5 1 1 31913
0 31915 7 1 2 91728 31914
0 31916 5 1 1 31915
0 31917 7 1 2 31879 31916
0 31918 7 1 2 31861 31917
0 31919 7 1 2 31826 31918
0 31920 7 1 2 31775 31919
0 31921 5 1 1 31920
0 31922 7 1 2 60599 31921
0 31923 5 1 1 31922
0 31924 7 1 2 80975 91218
0 31925 5 1 1 31924
0 31926 7 1 2 88135 89972
0 31927 7 1 2 89371 31926
0 31928 5 1 1 31927
0 31929 7 1 2 31925 31928
0 31930 5 1 1 31929
0 31931 7 1 2 86258 89906
0 31932 7 1 2 31930 31931
0 31933 5 1 1 31932
0 31934 7 1 2 31923 31933
0 31935 5 1 1 31934
0 31936 7 1 2 80031 31935
0 31937 5 1 1 31936
0 31938 7 1 2 31743 31937
0 31939 5 1 1 31938
0 31940 7 1 2 68241 31939
0 31941 5 1 1 31940
0 31942 7 1 2 66599 31941
0 31943 7 1 2 31677 31942
0 31944 5 1 1 31943
0 31945 7 1 2 68094 31944
0 31946 7 1 2 31214 31945
0 31947 5 1 1 31946
0 31948 7 1 2 60600 20221
0 31949 5 1 1 31948
0 31950 7 2 2 10746 31949
0 31951 7 1 2 83226 92639
0 31952 5 1 1 31951
0 31953 7 1 2 63046 31952
0 31954 5 1 1 31953
0 31955 7 1 2 9754 31954
0 31956 5 1 1 31955
0 31957 7 1 2 81338 31956
0 31958 5 1 1 31957
0 31959 7 1 2 58306 83908
0 31960 5 1 1 31959
0 31961 7 1 2 83347 31960
0 31962 5 1 1 31961
0 31963 7 1 2 82383 31962
0 31964 5 1 1 31963
0 31965 7 1 2 31958 31964
0 31966 5 1 1 31965
0 31967 7 1 2 64570 31966
0 31968 5 1 1 31967
0 31969 7 1 2 77697 80357
0 31970 5 1 1 31969
0 31971 7 1 2 63047 83909
0 31972 5 1 1 31971
0 31973 7 1 2 91854 31972
0 31974 7 1 2 31970 31973
0 31975 5 2 1 31974
0 31976 7 1 2 89524 92641
0 31977 5 1 1 31976
0 31978 7 1 2 31968 31977
0 31979 5 1 1 31978
0 31980 7 1 2 63321 31979
0 31981 5 1 1 31980
0 31982 7 1 2 61652 87823
0 31983 7 1 2 92642 31982
0 31984 5 1 1 31983
0 31985 7 1 2 31981 31984
0 31986 5 1 1 31985
0 31987 7 1 2 72746 31986
0 31988 5 1 1 31987
0 31989 7 2 2 66973 74591
0 31990 7 1 2 73349 92643
0 31991 5 1 1 31990
0 31992 7 2 2 62750 67055
0 31993 5 1 1 92645
0 31994 7 2 2 60391 92646
0 31995 5 1 1 92647
0 31996 7 1 2 71784 92648
0 31997 5 1 1 31996
0 31998 7 1 2 31991 31997
0 31999 5 1 1 31998
0 32000 7 1 2 80851 31999
0 32001 5 1 1 32000
0 32002 7 1 2 74001 79640
0 32003 7 1 2 92644 32002
0 32004 5 1 1 32003
0 32005 7 1 2 32001 32004
0 32006 5 1 1 32005
0 32007 7 1 2 61653 32006
0 32008 5 1 1 32007
0 32009 7 1 2 88964 91940
0 32010 5 1 1 32009
0 32011 7 2 2 60135 69165
0 32012 5 2 1 92649
0 32013 7 1 2 64348 92650
0 32014 5 1 1 32013
0 32015 7 1 2 32010 32014
0 32016 5 1 1 32015
0 32017 7 1 2 63048 32016
0 32018 5 1 1 32017
0 32019 7 1 2 58307 88965
0 32020 5 1 1 32019
0 32021 7 1 2 92651 32020
0 32022 5 1 1 32021
0 32023 7 1 2 77629 32022
0 32024 5 1 1 32023
0 32025 7 1 2 32018 32024
0 32026 5 1 1 32025
0 32027 7 1 2 88560 32026
0 32028 5 1 1 32027
0 32029 7 1 2 32008 32028
0 32030 5 1 1 32029
0 32031 7 1 2 63635 32030
0 32032 5 1 1 32031
0 32033 7 1 2 68242 87447
0 32034 5 1 1 32033
0 32035 7 1 2 83724 88014
0 32036 5 1 1 32035
0 32037 7 1 2 32034 32036
0 32038 5 1 1 32037
0 32039 7 1 2 62751 32038
0 32040 5 1 1 32039
0 32041 7 1 2 26871 32040
0 32042 5 1 1 32041
0 32043 7 1 2 74097 91526
0 32044 7 1 2 32042 32043
0 32045 5 1 1 32044
0 32046 7 1 2 32032 32045
0 32047 5 1 1 32046
0 32048 7 1 2 68866 32047
0 32049 5 1 1 32048
0 32050 7 1 2 62752 15315
0 32051 5 1 1 32050
0 32052 7 1 2 79684 32051
0 32053 5 1 1 32052
0 32054 7 1 2 57711 88439
0 32055 5 1 1 32054
0 32056 7 1 2 32053 32055
0 32057 5 1 1 32056
0 32058 7 1 2 61654 90824
0 32059 7 1 2 32057 32058
0 32060 5 1 1 32059
0 32061 7 1 2 88443 87980
0 32062 7 1 2 88441 32061
0 32063 5 1 1 32062
0 32064 7 1 2 75547 81558
0 32065 7 1 2 32063 32064
0 32066 5 1 1 32065
0 32067 7 1 2 32060 32066
0 32068 5 1 1 32067
0 32069 7 1 2 84224 32068
0 32070 5 1 1 32069
0 32071 7 1 2 32049 32070
0 32072 7 1 2 31988 32071
0 32073 5 1 1 32072
0 32074 7 1 2 66709 32073
0 32075 5 1 1 32074
0 32076 7 4 2 66272 67754
0 32077 7 1 2 75548 92653
0 32078 5 1 1 32077
0 32079 7 1 2 26809 32078
0 32080 5 1 1 32079
0 32081 7 1 2 68867 91974
0 32082 7 2 2 32080 32081
0 32083 7 1 2 69487 92657
0 32084 5 1 1 32083
0 32085 7 1 2 58308 19688
0 32086 5 1 1 32085
0 32087 7 1 2 88015 32086
0 32088 5 1 1 32087
0 32089 7 1 2 70649 84345
0 32090 7 1 2 80374 32089
0 32091 5 1 1 32090
0 32092 7 2 2 58309 83033
0 32093 7 1 2 83234 92659
0 32094 7 1 2 32091 32093
0 32095 5 1 1 32094
0 32096 7 1 2 87448 32095
0 32097 5 1 1 32096
0 32098 7 1 2 32088 32097
0 32099 5 1 1 32098
0 32100 7 1 2 64349 32099
0 32101 5 1 1 32100
0 32102 7 1 2 63049 6781
0 32103 5 1 1 32102
0 32104 7 1 2 78163 87261
0 32105 7 1 2 32103 32104
0 32106 5 1 1 32105
0 32107 7 1 2 32101 32106
0 32108 5 1 1 32107
0 32109 7 2 2 67480 32108
0 32110 5 1 1 92661
0 32111 7 1 2 67930 92662
0 32112 5 1 1 32111
0 32113 7 1 2 32084 32112
0 32114 7 1 2 32075 32113
0 32115 5 1 1 32114
0 32116 7 1 2 64903 32115
0 32117 5 1 1 32116
0 32118 7 1 2 64350 92658
0 32119 5 1 1 32118
0 32120 7 1 2 32110 32119
0 32121 5 2 1 32120
0 32122 7 1 2 87863 92663
0 32123 5 1 1 32122
0 32124 7 1 2 32117 32123
0 32125 5 1 1 32124
0 32126 7 1 2 63731 32125
0 32127 5 1 1 32126
0 32128 7 1 2 88095 92664
0 32129 5 1 1 32128
0 32130 7 1 2 32127 32129
0 32131 5 1 1 32130
0 32132 7 1 2 61851 32131
0 32133 5 1 1 32132
0 32134 7 1 2 58048 72693
0 32135 5 1 1 32134
0 32136 7 1 2 10361 32135
0 32137 5 1 1 32136
0 32138 7 1 2 64904 32137
0 32139 5 1 1 32138
0 32140 7 1 2 87864 91357
0 32141 5 1 1 32140
0 32142 7 1 2 32139 32141
0 32143 5 1 1 32142
0 32144 7 1 2 63732 32143
0 32145 5 1 1 32144
0 32146 7 1 2 69555 88864
0 32147 7 1 2 89306 32146
0 32148 5 1 1 32147
0 32149 7 1 2 32145 32148
0 32150 5 1 1 32149
0 32151 7 1 2 68623 32150
0 32152 5 1 1 32151
0 32153 7 1 2 88865 91298
0 32154 7 1 2 72694 32153
0 32155 5 1 1 32154
0 32156 7 1 2 32152 32155
0 32157 5 1 1 32156
0 32158 7 1 2 65273 32157
0 32159 5 1 1 32158
0 32160 7 2 2 70872 79794
0 32161 5 1 1 92665
0 32162 7 1 2 63050 32161
0 32163 5 1 1 32162
0 32164 7 1 2 72747 32163
0 32165 5 1 1 32164
0 32166 7 2 2 68779 71061
0 32167 7 1 2 88966 92667
0 32168 5 1 1 32167
0 32169 7 1 2 32165 32168
0 32170 5 1 1 32169
0 32171 7 1 2 88149 32170
0 32172 5 1 1 32171
0 32173 7 1 2 32159 32172
0 32174 5 1 1 32173
0 32175 7 1 2 73725 32174
0 32176 5 1 1 32175
0 32177 7 2 2 82157 66974
0 32178 7 1 2 60601 92669
0 32179 5 1 1 32178
0 32180 7 1 2 67084 32179
0 32181 5 1 1 32180
0 32182 7 1 2 63636 32181
0 32183 5 1 1 32182
0 32184 7 1 2 84772 32183
0 32185 5 1 1 32184
0 32186 7 2 2 88368 32185
0 32187 7 1 2 63733 79662
0 32188 7 1 2 92671 32187
0 32189 5 1 1 32188
0 32190 7 1 2 32176 32189
0 32191 5 1 1 32190
0 32192 7 1 2 63322 32191
0 32193 5 1 1 32192
0 32194 7 1 2 77823 92624
0 32195 7 1 2 92672 32194
0 32196 5 1 1 32195
0 32197 7 1 2 32193 32196
0 32198 5 1 1 32197
0 32199 7 1 2 61852 32198
0 32200 5 1 1 32199
0 32201 7 1 2 73405 70554
0 32202 5 1 1 32201
0 32203 7 1 2 74517 71088
0 32204 5 1 1 32203
0 32205 7 1 2 32202 32204
0 32206 5 1 1 32205
0 32207 7 1 2 91744 91971
0 32208 7 1 2 32206 32207
0 32209 5 1 1 32208
0 32210 7 1 2 32200 32209
0 32211 5 1 1 32210
0 32212 7 1 2 61655 32211
0 32213 5 1 1 32212
0 32214 7 3 2 66273 80814
0 32215 7 1 2 88830 91116
0 32216 7 1 2 92622 32215
0 32217 7 1 2 92673 32216
0 32218 7 1 2 72695 32217
0 32219 5 1 1 32218
0 32220 7 1 2 32213 32219
0 32221 5 1 1 32220
0 32222 7 1 2 68378 32221
0 32223 5 1 1 32222
0 32224 7 1 2 65274 82238
0 32225 5 1 1 32224
0 32226 7 1 2 75131 32225
0 32227 5 1 1 32226
0 32228 7 1 2 73413 83805
0 32229 5 1 1 32228
0 32230 7 1 2 59132 32229
0 32231 5 1 1 32230
0 32232 7 1 2 92284 32231
0 32233 7 1 2 32227 32232
0 32234 5 1 1 32233
0 32235 7 1 2 70085 80109
0 32236 5 1 1 32235
0 32237 7 1 2 71601 32236
0 32238 5 1 1 32237
0 32239 7 1 2 78529 89385
0 32240 7 1 2 32238 32239
0 32241 5 1 1 32240
0 32242 7 1 2 32234 32241
0 32243 5 1 1 32242
0 32244 7 1 2 71076 32243
0 32245 5 1 1 32244
0 32246 7 2 2 78601 84166
0 32247 7 1 2 60136 89973
0 32248 7 1 2 92676 32247
0 32249 5 1 1 32248
0 32250 7 1 2 32245 32249
0 32251 5 1 1 32250
0 32252 7 1 2 63637 32251
0 32253 5 1 1 32252
0 32254 7 1 2 70457 89974
0 32255 7 1 2 92677 32254
0 32256 5 1 1 32255
0 32257 7 1 2 32253 32256
0 32258 5 1 1 32257
0 32259 7 1 2 91972 32258
0 32260 5 1 1 32259
0 32261 7 1 2 32223 32260
0 32262 7 1 2 32133 32261
0 32263 5 1 1 32262
0 32264 7 1 2 66919 32263
0 32265 5 1 1 32264
0 32266 7 2 2 66485 84078
0 32267 7 1 2 88016 92678
0 32268 5 1 1 32267
0 32269 7 1 2 74376 91256
0 32270 5 1 1 32269
0 32271 7 1 2 32268 32270
0 32272 5 1 1 32271
0 32273 7 1 2 77673 32272
0 32274 5 1 1 32273
0 32275 7 1 2 67755 84327
0 32276 5 1 1 32275
0 32277 7 1 2 69396 70650
0 32278 5 1 1 32277
0 32279 7 1 2 58310 32278
0 32280 7 1 2 32276 32279
0 32281 5 1 1 32280
0 32282 7 1 2 91257 32281
0 32283 5 1 1 32282
0 32284 7 1 2 58049 81959
0 32285 5 1 1 32284
0 32286 7 1 2 88017 92259
0 32287 7 1 2 32285 32286
0 32288 5 1 1 32287
0 32289 7 1 2 32283 32288
0 32290 7 1 2 32274 32289
0 32291 5 1 1 32290
0 32292 7 1 2 64351 32291
0 32293 5 1 1 32292
0 32294 7 1 2 84062 89059
0 32295 5 1 1 32294
0 32296 7 1 2 32293 32295
0 32297 5 1 1 32296
0 32298 7 1 2 91301 32297
0 32299 5 1 1 32298
0 32300 7 1 2 63780 89736
0 32301 5 1 1 32300
0 32302 7 1 2 89745 32301
0 32303 5 2 1 32302
0 32304 7 1 2 58571 92680
0 32305 5 1 1 32304
0 32306 7 1 2 86832 89730
0 32307 5 1 1 32306
0 32308 7 1 2 32305 32307
0 32309 5 1 1 32308
0 32310 7 1 2 62222 32309
0 32311 5 1 1 32310
0 32312 7 1 2 84520 90895
0 32313 5 1 1 32312
0 32314 7 1 2 32311 32313
0 32315 5 1 1 32314
0 32316 7 1 2 84559 87944
0 32317 7 1 2 32315 32316
0 32318 5 1 1 32317
0 32319 7 1 2 89854 92681
0 32320 5 1 1 32319
0 32321 7 1 2 78083 89652
0 32322 7 1 2 92329 32321
0 32323 5 1 1 32322
0 32324 7 1 2 21821 32323
0 32325 7 1 2 32320 32324
0 32326 5 1 1 32325
0 32327 7 1 2 65275 87960
0 32328 7 1 2 32326 32327
0 32329 5 1 1 32328
0 32330 7 1 2 32318 32329
0 32331 5 1 1 32330
0 32332 7 1 2 60392 32331
0 32333 5 1 1 32332
0 32334 7 2 2 76649 69874
0 32335 7 1 2 89888 92682
0 32336 5 2 1 32335
0 32337 7 2 2 88797 91343
0 32338 7 1 2 87786 87961
0 32339 7 1 2 92686 32338
0 32340 5 1 1 32339
0 32341 7 1 2 92684 32340
0 32342 5 1 1 32341
0 32343 7 1 2 58982 32342
0 32344 5 1 1 32343
0 32345 7 2 2 77361 81339
0 32346 5 1 1 92688
0 32347 7 1 2 63903 88798
0 32348 7 2 2 92689 32347
0 32349 7 1 2 91573 92690
0 32350 5 1 1 32349
0 32351 7 1 2 70817 82564
0 32352 7 1 2 89876 32351
0 32353 5 1 1 32352
0 32354 7 1 2 32350 32353
0 32355 5 1 1 32354
0 32356 7 1 2 58050 32355
0 32357 5 1 1 32356
0 32358 7 1 2 74594 92330
0 32359 7 1 2 92687 32358
0 32360 5 1 1 32359
0 32361 7 1 2 92685 32360
0 32362 5 1 1 32361
0 32363 7 1 2 57428 32362
0 32364 5 1 1 32363
0 32365 7 1 2 32357 32364
0 32366 7 1 2 32344 32365
0 32367 7 1 2 32333 32366
0 32368 5 1 1 32367
0 32369 7 1 2 62474 32368
0 32370 5 1 1 32369
0 32371 7 1 2 58051 91584
0 32372 5 1 1 32371
0 32373 7 1 2 89234 92013
0 32374 5 3 1 32373
0 32375 7 1 2 32372 92692
0 32376 5 1 1 32375
0 32377 7 1 2 71183 32376
0 32378 5 1 1 32377
0 32379 7 1 2 88572 92603
0 32380 5 1 1 32379
0 32381 7 1 2 32378 32380
0 32382 5 1 1 32381
0 32383 7 1 2 68868 32382
0 32384 5 1 1 32383
0 32385 7 1 2 66486 88505
0 32386 7 1 2 92301 32385
0 32387 7 1 2 90825 32386
0 32388 5 1 1 32387
0 32389 7 1 2 32384 32388
0 32390 5 1 1 32389
0 32391 7 1 2 61656 32390
0 32392 5 1 1 32391
0 32393 7 1 2 61853 92285
0 32394 7 1 2 88574 32393
0 32395 5 1 1 32394
0 32396 7 1 2 32392 32395
0 32397 5 1 1 32396
0 32398 7 1 2 74592 32397
0 32399 5 1 1 32398
0 32400 7 1 2 76459 90191
0 32401 5 1 1 32400
0 32402 7 1 2 77549 91161
0 32403 5 1 1 32402
0 32404 7 1 2 32401 32403
0 32405 5 1 1 32404
0 32406 7 1 2 76755 32405
0 32407 5 1 1 32406
0 32408 7 1 2 89848 90896
0 32409 5 1 1 32408
0 32410 7 1 2 77785 81695
0 32411 7 1 2 91271 32410
0 32412 5 1 1 32411
0 32413 7 1 2 32409 32412
0 32414 5 1 1 32413
0 32415 7 1 2 57429 32414
0 32416 5 1 1 32415
0 32417 7 1 2 10522 84072
0 32418 5 1 1 32417
0 32419 7 1 2 89060 32418
0 32420 5 1 1 32419
0 32421 7 1 2 32416 32420
0 32422 7 1 2 32407 32421
0 32423 5 1 1 32422
0 32424 7 1 2 71895 32423
0 32425 5 1 1 32424
0 32426 7 1 2 63051 87521
0 32427 7 1 2 92691 32426
0 32428 5 1 1 32427
0 32429 7 1 2 32425 32428
0 32430 5 1 1 32429
0 32431 7 1 2 87984 32430
0 32432 5 1 1 32431
0 32433 7 1 2 32399 32432
0 32434 7 1 2 32370 32433
0 32435 5 1 1 32434
0 32436 7 1 2 66785 88136
0 32437 7 1 2 69273 32436
0 32438 7 1 2 32435 32437
0 32439 5 1 1 32438
0 32440 7 1 2 32299 32439
0 32441 5 1 1 32440
0 32442 7 1 2 66600 32441
0 32443 5 1 1 32442
0 32444 7 2 2 80815 90632
0 32445 7 1 2 91911 92695
0 32446 5 1 1 32445
0 32447 7 2 2 69820 89204
0 32448 7 1 2 58572 74222
0 32449 7 1 2 89883 32448
0 32450 7 1 2 92697 32449
0 32451 5 1 1 32450
0 32452 7 1 2 32446 32451
0 32453 5 1 1 32452
0 32454 7 2 2 88407 88150
0 32455 7 1 2 32453 92699
0 32456 5 1 1 32455
0 32457 7 1 2 59604 91213
0 32458 5 1 1 32457
0 32459 7 1 2 82998 88096
0 32460 5 1 1 32459
0 32461 7 1 2 32458 32460
0 32462 5 1 1 32461
0 32463 7 1 2 61854 91889
0 32464 5 1 1 32463
0 32465 7 2 2 89653 92304
0 32466 5 1 1 92701
0 32467 7 1 2 83684 92702
0 32468 5 1 1 32467
0 32469 7 1 2 32464 32468
0 32470 5 1 1 32469
0 32471 7 1 2 83147 32470
0 32472 7 1 2 32462 32471
0 32473 5 1 1 32472
0 32474 7 1 2 32456 32473
0 32475 5 1 1 32474
0 32476 7 1 2 67862 32475
0 32477 5 1 1 32476
0 32478 7 1 2 83512 88806
0 32479 5 1 1 32478
0 32480 7 1 2 58311 32479
0 32481 5 1 1 32480
0 32482 7 1 2 86378 32481
0 32483 5 1 1 32482
0 32484 7 1 2 91134 32483
0 32485 5 1 1 32484
0 32486 7 1 2 60602 89924
0 32487 7 1 2 87100 32486
0 32488 5 1 1 32487
0 32489 7 1 2 32485 32488
0 32490 5 1 1 32489
0 32491 7 1 2 76756 32490
0 32492 5 1 1 32491
0 32493 7 2 2 57430 80110
0 32494 5 1 1 92703
0 32495 7 1 2 91930 92704
0 32496 5 1 1 32495
0 32497 7 1 2 74455 81559
0 32498 5 1 1 32497
0 32499 7 1 2 32496 32498
0 32500 5 1 1 32499
0 32501 7 1 2 68998 32500
0 32502 5 1 1 32501
0 32503 7 1 2 78530 81431
0 32504 5 1 1 32503
0 32505 7 1 2 90439 32504
0 32506 5 1 1 32505
0 32507 7 1 2 58052 32506
0 32508 5 1 1 32507
0 32509 7 1 2 70709 73209
0 32510 7 1 2 84129 32509
0 32511 5 1 1 32510
0 32512 7 1 2 32508 32511
0 32513 7 1 2 32502 32512
0 32514 5 1 1 32513
0 32515 7 1 2 89093 32514
0 32516 5 1 1 32515
0 32517 7 1 2 88807 92640
0 32518 5 1 1 32517
0 32519 7 1 2 63052 32518
0 32520 5 1 1 32519
0 32521 7 4 2 68243 70093
0 32522 5 1 1 92705
0 32523 7 1 2 75360 92706
0 32524 5 1 1 32523
0 32525 7 1 2 32520 32524
0 32526 5 1 1 32525
0 32527 7 1 2 81340 32526
0 32528 5 1 1 32527
0 32529 7 1 2 83927 81284
0 32530 7 1 2 32494 32529
0 32531 5 1 1 32530
0 32532 7 1 2 82384 32531
0 32533 5 1 1 32532
0 32534 7 1 2 32528 32533
0 32535 5 1 1 32534
0 32536 7 1 2 89061 32535
0 32537 5 1 1 32536
0 32538 7 1 2 32516 32537
0 32539 7 1 2 32492 32538
0 32540 5 1 1 32539
0 32541 7 1 2 92700 32540
0 32542 5 1 1 32541
0 32543 7 1 2 32477 32542
0 32544 7 1 2 32443 32543
0 32545 7 1 2 75172 90897
0 32546 5 1 1 32545
0 32547 7 1 2 58053 89737
0 32548 5 1 1 32547
0 32549 7 1 2 32546 32548
0 32550 5 1 1 32549
0 32551 7 1 2 63323 32550
0 32552 5 1 1 32551
0 32553 7 1 2 82594 87438
0 32554 5 3 1 32553
0 32555 7 2 2 58573 92709
0 32556 5 1 1 92712
0 32557 7 3 2 65053 61855
0 32558 7 2 2 57431 82565
0 32559 5 4 1 92717
0 32560 7 1 2 63781 92719
0 32561 5 1 1 32560
0 32562 7 1 2 92714 32561
0 32563 7 1 2 92713 32562
0 32564 5 1 1 32563
0 32565 7 1 2 32552 32564
0 32566 5 1 1 32565
0 32567 7 1 2 91303 32566
0 32568 5 1 1 32567
0 32569 7 1 2 89205 90361
0 32570 5 1 1 32569
0 32571 7 2 2 58574 87338
0 32572 5 3 1 92723
0 32573 7 1 2 77363 25651
0 32574 7 1 2 92724 32573
0 32575 5 1 1 32574
0 32576 7 1 2 32570 32575
0 32577 5 1 1 32576
0 32578 7 1 2 72821 88151
0 32579 7 1 2 32577 32578
0 32580 7 1 2 92098 32579
0 32581 5 1 1 32580
0 32582 7 1 2 32568 32581
0 32583 5 1 1 32582
0 32584 7 1 2 65276 32583
0 32585 5 1 1 32584
0 32586 7 1 2 76757 81473
0 32587 5 1 1 32586
0 32588 7 1 2 89364 32587
0 32589 5 1 1 32588
0 32590 7 1 2 61856 32589
0 32591 5 1 1 32590
0 32592 7 2 2 77362 89654
0 32593 5 1 1 92728
0 32594 7 1 2 89930 92729
0 32595 5 1 1 32594
0 32596 7 1 2 32591 32595
0 32597 5 1 1 32596
0 32598 7 1 2 58312 32597
0 32599 5 1 1 32598
0 32600 7 1 2 70722 86847
0 32601 7 6 2 58983 61657
0 32602 7 1 2 89235 92730
0 32603 7 1 2 32600 32602
0 32604 5 1 1 32603
0 32605 7 1 2 32599 32604
0 32606 5 1 1 32605
0 32607 7 1 2 88408 32606
0 32608 5 1 1 32607
0 32609 7 1 2 74908 84313
0 32610 7 1 2 82992 32609
0 32611 7 1 2 89209 88079
0 32612 7 1 2 32610 32611
0 32613 5 1 1 32612
0 32614 7 1 2 32608 32613
0 32615 5 1 1 32614
0 32616 7 1 2 88152 32615
0 32617 5 1 1 32616
0 32618 7 1 2 32585 32617
0 32619 5 1 1 32618
0 32620 7 1 2 59605 32619
0 32621 5 1 1 32620
0 32622 7 1 2 89746 32593
0 32623 5 1 1 32622
0 32624 7 1 2 58575 32623
0 32625 5 1 1 32624
0 32626 7 1 2 85251 89655
0 32627 5 1 1 32626
0 32628 7 1 2 32625 32627
0 32629 5 1 1 32628
0 32630 7 2 2 66710 68709
0 32631 7 1 2 92575 92736
0 32632 7 1 2 86070 32631
0 32633 7 1 2 32629 32632
0 32634 5 1 1 32633
0 32635 7 1 2 32621 32634
0 32636 5 1 1 32635
0 32637 7 1 2 68379 32636
0 32638 5 1 1 32637
0 32639 7 1 2 80350 89094
0 32640 7 1 2 91304 32639
0 32641 5 1 1 32640
0 32642 7 1 2 76650 77652
0 32643 7 1 2 88153 32642
0 32644 7 1 2 92099 32643
0 32645 5 1 1 32644
0 32646 7 1 2 32641 32645
0 32647 5 1 1 32646
0 32648 7 1 2 65277 32647
0 32649 5 1 1 32648
0 32650 7 1 2 67665 86313
0 32651 7 1 2 90416 32650
0 32652 7 1 2 92428 32651
0 32653 5 1 1 32652
0 32654 7 1 2 32649 32653
0 32655 5 1 1 32654
0 32656 7 1 2 82385 32655
0 32657 5 1 1 32656
0 32658 7 1 2 64905 73979
0 32659 7 1 2 87236 80661
0 32660 7 1 2 32658 32659
0 32661 7 1 2 92625 32660
0 32662 7 1 2 91292 32661
0 32663 5 1 1 32662
0 32664 7 1 2 32657 32663
0 32665 5 1 1 32664
0 32666 7 1 2 71741 32665
0 32667 5 1 1 32666
0 32668 7 1 2 32638 32667
0 32669 7 1 2 32544 32668
0 32670 7 1 2 32265 32669
0 32671 5 1 1 32670
0 32672 7 1 2 85506 5514
0 32673 7 1 2 32671 32672
0 32674 5 1 1 32673
0 32675 7 1 2 31947 32674
0 32676 7 1 2 29963 32675
0 32677 7 1 2 27758 32676
0 32678 7 1 2 23930 32677
0 32679 7 1 2 21113 32678
0 32680 7 1 2 18676 32679
0 32681 7 1 2 18548 32680
0 32682 5 1 1 32681
0 32683 7 1 2 51 32682
0 32684 5 1 1 32683
0 32685 7 1 2 78834 78859
0 32686 5 1 1 32685
0 32687 7 2 2 79674 32686
0 32688 5 2 1 92738
0 32689 7 1 2 85569 92740
0 32690 5 1 1 32689
0 32691 7 1 2 67015 84109
0 32692 5 2 1 32691
0 32693 7 1 2 82124 92742
0 32694 5 1 1 32693
0 32695 7 1 2 32690 32694
0 32696 5 1 1 32695
0 32697 7 1 2 92438 32696
0 32698 5 1 1 32697
0 32699 7 2 2 70818 87122
0 32700 5 1 1 92744
0 32701 7 1 2 62475 79124
0 32702 5 2 1 32701
0 32703 7 1 2 32700 92746
0 32704 5 2 1 32703
0 32705 7 1 2 68095 92748
0 32706 5 1 1 32705
0 32707 7 2 2 81839 72193
0 32708 5 5 1 92750
0 32709 7 1 2 67326 92752
0 32710 7 1 2 32706 32709
0 32711 5 2 1 32710
0 32712 7 1 2 62223 92757
0 32713 5 1 1 32712
0 32714 7 3 2 72245 73898
0 32715 5 1 1 92759
0 32716 7 2 2 67327 78317
0 32717 5 1 1 92762
0 32718 7 1 2 32715 32717
0 32719 5 1 1 32718
0 32720 7 1 2 80208 84544
0 32721 5 7 1 32720
0 32722 7 1 2 78213 92764
0 32723 5 1 1 32722
0 32724 7 2 2 32719 32723
0 32725 7 3 2 57712 79795
0 32726 7 2 2 69973 69875
0 32727 7 1 2 92773 92776
0 32728 5 2 1 32727
0 32729 7 1 2 64352 92778
0 32730 5 1 1 32729
0 32731 7 1 2 92771 32730
0 32732 7 1 2 32713 32731
0 32733 5 1 1 32732
0 32734 7 1 2 60971 32733
0 32735 5 1 1 32734
0 32736 7 1 2 68096 79055
0 32737 5 3 1 32736
0 32738 7 1 2 73580 92780
0 32739 5 1 1 32738
0 32740 7 1 2 68244 32739
0 32741 5 1 1 32740
0 32742 7 1 2 72526 32741
0 32743 5 1 1 32742
0 32744 7 1 2 60603 32743
0 32745 5 1 1 32744
0 32746 7 1 2 65278 68206
0 32747 5 3 1 32746
0 32748 7 2 2 73294 92783
0 32749 5 1 1 92786
0 32750 7 1 2 73598 92787
0 32751 5 1 1 32750
0 32752 7 4 2 62224 68097
0 32753 5 2 1 92788
0 32754 7 1 2 64353 92789
0 32755 5 1 1 32754
0 32756 7 1 2 32751 32755
0 32757 5 1 1 32756
0 32758 7 1 2 69038 32757
0 32759 5 1 1 32758
0 32760 7 1 2 73599 72335
0 32761 5 1 1 32760
0 32762 7 1 2 72527 32761
0 32763 5 1 1 32762
0 32764 7 1 2 87990 32763
0 32765 5 1 1 32764
0 32766 7 1 2 87691 84398
0 32767 5 1 1 32766
0 32768 7 1 2 77914 32767
0 32769 7 1 2 32765 32768
0 32770 7 1 2 32759 32769
0 32771 7 1 2 32745 32770
0 32772 7 1 2 32735 32771
0 32773 5 1 1 32772
0 32774 7 1 2 79553 32773
0 32775 5 1 1 32774
0 32776 7 4 2 71686 79671
0 32777 5 2 1 92794
0 32778 7 1 2 90086 92795
0 32779 5 1 1 32778
0 32780 7 1 2 79563 32779
0 32781 5 1 1 32780
0 32782 7 5 2 62225 64354
0 32783 5 1 1 92800
0 32784 7 1 2 60972 92801
0 32785 7 1 2 32781 32784
0 32786 5 1 1 32785
0 32787 7 1 2 32775 32786
0 32788 5 1 1 32787
0 32789 7 1 2 61342 32788
0 32790 5 1 1 32789
0 32791 7 1 2 32698 32790
0 32792 5 1 1 32791
0 32793 7 1 2 63053 32792
0 32794 5 1 1 32793
0 32795 7 3 2 58754 73364
0 32796 5 1 1 92805
0 32797 7 1 2 73124 79083
0 32798 5 1 1 32797
0 32799 7 1 2 73125 76355
0 32800 5 2 1 32799
0 32801 7 1 2 57432 92808
0 32802 5 1 1 32801
0 32803 7 2 2 71687 75088
0 32804 5 2 1 92810
0 32805 7 1 2 73175 92812
0 32806 5 3 1 32805
0 32807 7 1 2 63904 92814
0 32808 7 1 2 32802 32807
0 32809 5 1 1 32808
0 32810 7 1 2 32798 32809
0 32811 5 1 1 32810
0 32812 7 1 2 62476 32811
0 32813 5 1 1 32812
0 32814 7 1 2 62226 81627
0 32815 5 2 1 32814
0 32816 7 2 2 81597 92817
0 32817 5 5 1 92819
0 32818 7 1 2 73126 92821
0 32819 5 1 1 32818
0 32820 7 2 2 32813 32819
0 32821 5 2 1 92826
0 32822 7 1 2 64355 92828
0 32823 5 2 1 32822
0 32824 7 2 2 2412 91070
0 32825 5 1 1 92832
0 32826 7 1 2 75200 3702
0 32827 7 1 2 92833 32826
0 32828 5 1 1 32827
0 32829 7 1 2 63905 32828
0 32830 5 1 1 32829
0 32831 7 1 2 65616 78411
0 32832 5 1 1 32831
0 32833 7 1 2 70210 87397
0 32834 7 1 2 32832 32833
0 32835 5 1 1 32834
0 32836 7 1 2 32830 32835
0 32837 5 1 1 32836
0 32838 7 1 2 62477 32837
0 32839 5 1 1 32838
0 32840 7 1 2 60973 86766
0 32841 5 1 1 32840
0 32842 7 1 2 73176 77530
0 32843 5 1 1 32842
0 32844 7 1 2 75089 32843
0 32845 5 1 1 32844
0 32846 7 1 2 32841 32845
0 32847 7 1 2 32839 32846
0 32848 5 1 1 32847
0 32849 7 1 2 64356 32848
0 32850 5 1 1 32849
0 32851 7 1 2 76801 90499
0 32852 5 2 1 32851
0 32853 7 1 2 32850 92834
0 32854 5 1 1 32853
0 32855 7 1 2 62753 32854
0 32856 5 1 1 32855
0 32857 7 1 2 92830 32856
0 32858 5 1 1 32857
0 32859 7 1 2 92806 32858
0 32860 5 1 1 32859
0 32861 7 1 2 32794 32860
0 32862 5 1 1 32861
0 32863 7 1 2 63324 32862
0 32864 5 1 1 32863
0 32865 7 1 2 71825 71688
0 32866 5 1 1 32865
0 32867 7 1 2 62478 92745
0 32868 5 1 1 32867
0 32869 7 2 2 32866 32868
0 32870 5 1 1 92836
0 32871 7 1 2 65962 92837
0 32872 5 1 1 32871
0 32873 7 1 2 62754 32872
0 32874 5 1 1 32873
0 32875 7 1 2 4136 32874
0 32876 5 1 1 32875
0 32877 7 1 2 85152 32876
0 32878 5 1 1 32877
0 32879 7 1 2 75132 81159
0 32880 5 1 1 32879
0 32881 7 1 2 85130 32880
0 32882 5 1 1 32881
0 32883 7 1 2 63325 67756
0 32884 5 1 1 32883
0 32885 7 1 2 57433 84322
0 32886 7 1 2 32884 32885
0 32887 5 1 1 32886
0 32888 7 1 2 32882 32887
0 32889 5 1 1 32888
0 32890 7 1 2 67328 92781
0 32891 5 2 1 32890
0 32892 7 1 2 81167 92838
0 32893 5 1 1 32892
0 32894 7 1 2 86021 32893
0 32895 7 1 2 32889 32894
0 32896 5 1 1 32895
0 32897 7 1 2 61343 32896
0 32898 5 1 1 32897
0 32899 7 2 2 72194 81656
0 32900 5 1 1 92840
0 32901 7 1 2 83913 92841
0 32902 5 1 1 32901
0 32903 7 5 2 71689 78243
0 32904 5 1 1 92842
0 32905 7 1 2 84320 92843
0 32906 5 1 1 32905
0 32907 7 1 2 32902 32906
0 32908 7 1 2 32898 32907
0 32909 5 1 1 32908
0 32910 7 1 2 60974 32909
0 32911 5 1 1 32910
0 32912 7 1 2 63326 73414
0 32913 5 1 1 32912
0 32914 7 2 2 60604 80703
0 32915 5 1 1 92847
0 32916 7 1 2 90577 92848
0 32917 5 1 1 32916
0 32918 7 1 2 32913 32917
0 32919 5 1 1 32918
0 32920 7 1 2 71290 32919
0 32921 5 1 1 32920
0 32922 7 1 2 32911 32921
0 32923 7 1 2 32878 32922
0 32924 5 1 1 32923
0 32925 7 1 2 70211 32924
0 32926 5 1 1 32925
0 32927 7 1 2 82922 70212
0 32928 5 2 1 32927
0 32929 7 1 2 91622 92849
0 32930 5 1 1 32929
0 32931 7 1 2 62227 32930
0 32932 5 1 1 32931
0 32933 7 1 2 21009 26107
0 32934 5 1 1 32933
0 32935 7 1 2 71291 32934
0 32936 5 1 1 32935
0 32937 7 2 2 85153 92790
0 32938 5 1 1 92851
0 32939 7 1 2 73882 92852
0 32940 5 1 1 32939
0 32941 7 1 2 32936 32940
0 32942 5 1 1 32941
0 32943 7 1 2 81086 32942
0 32944 5 1 1 32943
0 32945 7 4 2 61344 85482
0 32946 5 1 1 92853
0 32947 7 1 2 62479 92784
0 32948 5 2 1 32947
0 32949 7 1 2 72058 32938
0 32950 7 1 2 92857 32949
0 32951 5 1 1 32950
0 32952 7 1 2 92854 32951
0 32953 5 1 1 32952
0 32954 7 1 2 32944 32953
0 32955 7 1 2 32932 32954
0 32956 5 1 1 32955
0 32957 7 1 2 69039 32956
0 32958 5 1 1 32957
0 32959 7 1 2 65963 89419
0 32960 5 1 1 32959
0 32961 7 1 2 63327 32960
0 32962 5 1 1 32961
0 32963 7 1 2 58054 11078
0 32964 5 1 1 32963
0 32965 7 2 2 63906 61345
0 32966 7 1 2 91554 92859
0 32967 5 1 1 32966
0 32968 7 1 2 58576 32967
0 32969 5 1 1 32968
0 32970 7 1 2 60605 32969
0 32971 7 1 2 32964 32970
0 32972 5 1 1 32971
0 32973 7 1 2 32962 32972
0 32974 5 1 1 32973
0 32975 7 1 2 78659 32974
0 32976 5 1 1 32975
0 32977 7 1 2 75467 72336
0 32978 5 1 1 32977
0 32979 7 1 2 84879 32978
0 32980 5 1 1 32979
0 32981 7 1 2 81144 32980
0 32982 5 1 1 32981
0 32983 7 1 2 85154 85836
0 32984 5 1 1 32983
0 32985 7 1 2 32984 92850
0 32986 7 1 2 32982 32985
0 32987 7 1 2 62228 78485
0 32988 5 2 1 32987
0 32989 7 1 2 77434 92861
0 32990 5 1 1 32989
0 32991 7 1 2 90858 32990
0 32992 5 1 1 32991
0 32993 7 1 2 72337 90056
0 32994 7 1 2 90846 32993
0 32995 5 1 1 32994
0 32996 7 1 2 32992 32995
0 32997 7 1 2 32986 32996
0 32998 5 1 1 32997
0 32999 7 1 2 87991 32998
0 33000 5 1 1 32999
0 33001 7 1 2 61346 92368
0 33002 5 1 1 33001
0 33003 7 1 2 78576 33002
0 33004 5 1 1 33003
0 33005 7 1 2 73127 33004
0 33006 5 1 1 33005
0 33007 7 1 2 21960 33006
0 33008 5 1 1 33007
0 33009 7 1 2 77674 33008
0 33010 5 1 1 33009
0 33011 7 1 2 89417 92855
0 33012 5 1 1 33011
0 33013 7 1 2 78486 77675
0 33014 5 1 1 33013
0 33015 7 1 2 58577 33014
0 33016 5 1 1 33015
0 33017 7 1 2 91589 33016
0 33018 5 1 1 33017
0 33019 7 1 2 33012 33018
0 33020 7 1 2 33010 33019
0 33021 7 1 2 33000 33020
0 33022 7 1 2 32976 33021
0 33023 7 1 2 32958 33022
0 33024 7 2 2 32926 33023
0 33025 5 1 1 92863
0 33026 7 1 2 59848 92864
0 33027 5 1 1 33026
0 33028 7 1 2 72904 83814
0 33029 5 1 1 33028
0 33030 7 1 2 85409 33029
0 33031 5 1 1 33030
0 33032 7 1 2 65617 33031
0 33033 5 1 1 33032
0 33034 7 2 2 59133 73314
0 33035 5 1 1 92865
0 33036 7 1 2 74147 85410
0 33037 7 1 2 33035 33036
0 33038 5 1 1 33037
0 33039 7 1 2 81582 33038
0 33040 5 1 1 33039
0 33041 7 1 2 72905 69128
0 33042 5 1 1 33041
0 33043 7 1 2 73331 33042
0 33044 5 1 1 33043
0 33045 7 1 2 57713 33044
0 33046 5 1 1 33045
0 33047 7 1 2 58984 73315
0 33048 5 2 1 33047
0 33049 7 1 2 65054 73232
0 33050 5 1 1 33049
0 33051 7 1 2 92867 33050
0 33052 5 1 1 33051
0 33053 7 1 2 57434 33052
0 33054 5 1 1 33053
0 33055 7 1 2 33046 33054
0 33056 7 1 2 33040 33055
0 33057 5 1 1 33056
0 33058 7 1 2 65279 33057
0 33059 5 1 1 33058
0 33060 7 1 2 33033 33059
0 33061 5 1 1 33060
0 33062 7 1 2 63328 33061
0 33063 5 1 1 33062
0 33064 7 1 2 68431 87721
0 33065 5 1 1 33064
0 33066 7 1 2 67757 77045
0 33067 5 2 1 33066
0 33068 7 1 2 90754 92869
0 33069 5 1 1 33068
0 33070 7 1 2 73666 33069
0 33071 5 1 1 33070
0 33072 7 1 2 33065 33071
0 33073 5 1 1 33072
0 33074 7 1 2 62229 33073
0 33075 5 1 1 33074
0 33076 7 1 2 86246 77009
0 33077 5 1 1 33076
0 33078 7 1 2 33075 33077
0 33079 5 1 1 33078
0 33080 7 1 2 69040 33079
0 33081 5 1 1 33080
0 33082 7 1 2 68245 78648
0 33083 5 4 1 33082
0 33084 7 2 2 65280 92871
0 33085 5 1 1 92875
0 33086 7 1 2 60975 33085
0 33087 5 1 1 33086
0 33088 7 1 2 78172 80480
0 33089 5 12 1 33088
0 33090 7 3 2 67329 92877
0 33091 5 1 1 92889
0 33092 7 1 2 33087 92890
0 33093 5 1 1 33092
0 33094 7 1 2 78813 80506
0 33095 5 1 1 33094
0 33096 7 1 2 68098 87722
0 33097 7 1 2 33095 33096
0 33098 5 1 1 33097
0 33099 7 1 2 78487 89457
0 33100 7 1 2 87992 33099
0 33101 5 1 1 33100
0 33102 7 3 2 60393 77493
0 33103 5 2 1 92892
0 33104 7 1 2 73781 92893
0 33105 7 1 2 89714 33104
0 33106 5 1 1 33105
0 33107 7 1 2 64571 87031
0 33108 7 1 2 33106 33107
0 33109 7 1 2 33101 33108
0 33110 7 1 2 33098 33109
0 33111 7 1 2 33093 33110
0 33112 7 1 2 80563 81619
0 33113 5 1 1 33112
0 33114 7 3 2 65964 89715
0 33115 5 1 1 92897
0 33116 7 1 2 81628 92898
0 33117 5 1 1 33116
0 33118 7 1 2 33113 33117
0 33119 5 1 1 33118
0 33120 7 1 2 62480 33119
0 33121 5 1 1 33120
0 33122 7 5 2 58985 73464
0 33123 5 2 1 92900
0 33124 7 1 2 80579 92905
0 33125 5 1 1 33124
0 33126 7 1 2 72704 33125
0 33127 5 1 1 33126
0 33128 7 1 2 72059 87084
0 33129 5 1 1 33128
0 33130 7 1 2 72873 33129
0 33131 7 1 2 33127 33130
0 33132 5 1 1 33131
0 33133 7 1 2 70410 85878
0 33134 7 1 2 33132 33133
0 33135 5 1 1 33134
0 33136 7 1 2 33121 33135
0 33137 7 1 2 33111 33136
0 33138 7 1 2 33081 33137
0 33139 7 1 2 33063 33138
0 33140 7 1 2 80564 83358
0 33141 5 1 1 33140
0 33142 7 1 2 67758 82489
0 33143 5 2 1 33142
0 33144 7 4 2 67330 92907
0 33145 5 1 1 92909
0 33146 7 1 2 58313 92910
0 33147 5 2 1 33146
0 33148 7 1 2 78860 92913
0 33149 5 1 1 33148
0 33150 7 1 2 80238 80922
0 33151 5 1 1 33150
0 33152 7 1 2 62755 33151
0 33153 5 1 1 33152
0 33154 7 1 2 87601 33153
0 33155 7 1 2 33149 33154
0 33156 5 1 1 33155
0 33157 7 1 2 73667 33156
0 33158 5 1 1 33157
0 33159 7 1 2 33141 33158
0 33160 5 1 1 33159
0 33161 7 1 2 60976 33160
0 33162 5 1 1 33161
0 33163 7 1 2 68999 73449
0 33164 5 1 1 33163
0 33165 7 1 2 73787 33164
0 33166 5 1 1 33165
0 33167 7 1 2 57714 33166
0 33168 5 1 1 33167
0 33169 7 1 2 73531 69129
0 33170 5 2 1 33169
0 33171 7 1 2 33168 92915
0 33172 5 1 1 33171
0 33173 7 1 2 67331 33172
0 33174 5 1 1 33173
0 33175 7 1 2 76328 75890
0 33176 5 1 1 33175
0 33177 7 1 2 78861 33176
0 33178 5 1 1 33177
0 33179 7 2 2 67759 83949
0 33180 5 2 1 92917
0 33181 7 3 2 73934 92919
0 33182 7 2 2 60606 68432
0 33183 5 1 1 92924
0 33184 7 1 2 58314 33183
0 33185 7 1 2 92921 33184
0 33186 7 1 2 33178 33185
0 33187 5 2 1 33186
0 33188 7 1 2 58578 92926
0 33189 5 1 1 33188
0 33190 7 1 2 84431 33189
0 33191 7 1 2 33174 33190
0 33192 5 1 1 33191
0 33193 7 1 2 64357 33192
0 33194 5 1 1 33193
0 33195 7 1 2 33162 33194
0 33196 7 1 2 33139 33195
0 33197 5 1 1 33196
0 33198 7 1 2 63503 33197
0 33199 7 1 2 33027 33198
0 33200 5 1 1 33199
0 33201 7 1 2 85609 79465
0 33202 7 1 2 86870 33201
0 33203 5 1 1 33202
0 33204 7 1 2 33200 33203
0 33205 7 1 2 32864 33204
0 33206 5 1 1 33205
0 33207 7 1 2 61857 33206
0 33208 5 1 1 33207
0 33209 7 2 2 60607 89075
0 33210 5 1 1 92928
0 33211 7 1 2 84372 92929
0 33212 5 1 1 33211
0 33213 7 1 2 71690 90727
0 33214 5 1 1 33213
0 33215 7 1 2 67332 33214
0 33216 5 1 1 33215
0 33217 7 1 2 62230 33216
0 33218 5 2 1 33217
0 33219 7 1 2 67203 74817
0 33220 5 1 1 33219
0 33221 7 1 2 92930 33220
0 33222 5 1 1 33221
0 33223 7 1 2 70819 33222
0 33224 5 1 1 33223
0 33225 7 1 2 91057 92765
0 33226 5 1 1 33225
0 33227 7 1 2 67333 83934
0 33228 5 1 1 33227
0 33229 7 1 2 70045 33228
0 33230 5 1 1 33229
0 33231 7 1 2 71503 33230
0 33232 5 1 1 33231
0 33233 7 1 2 68099 33232
0 33234 5 1 1 33233
0 33235 7 1 2 33226 33234
0 33236 7 1 2 33224 33235
0 33237 5 1 1 33236
0 33238 7 1 2 78047 33237
0 33239 5 1 1 33238
0 33240 7 1 2 33212 33239
0 33241 5 1 1 33240
0 33242 7 1 2 61347 33241
0 33243 5 1 1 33242
0 33244 7 1 2 64089 88930
0 33245 5 1 1 33244
0 33246 7 1 2 92931 33245
0 33247 5 1 1 33246
0 33248 7 1 2 70820 33247
0 33249 5 1 1 33248
0 33250 7 1 2 78349 92766
0 33251 5 1 1 33250
0 33252 7 1 2 33249 33251
0 33253 5 1 1 33252
0 33254 7 1 2 60977 33253
0 33255 5 1 1 33254
0 33256 7 1 2 90750 92477
0 33257 5 1 1 33256
0 33258 7 2 2 67760 85363
0 33259 5 1 1 92932
0 33260 7 1 2 80378 33259
0 33261 7 1 2 81197 33260
0 33262 5 1 1 33261
0 33263 7 1 2 81075 33262
0 33264 5 1 1 33263
0 33265 7 1 2 67334 33264
0 33266 5 1 1 33265
0 33267 7 1 2 61348 33266
0 33268 5 1 1 33267
0 33269 7 1 2 33257 33268
0 33270 7 1 2 33255 33269
0 33271 5 1 1 33270
0 33272 7 1 2 71433 33271
0 33273 5 1 1 33272
0 33274 7 1 2 84201 85813
0 33275 5 2 1 33274
0 33276 7 1 2 58315 87700
0 33277 5 1 1 33276
0 33278 7 2 2 92934 33277
0 33279 7 1 2 67204 92936
0 33280 5 1 1 33279
0 33281 7 1 2 91445 33280
0 33282 5 1 1 33281
0 33283 7 1 2 57715 77041
0 33284 5 3 1 33283
0 33285 7 1 2 80583 92938
0 33286 7 1 2 33282 33285
0 33287 5 1 1 33286
0 33288 7 1 2 33273 33287
0 33289 7 1 2 33243 33288
0 33290 5 1 1 33289
0 33291 7 16 2 63504 66487
0 33292 7 1 2 75549 92941
0 33293 7 1 2 33290 33292
0 33294 5 1 1 33293
0 33295 7 1 2 60011 33294
0 33296 7 1 2 33208 33295
0 33297 5 1 1 33296
0 33298 7 1 2 63054 78835
0 33299 5 1 1 33298
0 33300 7 1 2 90376 33299
0 33301 5 1 1 33300
0 33302 7 1 2 68521 33301
0 33303 5 1 1 33302
0 33304 7 1 2 63055 80941
0 33305 5 1 1 33304
0 33306 7 1 2 33303 33305
0 33307 5 1 1 33306
0 33308 7 1 2 68100 33307
0 33309 5 1 1 33308
0 33310 7 1 2 13641 33309
0 33311 5 1 1 33310
0 33312 7 1 2 82803 33311
0 33313 5 1 1 33312
0 33314 7 1 2 76923 87247
0 33315 5 1 1 33314
0 33316 7 1 2 82804 84373
0 33317 5 2 1 33316
0 33318 7 1 2 65281 76924
0 33319 5 1 1 33318
0 33320 7 1 2 92957 33319
0 33321 5 1 1 33320
0 33322 7 1 2 76959 33321
0 33323 5 1 1 33322
0 33324 7 1 2 33315 33323
0 33325 7 1 2 33313 33324
0 33326 5 1 1 33325
0 33327 7 1 2 60394 33326
0 33328 5 1 1 33327
0 33329 7 1 2 86168 83136
0 33330 5 1 1 33329
0 33331 7 1 2 30594 92958
0 33332 5 1 1 33331
0 33333 7 1 2 33330 33332
0 33334 5 1 1 33333
0 33335 7 1 2 69424 76925
0 33336 5 1 1 33335
0 33337 7 1 2 71504 84829
0 33338 5 1 1 33337
0 33339 7 1 2 71292 82805
0 33340 7 1 2 33338 33339
0 33341 5 1 1 33340
0 33342 7 1 2 33336 33341
0 33343 5 1 1 33342
0 33344 7 1 2 68101 33343
0 33345 5 1 1 33344
0 33346 7 1 2 33334 33345
0 33347 7 1 2 33328 33346
0 33348 5 1 1 33347
0 33349 7 1 2 66488 33348
0 33350 5 1 1 33349
0 33351 7 2 2 61858 91826
0 33352 7 1 2 68007 79597
0 33353 5 2 1 33352
0 33354 7 1 2 92959 92961
0 33355 5 1 1 33354
0 33356 7 1 2 87248 92942
0 33357 5 1 1 33356
0 33358 7 2 2 69192 88733
0 33359 7 4 2 58579 59134
0 33360 7 1 2 76865 92965
0 33361 7 1 2 92963 33360
0 33362 5 1 1 33361
0 33363 7 1 2 33357 33362
0 33364 5 1 1 33363
0 33365 7 1 2 91915 33364
0 33366 5 1 1 33365
0 33367 7 1 2 33355 33366
0 33368 7 1 2 33350 33367
0 33369 5 1 1 33368
0 33370 7 1 2 60978 33369
0 33371 5 1 1 33370
0 33372 7 1 2 74829 92605
0 33373 5 1 1 33372
0 33374 7 1 2 65055 86187
0 33375 5 2 1 33374
0 33376 7 1 2 68380 75201
0 33377 5 2 1 33376
0 33378 7 1 2 92969 92971
0 33379 5 1 1 33378
0 33380 7 1 2 92943 33379
0 33381 5 1 1 33380
0 33382 7 14 2 58755 61859
0 33383 5 4 1 92973
0 33384 7 1 2 57435 92944
0 33385 5 1 1 33384
0 33386 7 1 2 92987 33385
0 33387 5 2 1 33386
0 33388 7 1 2 81583 92991
0 33389 5 1 1 33388
0 33390 7 1 2 82784 92715
0 33391 5 1 1 33390
0 33392 7 1 2 79515 92945
0 33393 5 1 1 33392
0 33394 7 1 2 33391 33393
0 33395 7 1 2 33389 33394
0 33396 5 1 1 33395
0 33397 7 1 2 65282 33396
0 33398 5 1 1 33397
0 33399 7 1 2 58756 89496
0 33400 5 1 1 33399
0 33401 7 1 2 33398 33400
0 33402 7 1 2 33381 33401
0 33403 5 1 1 33402
0 33404 7 1 2 58316 33403
0 33405 5 1 1 33404
0 33406 7 1 2 33373 33405
0 33407 5 1 1 33406
0 33408 7 1 2 67335 33407
0 33409 5 1 1 33408
0 33410 7 1 2 71032 89816
0 33411 5 1 1 33410
0 33412 7 1 2 70411 33411
0 33413 5 1 1 33412
0 33414 7 1 2 70821 84924
0 33415 7 1 2 33413 33414
0 33416 5 1 1 33415
0 33417 7 1 2 81862 17889
0 33418 5 2 1 33417
0 33419 7 1 2 78350 92993
0 33420 5 1 1 33419
0 33421 7 2 2 63056 92767
0 33422 5 1 1 92995
0 33423 7 1 2 33420 33422
0 33424 7 1 2 33416 33423
0 33425 5 2 1 33424
0 33426 7 1 2 82806 92997
0 33427 5 1 1 33426
0 33428 7 1 2 86251 76013
0 33429 5 1 1 33428
0 33430 7 1 2 33427 33429
0 33431 5 1 1 33430
0 33432 7 1 2 66489 33431
0 33433 5 1 1 33432
0 33434 7 1 2 81598 92974
0 33435 5 1 1 33434
0 33436 7 2 2 65283 92946
0 33437 7 1 2 59135 92999
0 33438 5 1 1 33437
0 33439 7 1 2 33435 33438
0 33440 5 1 1 33439
0 33441 7 1 2 57716 33440
0 33442 5 1 1 33441
0 33443 7 1 2 80048 92975
0 33444 5 1 1 33443
0 33445 7 1 2 72390 92947
0 33446 7 1 2 76075 33445
0 33447 5 1 1 33446
0 33448 7 1 2 33444 33447
0 33449 7 1 2 33442 33448
0 33450 5 1 1 33449
0 33451 7 1 2 65618 33450
0 33452 5 1 1 33451
0 33453 7 1 2 63782 82790
0 33454 5 1 1 33453
0 33455 7 1 2 65284 33454
0 33456 7 1 2 92992 33455
0 33457 5 1 1 33456
0 33458 7 4 2 65619 92948
0 33459 7 1 2 58986 93001
0 33460 5 1 1 33459
0 33461 7 1 2 33457 33460
0 33462 5 1 1 33461
0 33463 7 1 2 72379 33462
0 33464 5 1 1 33463
0 33465 7 1 2 33452 33464
0 33466 5 1 1 33465
0 33467 7 1 2 70412 33466
0 33468 5 1 1 33467
0 33469 7 2 2 68008 92976
0 33470 5 1 1 93005
0 33471 7 1 2 58317 93006
0 33472 5 1 1 33471
0 33473 7 1 2 33468 33472
0 33474 7 1 2 33433 33473
0 33475 7 1 2 33409 33474
0 33476 5 1 1 33475
0 33477 7 1 2 64358 33476
0 33478 5 1 1 33477
0 33479 7 2 2 78719 92949
0 33480 5 2 1 93007
0 33481 7 1 2 57436 93009
0 33482 5 1 1 33481
0 33483 7 1 2 92988 93010
0 33484 5 2 1 33483
0 33485 7 1 2 68102 93011
0 33486 7 1 2 33482 33485
0 33487 5 1 1 33486
0 33488 7 1 2 71826 92977
0 33489 5 1 1 33488
0 33490 7 1 2 92978 92785
0 33491 5 1 1 33490
0 33492 7 1 2 71827 93002
0 33493 5 2 1 33492
0 33494 7 1 2 33491 93013
0 33495 5 1 1 33494
0 33496 7 1 2 62481 33495
0 33497 5 1 1 33496
0 33498 7 1 2 33489 33497
0 33499 7 1 2 33487 33498
0 33500 5 1 1 33499
0 33501 7 1 2 58580 33500
0 33502 5 1 1 33501
0 33503 7 2 2 58757 84413
0 33504 7 1 2 64090 80816
0 33505 7 1 2 89860 33504
0 33506 7 1 2 93015 33505
0 33507 5 1 1 33506
0 33508 7 1 2 33502 33507
0 33509 5 1 1 33508
0 33510 7 1 2 69041 33509
0 33511 5 1 1 33510
0 33512 7 1 2 84925 93003
0 33513 5 1 1 33512
0 33514 7 1 2 92989 33513
0 33515 5 1 1 33514
0 33516 7 1 2 68103 33515
0 33517 5 1 1 33516
0 33518 7 1 2 80934 93008
0 33519 5 1 1 33518
0 33520 7 1 2 33517 33519
0 33521 5 1 1 33520
0 33522 7 1 2 58581 33521
0 33523 5 1 1 33522
0 33524 7 1 2 86423 91353
0 33525 7 1 2 83995 33524
0 33526 5 1 1 33525
0 33527 7 1 2 33523 33526
0 33528 5 1 1 33527
0 33529 7 1 2 70822 33528
0 33530 5 1 1 33529
0 33531 7 2 2 59374 76317
0 33532 5 3 1 93017
0 33533 7 1 2 92960 93019
0 33534 5 1 1 33533
0 33535 7 1 2 63505 80587
0 33536 5 1 1 33535
0 33537 7 2 2 71828 76886
0 33538 5 1 1 93022
0 33539 7 1 2 82807 93023
0 33540 5 1 1 33539
0 33541 7 1 2 33536 33540
0 33542 5 1 1 33541
0 33543 7 1 2 87114 92618
0 33544 7 1 2 33542 33543
0 33545 5 1 1 33544
0 33546 7 1 2 33534 33545
0 33547 5 1 1 33546
0 33548 7 1 2 78296 33547
0 33549 5 1 1 33548
0 33550 7 1 2 81620 72365
0 33551 5 1 1 33550
0 33552 7 1 2 76150 33551
0 33553 5 1 1 33552
0 33554 7 1 2 92979 33553
0 33555 5 1 1 33554
0 33556 7 1 2 81853 84545
0 33557 5 1 1 33556
0 33558 7 1 2 60979 80386
0 33559 5 2 1 33558
0 33560 7 1 2 92950 93024
0 33561 7 1 2 33557 33560
0 33562 5 1 1 33561
0 33563 7 1 2 33555 33562
0 33564 5 1 1 33563
0 33565 7 1 2 58582 33564
0 33566 5 1 1 33565
0 33567 7 1 2 61349 33566
0 33568 7 1 2 33549 33567
0 33569 7 1 2 33530 33568
0 33570 7 1 2 33511 33569
0 33571 7 1 2 33478 33570
0 33572 7 1 2 33371 33571
0 33573 5 1 1 33572
0 33574 7 1 2 83815 92980
0 33575 5 1 1 33574
0 33576 7 1 2 77216 90184
0 33577 7 1 2 74556 33576
0 33578 5 1 1 33577
0 33579 7 1 2 33575 33578
0 33580 5 1 1 33579
0 33581 7 1 2 67336 33580
0 33582 5 1 1 33581
0 33583 7 2 2 58583 79606
0 33584 5 2 1 93026
0 33585 7 1 2 70413 82158
0 33586 5 1 1 33585
0 33587 7 1 2 93028 33586
0 33588 5 1 1 33587
0 33589 7 1 2 92951 33588
0 33590 5 1 1 33589
0 33591 7 1 2 33582 33590
0 33592 5 1 1 33591
0 33593 7 1 2 64359 33592
0 33594 5 1 1 33593
0 33595 7 4 2 58758 89871
0 33596 5 2 1 93030
0 33597 7 1 2 81453 92452
0 33598 5 1 1 33597
0 33599 7 1 2 93034 33598
0 33600 5 1 1 33599
0 33601 7 1 2 76205 33600
0 33602 5 1 1 33601
0 33603 7 1 2 66490 78120
0 33604 7 1 2 75369 33603
0 33605 5 1 1 33604
0 33606 7 1 2 62231 83637
0 33607 7 1 2 89443 33606
0 33608 5 1 1 33607
0 33609 7 1 2 33605 33608
0 33610 5 1 1 33609
0 33611 7 1 2 69042 33610
0 33612 5 1 1 33611
0 33613 7 1 2 62232 92453
0 33614 5 1 1 33613
0 33615 7 1 2 93035 33614
0 33616 5 1 1 33615
0 33617 7 1 2 83871 33616
0 33618 5 1 1 33617
0 33619 7 1 2 33612 33618
0 33620 5 1 1 33619
0 33621 7 1 2 68104 33620
0 33622 5 1 1 33621
0 33623 7 1 2 33602 33622
0 33624 7 1 2 33594 33623
0 33625 5 1 1 33624
0 33626 7 1 2 60608 33625
0 33627 5 1 1 33626
0 33628 7 2 2 74929 88182
0 33629 5 1 1 93036
0 33630 7 1 2 5996 33629
0 33631 5 1 1 33630
0 33632 7 1 2 68105 33631
0 33633 5 1 1 33632
0 33634 7 1 2 76206 73760
0 33635 5 1 1 33634
0 33636 7 1 2 75454 33635
0 33637 5 2 1 33636
0 33638 7 1 2 83819 93038
0 33639 5 1 1 33638
0 33640 7 1 2 33633 33639
0 33641 5 1 1 33640
0 33642 7 1 2 92952 33641
0 33643 5 1 1 33642
0 33644 7 1 2 62233 93000
0 33645 5 1 1 33644
0 33646 7 1 2 92990 33645
0 33647 5 1 1 33646
0 33648 7 1 2 89716 33647
0 33649 5 1 1 33648
0 33650 7 1 2 66491 89458
0 33651 7 1 2 90303 33650
0 33652 5 1 1 33651
0 33653 7 1 2 33649 33652
0 33654 5 1 1 33653
0 33655 7 1 2 87993 33654
0 33656 5 1 1 33655
0 33657 7 1 2 76151 88816
0 33658 5 7 1 33657
0 33659 7 1 2 78840 93040
0 33660 5 1 1 33659
0 33661 7 1 2 68106 89418
0 33662 5 1 1 33661
0 33663 7 1 2 70414 33662
0 33664 7 1 2 33660 33663
0 33665 5 1 1 33664
0 33666 7 1 2 93031 33665
0 33667 5 1 1 33666
0 33668 7 1 2 33656 33667
0 33669 7 1 2 33643 33668
0 33670 7 1 2 33627 33669
0 33671 5 1 1 33670
0 33672 7 1 2 60980 33671
0 33673 5 1 1 33672
0 33674 7 1 2 78569 93012
0 33675 5 1 1 33674
0 33676 7 1 2 91467 92981
0 33677 5 1 1 33676
0 33678 7 1 2 70371 93004
0 33679 5 1 1 33678
0 33680 7 1 2 33677 33679
0 33681 5 1 1 33680
0 33682 7 1 2 59606 33681
0 33683 5 1 1 33682
0 33684 7 1 2 72510 92454
0 33685 5 1 1 33684
0 33686 7 1 2 33683 33685
0 33687 5 1 1 33686
0 33688 7 1 2 70823 33687
0 33689 5 1 1 33688
0 33690 7 1 2 33675 33689
0 33691 5 1 1 33690
0 33692 7 1 2 78862 33691
0 33693 5 1 1 33692
0 33694 7 1 2 78863 87115
0 33695 5 1 1 33694
0 33696 7 1 2 92760 33695
0 33697 5 1 1 33696
0 33698 7 2 2 90989 92953
0 33699 7 1 2 62482 93047
0 33700 5 1 1 33699
0 33701 7 1 2 63057 93032
0 33702 5 1 1 33701
0 33703 7 1 2 33700 33702
0 33704 5 1 1 33703
0 33705 7 1 2 33697 33704
0 33706 5 1 1 33705
0 33707 7 1 2 62756 93048
0 33708 5 1 1 33707
0 33709 7 1 2 75381 91629
0 33710 5 1 1 33709
0 33711 7 1 2 33708 33710
0 33712 5 1 1 33711
0 33713 7 1 2 75903 33712
0 33714 5 1 1 33713
0 33715 7 1 2 77471 93033
0 33716 5 1 1 33715
0 33717 7 1 2 64360 92455
0 33718 5 1 1 33717
0 33719 7 1 2 33716 33718
0 33720 5 1 1 33719
0 33721 7 1 2 81857 33720
0 33722 5 1 1 33721
0 33723 7 1 2 62757 92982
0 33724 5 1 1 33723
0 33725 7 1 2 93014 33724
0 33726 5 1 1 33725
0 33727 7 1 2 92192 33726
0 33728 5 1 1 33727
0 33729 7 1 2 65965 33728
0 33730 7 1 2 33722 33729
0 33731 7 1 2 33714 33730
0 33732 7 1 2 33706 33731
0 33733 7 1 2 33693 33732
0 33734 7 1 2 33673 33733
0 33735 5 1 1 33734
0 33736 7 1 2 33573 33735
0 33737 5 1 1 33736
0 33738 7 1 2 74341 75329
0 33739 5 2 1 33738
0 33740 7 1 2 61350 93049
0 33741 5 1 1 33740
0 33742 7 1 2 58987 33741
0 33743 5 1 1 33742
0 33744 7 3 2 69452 68381
0 33745 5 1 1 93051
0 33746 7 1 2 67337 93052
0 33747 5 1 1 33746
0 33748 7 1 2 33743 33747
0 33749 5 1 1 33748
0 33750 7 1 2 57437 33749
0 33751 5 1 1 33750
0 33752 7 1 2 65056 67893
0 33753 5 1 1 33752
0 33754 7 1 2 58318 85814
0 33755 5 1 1 33754
0 33756 7 1 2 33753 33755
0 33757 7 1 2 33751 33756
0 33758 5 1 1 33757
0 33759 7 1 2 59607 33758
0 33760 5 1 1 33759
0 33761 7 1 2 78737 83734
0 33762 5 1 1 33761
0 33763 7 1 2 65057 85403
0 33764 7 1 2 33762 33763
0 33765 5 1 1 33764
0 33766 7 1 2 33760 33765
0 33767 5 1 1 33766
0 33768 7 1 2 63506 33767
0 33769 5 1 1 33768
0 33770 7 1 2 62483 92822
0 33771 5 2 1 33770
0 33772 7 3 2 85122 93054
0 33773 5 3 1 93056
0 33774 7 1 2 60981 93059
0 33775 5 1 1 33774
0 33776 7 1 2 76360 81798
0 33777 5 1 1 33776
0 33778 7 1 2 60982 77540
0 33779 5 2 1 33778
0 33780 7 1 2 68780 93062
0 33781 5 1 1 33780
0 33782 7 1 2 62484 89616
0 33783 7 1 2 33781 33782
0 33784 5 1 1 33783
0 33785 7 1 2 70969 93063
0 33786 5 1 1 33785
0 33787 7 1 2 62234 92906
0 33788 7 1 2 33786 33787
0 33789 5 1 1 33788
0 33790 7 2 2 33784 33789
0 33791 7 1 2 33777 93064
0 33792 5 1 1 33791
0 33793 7 1 2 67205 33792
0 33794 5 1 1 33793
0 33795 7 1 2 33775 33794
0 33796 5 1 1 33795
0 33797 7 1 2 72511 75382
0 33798 7 1 2 33796 33797
0 33799 5 1 1 33798
0 33800 7 1 2 33769 33799
0 33801 5 1 1 33800
0 33802 7 1 2 66492 33801
0 33803 5 1 1 33802
0 33804 7 1 2 65620 80056
0 33805 5 2 1 33804
0 33806 7 1 2 65621 81599
0 33807 5 1 1 33806
0 33808 7 1 2 76248 33807
0 33809 5 1 1 33808
0 33810 7 1 2 67338 33809
0 33811 5 1 1 33810
0 33812 7 3 2 65285 70415
0 33813 5 2 1 93068
0 33814 7 3 2 16566 93071
0 33815 5 1 1 93073
0 33816 7 1 2 33811 93074
0 33817 7 1 2 93066 33816
0 33818 5 1 1 33817
0 33819 7 1 2 92954 33818
0 33820 5 1 1 33819
0 33821 7 1 2 33470 33820
0 33822 5 1 1 33821
0 33823 7 1 2 72906 33822
0 33824 5 1 1 33823
0 33825 7 1 2 79804 80717
0 33826 5 1 1 33825
0 33827 7 1 2 68382 33826
0 33828 5 1 1 33827
0 33829 7 3 2 72029 72391
0 33830 5 3 1 93076
0 33831 7 2 2 33828 93079
0 33832 5 1 1 93082
0 33833 7 1 2 75330 84357
0 33834 5 1 1 33833
0 33835 7 1 2 78998 33834
0 33836 7 1 2 93083 33835
0 33837 5 1 1 33836
0 33838 7 1 2 14596 92983
0 33839 7 1 2 33837 33838
0 33840 5 1 1 33839
0 33841 7 1 2 33824 33840
0 33842 7 1 2 33803 33841
0 33843 5 1 1 33842
0 33844 7 1 2 63329 33843
0 33845 5 1 1 33844
0 33846 7 1 2 79455 89446
0 33847 7 1 2 92927 33846
0 33848 5 1 1 33847
0 33849 7 1 2 64572 33848
0 33850 7 1 2 33845 33849
0 33851 7 1 2 33737 33850
0 33852 5 1 1 33851
0 33853 7 1 2 73629 78760
0 33854 5 1 1 33853
0 33855 7 2 2 64361 84079
0 33856 5 1 1 93084
0 33857 7 1 2 68522 79361
0 33858 5 2 1 33857
0 33859 7 1 2 33856 93086
0 33860 5 1 1 33859
0 33861 7 1 2 65966 33860
0 33862 5 1 1 33861
0 33863 7 1 2 33854 33862
0 33864 5 1 1 33863
0 33865 7 1 2 63330 33864
0 33866 5 1 1 33865
0 33867 7 1 2 69743 78761
0 33868 5 1 1 33867
0 33869 7 1 2 74541 80485
0 33870 5 1 1 33869
0 33871 7 1 2 33868 33870
0 33872 5 2 1 33871
0 33873 7 1 2 61351 93088
0 33874 5 1 1 33873
0 33875 7 1 2 79056 75419
0 33876 5 1 1 33875
0 33877 7 1 2 58584 33876
0 33878 5 1 1 33877
0 33879 7 1 2 65967 84080
0 33880 7 1 2 33878 33879
0 33881 5 1 1 33880
0 33882 7 1 2 33874 33881
0 33883 5 1 1 33882
0 33884 7 1 2 63058 33883
0 33885 5 1 1 33884
0 33886 7 1 2 33866 33885
0 33887 5 1 1 33886
0 33888 7 1 2 67761 33887
0 33889 5 1 1 33888
0 33890 7 1 2 80430 74602
0 33891 5 1 1 33890
0 33892 7 1 2 27205 33891
0 33893 5 1 1 33892
0 33894 7 1 2 68869 33893
0 33895 5 1 1 33894
0 33896 7 1 2 65968 92398
0 33897 5 1 1 33896
0 33898 7 1 2 33895 33897
0 33899 5 1 1 33898
0 33900 7 1 2 60609 33899
0 33901 5 1 1 33900
0 33902 7 5 2 61352 68523
0 33903 5 1 1 93090
0 33904 7 2 2 74989 93091
0 33905 5 1 1 93095
0 33906 7 1 2 65286 93096
0 33907 5 1 1 33906
0 33908 7 1 2 86739 33907
0 33909 5 1 1 33908
0 33910 7 1 2 68246 33909
0 33911 5 1 1 33910
0 33912 7 1 2 6193 33911
0 33913 7 1 2 33901 33912
0 33914 5 1 1 33913
0 33915 7 1 2 71293 33914
0 33916 5 1 1 33915
0 33917 7 2 2 61353 78144
0 33918 7 1 2 79383 93097
0 33919 5 1 1 33918
0 33920 7 1 2 65969 68383
0 33921 5 2 1 33920
0 33922 7 1 2 85507 93099
0 33923 7 1 2 79084 33922
0 33924 5 1 1 33923
0 33925 7 1 2 33919 33924
0 33926 5 1 1 33925
0 33927 7 1 2 85155 33926
0 33928 5 1 1 33927
0 33929 7 2 2 70300 78504
0 33930 5 1 1 93101
0 33931 7 1 2 75487 92860
0 33932 7 1 2 93102 33931
0 33933 5 1 1 33932
0 33934 7 1 2 33928 33933
0 33935 7 1 2 33916 33934
0 33936 7 1 2 33889 33935
0 33937 5 1 1 33936
0 33938 7 1 2 68107 33937
0 33939 5 1 1 33938
0 33940 7 1 2 65970 89410
0 33941 5 1 1 33940
0 33942 7 1 2 85416 33941
0 33943 5 1 1 33942
0 33944 7 1 2 69043 33943
0 33945 5 1 1 33944
0 33946 7 1 2 63783 91723
0 33947 5 1 1 33946
0 33948 7 1 2 75031 92544
0 33949 5 1 1 33948
0 33950 7 1 2 33947 33949
0 33951 7 1 2 33945 33950
0 33952 5 1 1 33951
0 33953 7 1 2 60610 33952
0 33954 5 1 1 33953
0 33955 7 4 2 60395 73630
0 33956 5 1 1 93103
0 33957 7 1 2 64091 83904
0 33958 7 1 2 93104 33957
0 33959 5 1 1 33958
0 33960 7 1 2 33954 33959
0 33961 5 1 1 33960
0 33962 7 1 2 63907 33961
0 33963 5 1 1 33962
0 33964 7 1 2 85951 79678
0 33965 5 1 1 33964
0 33966 7 1 2 33963 33965
0 33967 5 1 1 33966
0 33968 7 1 2 62485 33967
0 33969 5 1 1 33968
0 33970 7 1 2 61354 3676
0 33971 5 1 1 33970
0 33972 7 1 2 85555 76960
0 33973 7 1 2 33971 33972
0 33974 5 1 1 33973
0 33975 7 1 2 31139 33974
0 33976 5 1 1 33975
0 33977 7 1 2 60396 33976
0 33978 5 1 1 33977
0 33979 7 1 2 85556 85815
0 33980 7 1 2 87597 33979
0 33981 7 1 2 81200 33980
0 33982 5 1 1 33981
0 33983 7 1 2 33978 33982
0 33984 5 1 1 33983
0 33985 7 1 2 60983 33984
0 33986 5 1 1 33985
0 33987 7 2 2 63331 79371
0 33988 5 1 1 93107
0 33989 7 1 2 61355 93108
0 33990 5 1 1 33989
0 33991 7 1 2 14554 86740
0 33992 5 1 1 33991
0 33993 7 1 2 67206 33992
0 33994 5 1 1 33993
0 33995 7 1 2 33990 33994
0 33996 7 1 2 33986 33995
0 33997 7 1 2 33969 33996
0 33998 5 1 1 33997
0 33999 7 1 2 71294 33998
0 34000 5 1 1 33999
0 34001 7 2 2 33939 34000
0 34002 7 1 2 74483 88933
0 34003 5 1 1 34002
0 34004 7 1 2 65622 92140
0 34005 5 1 1 34004
0 34006 7 1 2 34003 34005
0 34007 5 1 1 34006
0 34008 7 1 2 60611 34007
0 34009 5 1 1 34008
0 34010 7 1 2 72001 93092
0 34011 5 1 1 34010
0 34012 7 1 2 34009 34011
0 34013 5 1 1 34012
0 34014 7 1 2 63908 34013
0 34015 5 1 1 34014
0 34016 7 2 2 85801 83488
0 34017 5 1 1 93111
0 34018 7 1 2 72338 93112
0 34019 5 1 1 34018
0 34020 7 1 2 34015 34019
0 34021 5 1 1 34020
0 34022 7 1 2 62486 34021
0 34023 5 1 1 34022
0 34024 7 1 2 13232 73631
0 34025 5 1 1 34024
0 34026 7 1 2 81198 600
0 34027 5 1 1 34026
0 34028 7 1 2 85802 76974
0 34029 5 1 1 34028
0 34030 7 1 2 60984 85411
0 34031 7 1 2 34029 34030
0 34032 7 1 2 34027 34031
0 34033 5 1 1 34032
0 34034 7 1 2 34025 34033
0 34035 7 1 2 34023 34034
0 34036 5 1 1 34035
0 34037 7 1 2 85156 34036
0 34038 5 1 1 34037
0 34039 7 1 2 60985 86907
0 34040 5 1 1 34039
0 34041 7 1 2 86973 34040
0 34042 5 1 1 34041
0 34043 7 1 2 63059 34042
0 34044 5 1 1 34043
0 34045 7 2 2 34038 34044
0 34046 7 2 2 78488 86635
0 34047 7 1 2 32900 93115
0 34048 5 1 1 34047
0 34049 7 1 2 93113 34048
0 34050 7 1 2 93109 34049
0 34051 5 1 1 34050
0 34052 7 1 2 66493 34051
0 34053 5 1 1 34052
0 34054 7 2 2 63332 69397
0 34055 7 1 2 90963 93117
0 34056 5 2 1 34055
0 34057 7 3 2 58319 72989
0 34058 7 1 2 69118 92964
0 34059 7 1 2 93121 34058
0 34060 5 1 1 34059
0 34061 7 1 2 93119 34060
0 34062 5 1 1 34061
0 34063 7 1 2 57438 34062
0 34064 5 1 1 34063
0 34065 7 1 2 65971 74038
0 34066 5 1 1 34065
0 34067 7 2 2 69876 72409
0 34068 5 2 1 93124
0 34069 7 1 2 34066 93126
0 34070 5 1 1 34069
0 34071 7 1 2 57717 34070
0 34072 5 1 1 34071
0 34073 7 1 2 69000 73953
0 34074 5 2 1 34073
0 34075 7 1 2 34072 93128
0 34076 5 1 1 34075
0 34077 7 1 2 89447 34076
0 34078 5 1 1 34077
0 34079 7 1 2 93120 34078
0 34080 5 1 1 34079
0 34081 7 1 2 67339 34080
0 34082 5 1 1 34081
0 34083 7 1 2 34064 34082
0 34084 7 1 2 34053 34083
0 34085 5 1 1 34084
0 34086 7 1 2 63507 34085
0 34087 5 1 1 34086
0 34088 7 1 2 92984 33025
0 34089 5 1 1 34088
0 34090 7 1 2 59849 34089
0 34091 7 1 2 34087 34090
0 34092 5 1 1 34091
0 34093 7 1 2 33852 34092
0 34094 5 1 1 34093
0 34095 7 1 2 76152 87362
0 34096 5 1 1 34095
0 34097 7 2 2 78489 79496
0 34098 5 1 1 93130
0 34099 7 2 2 34096 93131
0 34100 7 1 2 90449 93132
0 34101 5 1 1 34100
0 34102 7 1 2 65058 92901
0 34103 5 2 1 34102
0 34104 7 1 2 72099 93134
0 34105 5 1 1 34104
0 34106 7 1 2 57718 34105
0 34107 5 2 1 34106
0 34108 7 1 2 74766 75159
0 34109 5 1 1 34108
0 34110 7 1 2 65623 34109
0 34111 5 1 1 34110
0 34112 7 1 2 80713 81584
0 34113 5 1 1 34112
0 34114 7 1 2 71295 73883
0 34115 7 1 2 34113 34114
0 34116 7 1 2 34111 34115
0 34117 7 1 2 93136 34116
0 34118 5 1 1 34117
0 34119 7 4 2 61356 71296
0 34120 5 3 1 93138
0 34121 7 1 2 61860 93142
0 34122 7 1 2 34118 34121
0 34123 5 1 1 34122
0 34124 7 1 2 34101 34123
0 34125 5 1 1 34124
0 34126 7 1 2 92036 34125
0 34127 5 1 1 34126
0 34128 7 1 2 64714 34127
0 34129 7 1 2 34094 34128
0 34130 5 1 1 34129
0 34131 7 1 2 61658 34130
0 34132 7 1 2 33297 34131
0 34133 5 1 1 34132
0 34134 7 1 2 68384 88164
0 34135 5 4 1 34134
0 34136 7 2 2 68108 93145
0 34137 5 1 1 93149
0 34138 7 1 2 87829 93150
0 34139 5 1 1 34138
0 34140 7 1 2 80855 90089
0 34141 7 1 2 34139 34140
0 34142 5 1 1 34141
0 34143 7 2 2 87711 34142
0 34144 7 1 2 88878 93151
0 34145 5 1 1 34144
0 34146 7 1 2 34133 34145
0 34147 5 1 1 34146
0 34148 7 1 2 66711 34147
0 34149 5 1 1 34148
0 34150 7 2 2 63909 92048
0 34151 5 1 1 93153
0 34152 7 2 2 60612 80157
0 34153 5 1 1 93155
0 34154 7 1 2 34151 34153
0 34155 5 1 1 34154
0 34156 7 1 2 62487 34155
0 34157 5 1 1 34156
0 34158 7 1 2 71829 80158
0 34159 5 1 1 34158
0 34160 7 1 2 34157 34159
0 34161 5 2 1 34160
0 34162 7 1 2 76678 93157
0 34163 5 1 1 34162
0 34164 7 2 2 59608 79860
0 34165 5 1 1 93159
0 34166 7 1 2 93146 93160
0 34167 5 1 1 34166
0 34168 7 1 2 34163 34167
0 34169 5 1 1 34168
0 34170 7 1 2 68109 34169
0 34171 5 1 1 34170
0 34172 7 1 2 69425 78841
0 34173 5 3 1 34172
0 34174 7 1 2 65287 87994
0 34175 5 1 1 34174
0 34176 7 1 2 93161 34175
0 34177 5 2 1 34176
0 34178 7 1 2 76679 93164
0 34179 5 1 1 34178
0 34180 7 1 2 34165 34179
0 34181 5 1 1 34180
0 34182 7 1 2 67207 34181
0 34183 5 1 1 34182
0 34184 7 1 2 34171 34183
0 34185 5 1 1 34184
0 34186 7 1 2 60986 34185
0 34187 5 1 1 34186
0 34188 7 1 2 76680 75032
0 34189 7 1 2 92741 34188
0 34190 5 1 1 34189
0 34191 7 1 2 63060 34190
0 34192 7 1 2 34187 34191
0 34193 5 1 1 34192
0 34194 7 1 2 60012 80774
0 34195 7 1 2 78726 34194
0 34196 7 1 2 34193 34195
0 34197 5 1 1 34196
0 34198 7 2 2 60013 76681
0 34199 7 3 2 62488 92791
0 34200 7 1 2 84641 93168
0 34201 5 1 1 34200
0 34202 7 1 2 80270 91468
0 34203 5 1 1 34202
0 34204 7 1 2 70416 34203
0 34205 5 1 1 34204
0 34206 7 1 2 65624 34205
0 34207 5 1 1 34206
0 34208 7 1 2 34201 34207
0 34209 5 1 1 34208
0 34210 7 1 2 70824 34209
0 34211 5 1 1 34210
0 34212 7 1 2 65625 91495
0 34213 5 1 1 34212
0 34214 7 1 2 91603 34213
0 34215 5 2 1 34214
0 34216 7 1 2 81858 93171
0 34217 5 1 1 34216
0 34218 7 1 2 65626 92409
0 34219 5 1 1 34218
0 34220 7 1 2 74943 84642
0 34221 5 1 1 34220
0 34222 7 1 2 34219 34221
0 34223 5 1 1 34222
0 34224 7 1 2 75904 34223
0 34225 5 1 1 34224
0 34226 7 2 2 67666 77117
0 34227 5 1 1 93173
0 34228 7 1 2 76207 34227
0 34229 5 1 1 34228
0 34230 7 1 2 72268 85364
0 34231 5 1 1 34230
0 34232 7 1 2 70417 34231
0 34233 7 2 2 34229 34232
0 34234 5 1 1 93175
0 34235 7 1 2 72148 34234
0 34236 5 1 1 34235
0 34237 7 1 2 67208 75145
0 34238 5 3 1 34237
0 34239 7 1 2 34236 93177
0 34240 7 1 2 34225 34239
0 34241 7 1 2 34217 34240
0 34242 7 1 2 34211 34241
0 34243 5 1 1 34242
0 34244 7 1 2 93166 34243
0 34245 5 1 1 34244
0 34246 7 2 2 79100 72060
0 34247 5 1 1 93180
0 34248 7 1 2 93137 34247
0 34249 5 1 1 34248
0 34250 7 1 2 57439 34249
0 34251 5 1 1 34250
0 34252 7 1 2 71972 34251
0 34253 5 4 1 34252
0 34254 7 1 2 70418 79827
0 34255 7 1 2 93182 34254
0 34256 5 1 1 34255
0 34257 7 1 2 34245 34256
0 34258 5 1 1 34257
0 34259 7 1 2 64362 34258
0 34260 5 1 1 34259
0 34261 7 1 2 77118 74884
0 34262 7 1 2 78516 34261
0 34263 5 1 1 34262
0 34264 7 1 2 80147 34263
0 34265 5 1 1 34264
0 34266 7 1 2 68009 71042
0 34267 5 2 1 34266
0 34268 7 1 2 70825 93186
0 34269 5 1 1 34268
0 34270 7 1 2 73874 34269
0 34271 7 1 2 34265 34270
0 34272 5 1 1 34271
0 34273 7 1 2 68010 93174
0 34274 5 2 1 34273
0 34275 7 1 2 65288 93188
0 34276 5 1 1 34275
0 34277 7 1 2 60987 80164
0 34278 7 1 2 76823 34277
0 34279 7 1 2 34276 34278
0 34280 5 1 1 34279
0 34281 7 1 2 87174 34280
0 34282 7 1 2 34272 34281
0 34283 5 1 1 34282
0 34284 7 1 2 34260 34283
0 34285 7 1 2 34197 34284
0 34286 5 1 1 34285
0 34287 7 1 2 63508 34286
0 34288 5 1 1 34287
0 34289 7 1 2 58320 83919
0 34290 5 1 1 34289
0 34291 7 1 2 87021 34290
0 34292 5 2 1 34291
0 34293 7 1 2 79037 93190
0 34294 5 1 1 34293
0 34295 7 1 2 82923 92178
0 34296 5 1 1 34295
0 34297 7 1 2 34294 34296
0 34298 5 1 1 34297
0 34299 7 1 2 70323 34298
0 34300 5 1 1 34299
0 34301 7 1 2 74201 33930
0 34302 5 1 1 34301
0 34303 7 1 2 67209 34302
0 34304 5 2 1 34303
0 34305 7 3 2 60613 78145
0 34306 5 1 1 93194
0 34307 7 1 2 77406 90555
0 34308 5 1 1 34307
0 34309 7 1 2 93195 34308
0 34310 5 1 1 34309
0 34311 7 1 2 67762 83199
0 34312 5 2 1 34311
0 34313 7 1 2 70324 77104
0 34314 7 1 2 81233 34313
0 34315 5 2 1 34314
0 34316 7 1 2 78146 84583
0 34317 5 1 1 34316
0 34318 7 1 2 93199 34317
0 34319 7 2 2 93197 34318
0 34320 7 1 2 34310 93201
0 34321 5 1 1 34320
0 34322 7 1 2 63333 34321
0 34323 5 1 1 34322
0 34324 7 1 2 93192 34323
0 34325 5 1 1 34324
0 34326 7 1 2 64573 34325
0 34327 5 1 1 34326
0 34328 7 1 2 68524 86407
0 34329 5 1 1 34328
0 34330 7 1 2 69758 34329
0 34331 5 1 1 34330
0 34332 7 1 2 76682 34331
0 34333 5 1 1 34332
0 34334 7 2 2 70301 77105
0 34335 5 1 1 93203
0 34336 7 1 2 73726 93204
0 34337 5 1 1 34336
0 34338 7 1 2 34333 34337
0 34339 5 1 1 34338
0 34340 7 1 2 63061 34339
0 34341 5 1 1 34340
0 34342 7 2 2 60988 92412
0 34343 7 1 2 64363 80159
0 34344 7 1 2 93205 34343
0 34345 5 1 1 34344
0 34346 7 1 2 78399 34345
0 34347 7 1 2 34341 34346
0 34348 5 1 1 34347
0 34349 7 1 2 67763 34348
0 34350 5 1 1 34349
0 34351 7 2 2 72477 78847
0 34352 5 2 1 93207
0 34353 7 2 2 70325 93209
0 34354 7 1 2 80782 93211
0 34355 5 1 1 34354
0 34356 7 1 2 71297 84243
0 34357 7 1 2 93154 34356
0 34358 5 1 1 34357
0 34359 7 1 2 34355 34358
0 34360 5 1 1 34359
0 34361 7 1 2 76683 34360
0 34362 5 1 1 34361
0 34363 7 2 2 62489 81657
0 34364 5 2 1 93213
0 34365 7 1 2 78531 79984
0 34366 7 1 2 93214 34365
0 34367 5 1 1 34366
0 34368 7 1 2 34362 34367
0 34369 7 1 2 34350 34368
0 34370 5 1 1 34369
0 34371 7 1 2 68110 34370
0 34372 5 1 1 34371
0 34373 7 2 2 75055 93202
0 34374 5 1 1 93217
0 34375 7 1 2 84374 34374
0 34376 5 1 1 34375
0 34377 7 1 2 75146 75058
0 34378 5 3 1 34377
0 34379 7 1 2 34376 93219
0 34380 5 1 1 34379
0 34381 7 1 2 76684 34380
0 34382 5 1 1 34381
0 34383 7 2 2 34372 34382
0 34384 7 1 2 34327 93222
0 34385 5 1 1 34384
0 34386 7 1 2 79432 34385
0 34387 5 1 1 34386
0 34388 7 1 2 34300 34387
0 34389 7 1 2 34288 34388
0 34390 5 1 1 34389
0 34391 7 1 2 61357 34390
0 34392 5 1 1 34391
0 34393 7 2 2 58988 73227
0 34394 7 1 2 87428 93224
0 34395 5 1 1 34394
0 34396 7 1 2 87315 34395
0 34397 5 1 1 34396
0 34398 7 1 2 58321 34397
0 34399 5 1 1 34398
0 34400 7 1 2 85398 69086
0 34401 5 1 1 34400
0 34402 7 1 2 78173 34401
0 34403 5 1 1 34402
0 34404 7 1 2 59850 34403
0 34405 5 1 1 34404
0 34406 7 1 2 34399 34405
0 34407 5 1 1 34406
0 34408 7 1 2 57719 34407
0 34409 5 1 1 34408
0 34410 7 4 2 59851 92878
0 34411 5 1 1 93226
0 34412 7 1 2 74039 93227
0 34413 5 1 1 34412
0 34414 7 1 2 34409 34413
0 34415 5 1 1 34414
0 34416 7 1 2 57440 34415
0 34417 5 1 1 34416
0 34418 7 1 2 79516 93228
0 34419 5 1 1 34418
0 34420 7 1 2 34417 34419
0 34421 5 1 1 34420
0 34422 7 1 2 65289 34421
0 34423 5 1 1 34422
0 34424 7 2 2 65627 78744
0 34425 5 1 1 93230
0 34426 7 1 2 64574 93231
0 34427 5 1 1 34426
0 34428 7 1 2 61358 90611
0 34429 5 1 1 34428
0 34430 7 1 2 34427 34429
0 34431 5 1 1 34430
0 34432 7 1 2 58585 34431
0 34433 5 1 1 34432
0 34434 7 2 2 65628 71113
0 34435 5 1 1 93232
0 34436 7 1 2 93229 93233
0 34437 5 1 1 34436
0 34438 7 1 2 34433 34437
0 34439 7 1 2 34423 34438
0 34440 5 1 1 34439
0 34441 7 1 2 64715 34440
0 34442 5 1 1 34441
0 34443 7 1 2 85114 85983
0 34444 5 1 1 34443
0 34445 7 1 2 34442 34444
0 34446 5 1 1 34445
0 34447 7 1 2 63509 34446
0 34448 5 1 1 34447
0 34449 7 1 2 70302 74655
0 34450 7 1 2 89198 34449
0 34451 5 1 1 34450
0 34452 7 1 2 34448 34451
0 34453 5 1 1 34452
0 34454 7 1 2 67340 34453
0 34455 5 1 1 34454
0 34456 7 1 2 58322 77882
0 34457 5 2 1 34456
0 34458 7 1 2 19292 93234
0 34459 5 1 1 34458
0 34460 7 1 2 70326 34459
0 34461 5 1 1 34460
0 34462 7 2 2 64575 78921
0 34463 5 1 1 93236
0 34464 7 1 2 76685 34463
0 34465 7 1 2 93183 34464
0 34466 5 1 1 34465
0 34467 7 1 2 34461 34466
0 34468 5 1 1 34467
0 34469 7 1 2 82999 34468
0 34470 5 1 1 34469
0 34471 7 1 2 34455 34470
0 34472 7 1 2 34392 34471
0 34473 5 1 1 34472
0 34474 7 1 2 90675 34473
0 34475 5 1 1 34474
0 34476 7 1 2 70213 80051
0 34477 5 1 1 34476
0 34478 7 2 2 73177 34477
0 34479 5 1 1 93238
0 34480 7 1 2 69001 84899
0 34481 5 1 1 34480
0 34482 7 1 2 72100 75905
0 34483 7 1 2 34481 34482
0 34484 5 1 1 34483
0 34485 7 1 2 57720 34484
0 34486 5 1 1 34485
0 34487 7 2 2 34479 34486
0 34488 5 1 1 93240
0 34489 7 1 2 58055 34488
0 34490 5 1 1 34489
0 34491 7 1 2 81096 87085
0 34492 5 1 1 34491
0 34493 7 1 2 81540 34492
0 34494 7 1 2 34490 34493
0 34495 5 1 1 34494
0 34496 7 1 2 80757 34495
0 34497 5 1 1 34496
0 34498 7 1 2 68011 19001
0 34499 5 2 1 34498
0 34500 7 1 2 71434 93242
0 34501 5 1 1 34500
0 34502 7 4 2 71298 85360
0 34503 5 1 1 93244
0 34504 7 1 2 75331 77150
0 34505 5 1 1 34504
0 34506 7 1 2 60614 34505
0 34507 7 1 2 93245 34506
0 34508 5 1 1 34507
0 34509 7 1 2 34501 34508
0 34510 5 2 1 34509
0 34511 7 1 2 74656 72313
0 34512 7 1 2 83666 34511
0 34513 7 1 2 93248 34512
0 34514 5 1 1 34513
0 34515 7 1 2 34497 34514
0 34516 5 1 1 34515
0 34517 7 1 2 59852 34516
0 34518 5 1 1 34517
0 34519 7 3 2 79541 92939
0 34520 7 1 2 76686 93250
0 34521 5 1 1 34520
0 34522 7 1 2 58586 79291
0 34523 5 1 1 34522
0 34524 7 1 2 34521 34523
0 34525 5 1 1 34524
0 34526 7 1 2 85471 34525
0 34527 5 1 1 34526
0 34528 7 2 2 84202 73454
0 34529 5 1 1 93253
0 34530 7 1 2 62490 79542
0 34531 5 1 1 34530
0 34532 7 1 2 34529 34531
0 34533 5 1 1 34532
0 34534 7 2 2 64576 84985
0 34535 5 1 1 93255
0 34536 7 1 2 34533 93256
0 34537 5 1 1 34536
0 34538 7 2 2 67563 77034
0 34539 5 3 1 93257
0 34540 7 1 2 90808 93258
0 34541 5 1 1 34540
0 34542 7 1 2 84346 90790
0 34543 5 1 1 34542
0 34544 7 1 2 34541 34543
0 34545 5 1 1 34544
0 34546 7 5 2 68111 76687
0 34547 5 2 1 93262
0 34548 7 1 2 85425 93263
0 34549 7 1 2 34545 34548
0 34550 5 1 1 34549
0 34551 7 1 2 84884 93251
0 34552 5 1 1 34551
0 34553 7 1 2 34550 34552
0 34554 7 1 2 34537 34553
0 34555 7 1 2 34527 34554
0 34556 5 1 1 34555
0 34557 7 1 2 78864 34556
0 34558 5 1 1 34557
0 34559 7 1 2 70419 92870
0 34560 5 1 1 34559
0 34561 7 1 2 76979 34560
0 34562 5 1 1 34561
0 34563 7 1 2 63062 88420
0 34564 5 2 1 34563
0 34565 7 1 2 63334 93269
0 34566 5 1 1 34565
0 34567 7 1 2 34562 34566
0 34568 5 1 1 34567
0 34569 7 1 2 64577 34568
0 34570 5 1 1 34569
0 34571 7 1 2 65629 92996
0 34572 5 1 1 34571
0 34573 7 1 2 34570 34572
0 34574 5 1 1 34573
0 34575 7 1 2 85209 34574
0 34576 5 1 1 34575
0 34577 7 1 2 84986 93254
0 34578 5 1 1 34577
0 34579 7 5 2 63335 68112
0 34580 5 1 1 93271
0 34581 7 1 2 87751 93272
0 34582 5 1 1 34581
0 34583 7 1 2 34578 34582
0 34584 5 1 1 34583
0 34585 7 1 2 64578 34584
0 34586 5 1 1 34585
0 34587 7 1 2 87759 89978
0 34588 5 1 1 34587
0 34589 7 2 2 63063 70327
0 34590 5 1 1 93276
0 34591 7 2 2 70826 83950
0 34592 5 1 1 93278
0 34593 7 1 2 93277 93279
0 34594 5 1 1 34593
0 34595 7 1 2 69925 78784
0 34596 5 1 1 34595
0 34597 7 1 2 34594 34596
0 34598 5 1 1 34597
0 34599 7 1 2 85210 34598
0 34600 5 1 1 34599
0 34601 7 1 2 34588 34600
0 34602 7 1 2 34586 34601
0 34603 5 1 1 34602
0 34604 7 1 2 62491 34603
0 34605 5 1 1 34604
0 34606 7 2 2 60989 87116
0 34607 7 1 2 58587 33538
0 34608 5 1 1 34607
0 34609 7 1 2 93280 34608
0 34610 5 1 1 34609
0 34611 7 1 2 80824 34610
0 34612 5 1 1 34611
0 34613 7 1 2 59609 34612
0 34614 5 1 1 34613
0 34615 7 1 2 74192 92768
0 34616 5 1 1 34615
0 34617 7 1 2 34614 34616
0 34618 5 1 1 34617
0 34619 7 1 2 64579 34618
0 34620 5 1 1 34619
0 34621 7 1 2 34605 34620
0 34622 7 1 2 34576 34621
0 34623 7 1 2 34558 34622
0 34624 5 1 1 34623
0 34625 7 1 2 61359 74307
0 34626 7 1 2 34624 34625
0 34627 5 1 1 34626
0 34628 7 1 2 34518 34627
0 34629 5 1 1 34628
0 34630 7 1 2 66494 34629
0 34631 5 1 1 34630
0 34632 7 1 2 67210 85033
0 34633 5 1 1 34632
0 34634 7 1 2 34335 34633
0 34635 5 1 1 34634
0 34636 7 1 2 67879 34635
0 34637 5 1 1 34636
0 34638 7 3 2 85570 78624
0 34639 7 1 2 79085 93282
0 34640 5 1 1 34639
0 34641 7 2 2 73128 84414
0 34642 5 4 1 93285
0 34643 7 1 2 34640 93287
0 34644 7 1 2 34637 34643
0 34645 5 1 1 34644
0 34646 7 1 2 80790 34645
0 34647 5 1 1 34646
0 34648 7 1 2 71742 84338
0 34649 5 1 1 34648
0 34650 7 1 2 80924 34649
0 34651 5 1 1 34650
0 34652 7 1 2 91861 34651
0 34653 5 2 1 34652
0 34654 7 1 2 83951 93291
0 34655 5 1 1 34654
0 34656 7 1 2 90985 34655
0 34657 7 1 2 93057 34656
0 34658 5 1 1 34657
0 34659 7 1 2 80979 34658
0 34660 5 1 1 34659
0 34661 7 2 2 34647 34660
0 34662 5 1 1 93293
0 34663 7 2 2 66712 34662
0 34664 7 1 2 92510 93295
0 34665 5 1 1 34664
0 34666 7 1 2 57721 81600
0 34667 5 2 1 34666
0 34668 7 2 2 81799 93297
0 34669 5 2 1 93299
0 34670 7 1 2 72492 87587
0 34671 7 1 2 72623 34670
0 34672 7 1 2 93300 34671
0 34673 5 1 1 34672
0 34674 7 6 2 71184 76651
0 34675 5 2 1 93303
0 34676 7 1 2 62111 88674
0 34677 7 1 2 93304 34676
0 34678 7 1 2 34673 34677
0 34679 5 1 1 34678
0 34680 7 1 2 34665 34679
0 34681 5 1 1 34680
0 34682 7 1 2 58759 34681
0 34683 5 1 1 34682
0 34684 7 2 2 71656 79512
0 34685 7 1 2 79194 93311
0 34686 5 1 1 34685
0 34687 7 1 2 67341 83574
0 34688 5 2 1 34687
0 34689 7 1 2 71299 93313
0 34690 5 1 1 34689
0 34691 7 1 2 12904 79393
0 34692 5 1 1 34691
0 34693 7 1 2 34690 34692
0 34694 5 1 1 34693
0 34695 7 1 2 67764 34694
0 34696 5 1 1 34695
0 34697 7 1 2 68113 92707
0 34698 5 1 1 34697
0 34699 7 1 2 67211 78762
0 34700 5 1 1 34699
0 34701 7 3 2 60990 68433
0 34702 5 3 1 93315
0 34703 7 1 2 34700 93318
0 34704 7 1 2 34698 34703
0 34705 5 1 1 34704
0 34706 7 1 2 71300 34705
0 34707 5 1 1 34706
0 34708 7 1 2 62758 77759
0 34709 7 1 2 90982 34708
0 34710 5 1 1 34709
0 34711 7 1 2 71435 78763
0 34712 5 2 1 34711
0 34713 7 1 2 34710 93321
0 34714 7 1 2 34707 34713
0 34715 7 1 2 34696 34714
0 34716 5 1 1 34715
0 34717 7 1 2 64580 34716
0 34718 5 1 1 34717
0 34719 7 1 2 34686 34718
0 34720 5 1 1 34719
0 34721 7 1 2 63336 34720
0 34722 5 1 1 34721
0 34723 7 1 2 77167 84415
0 34724 7 1 2 80791 34723
0 34725 5 1 1 34724
0 34726 7 1 2 80981 34725
0 34727 5 1 1 34726
0 34728 7 1 2 88161 34727
0 34729 5 1 1 34728
0 34730 7 1 2 9247 86793
0 34731 5 2 1 34730
0 34732 7 1 2 71505 93323
0 34733 5 2 1 34732
0 34734 7 1 2 75550 93325
0 34735 5 1 1 34734
0 34736 7 1 2 34729 34735
0 34737 5 1 1 34736
0 34738 7 1 2 70214 34737
0 34739 5 1 1 34738
0 34740 7 1 2 62759 83301
0 34741 5 1 1 34740
0 34742 7 1 2 87072 34741
0 34743 5 1 1 34742
0 34744 7 1 2 60615 34743
0 34745 5 2 1 34744
0 34746 7 1 2 67819 77106
0 34747 5 1 1 34746
0 34748 7 1 2 93327 34747
0 34749 5 1 1 34748
0 34750 7 1 2 75575 86443
0 34751 5 1 1 34750
0 34752 7 2 2 76688 34751
0 34753 7 1 2 63064 93329
0 34754 5 1 1 34753
0 34755 7 1 2 64581 91618
0 34756 5 1 1 34755
0 34757 7 1 2 34754 34756
0 34758 5 1 1 34757
0 34759 7 1 2 34749 34758
0 34760 5 1 1 34759
0 34761 7 1 2 85640 93312
0 34762 5 1 1 34761
0 34763 7 1 2 34760 34762
0 34764 7 1 2 34739 34763
0 34765 7 1 2 34722 34764
0 34766 5 1 1 34765
0 34767 7 1 2 88666 34766
0 34768 5 1 1 34767
0 34769 7 1 2 59610 92998
0 34770 5 1 1 34769
0 34771 7 2 2 68385 88778
0 34772 5 1 1 93331
0 34773 7 1 2 60616 74010
0 34774 5 1 1 34773
0 34775 7 3 2 93332 34774
0 34776 7 1 2 63337 93333
0 34777 5 1 1 34776
0 34778 7 1 2 34770 34777
0 34779 5 1 1 34778
0 34780 7 1 2 65630 34779
0 34781 5 1 1 34780
0 34782 7 2 2 58588 83837
0 34783 5 1 1 93336
0 34784 7 1 2 74342 81672
0 34785 5 1 1 34784
0 34786 7 1 2 83952 34785
0 34787 5 1 1 34786
0 34788 7 1 2 92376 34787
0 34789 5 1 1 34788
0 34790 7 1 2 67765 34789
0 34791 5 1 1 34790
0 34792 7 2 2 76329 70121
0 34793 5 4 1 93338
0 34794 7 1 2 84328 93340
0 34795 5 1 1 34794
0 34796 7 1 2 68434 77073
0 34797 5 1 1 34796
0 34798 7 1 2 34795 34797
0 34799 7 1 2 34791 34798
0 34800 5 1 1 34799
0 34801 7 1 2 64364 34800
0 34802 5 1 1 34801
0 34803 7 1 2 86817 34802
0 34804 5 1 1 34803
0 34805 7 1 2 93337 34804
0 34806 5 2 1 34805
0 34807 7 1 2 82473 87522
0 34808 5 1 1 34807
0 34809 7 1 2 76208 81201
0 34810 5 1 1 34809
0 34811 7 1 2 71615 88809
0 34812 5 1 1 34811
0 34813 7 1 2 70420 34812
0 34814 7 1 2 34810 34813
0 34815 5 1 1 34814
0 34816 7 1 2 74542 34815
0 34817 5 2 1 34816
0 34818 7 1 2 34808 93346
0 34819 5 1 1 34818
0 34820 7 1 2 65059 34819
0 34821 5 1 1 34820
0 34822 7 1 2 63338 6526
0 34823 5 1 1 34822
0 34824 7 1 2 68525 88810
0 34825 5 1 1 34824
0 34826 7 1 2 70421 78469
0 34827 7 1 2 34825 34826
0 34828 5 1 1 34827
0 34829 7 1 2 72149 5721
0 34830 7 1 2 34828 34829
0 34831 5 1 1 34830
0 34832 7 1 2 34823 34831
0 34833 5 1 1 34832
0 34834 7 1 2 59611 34833
0 34835 5 1 1 34834
0 34836 7 1 2 79362 69776
0 34837 5 1 1 34836
0 34838 7 1 2 83685 34837
0 34839 5 2 1 34838
0 34840 7 1 2 70422 93348
0 34841 5 1 1 34840
0 34842 7 1 2 59853 34841
0 34843 7 1 2 34835 34842
0 34844 7 1 2 34821 34843
0 34845 7 1 2 93344 34844
0 34846 7 1 2 34781 34845
0 34847 5 1 1 34846
0 34848 7 1 2 82949 93184
0 34849 5 1 1 34848
0 34850 7 1 2 64582 84486
0 34851 7 1 2 34849 34850
0 34852 5 1 1 34851
0 34853 7 1 2 34847 34852
0 34854 5 1 1 34853
0 34855 7 1 2 63339 69426
0 34856 5 2 1 34855
0 34857 7 1 2 74624 75420
0 34858 5 1 1 34857
0 34859 7 1 2 93350 34858
0 34860 5 1 1 34859
0 34861 7 1 2 59854 34860
0 34862 5 1 1 34861
0 34863 7 9 2 64583 82950
0 34864 5 1 1 93352
0 34865 7 1 2 72353 93353
0 34866 5 1 1 34865
0 34867 7 1 2 34862 34866
0 34868 5 1 1 34867
0 34869 7 1 2 59136 34868
0 34870 5 1 1 34869
0 34871 7 1 2 76763 79644
0 34872 5 5 1 34871
0 34873 7 1 2 80094 93361
0 34874 5 1 1 34873
0 34875 7 1 2 34870 34874
0 34876 5 1 1 34875
0 34877 7 1 2 57722 34876
0 34878 5 1 1 34877
0 34879 7 1 2 78931 79380
0 34880 5 1 1 34879
0 34881 7 1 2 78174 34880
0 34882 5 2 1 34881
0 34883 7 1 2 59855 93366
0 34884 5 2 1 34883
0 34885 7 1 2 71896 75202
0 34886 5 2 1 34885
0 34887 7 1 2 73991 93370
0 34888 5 1 1 34887
0 34889 7 1 2 93362 34888
0 34890 5 1 1 34889
0 34891 7 1 2 93368 34890
0 34892 7 1 2 34878 34891
0 34893 5 1 1 34892
0 34894 7 1 2 67342 34893
0 34895 5 1 1 34894
0 34896 7 1 2 65290 79645
0 34897 5 1 1 34896
0 34898 7 1 2 78084 74990
0 34899 5 2 1 34898
0 34900 7 1 2 79421 93372
0 34901 5 2 1 34900
0 34902 7 1 2 68012 93374
0 34903 7 1 2 34897 34902
0 34904 5 1 1 34903
0 34905 7 1 2 93369 34904
0 34906 5 1 1 34905
0 34907 7 1 2 71114 34906
0 34908 5 1 1 34907
0 34909 7 2 2 64584 83648
0 34910 5 1 1 93376
0 34911 7 1 2 76689 34910
0 34912 7 1 2 33815 34911
0 34913 5 1 1 34912
0 34914 7 1 2 64716 34913
0 34915 7 1 2 34908 34914
0 34916 7 1 2 34895 34915
0 34917 7 1 2 34854 34916
0 34918 5 1 1 34917
0 34919 7 1 2 60014 93294
0 34920 5 1 1 34919
0 34921 7 1 2 61861 34920
0 34922 7 1 2 34918 34921
0 34923 5 1 1 34922
0 34924 7 1 2 34768 34923
0 34925 5 1 1 34924
0 34926 7 1 2 79942 34925
0 34927 5 1 1 34926
0 34928 7 1 2 34683 34927
0 34929 5 1 1 34928
0 34930 7 1 2 65972 34929
0 34931 5 1 1 34930
0 34932 7 1 2 34631 34931
0 34933 7 1 2 34475 34932
0 34934 5 1 1 34933
0 34935 7 1 2 66274 34934
0 34936 5 1 1 34935
0 34937 7 1 2 72990 79265
0 34938 7 4 2 58760 65973
0 34939 7 1 2 87815 93378
0 34940 7 1 2 34937 34939
0 34941 7 1 2 86322 34940
0 34942 7 1 2 93125 34941
0 34943 5 1 1 34942
0 34944 7 1 2 34936 34943
0 34945 7 1 2 34149 34944
0 34946 5 1 1 34945
0 34947 7 1 2 60137 34946
0 34948 5 1 1 34947
0 34949 7 1 2 62492 87117
0 34950 5 2 1 34949
0 34951 7 1 2 92761 93382
0 34952 5 3 1 34951
0 34953 7 1 2 78865 93384
0 34954 5 1 1 34953
0 34955 7 2 2 92908 34954
0 34956 7 2 2 67343 93387
0 34957 5 1 1 93389
0 34958 7 1 2 58589 34957
0 34959 5 2 1 34958
0 34960 7 1 2 57723 81797
0 34961 5 1 1 34960
0 34962 7 1 2 63065 34961
0 34963 5 1 1 34962
0 34964 7 1 2 83920 34963
0 34965 5 1 1 34964
0 34966 7 1 2 93391 34965
0 34967 5 1 1 34966
0 34968 7 1 2 61360 34967
0 34969 5 1 1 34968
0 34970 7 1 2 69890 91392
0 34971 5 1 1 34970
0 34972 7 1 2 68114 83085
0 34973 7 1 2 73824 8626
0 34974 7 2 2 34972 34973
0 34975 5 1 1 93393
0 34976 7 1 2 34971 34975
0 34977 5 1 1 34976
0 34978 7 1 2 63066 34977
0 34979 5 1 1 34978
0 34980 7 3 2 68247 76209
0 34981 5 1 1 93395
0 34982 7 2 2 70423 34981
0 34983 5 2 1 93398
0 34984 7 2 2 60617 93400
0 34985 5 1 1 93402
0 34986 7 1 2 83310 77151
0 34987 5 1 1 34986
0 34988 7 1 2 93403 34987
0 34989 5 1 1 34988
0 34990 7 1 2 34979 34989
0 34991 5 1 1 34990
0 34992 7 1 2 73668 34991
0 34993 5 1 1 34992
0 34994 7 2 2 71185 85935
0 34995 7 1 2 75715 93404
0 34996 5 3 1 34995
0 34997 7 1 2 71506 93406
0 34998 5 1 1 34997
0 34999 7 1 2 60397 67894
0 35000 5 1 1 34999
0 35001 7 1 2 83501 35000
0 35002 7 2 2 34998 35001
0 35003 5 1 1 93409
0 35004 7 1 2 65974 35003
0 35005 5 1 1 35004
0 35006 7 1 2 59612 85852
0 35007 5 1 1 35006
0 35008 7 1 2 35005 35007
0 35009 5 1 1 35008
0 35010 7 1 2 63340 35009
0 35011 5 1 1 35010
0 35012 7 1 2 34993 35011
0 35013 7 1 2 34969 35012
0 35014 5 1 1 35013
0 35015 7 1 2 66275 35014
0 35016 5 1 1 35015
0 35017 7 2 2 58590 86488
0 35018 5 4 1 93411
0 35019 7 1 2 69453 93412
0 35020 5 3 1 35019
0 35021 7 1 2 69454 80477
0 35022 5 3 1 35021
0 35023 7 1 2 69455 73053
0 35024 5 3 1 35023
0 35025 7 1 2 69827 80507
0 35026 5 1 1 35025
0 35027 7 1 2 75233 35026
0 35028 5 3 1 35027
0 35029 7 1 2 65975 93426
0 35030 5 1 1 35029
0 35031 7 1 2 93423 35030
0 35032 5 1 1 35031
0 35033 7 1 2 63341 35032
0 35034 5 1 1 35033
0 35035 7 1 2 93420 35034
0 35036 5 1 1 35035
0 35037 7 1 2 66276 35036
0 35038 5 1 1 35037
0 35039 7 1 2 93417 35038
0 35040 5 1 1 35039
0 35041 7 1 2 75332 35040
0 35042 5 1 1 35041
0 35043 7 1 2 83041 35042
0 35044 7 1 2 35016 35043
0 35045 5 1 1 35044
0 35046 7 1 2 65631 35045
0 35047 5 1 1 35046
0 35048 7 1 2 63342 16841
0 35049 5 1 1 35048
0 35050 7 2 2 64365 85853
0 35051 5 4 1 93429
0 35052 7 1 2 35049 93431
0 35053 5 1 1 35052
0 35054 7 1 2 66277 35053
0 35055 5 1 1 35054
0 35056 7 1 2 93413 35055
0 35057 5 1 1 35056
0 35058 7 1 2 93077 35057
0 35059 5 1 1 35058
0 35060 7 1 2 68115 82908
0 35061 5 2 1 35060
0 35062 7 2 2 85907 93435
0 35063 5 2 1 93437
0 35064 7 1 2 75455 93439
0 35065 5 3 1 35064
0 35066 7 1 2 84668 93441
0 35067 5 1 1 35066
0 35068 7 1 2 83042 35067
0 35069 7 1 2 35059 35068
0 35070 5 2 1 35069
0 35071 7 1 2 68386 93444
0 35072 5 1 1 35071
0 35073 7 1 2 85854 89187
0 35074 5 1 1 35073
0 35075 7 2 2 65291 84502
0 35076 5 1 1 93446
0 35077 7 1 2 60991 90334
0 35078 7 1 2 93447 35077
0 35079 5 1 1 35078
0 35080 7 1 2 35074 35079
0 35081 5 1 1 35080
0 35082 7 1 2 59613 35081
0 35083 5 1 1 35082
0 35084 7 1 2 80665 93069
0 35085 5 1 1 35084
0 35086 7 1 2 78932 74051
0 35087 7 1 2 79796 35086
0 35088 5 1 1 35087
0 35089 7 1 2 35085 35088
0 35090 7 1 2 35083 35089
0 35091 5 1 1 35090
0 35092 7 1 2 65060 35091
0 35093 5 1 1 35092
0 35094 7 1 2 78906 85999
0 35095 5 1 1 35094
0 35096 7 1 2 61361 93070
0 35097 5 1 1 35096
0 35098 7 1 2 5693 35097
0 35099 5 1 1 35098
0 35100 7 1 2 78164 35099
0 35101 5 1 1 35100
0 35102 7 1 2 35095 35101
0 35103 7 1 2 35093 35102
0 35104 5 1 1 35103
0 35105 7 1 2 66278 35104
0 35106 5 1 1 35105
0 35107 7 1 2 35072 35106
0 35108 7 1 2 35047 35107
0 35109 7 1 2 60992 93243
0 35110 5 1 1 35109
0 35111 7 1 2 58323 35110
0 35112 5 1 1 35111
0 35113 7 1 2 84669 35112
0 35114 5 1 1 35113
0 35115 7 1 2 81432 92862
0 35116 5 1 1 35115
0 35117 7 1 2 35114 35116
0 35118 5 1 1 35117
0 35119 7 1 2 59614 35118
0 35120 5 1 1 35119
0 35121 7 2 2 58056 70980
0 35122 5 1 1 93448
0 35123 7 1 2 86762 93449
0 35124 5 1 1 35123
0 35125 7 1 2 60993 35124
0 35126 5 1 1 35125
0 35127 7 1 2 88165 92858
0 35128 5 1 1 35127
0 35129 7 1 2 68116 35128
0 35130 5 1 1 35129
0 35131 7 2 2 76210 74229
0 35132 5 1 1 93450
0 35133 7 2 2 90336 35132
0 35134 5 1 1 93452
0 35135 7 1 2 80235 92753
0 35136 7 1 2 93453 35135
0 35137 7 1 2 35130 35136
0 35138 7 1 2 35126 35137
0 35139 5 1 1 35138
0 35140 7 1 2 88071 35139
0 35141 5 1 1 35140
0 35142 7 1 2 74697 35141
0 35143 5 1 1 35142
0 35144 7 1 2 64366 35143
0 35145 5 1 1 35144
0 35146 7 1 2 60618 72512
0 35147 5 1 1 35146
0 35148 7 1 2 85695 70445
0 35149 5 1 1 35148
0 35150 7 1 2 65976 35149
0 35151 7 1 2 35147 35150
0 35152 5 1 1 35151
0 35153 7 1 2 61362 84253
0 35154 5 1 1 35153
0 35155 7 1 2 79115 35154
0 35156 7 1 2 35152 35155
0 35157 5 1 1 35156
0 35158 7 1 2 35145 35157
0 35159 7 1 2 60994 72339
0 35160 5 1 1 35159
0 35161 7 1 2 59615 35160
0 35162 5 2 1 35161
0 35163 7 1 2 93041 93454
0 35164 5 1 1 35163
0 35165 7 1 2 82474 84552
0 35166 5 1 1 35165
0 35167 7 1 2 92802 35166
0 35168 5 1 1 35167
0 35169 7 1 2 35164 35168
0 35170 5 1 1 35169
0 35171 7 1 2 65977 35170
0 35172 5 2 1 35171
0 35173 7 1 2 79525 92545
0 35174 5 1 1 35173
0 35175 7 1 2 93456 35174
0 35176 5 1 1 35175
0 35177 7 1 2 69044 35176
0 35178 5 1 1 35177
0 35179 7 2 2 80399 69799
0 35180 5 1 1 93458
0 35181 7 2 2 58324 92754
0 35182 5 3 1 93460
0 35183 7 1 2 62760 93462
0 35184 5 2 1 35183
0 35185 7 1 2 64092 93463
0 35186 5 2 1 35185
0 35187 7 1 2 77497 88779
0 35188 5 1 1 35187
0 35189 7 1 2 89817 35188
0 35190 5 2 1 35189
0 35191 7 1 2 67564 76211
0 35192 5 1 1 35191
0 35193 7 1 2 93469 35192
0 35194 7 1 2 93467 35193
0 35195 7 1 2 93465 35194
0 35196 5 1 1 35195
0 35197 7 1 2 65978 35196
0 35198 5 1 1 35197
0 35199 7 1 2 35180 35198
0 35200 5 1 1 35199
0 35201 7 1 2 60995 35200
0 35202 5 1 1 35201
0 35203 7 1 2 35178 35202
0 35204 7 1 2 35158 35203
0 35205 5 1 1 35204
0 35206 7 1 2 66279 35205
0 35207 5 1 1 35206
0 35208 7 1 2 35120 35207
0 35209 5 1 1 35208
0 35210 7 1 2 58591 35209
0 35211 5 1 1 35210
0 35212 7 1 2 65979 76399
0 35213 5 1 1 35212
0 35214 7 1 2 76366 73054
0 35215 5 1 1 35214
0 35216 7 1 2 35213 35215
0 35217 5 1 1 35216
0 35218 7 1 2 63343 35217
0 35219 5 1 1 35218
0 35220 7 1 2 76367 80478
0 35221 5 1 1 35220
0 35222 7 1 2 35219 35221
0 35223 5 1 1 35222
0 35224 7 1 2 66280 35223
0 35225 5 1 1 35224
0 35226 7 1 2 76368 86946
0 35227 5 1 1 35226
0 35228 7 1 2 35225 35227
0 35229 5 2 1 35228
0 35230 7 1 2 68387 93471
0 35231 5 1 1 35230
0 35232 7 1 2 76566 87006
0 35233 5 1 1 35232
0 35234 7 1 2 93424 35233
0 35235 5 1 1 35234
0 35236 7 1 2 63344 35235
0 35237 5 1 1 35236
0 35238 7 1 2 93421 35237
0 35239 5 1 1 35238
0 35240 7 1 2 66281 35239
0 35241 5 1 1 35240
0 35242 7 1 2 93418 35241
0 35243 5 1 1 35242
0 35244 7 1 2 67667 35243
0 35245 5 1 1 35244
0 35246 7 1 2 86692 84073
0 35247 5 1 1 35246
0 35248 7 1 2 58592 35247
0 35249 5 1 1 35248
0 35250 7 1 2 82880 74675
0 35251 5 1 1 35250
0 35252 7 1 2 35249 35251
0 35253 7 1 2 35245 35252
0 35254 7 1 2 35231 35253
0 35255 5 1 1 35254
0 35256 7 1 2 67344 35255
0 35257 5 1 1 35256
0 35258 7 1 2 35211 35257
0 35259 7 1 2 35108 35258
0 35260 5 1 1 35259
0 35261 7 1 2 59856 35260
0 35262 5 1 1 35261
0 35263 7 1 2 70111 10693
0 35264 5 1 1 35263
0 35265 7 2 2 67345 35264
0 35266 5 1 1 93473
0 35267 7 1 2 68013 76567
0 35268 5 1 1 35267
0 35269 7 1 2 35266 35268
0 35270 5 1 1 35269
0 35271 7 1 2 57441 35270
0 35272 5 1 1 35271
0 35273 7 1 2 68435 35272
0 35274 5 2 1 35273
0 35275 7 1 2 71186 93475
0 35276 5 1 1 35275
0 35277 7 1 2 57442 93474
0 35278 5 2 1 35277
0 35279 7 1 2 71301 93477
0 35280 5 1 1 35279
0 35281 7 1 2 58593 35280
0 35282 5 1 1 35281
0 35283 7 1 2 60996 35282
0 35284 7 1 2 35276 35283
0 35285 5 1 1 35284
0 35286 7 1 2 85348 76768
0 35287 5 1 1 35286
0 35288 7 1 2 69846 35287
0 35289 5 1 1 35288
0 35290 7 1 2 68117 78417
0 35291 5 1 1 35290
0 35292 7 1 2 67346 74377
0 35293 7 1 2 35291 35292
0 35294 5 1 1 35293
0 35295 7 1 2 85131 93407
0 35296 5 1 1 35295
0 35297 7 1 2 81219 72537
0 35298 5 1 1 35297
0 35299 7 1 2 67347 35298
0 35300 5 1 1 35299
0 35301 7 1 2 74518 79598
0 35302 5 1 1 35301
0 35303 7 2 2 35300 35302
0 35304 5 1 1 93479
0 35305 7 1 2 35296 93480
0 35306 7 1 2 35294 35305
0 35307 7 1 2 35289 35306
0 35308 5 1 1 35307
0 35309 7 1 2 82951 35308
0 35310 5 1 1 35309
0 35311 7 1 2 83137 93442
0 35312 5 1 1 35311
0 35313 7 1 2 9014 35312
0 35314 5 1 1 35313
0 35315 7 1 2 74343 35314
0 35316 5 1 1 35315
0 35317 7 1 2 65632 35316
0 35318 7 1 2 35310 35317
0 35319 5 1 1 35318
0 35320 7 1 2 65980 35319
0 35321 7 1 2 35285 35320
0 35322 5 1 1 35321
0 35323 7 2 2 76436 92774
0 35324 5 1 1 93481
0 35325 7 1 2 63345 35324
0 35326 5 1 1 35325
0 35327 7 1 2 71897 35326
0 35328 5 1 1 35327
0 35329 7 1 2 63346 84914
0 35330 5 1 1 35329
0 35331 7 2 2 58594 82129
0 35332 5 1 1 93483
0 35333 7 1 2 78304 35332
0 35334 5 1 1 35333
0 35335 7 1 2 35330 35334
0 35336 5 1 1 35335
0 35337 7 1 2 35328 35336
0 35338 5 1 1 35337
0 35339 7 1 2 74755 35338
0 35340 5 1 1 35339
0 35341 7 1 2 35322 35340
0 35342 5 2 1 35341
0 35343 7 1 2 82209 93485
0 35344 5 1 1 35343
0 35345 7 1 2 35262 35344
0 35346 5 1 1 35345
0 35347 7 1 2 66495 35346
0 35348 5 1 1 35347
0 35349 7 5 2 86291 90898
0 35350 7 1 2 80052 93298
0 35351 5 3 1 35350
0 35352 7 1 2 65981 93492
0 35353 5 2 1 35352
0 35354 7 1 2 61363 82086
0 35355 5 3 1 35354
0 35356 7 1 2 58057 93497
0 35357 5 1 1 35356
0 35358 7 1 2 93495 35357
0 35359 5 1 1 35358
0 35360 7 1 2 57443 35359
0 35361 5 1 1 35360
0 35362 7 1 2 65982 77702
0 35363 5 1 1 35362
0 35364 7 1 2 35361 35363
0 35365 5 1 1 35364
0 35366 7 1 2 73178 35365
0 35367 5 1 1 35366
0 35368 7 2 2 70927 78564
0 35369 5 1 1 93500
0 35370 7 1 2 87052 35369
0 35371 5 1 1 35370
0 35372 7 1 2 69002 73899
0 35373 5 2 1 35372
0 35374 7 1 2 74874 93502
0 35375 5 1 1 35374
0 35376 7 1 2 57724 35375
0 35377 5 1 1 35376
0 35378 7 1 2 79101 74861
0 35379 5 1 1 35378
0 35380 7 1 2 35377 35379
0 35381 5 1 1 35380
0 35382 7 1 2 57444 35381
0 35383 5 1 1 35382
0 35384 7 1 2 87091 35383
0 35385 5 1 1 35384
0 35386 7 1 2 72934 35385
0 35387 5 1 1 35386
0 35388 7 1 2 35371 35387
0 35389 7 1 2 35367 35388
0 35390 5 1 1 35389
0 35391 7 1 2 93487 35390
0 35392 5 1 1 35391
0 35393 7 1 2 35348 35392
0 35394 5 1 1 35393
0 35395 7 1 2 60015 35394
0 35396 5 1 1 35395
0 35397 7 1 2 65983 93476
0 35398 5 1 1 35397
0 35399 7 1 2 87462 73903
0 35400 5 1 1 35399
0 35401 7 1 2 81062 35400
0 35402 5 1 1 35401
0 35403 7 1 2 78318 35402
0 35404 5 1 1 35403
0 35405 7 1 2 65984 80327
0 35406 5 1 1 35405
0 35407 7 1 2 84926 70942
0 35408 5 1 1 35407
0 35409 7 1 2 65985 35408
0 35410 5 1 1 35409
0 35411 7 1 2 68014 88256
0 35412 5 1 1 35411
0 35413 7 1 2 35410 35412
0 35414 5 1 1 35413
0 35415 7 1 2 71898 35414
0 35416 5 1 1 35415
0 35417 7 1 2 35406 35416
0 35418 7 1 2 35404 35417
0 35419 5 1 1 35418
0 35420 7 1 2 65633 35419
0 35421 5 1 1 35420
0 35422 7 1 2 35398 35421
0 35423 5 2 1 35422
0 35424 7 2 2 86292 89427
0 35425 7 1 2 87533 93506
0 35426 7 1 2 93504 35425
0 35427 5 1 1 35426
0 35428 7 1 2 63510 35427
0 35429 7 1 2 35396 35428
0 35430 5 1 1 35429
0 35431 7 1 2 59857 93472
0 35432 5 1 1 35431
0 35433 7 3 2 86565 93354
0 35434 7 1 2 76400 93508
0 35435 5 1 1 35434
0 35436 7 1 2 35432 35435
0 35437 5 1 1 35436
0 35438 7 1 2 66496 35437
0 35439 5 1 1 35438
0 35440 7 1 2 58595 91990
0 35441 7 1 2 80095 35440
0 35442 5 1 1 35441
0 35443 7 1 2 35439 35442
0 35444 5 1 1 35443
0 35445 7 1 2 67348 35444
0 35446 5 1 1 35445
0 35447 7 1 2 59858 93445
0 35448 5 1 1 35447
0 35449 7 1 2 87463 93438
0 35450 5 1 1 35449
0 35451 7 2 2 78907 73055
0 35452 5 2 1 93511
0 35453 7 1 2 35450 93513
0 35454 5 1 1 35453
0 35455 7 1 2 93078 35454
0 35456 5 1 1 35455
0 35457 7 1 2 83975 87671
0 35458 5 1 1 35457
0 35459 7 1 2 4506 74678
0 35460 5 1 1 35459
0 35461 7 1 2 58596 35460
0 35462 5 1 1 35461
0 35463 7 1 2 35458 35462
0 35464 7 1 2 35456 35463
0 35465 5 1 1 35464
0 35466 7 1 2 82210 35465
0 35467 5 1 1 35466
0 35468 7 1 2 35448 35467
0 35469 5 1 1 35468
0 35470 7 1 2 66497 35469
0 35471 5 1 1 35470
0 35472 7 2 2 65634 85842
0 35473 5 1 1 93515
0 35474 7 1 2 69476 93516
0 35475 5 1 1 35474
0 35476 7 1 2 73808 35475
0 35477 5 1 1 35476
0 35478 7 1 2 35477 93488
0 35479 5 1 1 35478
0 35480 7 1 2 35471 35479
0 35481 7 1 2 35446 35480
0 35482 5 1 1 35481
0 35483 7 1 2 68388 35482
0 35484 5 1 1 35483
0 35485 7 3 2 75851 88166
0 35486 7 1 2 71115 76387
0 35487 7 1 2 93517 35486
0 35488 5 1 1 35487
0 35489 7 1 2 68118 35488
0 35490 5 1 1 35489
0 35491 7 1 2 71691 70827
0 35492 5 1 1 35491
0 35493 7 1 2 76829 35492
0 35494 7 1 2 92747 35493
0 35495 5 1 1 35494
0 35496 7 1 2 60997 35495
0 35497 5 1 1 35496
0 35498 7 1 2 92798 35497
0 35499 7 1 2 35490 35498
0 35500 5 1 1 35499
0 35501 7 1 2 64367 35500
0 35502 5 1 1 35501
0 35503 7 1 2 59616 93461
0 35504 5 2 1 35503
0 35505 7 1 2 82295 93520
0 35506 5 1 1 35505
0 35507 7 1 2 59617 90557
0 35508 5 1 1 35507
0 35509 7 1 2 72340 35508
0 35510 5 1 1 35509
0 35511 7 1 2 90377 35510
0 35512 5 1 1 35511
0 35513 7 1 2 69045 35512
0 35514 5 1 1 35513
0 35515 7 1 2 35506 35514
0 35516 5 1 1 35515
0 35517 7 1 2 68119 35516
0 35518 5 1 1 35517
0 35519 7 1 2 76249 80998
0 35520 5 1 1 35519
0 35521 7 1 2 60998 77046
0 35522 5 1 1 35521
0 35523 7 1 2 35520 35522
0 35524 5 1 1 35523
0 35525 7 1 2 62235 35524
0 35526 5 1 1 35525
0 35527 7 1 2 85476 35526
0 35528 5 1 1 35527
0 35529 7 1 2 69046 35528
0 35530 5 1 1 35529
0 35531 7 3 2 68389 81616
0 35532 5 1 1 93522
0 35533 7 1 2 93518 93523
0 35534 5 1 1 35533
0 35535 7 1 2 80305 35534
0 35536 5 1 1 35535
0 35537 7 1 2 64368 35134
0 35538 5 2 1 35537
0 35539 7 1 2 35536 93525
0 35540 7 1 2 35530 35539
0 35541 7 1 2 35518 35540
0 35542 7 1 2 35502 35541
0 35543 5 1 1 35542
0 35544 7 1 2 58597 35543
0 35545 5 1 1 35544
0 35546 7 1 2 58325 83252
0 35547 7 1 2 90860 35546
0 35548 5 1 1 35547
0 35549 7 1 2 35545 35548
0 35550 5 1 1 35549
0 35551 7 1 2 59859 35550
0 35552 5 1 1 35551
0 35553 7 1 2 80271 75052
0 35554 5 1 1 35553
0 35555 7 1 2 68526 88221
0 35556 5 1 1 35555
0 35557 7 1 2 35554 35556
0 35558 5 1 1 35557
0 35559 7 1 2 90335 35558
0 35560 5 1 1 35559
0 35561 7 2 2 62761 89029
0 35562 5 1 1 93527
0 35563 7 1 2 76080 81194
0 35564 5 1 1 35563
0 35565 7 2 2 62493 89468
0 35566 5 2 1 93529
0 35567 7 1 2 83847 93531
0 35568 7 2 2 35564 35567
0 35569 5 1 1 93533
0 35570 7 1 2 35562 93534
0 35571 5 1 1 35570
0 35572 7 3 2 68120 75147
0 35573 7 1 2 35571 93535
0 35574 5 1 1 35573
0 35575 7 1 2 35560 35574
0 35576 5 2 1 35575
0 35577 7 1 2 59860 93538
0 35578 5 1 1 35577
0 35579 7 1 2 82003 81224
0 35580 5 1 1 35579
0 35581 7 2 2 60999 83269
0 35582 5 2 1 93540
0 35583 7 1 2 58326 82008
0 35584 7 1 2 93542 35583
0 35585 5 1 1 35584
0 35586 7 1 2 35580 35585
0 35587 5 1 1 35586
0 35588 7 1 2 88414 35587
0 35589 5 1 1 35588
0 35590 7 2 2 58327 83357
0 35591 5 3 1 93544
0 35592 7 1 2 65635 93545
0 35593 5 1 1 35592
0 35594 7 1 2 77883 70912
0 35595 7 1 2 35593 35594
0 35596 5 1 1 35595
0 35597 7 1 2 35589 35596
0 35598 7 1 2 35578 35597
0 35599 5 1 1 35598
0 35600 7 1 2 59618 35599
0 35601 5 1 1 35600
0 35602 7 1 2 77232 69877
0 35603 7 1 2 82830 35602
0 35604 5 1 1 35603
0 35605 7 1 2 74378 76758
0 35606 5 1 1 35605
0 35607 7 1 2 35604 35606
0 35608 5 1 1 35607
0 35609 7 1 2 65636 35608
0 35610 5 1 1 35609
0 35611 7 1 2 77804 88222
0 35612 5 1 1 35611
0 35613 7 1 2 35610 35612
0 35614 5 1 1 35613
0 35615 7 1 2 68015 35614
0 35616 5 1 1 35615
0 35617 7 2 2 58598 73546
0 35618 5 1 1 93549
0 35619 7 1 2 78933 93550
0 35620 5 1 1 35619
0 35621 7 1 2 65986 35620
0 35622 7 1 2 35616 35621
0 35623 7 1 2 35601 35622
0 35624 7 1 2 35552 35623
0 35625 5 1 1 35624
0 35626 7 1 2 93440 93392
0 35627 5 1 1 35626
0 35628 7 1 2 65637 35627
0 35629 5 1 1 35628
0 35630 7 1 2 59619 87118
0 35631 5 1 1 35630
0 35632 7 2 2 70112 80272
0 35633 5 3 1 93551
0 35634 7 1 2 79690 93553
0 35635 7 1 2 35631 35634
0 35636 5 1 1 35635
0 35637 7 1 2 61000 84203
0 35638 7 1 2 35636 35637
0 35639 5 1 1 35638
0 35640 7 1 2 87931 92062
0 35641 7 1 2 35639 35640
0 35642 5 1 1 35641
0 35643 7 1 2 58599 35642
0 35644 5 1 1 35643
0 35645 7 1 2 35629 35644
0 35646 5 1 1 35645
0 35647 7 1 2 59861 35646
0 35648 5 1 1 35647
0 35649 7 1 2 59862 85908
0 35650 5 1 1 35649
0 35651 7 1 2 75214 79426
0 35652 5 1 1 35651
0 35653 7 1 2 35650 35652
0 35654 5 1 1 35653
0 35655 7 1 2 68016 35654
0 35656 5 1 1 35655
0 35657 7 1 2 85242 35656
0 35658 5 1 1 35657
0 35659 7 1 2 69456 35658
0 35660 5 1 1 35659
0 35661 7 1 2 80588 79641
0 35662 5 2 1 35661
0 35663 7 1 2 61364 93556
0 35664 7 1 2 35660 35663
0 35665 7 1 2 35648 35664
0 35666 5 1 1 35665
0 35667 7 1 2 66282 35666
0 35668 7 1 2 35625 35667
0 35669 5 1 1 35668
0 35670 7 1 2 62236 87712
0 35671 5 1 1 35670
0 35672 7 2 2 58328 81258
0 35673 5 2 1 93558
0 35674 7 1 2 73836 93559
0 35675 7 1 2 35671 35674
0 35676 5 1 1 35675
0 35677 7 1 2 35669 35676
0 35678 5 1 1 35677
0 35679 7 1 2 66498 35678
0 35680 5 1 1 35679
0 35681 7 2 2 72048 93543
0 35682 7 1 2 65987 93562
0 35683 5 1 1 35682
0 35684 7 1 2 93425 35683
0 35685 5 1 1 35684
0 35686 7 1 2 63347 35685
0 35687 5 1 1 35686
0 35688 7 1 2 93422 35687
0 35689 5 1 1 35688
0 35690 7 1 2 66283 35689
0 35691 5 1 1 35690
0 35692 7 1 2 35691 93419
0 35693 5 1 1 35692
0 35694 7 1 2 59863 35693
0 35695 5 1 1 35694
0 35696 7 1 2 93509 93563
0 35697 5 1 1 35696
0 35698 7 1 2 35695 35697
0 35699 5 1 1 35698
0 35700 7 1 2 67668 35699
0 35701 5 1 1 35700
0 35702 7 1 2 82595 87459
0 35703 5 2 1 35702
0 35704 7 1 2 58600 93564
0 35705 5 1 1 35704
0 35706 7 1 2 61365 91882
0 35707 5 1 1 35706
0 35708 7 1 2 35705 35707
0 35709 5 1 1 35708
0 35710 7 1 2 71187 35709
0 35711 5 1 1 35710
0 35712 7 1 2 75447 91963
0 35713 5 1 1 35712
0 35714 7 1 2 35711 35713
0 35715 7 1 2 35701 35714
0 35716 5 1 1 35715
0 35717 7 1 2 66499 35716
0 35718 5 1 1 35717
0 35719 7 2 2 61366 93080
0 35720 5 4 1 93566
0 35721 7 1 2 57445 93568
0 35722 5 2 1 35721
0 35723 7 1 2 73572 93572
0 35724 5 1 1 35723
0 35725 7 1 2 89936 92017
0 35726 7 1 2 35724 35725
0 35727 5 1 1 35726
0 35728 7 1 2 35718 35727
0 35729 5 1 1 35728
0 35730 7 1 2 67349 35729
0 35731 5 1 1 35730
0 35732 7 1 2 67669 76369
0 35733 5 1 1 35732
0 35734 7 1 2 93567 35733
0 35735 5 1 1 35734
0 35736 7 1 2 57446 35735
0 35737 5 1 1 35736
0 35738 7 1 2 61367 76281
0 35739 5 5 1 35738
0 35740 7 1 2 65292 93574
0 35741 5 2 1 35740
0 35742 7 1 2 73332 93579
0 35743 7 1 2 35737 35742
0 35744 5 1 1 35743
0 35745 7 1 2 68017 35744
0 35746 5 1 1 35745
0 35747 7 2 2 72392 87464
0 35748 5 1 1 93581
0 35749 7 1 2 72030 93582
0 35750 5 1 1 35749
0 35751 7 1 2 35746 35750
0 35752 5 1 1 35751
0 35753 7 1 2 93489 35752
0 35754 5 1 1 35753
0 35755 7 1 2 64717 35754
0 35756 7 1 2 35731 35755
0 35757 7 1 2 35680 35756
0 35758 7 1 2 35484 35757
0 35759 5 1 1 35758
0 35760 7 2 2 77494 93169
0 35761 5 1 1 93583
0 35762 7 1 2 78470 35761
0 35763 5 1 1 35762
0 35764 7 1 2 81341 35763
0 35765 5 1 1 35764
0 35766 7 1 2 79607 81446
0 35767 5 1 1 35766
0 35768 7 1 2 35765 35767
0 35769 5 1 1 35768
0 35770 7 1 2 61001 35769
0 35771 5 1 1 35770
0 35772 7 2 2 68870 68436
0 35773 5 1 1 93585
0 35774 7 2 2 67876 35773
0 35775 5 1 1 93587
0 35776 7 1 2 81505 35775
0 35777 5 1 1 35776
0 35778 7 1 2 35771 35777
0 35779 5 1 1 35778
0 35780 7 1 2 58601 35779
0 35781 5 1 1 35780
0 35782 7 1 2 58602 93246
0 35783 5 1 1 35782
0 35784 7 1 2 91642 35783
0 35785 5 1 1 35784
0 35786 7 1 2 91461 35785
0 35787 5 1 1 35786
0 35788 7 2 2 82952 76815
0 35789 5 1 1 93589
0 35790 7 1 2 61659 93590
0 35791 5 1 1 35790
0 35792 7 1 2 61002 35791
0 35793 7 1 2 35787 35792
0 35794 5 1 1 35793
0 35795 7 2 2 61660 67766
0 35796 7 1 2 84521 93591
0 35797 5 1 1 35796
0 35798 7 1 2 85157 68437
0 35799 5 1 1 35798
0 35800 7 1 2 68248 78665
0 35801 5 1 1 35800
0 35802 7 1 2 35799 35801
0 35803 5 1 1 35802
0 35804 7 1 2 66284 35803
0 35805 5 1 1 35804
0 35806 7 1 2 35797 35805
0 35807 5 1 1 35806
0 35808 7 1 2 62237 35807
0 35809 5 1 1 35808
0 35810 7 1 2 85158 88116
0 35811 5 1 1 35810
0 35812 7 1 2 81269 35811
0 35813 5 1 1 35812
0 35814 7 1 2 68438 35813
0 35815 5 1 1 35814
0 35816 7 2 2 77472 79211
0 35817 5 1 1 93593
0 35818 7 1 2 90132 93594
0 35819 5 1 1 35818
0 35820 7 1 2 65638 35819
0 35821 7 1 2 35815 35820
0 35822 7 1 2 35809 35821
0 35823 5 1 1 35822
0 35824 7 1 2 60398 35823
0 35825 7 1 2 35794 35824
0 35826 5 1 1 35825
0 35827 7 1 2 68121 90791
0 35828 5 2 1 35827
0 35829 7 1 2 61003 85117
0 35830 5 1 1 35829
0 35831 7 1 2 93595 35830
0 35832 5 1 1 35831
0 35833 7 1 2 76961 35832
0 35834 5 1 1 35833
0 35835 7 1 2 59620 84632
0 35836 5 1 1 35835
0 35837 7 1 2 89941 35836
0 35838 5 1 1 35837
0 35839 7 1 2 63067 35838
0 35840 5 1 1 35839
0 35841 7 1 2 58603 77915
0 35842 5 1 1 35841
0 35843 7 1 2 65639 35842
0 35844 5 1 1 35843
0 35845 7 1 2 35840 35844
0 35846 5 1 1 35845
0 35847 7 1 2 76802 35846
0 35848 5 1 1 35847
0 35849 7 1 2 35834 35848
0 35850 5 1 1 35849
0 35851 7 1 2 66285 35850
0 35852 5 1 1 35851
0 35853 7 1 2 35826 35852
0 35854 7 1 2 35781 35853
0 35855 5 1 1 35854
0 35856 7 1 2 60619 35855
0 35857 5 1 1 35856
0 35858 7 1 2 62238 87995
0 35859 5 1 1 35858
0 35860 7 2 2 83816 35859
0 35861 5 6 1 93597
0 35862 7 1 2 65640 93599
0 35863 5 2 1 35862
0 35864 7 1 2 10264 93605
0 35865 5 1 1 35864
0 35866 7 1 2 61661 35865
0 35867 5 1 1 35866
0 35868 7 1 2 90437 35867
0 35869 5 1 1 35868
0 35870 7 1 2 58604 35869
0 35871 5 1 1 35870
0 35872 7 1 2 77178 90792
0 35873 5 1 1 35872
0 35874 7 1 2 30363 35873
0 35875 5 1 1 35874
0 35876 7 1 2 66286 35875
0 35877 5 1 1 35876
0 35878 7 1 2 35871 35877
0 35879 5 1 1 35878
0 35880 7 1 2 68122 35879
0 35881 5 1 1 35880
0 35882 7 1 2 78764 79805
0 35883 5 2 1 35882
0 35884 7 1 2 63910 93081
0 35885 5 1 1 35884
0 35886 7 1 2 57725 35885
0 35887 7 1 2 93607 35886
0 35888 5 1 1 35887
0 35889 7 1 2 86253 93127
0 35890 7 1 2 35888 35889
0 35891 5 1 1 35890
0 35892 7 1 2 68018 35891
0 35893 5 1 1 35892
0 35894 7 3 2 58989 72478
0 35895 5 2 1 93609
0 35896 7 1 2 65061 83055
0 35897 7 1 2 93610 35896
0 35898 5 1 1 35897
0 35899 7 1 2 61662 35898
0 35900 7 1 2 35893 35899
0 35901 5 1 1 35900
0 35902 7 1 2 80306 88447
0 35903 5 1 1 35902
0 35904 7 1 2 74025 79222
0 35905 5 2 1 35904
0 35906 7 1 2 63348 93614
0 35907 5 1 1 35906
0 35908 7 1 2 66287 93178
0 35909 7 1 2 35907 35908
0 35910 7 1 2 35903 35909
0 35911 5 1 1 35910
0 35912 7 1 2 64369 35911
0 35913 7 1 2 35901 35912
0 35914 5 1 1 35913
0 35915 7 1 2 78508 88632
0 35916 5 1 1 35915
0 35917 7 1 2 82881 35916
0 35918 5 1 1 35917
0 35919 7 1 2 65641 82895
0 35920 5 1 1 35919
0 35921 7 1 2 88448 89565
0 35922 5 1 1 35921
0 35923 7 1 2 35920 35922
0 35924 5 1 1 35923
0 35925 7 1 2 67212 35924
0 35926 5 1 1 35925
0 35927 7 1 2 58329 86880
0 35928 5 2 1 35927
0 35929 7 1 2 93025 93616
0 35930 5 1 1 35929
0 35931 7 2 2 67767 69427
0 35932 7 1 2 70094 93618
0 35933 5 1 1 35932
0 35934 7 1 2 80367 74604
0 35935 7 1 2 35933 35934
0 35936 5 1 1 35935
0 35937 7 1 2 61004 35936
0 35938 5 1 1 35937
0 35939 7 1 2 35930 35938
0 35940 5 1 1 35939
0 35941 7 1 2 81259 35940
0 35942 5 1 1 35941
0 35943 7 1 2 35926 35942
0 35944 7 1 2 35918 35943
0 35945 7 1 2 35914 35944
0 35946 7 1 2 35881 35945
0 35947 7 1 2 35857 35946
0 35948 5 1 1 35947
0 35949 7 1 2 61368 35948
0 35950 5 1 1 35949
0 35951 7 1 2 70424 79384
0 35952 5 1 1 35951
0 35953 7 1 2 76350 78134
0 35954 5 1 1 35953
0 35955 7 1 2 35952 35954
0 35956 5 1 1 35955
0 35957 7 1 2 61663 78165
0 35958 7 1 2 35956 35957
0 35959 5 1 1 35958
0 35960 7 1 2 35950 35959
0 35961 5 1 1 35960
0 35962 7 1 2 66500 35961
0 35963 5 1 1 35962
0 35964 7 1 2 79363 90031
0 35965 5 1 1 35964
0 35966 7 1 2 78745 91248
0 35967 5 1 1 35966
0 35968 7 1 2 35965 35967
0 35969 5 1 1 35968
0 35970 7 1 2 82953 35969
0 35971 5 1 1 35970
0 35972 7 1 2 78781 80100
0 35973 5 1 1 35972
0 35974 7 1 2 61664 92879
0 35975 7 1 2 35973 35974
0 35976 5 1 1 35975
0 35977 7 1 2 64370 86436
0 35978 5 1 1 35977
0 35979 7 1 2 35976 35978
0 35980 5 1 1 35979
0 35981 7 1 2 66501 35980
0 35982 5 1 1 35981
0 35983 7 1 2 35971 35982
0 35984 5 1 1 35983
0 35985 7 1 2 67350 35984
0 35986 5 1 1 35985
0 35987 7 1 2 58605 70328
0 35988 5 2 1 35987
0 35989 7 1 2 68019 93185
0 35990 5 1 1 35989
0 35991 7 1 2 93620 35990
0 35992 5 1 1 35991
0 35993 7 1 2 90192 35992
0 35994 5 1 1 35993
0 35995 7 1 2 35986 35994
0 35996 7 1 2 35963 35995
0 35997 5 1 1 35996
0 35998 7 1 2 64585 35997
0 35999 5 1 1 35998
0 36000 7 1 2 71302 84081
0 36001 5 1 1 36000
0 36002 7 1 2 93087 36001
0 36003 5 1 1 36002
0 36004 7 1 2 63349 36003
0 36005 5 1 1 36004
0 36006 7 3 2 62239 81013
0 36007 7 1 2 90587 93622
0 36008 5 1 1 36007
0 36009 7 1 2 36005 36008
0 36010 5 1 1 36009
0 36011 7 1 2 67768 36010
0 36012 5 1 1 36011
0 36013 7 1 2 77035 91339
0 36014 5 1 1 36013
0 36015 7 1 2 60399 82924
0 36016 5 1 1 36015
0 36017 7 1 2 36014 36016
0 36018 5 1 1 36017
0 36019 7 1 2 68871 36018
0 36020 5 1 1 36019
0 36021 7 1 2 74991 90383
0 36022 5 1 1 36021
0 36023 7 1 2 61005 83931
0 36024 5 1 1 36023
0 36025 7 1 2 30193 36024
0 36026 5 1 1 36025
0 36027 7 1 2 63350 36026
0 36028 5 1 1 36027
0 36029 7 1 2 36022 36028
0 36030 7 1 2 36020 36029
0 36031 5 1 1 36030
0 36032 7 1 2 60620 36031
0 36033 5 1 1 36032
0 36034 7 1 2 85159 86259
0 36035 5 1 1 36034
0 36036 7 1 2 82954 36035
0 36037 5 1 1 36036
0 36038 7 1 2 68249 36037
0 36039 5 1 1 36038
0 36040 7 1 2 87766 36039
0 36041 7 1 2 36033 36040
0 36042 7 1 2 36012 36041
0 36043 5 1 1 36042
0 36044 7 1 2 59864 36043
0 36045 5 1 1 36044
0 36046 7 1 2 86868 91377
0 36047 5 1 1 36046
0 36048 7 1 2 79504 90558
0 36049 5 1 1 36048
0 36050 7 1 2 60621 36049
0 36051 5 1 1 36050
0 36052 7 1 2 68624 79505
0 36053 5 1 1 36052
0 36054 7 1 2 67769 36053
0 36055 7 1 2 83838 36054
0 36056 5 1 1 36055
0 36057 7 1 2 36051 36056
0 36058 5 1 1 36057
0 36059 7 1 2 68872 36058
0 36060 5 1 1 36059
0 36061 7 1 2 70913 36060
0 36062 5 1 1 36061
0 36063 7 1 2 77824 36062
0 36064 5 1 1 36063
0 36065 7 1 2 36047 36064
0 36066 7 1 2 36045 36065
0 36067 5 1 1 36066
0 36068 7 1 2 68123 36067
0 36069 5 1 1 36068
0 36070 7 2 2 72269 78651
0 36071 5 2 1 93625
0 36072 7 1 2 59621 93627
0 36073 5 2 1 36072
0 36074 7 1 2 77805 93629
0 36075 5 1 1 36074
0 36076 7 1 2 77806 93600
0 36077 5 1 1 36076
0 36078 7 1 2 85316 78097
0 36079 7 1 2 86342 36078
0 36080 5 1 1 36079
0 36081 7 1 2 76759 79608
0 36082 5 1 1 36081
0 36083 7 1 2 24121 36082
0 36084 5 1 1 36083
0 36085 7 1 2 60622 36084
0 36086 5 1 1 36085
0 36087 7 1 2 36080 36086
0 36088 7 1 2 36077 36087
0 36089 5 1 1 36088
0 36090 7 1 2 61006 36089
0 36091 5 1 1 36090
0 36092 7 1 2 36075 36091
0 36093 5 1 1 36092
0 36094 7 1 2 76212 36093
0 36095 5 1 1 36094
0 36096 7 1 2 70949 77825
0 36097 7 1 2 78866 36096
0 36098 5 1 1 36097
0 36099 7 1 2 79065 93334
0 36100 5 1 1 36099
0 36101 7 1 2 61007 36100
0 36102 5 1 1 36101
0 36103 7 1 2 65642 71940
0 36104 5 1 1 36103
0 36105 7 2 2 76250 36104
0 36106 7 1 2 69047 93631
0 36107 5 1 1 36106
0 36108 7 1 2 92799 36107
0 36109 7 1 2 36102 36108
0 36110 5 1 1 36109
0 36111 7 1 2 59865 84987
0 36112 7 1 2 36110 36111
0 36113 5 1 1 36112
0 36114 7 1 2 36098 36113
0 36115 5 1 1 36114
0 36116 7 1 2 64371 36115
0 36117 5 1 1 36116
0 36118 7 1 2 90090 36117
0 36119 7 1 2 36095 36118
0 36120 7 1 2 36069 36119
0 36121 5 1 1 36120
0 36122 7 1 2 66502 36121
0 36123 5 1 1 36122
0 36124 7 1 2 62494 92994
0 36125 5 1 1 36124
0 36126 7 1 2 70828 70372
0 36127 5 1 1 36126
0 36128 7 1 2 36125 36127
0 36129 5 2 1 36128
0 36130 7 1 2 73727 92553
0 36131 7 1 2 93633 36130
0 36132 5 1 1 36131
0 36133 7 1 2 86854 89892
0 36134 5 1 1 36133
0 36135 7 2 2 63351 74344
0 36136 5 1 1 93635
0 36137 7 1 2 66503 92305
0 36138 7 1 2 93636 36137
0 36139 5 1 1 36138
0 36140 7 2 2 58606 69457
0 36141 7 1 2 89236 93637
0 36142 5 1 1 36141
0 36143 7 1 2 36139 36142
0 36144 5 2 1 36143
0 36145 7 1 2 68390 93639
0 36146 5 1 1 36145
0 36147 7 1 2 36134 36146
0 36148 7 1 2 36132 36147
0 36149 5 1 1 36148
0 36150 7 1 2 65643 36149
0 36151 5 1 1 36150
0 36152 7 1 2 73861 72403
0 36153 5 1 1 36152
0 36154 7 1 2 89095 36153
0 36155 5 1 1 36154
0 36156 7 1 2 58990 89242
0 36157 5 1 1 36156
0 36158 7 1 2 36155 36157
0 36159 5 1 1 36158
0 36160 7 1 2 65062 36159
0 36161 5 1 1 36160
0 36162 7 1 2 71899 89062
0 36163 5 2 1 36162
0 36164 7 1 2 36161 93641
0 36165 5 1 1 36164
0 36166 7 1 2 57726 36165
0 36167 5 1 1 36166
0 36168 7 1 2 59137 93640
0 36169 5 1 1 36168
0 36170 7 1 2 36167 36169
0 36171 5 1 1 36170
0 36172 7 1 2 67351 36171
0 36173 5 1 1 36172
0 36174 7 1 2 61665 36173
0 36175 7 1 2 36151 36174
0 36176 7 1 2 36123 36175
0 36177 5 1 1 36176
0 36178 7 1 2 60623 86348
0 36179 5 1 1 36178
0 36180 7 3 2 62240 61008
0 36181 5 2 1 93643
0 36182 7 1 2 90165 93646
0 36183 5 1 1 36182
0 36184 7 1 2 63784 36183
0 36185 5 1 1 36184
0 36186 7 1 2 74944 69891
0 36187 5 1 1 36186
0 36188 7 1 2 58058 68207
0 36189 5 1 1 36188
0 36190 7 1 2 64093 36189
0 36191 5 1 1 36190
0 36192 7 1 2 36187 36191
0 36193 7 1 2 36185 36192
0 36194 7 1 2 36179 36193
0 36195 5 1 1 36194
0 36196 7 1 2 62495 36195
0 36197 5 1 1 36196
0 36198 7 1 2 70028 70122
0 36199 5 1 1 36198
0 36200 7 1 2 61009 36199
0 36201 5 1 1 36200
0 36202 7 1 2 72246 76391
0 36203 7 1 2 59375 69795
0 36204 5 2 1 36203
0 36205 7 1 2 62241 93648
0 36206 5 1 1 36205
0 36207 7 1 2 81624 36206
0 36208 7 1 2 36202 36207
0 36209 5 1 1 36208
0 36210 7 1 2 62762 36209
0 36211 5 1 1 36210
0 36212 7 1 2 36201 36211
0 36213 7 1 2 36197 36212
0 36214 5 1 1 36213
0 36215 7 1 2 71303 36214
0 36216 5 1 1 36215
0 36217 7 1 2 73900 19112
0 36218 5 2 1 36217
0 36219 7 1 2 62496 93650
0 36220 5 1 1 36219
0 36221 7 1 2 73891 87123
0 36222 5 1 1 36221
0 36223 7 1 2 36220 36222
0 36224 5 1 1 36223
0 36225 7 2 2 73129 36224
0 36226 5 1 1 93652
0 36227 7 1 2 73406 80228
0 36228 5 2 1 36227
0 36229 7 1 2 71436 93654
0 36230 5 1 1 36229
0 36231 7 1 2 36226 36230
0 36232 7 1 2 36216 36231
0 36233 5 1 1 36232
0 36234 7 1 2 63352 36233
0 36235 5 1 1 36234
0 36236 7 3 2 62242 85160
0 36237 5 3 1 93656
0 36238 7 1 2 74715 93657
0 36239 5 1 1 36238
0 36240 7 1 2 63353 84273
0 36241 5 1 1 36240
0 36242 7 1 2 36239 36241
0 36243 5 1 1 36242
0 36244 7 1 2 62763 36243
0 36245 5 1 1 36244
0 36246 7 1 2 72341 91620
0 36247 5 1 1 36246
0 36248 7 1 2 64094 82925
0 36249 5 1 1 36248
0 36250 7 1 2 36247 36249
0 36251 7 1 2 36245 36250
0 36252 5 1 1 36251
0 36253 7 1 2 77676 36252
0 36254 5 1 1 36253
0 36255 7 1 2 6328 36254
0 36256 5 1 1 36255
0 36257 7 1 2 69048 36256
0 36258 5 1 1 36257
0 36259 7 1 2 63354 93326
0 36260 5 1 1 36259
0 36261 7 1 2 82926 83302
0 36262 5 1 1 36261
0 36263 7 1 2 80273 77473
0 36264 7 1 2 92422 36263
0 36265 5 1 1 36264
0 36266 7 1 2 36262 36265
0 36267 5 1 1 36266
0 36268 7 1 2 60624 36267
0 36269 5 1 1 36268
0 36270 7 1 2 36260 36269
0 36271 5 1 1 36270
0 36272 7 1 2 70215 36271
0 36273 5 1 1 36272
0 36274 7 1 2 71437 93653
0 36275 5 1 1 36274
0 36276 7 1 2 66504 36275
0 36277 7 1 2 36273 36276
0 36278 7 1 2 36258 36277
0 36279 7 1 2 36235 36278
0 36280 5 1 1 36279
0 36281 7 1 2 68020 5758
0 36282 5 1 1 36281
0 36283 7 1 2 63355 36282
0 36284 5 1 1 36283
0 36285 7 1 2 71188 36284
0 36286 5 1 1 36285
0 36287 7 1 2 73884 69485
0 36288 5 1 1 36287
0 36289 7 1 2 78623 36288
0 36290 5 1 1 36289
0 36291 7 1 2 73818 72362
0 36292 5 1 1 36291
0 36293 7 1 2 79628 36292
0 36294 7 1 2 36290 36293
0 36295 7 1 2 36286 36294
0 36296 5 1 1 36295
0 36297 7 1 2 82955 36296
0 36298 5 1 1 36297
0 36299 7 1 2 61862 36298
0 36300 5 1 1 36299
0 36301 7 1 2 64586 36300
0 36302 7 1 2 36280 36301
0 36303 5 1 1 36302
0 36304 7 1 2 87422 34783
0 36305 5 1 1 36304
0 36306 7 1 2 68873 36305
0 36307 5 2 1 36306
0 36308 7 1 2 60400 90990
0 36309 5 1 1 36308
0 36310 7 1 2 93662 36309
0 36311 5 1 1 36310
0 36312 7 1 2 67770 36311
0 36313 5 1 1 36312
0 36314 7 1 2 72150 78505
0 36315 5 1 1 36314
0 36316 7 1 2 79086 90991
0 36317 5 1 1 36316
0 36318 7 1 2 36315 36317
0 36319 7 1 2 36313 36318
0 36320 5 1 1 36319
0 36321 7 1 2 68124 36320
0 36322 5 1 1 36321
0 36323 7 1 2 74549 72806
0 36324 7 1 2 85696 36323
0 36325 7 1 2 93060 36324
0 36326 5 1 1 36325
0 36327 7 1 2 63068 85233
0 36328 5 1 1 36327
0 36329 7 1 2 63356 36328
0 36330 5 1 1 36329
0 36331 7 1 2 93347 36330
0 36332 5 1 1 36331
0 36333 7 1 2 65063 36332
0 36334 5 1 1 36333
0 36335 7 4 2 58059 72286
0 36336 5 1 1 93664
0 36337 7 1 2 83584 93665
0 36338 5 1 1 36337
0 36339 7 1 2 73980 79800
0 36340 5 1 1 36339
0 36341 7 1 2 36338 36340
0 36342 5 1 1 36341
0 36343 7 1 2 68391 36342
0 36344 5 1 1 36343
0 36345 7 1 2 73981 93053
0 36346 5 1 1 36345
0 36347 7 1 2 83441 90588
0 36348 5 1 1 36347
0 36349 7 1 2 36346 36348
0 36350 5 1 1 36349
0 36351 7 1 2 67352 36350
0 36352 5 1 1 36351
0 36353 7 1 2 93367 35817
0 36354 5 1 1 36353
0 36355 7 1 2 68021 93349
0 36356 5 1 1 36355
0 36357 7 1 2 36354 36356
0 36358 7 1 2 36352 36357
0 36359 7 1 2 36344 36358
0 36360 7 1 2 36334 36359
0 36361 7 1 2 36326 36360
0 36362 7 1 2 36322 36361
0 36363 5 1 1 36362
0 36364 7 1 2 89237 36363
0 36365 5 1 1 36364
0 36366 7 1 2 57727 84900
0 36367 5 1 1 36366
0 36368 7 1 2 77961 87756
0 36369 5 1 1 36368
0 36370 7 3 2 36367 36369
0 36371 5 1 1 93668
0 36372 7 1 2 62764 93669
0 36373 5 1 1 36372
0 36374 7 1 2 68250 81678
0 36375 5 2 1 36374
0 36376 7 1 2 36373 93671
0 36377 5 2 1 36376
0 36378 7 1 2 78867 93673
0 36379 5 1 1 36378
0 36380 7 1 2 84106 36379
0 36381 5 3 1 36380
0 36382 7 1 2 92696 93675
0 36383 5 1 1 36382
0 36384 7 1 2 66288 36383
0 36385 7 1 2 36365 36384
0 36386 7 1 2 36303 36385
0 36387 5 1 1 36386
0 36388 7 1 2 36177 36387
0 36389 5 1 1 36388
0 36390 7 1 2 76962 93039
0 36391 5 1 1 36390
0 36392 7 1 2 60625 84531
0 36393 5 1 1 36392
0 36394 7 1 2 77014 16921
0 36395 5 2 1 36394
0 36396 7 1 2 88811 93678
0 36397 5 1 1 36396
0 36398 7 1 2 36393 36397
0 36399 7 1 2 36391 36398
0 36400 5 1 1 36399
0 36401 7 1 2 60401 36400
0 36402 5 1 1 36401
0 36403 7 1 2 75448 88629
0 36404 5 1 1 36403
0 36405 7 1 2 36402 36404
0 36406 5 1 1 36405
0 36407 7 1 2 61010 36406
0 36408 5 1 1 36407
0 36409 7 2 2 11317 93075
0 36410 7 1 2 82927 93680
0 36411 5 1 1 36410
0 36412 7 1 2 75894 17450
0 36413 5 1 1 36412
0 36414 7 1 2 77991 36413
0 36415 5 1 1 36414
0 36416 7 1 2 84192 69926
0 36417 5 2 1 36416
0 36418 7 1 2 58607 93682
0 36419 7 1 2 36415 36418
0 36420 5 1 1 36419
0 36421 7 1 2 36411 36420
0 36422 5 1 1 36421
0 36423 7 1 2 80209 75456
0 36424 5 1 1 36423
0 36425 7 1 2 63069 36424
0 36426 5 1 1 36425
0 36427 7 1 2 68125 79685
0 36428 5 1 1 36427
0 36429 7 1 2 84546 36428
0 36430 7 1 2 36426 36429
0 36431 5 1 1 36430
0 36432 7 1 2 90992 36431
0 36433 5 1 1 36432
0 36434 7 1 2 36422 36433
0 36435 7 1 2 36408 36434
0 36436 5 1 1 36435
0 36437 7 1 2 89750 36436
0 36438 5 1 1 36437
0 36439 7 1 2 79364 83280
0 36440 5 1 1 36439
0 36441 7 1 2 83686 36440
0 36442 5 1 1 36441
0 36443 7 1 2 78814 36442
0 36444 5 1 1 36443
0 36445 7 1 2 79365 70443
0 36446 5 1 1 36445
0 36447 7 1 2 78175 36446
0 36448 5 1 1 36447
0 36449 7 1 2 57447 36448
0 36450 5 1 1 36449
0 36451 7 1 2 36444 36450
0 36452 5 1 1 36451
0 36453 7 1 2 89747 32466
0 36454 5 1 1 36453
0 36455 7 1 2 36452 36454
0 36456 5 1 1 36455
0 36457 7 1 2 65988 36456
0 36458 7 1 2 36438 36457
0 36459 7 1 2 36389 36458
0 36460 5 1 1 36459
0 36461 7 1 2 6940 90363
0 36462 5 2 1 36461
0 36463 7 1 2 60626 93684
0 36464 5 1 1 36463
0 36465 7 1 2 65064 93592
0 36466 5 1 1 36465
0 36467 7 1 2 36464 36466
0 36468 5 1 1 36467
0 36469 7 1 2 68874 36468
0 36470 5 1 1 36469
0 36471 7 1 2 65065 81087
0 36472 5 2 1 36471
0 36473 7 1 2 86357 93686
0 36474 5 1 1 36473
0 36475 7 1 2 61666 36474
0 36476 5 1 1 36475
0 36477 7 1 2 69857 82888
0 36478 5 1 1 36477
0 36479 7 1 2 76963 87241
0 36480 7 1 2 36478 36479
0 36481 5 1 1 36480
0 36482 7 1 2 36476 36481
0 36483 7 1 2 36470 36482
0 36484 5 1 1 36483
0 36485 7 1 2 61011 36484
0 36486 5 1 1 36485
0 36487 7 1 2 81506 93061
0 36488 5 1 1 36487
0 36489 7 1 2 36486 36488
0 36490 5 1 1 36489
0 36491 7 1 2 76213 36490
0 36492 5 1 1 36491
0 36493 7 1 2 61012 93351
0 36494 5 1 1 36493
0 36495 7 1 2 87780 36494
0 36496 5 1 1 36495
0 36497 7 1 2 36492 36496
0 36498 5 1 1 36497
0 36499 7 1 2 64372 36498
0 36500 5 1 1 36499
0 36501 7 1 2 65644 85244
0 36502 5 1 1 36501
0 36503 7 2 2 93198 36502
0 36504 7 1 2 77750 93688
0 36505 5 1 1 36504
0 36506 7 1 2 84724 36505
0 36507 5 1 1 36506
0 36508 7 1 2 33988 36507
0 36509 5 1 1 36508
0 36510 7 1 2 63070 36509
0 36511 5 1 1 36510
0 36512 7 1 2 80368 93687
0 36513 5 1 1 36512
0 36514 7 1 2 61013 36513
0 36515 5 1 1 36514
0 36516 7 1 2 61014 69860
0 36517 5 1 1 36516
0 36518 7 1 2 75036 36517
0 36519 5 1 1 36518
0 36520 7 1 2 63357 36519
0 36521 5 1 1 36520
0 36522 7 2 2 82467 75007
0 36523 7 1 2 68875 93690
0 36524 5 1 1 36523
0 36525 7 1 2 36521 36524
0 36526 7 1 2 36515 36525
0 36527 5 1 1 36526
0 36528 7 1 2 84988 36527
0 36529 5 1 1 36528
0 36530 7 1 2 36511 36529
0 36531 5 1 1 36530
0 36532 7 1 2 61667 36531
0 36533 5 1 1 36532
0 36534 7 1 2 84885 87789
0 36535 7 1 2 83303 36534
0 36536 5 1 1 36535
0 36537 7 1 2 36533 36536
0 36538 7 1 2 36500 36537
0 36539 5 1 1 36538
0 36540 7 1 2 66505 36539
0 36541 5 1 1 36540
0 36542 7 1 2 88638 90809
0 36543 5 1 1 36542
0 36544 7 1 2 68876 93685
0 36545 5 1 1 36544
0 36546 7 1 2 60627 16252
0 36547 7 1 2 36545 36546
0 36548 5 1 1 36547
0 36549 7 1 2 71304 87242
0 36550 7 1 2 85902 36549
0 36551 7 1 2 36548 36550
0 36552 5 1 1 36551
0 36553 7 1 2 36543 36552
0 36554 5 1 1 36553
0 36555 7 1 2 68251 36554
0 36556 5 1 1 36555
0 36557 7 1 2 85161 87305
0 36558 5 1 1 36557
0 36559 7 1 2 87807 36558
0 36560 7 1 2 36556 36559
0 36561 5 1 1 36560
0 36562 7 1 2 61015 36561
0 36563 5 1 1 36562
0 36564 7 1 2 61668 90793
0 36565 7 1 2 78425 36564
0 36566 5 1 1 36565
0 36567 7 1 2 36563 36566
0 36568 5 1 1 36567
0 36569 7 1 2 66506 36568
0 36570 5 1 1 36569
0 36571 7 1 2 91716 93212
0 36572 5 1 1 36571
0 36573 7 1 2 91162 92537
0 36574 5 1 1 36573
0 36575 7 1 2 91253 36574
0 36576 5 1 1 36575
0 36577 7 1 2 58608 36576
0 36578 5 1 1 36577
0 36579 7 1 2 63071 93089
0 36580 5 1 1 36579
0 36581 7 1 2 78765 74193
0 36582 5 1 1 36581
0 36583 7 1 2 36580 36582
0 36584 5 1 1 36583
0 36585 7 1 2 89656 36584
0 36586 5 1 1 36585
0 36587 7 1 2 36578 36586
0 36588 5 1 1 36587
0 36589 7 1 2 67771 36588
0 36590 5 1 1 36589
0 36591 7 1 2 36572 36590
0 36592 7 1 2 36570 36591
0 36593 5 1 1 36592
0 36594 7 1 2 68126 36593
0 36595 5 1 1 36594
0 36596 7 1 2 21819 91764
0 36597 5 1 1 36596
0 36598 7 1 2 75037 91604
0 36599 7 1 2 34590 36598
0 36600 7 1 2 93200 36599
0 36601 5 1 1 36600
0 36602 7 1 2 91717 36601
0 36603 5 1 1 36602
0 36604 7 1 2 70303 86875
0 36605 5 1 1 36604
0 36606 7 1 2 36605 93689
0 36607 7 1 2 36603 36606
0 36608 5 1 1 36607
0 36609 7 1 2 36597 36608
0 36610 5 1 1 36609
0 36611 7 1 2 76290 81534
0 36612 5 1 1 36611
0 36613 7 1 2 57728 36612
0 36614 5 1 1 36613
0 36615 7 1 2 59138 76153
0 36616 5 1 1 36615
0 36617 7 1 2 36614 36616
0 36618 5 1 1 36617
0 36619 7 1 2 57448 36618
0 36620 5 1 1 36619
0 36621 7 1 2 76292 36620
0 36622 5 1 1 36621
0 36623 7 1 2 65293 36622
0 36624 5 1 1 36623
0 36625 7 2 2 64095 76356
0 36626 5 1 1 93692
0 36627 7 1 2 58060 36626
0 36628 5 2 1 36627
0 36629 7 2 2 72393 68923
0 36630 5 1 1 93696
0 36631 7 1 2 93694 36630
0 36632 5 2 1 36631
0 36633 7 1 2 67670 93698
0 36634 5 1 1 36633
0 36635 7 1 2 76308 33745
0 36636 5 1 1 36635
0 36637 7 1 2 70425 36636
0 36638 5 1 1 36637
0 36639 7 1 2 36634 36638
0 36640 5 1 1 36639
0 36641 7 1 2 57449 36640
0 36642 5 1 1 36641
0 36643 7 1 2 59376 83056
0 36644 5 1 1 36643
0 36645 7 1 2 72218 69934
0 36646 5 1 1 36645
0 36647 7 1 2 58061 36646
0 36648 5 1 1 36647
0 36649 7 1 2 36644 36648
0 36650 7 1 2 36642 36649
0 36651 5 1 1 36650
0 36652 7 1 2 65645 36651
0 36653 5 1 1 36652
0 36654 7 1 2 36624 36653
0 36655 5 1 1 36654
0 36656 7 1 2 89674 36655
0 36657 5 1 1 36656
0 36658 7 1 2 36610 36657
0 36659 7 1 2 36595 36658
0 36660 7 1 2 36541 36659
0 36661 5 1 1 36660
0 36662 7 1 2 59866 36661
0 36663 5 1 1 36662
0 36664 7 1 2 78868 93252
0 36665 5 1 1 36664
0 36666 7 1 2 65294 87793
0 36667 5 1 1 36666
0 36668 7 1 2 36665 36667
0 36669 5 1 1 36668
0 36670 7 1 2 84375 36669
0 36671 5 2 1 36670
0 36672 7 1 2 93220 93700
0 36673 5 1 1 36672
0 36674 7 1 2 91761 36673
0 36675 5 1 1 36674
0 36676 7 2 2 68392 81960
0 36677 5 2 1 93702
0 36678 7 1 2 80762 89995
0 36679 7 1 2 93704 36678
0 36680 5 1 1 36679
0 36681 7 1 2 69744 67772
0 36682 7 1 2 92674 36681
0 36683 7 1 2 92679 36682
0 36684 5 1 1 36683
0 36685 7 1 2 36680 36684
0 36686 5 1 1 36685
0 36687 7 1 2 68127 36686
0 36688 5 1 1 36687
0 36689 7 1 2 61369 36688
0 36690 7 1 2 36675 36689
0 36691 7 1 2 36663 36690
0 36692 5 1 1 36691
0 36693 7 1 2 36460 36692
0 36694 5 1 1 36693
0 36695 7 1 2 57450 33832
0 36696 5 1 1 36695
0 36697 7 1 2 93681 36696
0 36698 5 1 1 36697
0 36699 7 1 2 82882 36698
0 36700 5 1 1 36699
0 36701 7 1 2 93560 36700
0 36702 5 1 1 36701
0 36703 7 1 2 59622 36702
0 36704 5 1 1 36703
0 36705 7 3 2 58609 58991
0 36706 7 2 2 67671 93706
0 36707 7 1 2 86237 81377
0 36708 7 1 2 93709 36707
0 36709 5 1 1 36708
0 36710 7 1 2 36704 36709
0 36711 5 1 1 36710
0 36712 7 1 2 89238 36711
0 36713 5 1 1 36712
0 36714 7 1 2 60016 36713
0 36715 7 1 2 36694 36714
0 36716 7 1 2 35999 36715
0 36717 5 1 1 36716
0 36718 7 1 2 35759 36717
0 36719 5 1 1 36718
0 36720 7 1 2 85765 80508
0 36721 5 1 1 36720
0 36722 7 1 2 75234 36721
0 36723 5 1 1 36722
0 36724 7 1 2 92446 36723
0 36725 5 1 1 36724
0 36726 7 1 2 61016 74230
0 36727 5 2 1 36726
0 36728 7 1 2 72354 80080
0 36729 7 2 2 93711 36728
0 36730 7 2 2 61863 93713
0 36731 7 2 2 11382 87168
0 36732 5 6 1 93717
0 36733 7 1 2 93715 93719
0 36734 5 1 1 36733
0 36735 7 1 2 36725 36734
0 36736 5 1 1 36735
0 36737 7 1 2 71189 36736
0 36738 5 1 1 36737
0 36739 7 1 2 88667 93427
0 36740 5 1 1 36739
0 36741 7 1 2 72355 88649
0 36742 5 1 1 36741
0 36743 7 1 2 36740 36742
0 36744 5 1 1 36743
0 36745 7 1 2 65646 36744
0 36746 5 1 1 36745
0 36747 7 4 2 60017 92716
0 36748 5 1 1 93725
0 36749 7 1 2 76540 93726
0 36750 5 1 1 36749
0 36751 7 1 2 36746 36750
0 36752 5 1 1 36751
0 36753 7 1 2 76760 36752
0 36754 5 1 1 36753
0 36755 7 1 2 36738 36754
0 36756 5 1 1 36755
0 36757 7 1 2 65989 36756
0 36758 5 1 1 36757
0 36759 7 2 2 60018 92880
0 36760 5 1 1 93729
0 36761 7 1 2 93716 93730
0 36762 5 1 1 36761
0 36763 7 2 2 69458 71507
0 36764 7 1 2 72663 73632
0 36765 7 1 2 88668 36764
0 36766 7 1 2 93731 36765
0 36767 5 1 1 36766
0 36768 7 1 2 36762 36767
0 36769 5 1 1 36768
0 36770 7 1 2 59867 36769
0 36771 5 1 1 36770
0 36772 7 1 2 66289 36771
0 36773 7 1 2 36758 36772
0 36774 5 1 1 36773
0 36775 7 1 2 92881 93608
0 36776 5 1 1 36775
0 36777 7 2 2 63358 73316
0 36778 5 3 1 93733
0 36779 7 1 2 69459 93734
0 36780 5 1 1 36779
0 36781 7 1 2 36776 36780
0 36782 5 1 1 36781
0 36783 7 1 2 89266 36782
0 36784 5 1 1 36783
0 36785 7 1 2 87499 89448
0 36786 7 1 2 76370 36785
0 36787 5 1 1 36786
0 36788 7 1 2 36784 36787
0 36789 5 1 1 36788
0 36790 7 1 2 60019 36789
0 36791 5 1 1 36790
0 36792 7 1 2 73382 82640
0 36793 7 1 2 90075 36792
0 36794 7 1 2 69460 36793
0 36795 5 1 1 36794
0 36796 7 1 2 61669 36795
0 36797 7 1 2 36791 36796
0 36798 5 1 1 36797
0 36799 7 1 2 75333 36798
0 36800 7 1 2 36774 36799
0 36801 5 1 1 36800
0 36802 7 1 2 58761 36801
0 36803 7 1 2 36719 36802
0 36804 5 1 1 36803
0 36805 7 1 2 69245 36804
0 36806 7 1 2 35430 36805
0 36807 5 1 1 36806
0 36808 7 1 2 34948 36807
0 36809 5 1 1 36808
0 36810 7 1 2 58864 36809
0 36811 5 1 1 36810
0 36812 7 2 2 70373 69745
0 36813 5 1 1 93738
0 36814 7 1 2 84851 93554
0 36815 5 1 1 36814
0 36816 7 1 2 93739 36815
0 36817 5 1 1 36816
0 36818 7 1 2 93701 36817
0 36819 5 1 1 36818
0 36820 7 1 2 61370 36819
0 36821 5 1 1 36820
0 36822 7 1 2 74728 93676
0 36823 5 1 1 36822
0 36824 7 1 2 36821 36823
0 36825 5 2 1 36824
0 36826 7 1 2 90104 93740
0 36827 5 1 1 36826
0 36828 7 1 2 70329 92918
0 36829 5 1 1 36828
0 36830 7 1 2 60628 78007
0 36831 7 1 2 93341 36830
0 36832 5 1 1 36831
0 36833 7 1 2 36829 36832
0 36834 5 1 1 36833
0 36835 7 1 2 92546 36834
0 36836 5 1 1 36835
0 36837 7 1 2 93457 36836
0 36838 5 1 1 36837
0 36839 7 1 2 69049 36838
0 36840 5 1 1 36839
0 36841 7 1 2 64373 93270
0 36842 5 2 1 36841
0 36843 7 2 2 78509 93742
0 36844 5 1 1 93744
0 36845 7 3 2 63911 72151
0 36846 5 1 1 93746
0 36847 7 1 2 71692 93747
0 36848 5 1 1 36847
0 36849 7 1 2 61371 75038
0 36850 7 1 2 36848 36849
0 36851 7 1 2 93745 36850
0 36852 5 1 1 36851
0 36853 7 1 2 64374 86764
0 36854 5 1 1 36853
0 36855 7 2 2 78244 77474
0 36856 5 1 1 93749
0 36857 7 1 2 93470 36856
0 36858 7 1 2 36854 36857
0 36859 5 1 1 36858
0 36860 7 1 2 61017 36859
0 36861 5 1 1 36860
0 36862 7 1 2 65990 93526
0 36863 7 1 2 36861 36862
0 36864 5 1 1 36863
0 36865 7 1 2 36852 36864
0 36866 5 1 1 36865
0 36867 7 1 2 64375 80517
0 36868 5 1 1 36867
0 36869 7 1 2 71693 77951
0 36870 5 1 1 36869
0 36871 7 1 2 36868 36870
0 36872 5 1 1 36871
0 36873 7 1 2 62497 36872
0 36874 5 1 1 36873
0 36875 7 1 2 76081 88774
0 36876 5 2 1 36875
0 36877 7 1 2 58330 93751
0 36878 5 1 1 36877
0 36879 7 1 2 64376 36878
0 36880 5 1 1 36879
0 36881 7 1 2 36874 36880
0 36882 5 1 1 36881
0 36883 7 1 2 65991 36882
0 36884 5 1 1 36883
0 36885 7 1 2 67565 73633
0 36886 5 1 1 36885
0 36887 7 1 2 36884 36886
0 36888 5 1 1 36887
0 36889 7 1 2 68128 36888
0 36890 5 1 1 36889
0 36891 7 1 2 86590 90012
0 36892 5 1 1 36891
0 36893 7 1 2 77495 90413
0 36894 5 1 1 36893
0 36895 7 1 2 36892 36894
0 36896 5 1 1 36895
0 36897 7 1 2 35122 36896
0 36898 5 1 1 36897
0 36899 7 3 2 79116 67024
0 36900 7 1 2 65992 72513
0 36901 5 1 1 36900
0 36902 7 1 2 86373 36901
0 36903 5 1 1 36902
0 36904 7 1 2 60629 36903
0 36905 5 1 1 36904
0 36906 7 2 2 62765 90931
0 36907 5 1 1 93756
0 36908 7 1 2 80447 93757
0 36909 5 1 1 36908
0 36910 7 1 2 61372 83457
0 36911 5 1 1 36910
0 36912 7 1 2 90904 36911
0 36913 7 1 2 36909 36912
0 36914 7 1 2 36905 36913
0 36915 5 1 1 36914
0 36916 7 1 2 93753 36915
0 36917 5 1 1 36916
0 36918 7 1 2 36898 36917
0 36919 7 1 2 36890 36918
0 36920 7 1 2 36866 36919
0 36921 7 1 2 36840 36920
0 36922 5 1 1 36921
0 36923 7 1 2 58610 36922
0 36924 5 1 1 36923
0 36925 7 1 2 72664 84906
0 36926 5 1 1 36925
0 36927 7 1 2 83945 86178
0 36928 5 1 1 36927
0 36929 7 1 2 82909 36928
0 36930 7 1 2 36926 36929
0 36931 5 1 1 36930
0 36932 7 1 2 78319 36931
0 36933 5 1 1 36932
0 36934 7 1 2 77520 88257
0 36935 5 1 1 36934
0 36936 7 1 2 78176 36935
0 36937 5 1 1 36936
0 36938 7 1 2 70256 36937
0 36939 5 1 1 36938
0 36940 7 1 2 72665 90978
0 36941 7 1 2 78221 36940
0 36942 5 1 1 36941
0 36943 7 4 2 59623 69003
0 36944 7 1 2 80651 93758
0 36945 5 1 1 36944
0 36946 7 1 2 86227 36945
0 36947 7 1 2 36942 36946
0 36948 7 1 2 36939 36947
0 36949 5 1 1 36948
0 36950 7 1 2 71900 36949
0 36951 5 1 1 36950
0 36952 7 1 2 69315 76330
0 36953 5 1 1 36952
0 36954 7 2 2 59624 78610
0 36955 5 1 1 93762
0 36956 7 1 2 63359 93763
0 36957 5 1 1 36956
0 36958 7 1 2 36953 36957
0 36959 5 1 1 36958
0 36960 7 1 2 58331 36959
0 36961 5 1 1 36960
0 36962 7 2 2 70174 79710
0 36963 5 1 1 93764
0 36964 7 1 2 63360 93765
0 36965 5 1 1 36964
0 36966 7 1 2 61373 36965
0 36967 7 1 2 36961 36966
0 36968 7 1 2 36951 36967
0 36969 7 1 2 36933 36968
0 36970 5 1 1 36969
0 36971 7 1 2 75334 93428
0 36972 5 1 1 36971
0 36973 7 1 2 76300 83281
0 36974 5 1 1 36973
0 36975 7 3 2 67353 80494
0 36976 7 1 2 74379 93766
0 36977 5 1 1 36976
0 36978 7 1 2 36974 36977
0 36979 5 1 1 36978
0 36980 7 1 2 68393 36979
0 36981 5 1 1 36980
0 36982 7 1 2 65647 36981
0 36983 7 1 2 36972 36982
0 36984 7 1 2 93410 36983
0 36985 5 1 1 36984
0 36986 7 1 2 84809 85321
0 36987 7 1 2 93478 36986
0 36988 5 1 1 36987
0 36989 7 1 2 63361 36988
0 36990 7 1 2 36985 36989
0 36991 5 1 1 36990
0 36992 7 1 2 59625 93539
0 36993 5 1 1 36992
0 36994 7 1 2 65993 36993
0 36995 7 1 2 36991 36994
0 36996 5 1 1 36995
0 36997 7 1 2 36970 36996
0 36998 5 1 1 36997
0 36999 7 1 2 36924 36998
0 37000 5 1 1 36999
0 37001 7 1 2 79901 37000
0 37002 5 1 1 37001
0 37003 7 1 2 80431 90105
0 37004 7 1 2 93249 37003
0 37005 5 1 1 37004
0 37006 7 1 2 59868 37005
0 37007 7 1 2 37002 37006
0 37008 5 1 1 37007
0 37009 7 2 2 80432 90810
0 37010 7 1 2 68252 93769
0 37011 5 1 1 37010
0 37012 7 2 2 85162 80448
0 37013 7 2 2 65994 87797
0 37014 5 3 1 93773
0 37015 7 1 2 93771 93775
0 37016 5 1 1 37015
0 37017 7 1 2 37011 37016
0 37018 5 1 1 37017
0 37019 7 1 2 60630 37018
0 37020 5 1 1 37019
0 37021 7 1 2 86247 90794
0 37022 5 1 1 37021
0 37023 7 1 2 37020 37022
0 37024 5 1 1 37023
0 37025 7 1 2 62243 37024
0 37026 5 1 1 37025
0 37027 7 1 2 73218 71651
0 37028 7 1 2 90784 37027
0 37029 5 1 1 37028
0 37030 7 1 2 37026 37029
0 37031 5 1 1 37030
0 37032 7 1 2 68129 37031
0 37033 5 1 1 37032
0 37034 7 1 2 60631 92390
0 37035 5 2 1 37034
0 37036 7 1 2 14606 86741
0 37037 5 2 1 37036
0 37038 7 1 2 67773 93780
0 37039 5 1 1 37038
0 37040 7 1 2 93778 37039
0 37041 5 1 1 37040
0 37042 7 1 2 61018 37041
0 37043 5 1 1 37042
0 37044 7 1 2 70950 90368
0 37045 5 1 1 37044
0 37046 7 1 2 37043 37045
0 37047 5 1 1 37046
0 37048 7 1 2 62244 37047
0 37049 5 1 1 37048
0 37050 7 1 2 86974 37049
0 37051 5 1 1 37050
0 37052 7 1 2 76214 37051
0 37053 5 1 1 37052
0 37054 7 2 2 62245 84989
0 37055 7 1 2 73076 74104
0 37056 5 1 1 37055
0 37057 7 1 2 61019 84347
0 37058 7 1 2 37056 37057
0 37059 5 1 1 37058
0 37060 7 1 2 14104 37059
0 37061 5 1 1 37060
0 37062 7 1 2 93782 37061
0 37063 5 1 1 37062
0 37064 7 3 2 80817 84612
0 37065 5 1 1 93784
0 37066 7 1 2 37063 37065
0 37067 7 1 2 37053 37066
0 37068 7 1 2 37033 37067
0 37069 5 1 1 37068
0 37070 7 1 2 69050 37069
0 37071 5 1 1 37070
0 37072 7 1 2 67213 87385
0 37073 5 2 1 37072
0 37074 7 1 2 78008 93787
0 37075 5 1 1 37074
0 37076 7 1 2 80818 37075
0 37077 5 1 1 37076
0 37078 7 1 2 77992 84990
0 37079 7 1 2 93754 37078
0 37080 5 1 1 37079
0 37081 7 1 2 65995 37080
0 37082 7 1 2 37077 37081
0 37083 5 1 1 37082
0 37084 7 2 2 61020 84991
0 37085 7 1 2 84204 70113
0 37086 7 1 2 93789 37085
0 37087 5 1 1 37086
0 37088 7 1 2 85163 84231
0 37089 5 1 1 37088
0 37090 7 1 2 37087 37089
0 37091 5 1 1 37090
0 37092 7 1 2 71694 37091
0 37093 5 1 1 37092
0 37094 7 1 2 63362 36844
0 37095 5 1 1 37094
0 37096 7 1 2 84205 67025
0 37097 7 2 2 84992 37096
0 37098 7 1 2 77036 93791
0 37099 5 1 1 37098
0 37100 7 1 2 61374 37099
0 37101 7 1 2 37095 37100
0 37102 7 1 2 37093 37101
0 37103 5 1 1 37102
0 37104 7 1 2 37083 37103
0 37105 5 1 1 37104
0 37106 7 1 2 62498 93781
0 37107 5 1 1 37106
0 37108 7 1 2 93779 37107
0 37109 5 1 1 37108
0 37110 7 1 2 79117 37109
0 37111 5 1 1 37110
0 37112 7 1 2 64377 93459
0 37113 5 1 1 37112
0 37114 7 1 2 37111 37113
0 37115 5 1 1 37114
0 37116 7 1 2 61021 37115
0 37117 5 1 1 37116
0 37118 7 1 2 86972 87386
0 37119 5 1 1 37118
0 37120 7 1 2 37117 37119
0 37121 5 1 1 37120
0 37122 7 1 2 76215 37121
0 37123 5 1 1 37122
0 37124 7 1 2 90795 93755
0 37125 5 1 1 37124
0 37126 7 1 2 30678 37125
0 37127 5 1 1 37126
0 37128 7 1 2 61375 37127
0 37129 5 1 1 37128
0 37130 7 1 2 60632 79118
0 37131 5 1 1 37130
0 37132 7 1 2 71508 71116
0 37133 7 1 2 88167 37132
0 37134 7 1 2 37131 37133
0 37135 5 1 1 37134
0 37136 7 1 2 90785 37135
0 37137 5 1 1 37136
0 37138 7 1 2 37129 37137
0 37139 5 1 1 37138
0 37140 7 1 2 68130 37139
0 37141 5 1 1 37140
0 37142 7 3 2 69791 77619
0 37143 5 1 1 93793
0 37144 7 1 2 63072 93794
0 37145 5 1 1 37144
0 37146 7 1 2 58611 37145
0 37147 5 1 1 37146
0 37148 7 1 2 73262 77610
0 37149 5 1 1 37148
0 37150 7 1 2 67566 76341
0 37151 7 1 2 92343 37150
0 37152 5 1 1 37151
0 37153 7 1 2 37149 37152
0 37154 5 1 1 37153
0 37155 7 1 2 37147 37154
0 37156 5 1 1 37155
0 37157 7 1 2 37141 37156
0 37158 7 1 2 58332 37143
0 37159 5 1 1 37158
0 37160 7 1 2 62766 90369
0 37161 5 1 1 37160
0 37162 7 1 2 61022 92391
0 37163 5 1 1 37162
0 37164 7 1 2 37161 37163
0 37165 5 1 1 37164
0 37166 7 1 2 67567 37165
0 37167 5 1 1 37166
0 37168 7 1 2 62767 80666
0 37169 5 1 1 37168
0 37170 7 1 2 37167 37169
0 37171 5 1 1 37170
0 37172 7 1 2 37159 37171
0 37173 5 1 1 37172
0 37174 7 1 2 62768 93770
0 37175 5 1 1 37174
0 37176 7 1 2 90787 37175
0 37177 5 1 1 37176
0 37178 7 1 2 67568 37177
0 37179 5 1 1 37178
0 37180 7 1 2 71305 80667
0 37181 5 1 1 37180
0 37182 7 1 2 67584 78805
0 37183 5 1 1 37182
0 37184 7 1 2 65996 75941
0 37185 5 2 1 37184
0 37186 7 1 2 37183 93796
0 37187 7 1 2 93772 37186
0 37188 5 1 1 37187
0 37189 7 1 2 37181 37188
0 37190 7 1 2 37179 37189
0 37191 5 1 1 37190
0 37192 7 1 2 69808 37191
0 37193 5 1 1 37192
0 37194 7 1 2 37173 37193
0 37195 7 1 2 37157 37194
0 37196 7 1 2 37123 37195
0 37197 7 1 2 37105 37196
0 37198 7 1 2 37071 37197
0 37199 5 1 1 37198
0 37200 7 1 2 66847 37199
0 37201 5 1 1 37200
0 37202 7 1 2 66920 93486
0 37203 5 1 1 37202
0 37204 7 1 2 64587 37203
0 37205 7 1 2 37201 37204
0 37206 5 1 1 37205
0 37207 7 1 2 37008 37206
0 37208 5 1 1 37207
0 37209 7 1 2 36827 37208
0 37210 5 1 1 37209
0 37211 7 1 2 60138 37210
0 37212 5 1 1 37211
0 37213 7 2 2 76652 85462
0 37214 5 1 1 93798
0 37215 7 1 2 71190 93799
0 37216 7 1 2 93505 37215
0 37217 5 1 1 37216
0 37218 7 1 2 37212 37217
0 37219 5 1 1 37218
0 37220 7 1 2 66290 37219
0 37221 5 1 1 37220
0 37222 7 1 2 90057 93644
0 37223 7 1 2 80316 37222
0 37224 5 1 1 37223
0 37225 7 1 2 71191 37224
0 37226 5 1 1 37225
0 37227 7 1 2 73885 78214
0 37228 5 1 1 37227
0 37229 7 1 2 71901 37228
0 37230 5 1 1 37229
0 37231 7 2 2 78320 73904
0 37232 5 1 1 93800
0 37233 7 1 2 73465 93801
0 37234 5 1 1 37233
0 37235 7 1 2 37230 37234
0 37236 5 1 1 37235
0 37237 7 1 2 65997 82130
0 37238 7 1 2 37236 37237
0 37239 5 1 1 37238
0 37240 7 1 2 37226 37239
0 37241 5 1 1 37240
0 37242 7 1 2 79902 37241
0 37243 5 1 1 37242
0 37244 7 1 2 58762 87150
0 37245 7 1 2 93133 37244
0 37246 5 1 1 37245
0 37247 7 1 2 37243 37246
0 37248 5 1 1 37247
0 37249 7 1 2 58612 37248
0 37250 5 1 1 37249
0 37251 7 1 2 63073 86871
0 37252 5 2 1 37251
0 37253 7 1 2 93116 93802
0 37254 5 1 1 37253
0 37255 7 1 2 93114 37254
0 37256 7 1 2 93110 37255
0 37257 5 1 1 37256
0 37258 7 1 2 66848 37257
0 37259 5 1 1 37258
0 37260 7 1 2 37250 37259
0 37261 5 1 1 37260
0 37262 7 1 2 59869 37261
0 37263 5 1 1 37262
0 37264 7 1 2 76361 87378
0 37265 5 1 1 37264
0 37266 7 1 2 76154 37265
0 37267 7 1 2 93065 37266
0 37268 5 1 1 37267
0 37269 7 1 2 64378 37268
0 37270 5 1 1 37269
0 37271 7 1 2 57729 84206
0 37272 5 1 1 37271
0 37273 7 1 2 79119 37272
0 37274 5 1 1 37273
0 37275 7 1 2 92895 37274
0 37276 5 1 1 37275
0 37277 7 1 2 93455 37276
0 37278 5 1 1 37277
0 37279 7 1 2 72628 79777
0 37280 5 1 1 37279
0 37281 7 1 2 32783 93259
0 37282 5 1 1 37281
0 37283 7 3 2 69051 84348
0 37284 5 1 1 93804
0 37285 7 1 2 37282 93805
0 37286 5 1 1 37285
0 37287 7 1 2 37280 37286
0 37288 7 1 2 37278 37287
0 37289 5 1 1 37288
0 37290 7 1 2 68131 37289
0 37291 5 1 1 37290
0 37292 7 2 2 64096 81454
0 37293 5 1 1 93807
0 37294 7 1 2 62769 93808
0 37295 5 3 1 37294
0 37296 7 2 2 81460 93809
0 37297 5 1 1 93812
0 37298 7 1 2 70304 37297
0 37299 5 1 1 37298
0 37300 7 1 2 58613 37299
0 37301 7 1 2 37291 37300
0 37302 7 1 2 37270 37301
0 37303 5 1 1 37302
0 37304 7 1 2 63363 93067
0 37305 5 1 1 37304
0 37306 7 1 2 65998 37305
0 37307 7 1 2 37303 37306
0 37308 5 1 1 37307
0 37309 7 1 2 70330 83953
0 37310 7 1 2 76964 37309
0 37311 5 1 1 37310
0 37312 7 1 2 4313 37311
0 37313 5 1 1 37312
0 37314 7 1 2 60402 37313
0 37315 5 1 1 37314
0 37316 7 1 2 81076 75008
0 37317 7 1 2 83144 37316
0 37318 5 1 1 37317
0 37319 7 1 2 68132 83603
0 37320 5 1 1 37319
0 37321 7 1 2 75039 37320
0 37322 7 1 2 37318 37321
0 37323 7 1 2 37315 37322
0 37324 5 1 1 37323
0 37325 7 1 2 58614 37324
0 37326 5 1 1 37325
0 37327 7 1 2 79372 93191
0 37328 5 2 1 37327
0 37329 7 1 2 83940 93339
0 37330 5 1 1 37329
0 37331 7 1 2 75187 37330
0 37332 5 1 1 37331
0 37333 7 1 2 92920 37332
0 37334 5 1 1 37333
0 37335 7 1 2 74992 35789
0 37336 5 1 1 37335
0 37337 7 1 2 63364 75009
0 37338 5 2 1 37337
0 37339 7 1 2 60633 93816
0 37340 7 1 2 37336 37339
0 37341 7 1 2 37334 37340
0 37342 5 1 1 37341
0 37343 7 1 2 93814 37342
0 37344 7 1 2 37326 37343
0 37345 5 1 1 37344
0 37346 7 1 2 61376 37345
0 37347 5 1 1 37346
0 37348 7 1 2 84622 4490
0 37349 5 1 1 37348
0 37350 7 1 2 57451 37349
0 37351 5 1 1 37350
0 37352 7 2 2 65648 75852
0 37353 5 1 1 93818
0 37354 7 2 2 76076 93819
0 37355 5 1 1 93820
0 37356 7 1 2 61377 93821
0 37357 5 1 1 37356
0 37358 7 1 2 37351 37357
0 37359 5 1 1 37358
0 37360 7 1 2 58992 37359
0 37361 5 1 1 37360
0 37362 7 1 2 67672 86028
0 37363 5 1 1 37362
0 37364 7 1 2 37361 37363
0 37365 5 1 1 37364
0 37366 7 1 2 64379 37365
0 37367 5 1 1 37366
0 37368 7 1 2 72960 83839
0 37369 5 1 1 37368
0 37370 7 1 2 63365 37369
0 37371 5 1 1 37370
0 37372 7 1 2 37367 37371
0 37373 5 1 1 37372
0 37374 7 1 2 70426 37373
0 37375 5 1 1 37374
0 37376 7 1 2 37347 37375
0 37377 7 1 2 37308 37376
0 37378 7 1 2 82956 79381
0 37379 5 1 1 37378
0 37380 7 2 2 57730 75203
0 37381 5 2 1 93822
0 37382 7 2 2 93371 93824
0 37383 7 1 2 73210 88780
0 37384 5 1 1 37383
0 37385 7 1 2 92970 37384
0 37386 7 1 2 93826 37385
0 37387 5 1 1 37386
0 37388 7 1 2 78934 37387
0 37389 5 1 1 37388
0 37390 7 1 2 37379 37389
0 37391 5 1 1 37390
0 37392 7 1 2 61378 37391
0 37393 5 1 1 37392
0 37394 7 1 2 79013 83703
0 37395 5 1 1 37394
0 37396 7 1 2 73956 81703
0 37397 5 1 1 37396
0 37398 7 1 2 57452 37397
0 37399 5 1 1 37398
0 37400 7 1 2 64380 80608
0 37401 5 4 1 37400
0 37402 7 1 2 59139 93828
0 37403 5 1 1 37402
0 37404 7 1 2 37399 37403
0 37405 5 1 1 37404
0 37406 7 1 2 65066 37405
0 37407 5 1 1 37406
0 37408 7 1 2 70781 72907
0 37409 5 2 1 37408
0 37410 7 1 2 85825 93832
0 37411 7 1 2 37407 37410
0 37412 5 1 1 37411
0 37413 7 1 2 63366 37412
0 37414 5 1 1 37413
0 37415 7 1 2 37395 37414
0 37416 5 1 1 37415
0 37417 7 1 2 57731 37416
0 37418 5 1 1 37417
0 37419 7 1 2 85823 81601
0 37420 5 1 1 37419
0 37421 7 1 2 79106 93759
0 37422 5 1 1 37421
0 37423 7 1 2 16686 82707
0 37424 5 1 1 37423
0 37425 7 1 2 73211 37424
0 37426 5 1 1 37425
0 37427 7 1 2 37422 37426
0 37428 7 1 2 37420 37427
0 37429 5 1 1 37428
0 37430 7 1 2 63367 37429
0 37431 5 1 1 37430
0 37432 7 1 2 37418 37431
0 37433 7 1 2 37393 37432
0 37434 5 1 1 37433
0 37435 7 1 2 67354 37434
0 37436 5 1 1 37435
0 37437 7 1 2 61379 82081
0 37438 5 1 1 37437
0 37439 7 1 2 57453 37438
0 37440 5 1 1 37439
0 37441 7 1 2 37440 37355
0 37442 5 1 1 37441
0 37443 7 1 2 58993 37442
0 37444 5 1 1 37443
0 37445 7 1 2 71973 78999
0 37446 7 1 2 37444 37445
0 37447 5 1 1 37446
0 37448 7 1 2 63368 37447
0 37449 5 1 1 37448
0 37450 7 1 2 62499 80072
0 37451 7 1 2 72424 37450
0 37452 5 1 1 37451
0 37453 7 1 2 36846 37452
0 37454 5 1 1 37453
0 37455 7 1 2 76216 37454
0 37456 5 1 1 37455
0 37457 7 3 2 65649 68133
0 37458 5 1 1 93834
0 37459 7 1 2 70114 77399
0 37460 7 1 2 93835 37459
0 37461 5 1 1 37460
0 37462 7 1 2 37456 37461
0 37463 5 1 1 37462
0 37464 7 1 2 69052 37463
0 37465 5 1 1 37464
0 37466 7 1 2 79120 75148
0 37467 5 1 1 37466
0 37468 7 1 2 80935 93748
0 37469 5 1 1 37468
0 37470 7 1 2 37467 37469
0 37471 5 1 1 37470
0 37472 7 1 2 62500 37471
0 37473 5 1 1 37472
0 37474 7 1 2 75149 92894
0 37475 5 1 1 37474
0 37476 7 1 2 37473 37475
0 37477 5 1 1 37476
0 37478 7 1 2 68134 37477
0 37479 5 1 1 37478
0 37480 7 1 2 80307 87965
0 37481 5 1 1 37480
0 37482 7 1 2 60634 93536
0 37483 5 1 1 37482
0 37484 7 1 2 37481 37483
0 37485 5 1 1 37484
0 37486 7 1 2 87996 37485
0 37487 5 1 1 37486
0 37488 7 2 2 7905 80073
0 37489 7 1 2 93396 93837
0 37490 5 1 1 37489
0 37491 7 1 2 93179 37490
0 37492 7 1 2 37487 37491
0 37493 7 1 2 37479 37492
0 37494 7 1 2 37465 37493
0 37495 5 1 1 37494
0 37496 7 1 2 65999 37495
0 37497 5 1 1 37496
0 37498 7 1 2 37449 37497
0 37499 5 1 1 37498
0 37500 7 1 2 59626 37499
0 37501 5 1 1 37500
0 37502 7 1 2 37436 37501
0 37503 7 1 2 37377 37502
0 37504 5 1 1 37503
0 37505 7 1 2 79570 37504
0 37506 5 1 1 37505
0 37507 7 1 2 37263 37506
0 37508 5 1 1 37507
0 37509 7 1 2 89567 37508
0 37510 5 1 1 37509
0 37511 7 1 2 37221 37510
0 37512 5 1 1 37511
0 37513 7 1 2 66507 37512
0 37514 5 1 1 37513
0 37515 7 1 2 87798 88817
0 37516 7 3 2 73935 37515
0 37517 5 2 1 93839
0 37518 7 1 2 92200 93840
0 37519 5 1 1 37518
0 37520 7 1 2 78686 91389
0 37521 5 1 1 37520
0 37522 7 1 2 65650 88485
0 37523 5 1 1 37522
0 37524 7 1 2 63074 75010
0 37525 7 1 2 37523 37524
0 37526 5 1 1 37525
0 37527 7 1 2 37521 37526
0 37528 5 1 1 37527
0 37529 7 1 2 75906 37528
0 37530 5 1 1 37529
0 37531 7 1 2 78687 88630
0 37532 5 1 1 37531
0 37533 7 1 2 62770 88493
0 37534 5 1 1 37533
0 37535 7 1 2 37532 37534
0 37536 5 1 1 37535
0 37537 7 1 2 81859 37536
0 37538 5 1 1 37537
0 37539 7 1 2 84927 93537
0 37540 5 1 1 37539
0 37541 7 2 2 91145 92475
0 37542 5 1 1 93844
0 37543 7 1 2 60403 9787
0 37544 5 2 1 37543
0 37545 7 1 2 76217 93846
0 37546 7 1 2 93845 37545
0 37547 5 1 1 37546
0 37548 7 1 2 37540 37547
0 37549 5 1 1 37548
0 37550 7 1 2 70829 37549
0 37551 5 1 1 37550
0 37552 7 1 2 72782 78127
0 37553 5 1 1 37552
0 37554 7 1 2 63369 77622
0 37555 5 1 1 37554
0 37556 7 1 2 37553 37555
0 37557 7 1 2 37551 37556
0 37558 7 1 2 37538 37557
0 37559 7 1 2 37530 37558
0 37560 5 1 1 37559
0 37561 7 1 2 59870 37560
0 37562 5 1 1 37561
0 37563 7 1 2 73936 77233
0 37564 5 1 1 37563
0 37565 7 1 2 77811 37564
0 37566 5 1 1 37565
0 37567 7 1 2 68394 37566
0 37568 5 1 1 37567
0 37569 7 1 2 77812 79321
0 37570 5 1 1 37569
0 37571 7 1 2 58062 37570
0 37572 5 1 1 37571
0 37573 7 1 2 93235 37572
0 37574 7 1 2 37568 37573
0 37575 7 1 2 37562 37574
0 37576 5 1 1 37575
0 37577 7 1 2 60020 37576
0 37578 5 1 1 37577
0 37579 7 1 2 37519 37578
0 37580 5 1 1 37579
0 37581 7 1 2 58763 37580
0 37582 5 1 1 37581
0 37583 7 5 2 86995 73966
0 37584 7 1 2 63511 93848
0 37585 7 1 2 93841 37584
0 37586 5 1 1 37585
0 37587 7 1 2 37582 37586
0 37588 5 1 1 37587
0 37589 7 1 2 59627 37588
0 37590 5 1 1 37589
0 37591 7 1 2 77826 85501
0 37592 5 1 1 37591
0 37593 7 1 2 76816 90589
0 37594 5 1 1 37593
0 37595 7 1 2 93817 37594
0 37596 5 1 1 37595
0 37597 7 1 2 70427 37596
0 37598 5 1 1 37597
0 37599 7 1 2 77923 90590
0 37600 5 1 1 37599
0 37601 7 1 2 78975 83720
0 37602 7 1 2 92972 37601
0 37603 5 1 1 37602
0 37604 7 1 2 63370 37603
0 37605 5 1 1 37604
0 37606 7 1 2 37600 37605
0 37607 5 1 1 37606
0 37608 7 1 2 67355 37607
0 37609 5 1 1 37608
0 37610 7 1 2 37598 37609
0 37611 7 1 2 93345 37610
0 37612 5 1 1 37611
0 37613 7 1 2 59871 37612
0 37614 5 1 1 37613
0 37615 7 1 2 37592 37614
0 37616 5 1 1 37615
0 37617 7 1 2 66849 37616
0 37618 5 1 1 37617
0 37619 7 1 2 37590 37618
0 37620 5 1 1 37619
0 37621 7 1 2 66000 37620
0 37622 5 1 1 37621
0 37623 7 2 2 61380 76980
0 37624 5 1 1 93853
0 37625 7 1 2 87249 80165
0 37626 5 1 1 37625
0 37627 7 1 2 93854 37626
0 37628 5 1 1 37627
0 37629 7 1 2 80148 78869
0 37630 5 1 1 37629
0 37631 7 1 2 86219 93383
0 37632 7 1 2 37630 37631
0 37633 5 1 1 37632
0 37634 7 1 2 80565 37633
0 37635 5 1 1 37634
0 37636 7 2 2 68135 91992
0 37637 5 1 1 93855
0 37638 7 1 2 92891 37637
0 37639 5 1 1 37638
0 37640 7 1 2 82910 37639
0 37641 7 1 2 37635 37640
0 37642 5 1 1 37641
0 37643 7 1 2 65651 37642
0 37644 5 1 1 37643
0 37645 7 1 2 37628 37644
0 37646 5 1 1 37645
0 37647 7 1 2 59872 37646
0 37648 5 1 1 37647
0 37649 7 1 2 93557 37648
0 37650 5 1 1 37649
0 37651 7 1 2 66850 37650
0 37652 5 1 1 37651
0 37653 7 1 2 37622 37652
0 37654 5 1 1 37653
0 37655 7 1 2 66291 37654
0 37656 5 1 1 37655
0 37657 7 4 2 60021 73317
0 37658 7 1 2 82785 93707
0 37659 7 1 2 93857 37658
0 37660 5 1 1 37659
0 37661 7 1 2 69004 66851
0 37662 7 1 2 85547 37661
0 37663 7 1 2 75335 37662
0 37664 5 1 1 37663
0 37665 7 1 2 37660 37664
0 37666 5 1 1 37665
0 37667 7 1 2 82566 37666
0 37668 5 1 1 37667
0 37669 7 1 2 70086 85843
0 37670 5 1 1 37669
0 37671 7 1 2 82451 37670
0 37672 5 1 1 37671
0 37673 7 1 2 65652 37672
0 37674 5 1 1 37673
0 37675 7 1 2 66001 67895
0 37676 5 1 1 37675
0 37677 7 2 2 37674 37676
0 37678 5 2 1 93861
0 37679 7 1 2 92203 93863
0 37680 5 1 1 37679
0 37681 7 1 2 85048 82452
0 37682 5 1 1 37681
0 37683 7 1 2 69005 37682
0 37684 5 1 1 37683
0 37685 7 1 2 76240 37684
0 37686 5 1 1 37685
0 37687 7 1 2 57454 37686
0 37688 5 1 1 37687
0 37689 7 1 2 76218 81077
0 37690 5 1 1 37689
0 37691 7 1 2 67673 37690
0 37692 5 1 1 37691
0 37693 7 1 2 78922 37692
0 37694 7 1 2 37688 37693
0 37695 5 1 1 37694
0 37696 7 1 2 64381 37695
0 37697 5 1 1 37696
0 37698 7 1 2 87022 37697
0 37699 5 1 1 37698
0 37700 7 1 2 61381 37699
0 37701 5 1 1 37700
0 37702 7 1 2 76965 92899
0 37703 5 1 1 37702
0 37704 7 1 2 58615 91284
0 37705 5 1 1 37704
0 37706 7 1 2 37703 37705
0 37707 5 1 1 37706
0 37708 7 1 2 60404 37707
0 37709 5 1 1 37708
0 37710 7 1 2 73669 93617
0 37711 5 1 1 37710
0 37712 7 1 2 80571 37711
0 37713 5 1 1 37712
0 37714 7 1 2 68022 29594
0 37715 5 1 1 37714
0 37716 7 1 2 37713 37715
0 37717 5 1 1 37716
0 37718 7 1 2 37709 37717
0 37719 5 1 1 37718
0 37720 7 1 2 61023 37719
0 37721 5 1 1 37720
0 37722 7 1 2 59628 75173
0 37723 5 1 1 37722
0 37724 7 1 2 34772 37723
0 37725 5 1 1 37724
0 37726 7 1 2 67356 37725
0 37727 5 1 1 37726
0 37728 7 1 2 70374 79621
0 37729 7 1 2 37727 37728
0 37730 5 1 1 37729
0 37731 7 1 2 86985 37730
0 37732 5 1 1 37731
0 37733 7 1 2 59873 37732
0 37734 7 1 2 37721 37733
0 37735 7 1 2 37701 37734
0 37736 5 1 1 37735
0 37737 7 1 2 63371 93862
0 37738 5 1 1 37737
0 37739 7 1 2 71192 37738
0 37740 5 1 1 37739
0 37741 7 1 2 79622 78819
0 37742 5 1 1 37741
0 37743 7 1 2 85548 37742
0 37744 5 1 1 37743
0 37745 7 1 2 64588 37744
0 37746 7 1 2 37740 37745
0 37747 5 1 1 37746
0 37748 7 1 2 60022 37747
0 37749 7 1 2 37736 37748
0 37750 5 1 1 37749
0 37751 7 1 2 37680 37750
0 37752 5 1 1 37751
0 37753 7 1 2 58764 37752
0 37754 5 1 1 37753
0 37755 7 2 2 74667 93849
0 37756 7 1 2 93864 93865
0 37757 5 1 1 37756
0 37758 7 1 2 71193 93720
0 37759 5 2 1 37758
0 37760 7 1 2 60023 76761
0 37761 5 1 1 37760
0 37762 7 1 2 93867 37761
0 37763 5 1 1 37762
0 37764 7 1 2 66002 37763
0 37765 5 1 1 37764
0 37766 7 1 2 73967 87147
0 37767 5 1 1 37766
0 37768 7 1 2 37765 37767
0 37769 5 1 1 37768
0 37770 7 1 2 58765 37769
0 37771 5 1 1 37770
0 37772 7 2 2 76926 87500
0 37773 7 1 2 82313 93869
0 37774 5 1 1 37773
0 37775 7 1 2 37771 37774
0 37776 5 1 1 37775
0 37777 7 1 2 75204 37776
0 37778 5 1 1 37777
0 37779 7 1 2 66852 74194
0 37780 7 1 2 73837 37779
0 37781 5 1 1 37780
0 37782 7 1 2 37778 37781
0 37783 5 1 1 37782
0 37784 7 1 2 75336 37783
0 37785 5 1 1 37784
0 37786 7 1 2 37757 37785
0 37787 7 1 2 37754 37786
0 37788 5 1 1 37787
0 37789 7 1 2 66292 37788
0 37790 5 1 1 37789
0 37791 7 1 2 37668 37790
0 37792 5 1 1 37791
0 37793 7 1 2 65295 37792
0 37794 5 1 1 37793
0 37795 7 1 2 87316 79422
0 37796 5 2 1 37795
0 37797 7 1 2 68023 93871
0 37798 5 3 1 37797
0 37799 7 1 2 59874 86986
0 37800 5 1 1 37799
0 37801 7 1 2 25925 37800
0 37802 7 2 2 92009 37801
0 37803 5 2 1 93876
0 37804 7 1 2 93873 93877
0 37805 5 1 1 37804
0 37806 7 2 2 65653 37805
0 37807 5 1 1 93880
0 37808 7 1 2 85404 93355
0 37809 5 1 1 37808
0 37810 7 1 2 37807 37809
0 37811 5 2 1 37810
0 37812 7 1 2 60024 93882
0 37813 5 1 1 37812
0 37814 7 4 2 72935 36907
0 37815 5 1 1 93884
0 37816 7 1 2 92204 93885
0 37817 5 1 1 37816
0 37818 7 1 2 37813 37817
0 37819 5 1 1 37818
0 37820 7 1 2 58766 37819
0 37821 5 1 1 37820
0 37822 7 1 2 93866 93886
0 37823 5 1 1 37822
0 37824 7 1 2 37821 37823
0 37825 5 1 1 37824
0 37826 7 1 2 86838 37825
0 37827 5 1 1 37826
0 37828 7 1 2 78611 86489
0 37829 7 1 2 92517 37828
0 37830 5 1 1 37829
0 37831 7 1 2 37827 37830
0 37832 5 1 1 37831
0 37833 7 1 2 93301 37832
0 37834 5 1 1 37833
0 37835 7 1 2 81433 92581
0 37836 5 1 1 37835
0 37837 7 1 2 4908 92167
0 37838 5 4 1 37837
0 37839 7 1 2 71194 93888
0 37840 5 1 1 37839
0 37841 7 1 2 86996 79554
0 37842 5 2 1 37841
0 37843 7 1 2 37840 93892
0 37844 5 1 1 37843
0 37845 7 1 2 86839 37844
0 37846 5 1 1 37845
0 37847 7 3 2 66853 89386
0 37848 5 1 1 93894
0 37849 7 1 2 37846 37848
0 37850 5 1 1 37849
0 37851 7 1 2 73875 37850
0 37852 5 1 1 37851
0 37853 7 1 2 86920 93889
0 37854 5 1 1 37853
0 37855 7 1 2 59875 90106
0 37856 5 1 1 37855
0 37857 7 1 2 37854 37856
0 37858 5 1 1 37857
0 37859 7 1 2 57455 81875
0 37860 7 1 2 37858 37859
0 37861 5 1 1 37860
0 37862 7 1 2 37852 37861
0 37863 5 1 1 37862
0 37864 7 1 2 93498 37863
0 37865 5 1 1 37864
0 37866 7 1 2 37836 37865
0 37867 7 1 2 37834 37866
0 37868 7 1 2 37794 37867
0 37869 7 1 2 37656 37868
0 37870 5 1 1 37869
0 37871 7 1 2 91321 37870
0 37872 5 1 1 37871
0 37873 7 1 2 37514 37872
0 37874 5 1 1 37873
0 37875 7 1 2 72562 37874
0 37876 5 1 1 37875
0 37877 7 1 2 36811 37876
0 37878 5 1 1 37877
0 37879 7 1 2 66601 37878
0 37880 5 1 1 37879
0 37881 7 2 2 79529 90032
0 37882 5 1 1 93897
0 37883 7 1 2 65654 83767
0 37884 5 1 1 37883
0 37885 7 1 2 73466 75174
0 37886 5 2 1 37885
0 37887 7 1 2 37884 93899
0 37888 5 1 1 37887
0 37889 7 1 2 57732 37888
0 37890 5 1 1 37889
0 37891 7 1 2 4556 37890
0 37892 5 2 1 37891
0 37893 7 1 2 66003 93901
0 37894 5 1 1 37893
0 37895 7 1 2 93621 37894
0 37896 5 1 1 37895
0 37897 7 1 2 89596 37896
0 37898 5 1 1 37897
0 37899 7 1 2 37882 37898
0 37900 5 1 1 37899
0 37901 7 1 2 64589 37900
0 37902 5 1 1 37901
0 37903 7 1 2 90005 37902
0 37904 5 1 1 37903
0 37905 7 1 2 66602 37904
0 37906 5 1 1 37905
0 37907 7 1 2 77152 82475
0 37908 5 2 1 37907
0 37909 7 1 2 81234 81455
0 37910 7 1 2 93903 37909
0 37911 5 1 1 37910
0 37912 7 2 2 90625 37911
0 37913 7 1 2 76653 93905
0 37914 5 1 1 37913
0 37915 7 1 2 37906 37914
0 37916 5 1 1 37915
0 37917 7 1 2 64718 37916
0 37918 5 1 1 37917
0 37919 7 1 2 76243 89267
0 37920 5 1 1 37919
0 37921 7 1 2 73467 89243
0 37922 5 2 1 37921
0 37923 7 1 2 66508 73547
0 37924 5 1 1 37923
0 37925 7 1 2 92693 37924
0 37926 5 1 1 37925
0 37927 7 1 2 71902 37926
0 37928 5 1 1 37927
0 37929 7 1 2 93907 37928
0 37930 7 1 2 37920 37929
0 37931 5 1 1 37930
0 37932 7 1 2 75285 37931
0 37933 5 1 1 37932
0 37934 7 1 2 72101 80689
0 37935 5 1 1 37934
0 37936 7 2 2 66509 37935
0 37937 7 1 2 64590 93909
0 37938 5 1 1 37937
0 37939 7 1 2 93908 37938
0 37940 5 1 1 37939
0 37941 7 1 2 57733 37940
0 37942 5 1 1 37941
0 37943 7 7 2 59140 64591
0 37944 7 1 2 88799 93911
0 37945 5 1 1 37944
0 37946 7 1 2 93642 37945
0 37947 5 1 1 37946
0 37948 7 1 2 65655 37947
0 37949 5 1 1 37948
0 37950 7 1 2 37942 37949
0 37951 7 1 2 37933 37950
0 37952 5 1 1 37951
0 37953 7 1 2 86566 37952
0 37954 5 1 1 37953
0 37955 7 1 2 61670 89008
0 37956 5 1 1 37955
0 37957 7 1 2 37954 37956
0 37958 5 1 1 37957
0 37959 7 1 2 75960 37958
0 37960 5 1 1 37959
0 37961 7 1 2 37918 37960
0 37962 5 1 1 37961
0 37963 7 1 2 63512 37962
0 37964 5 1 1 37963
0 37965 7 1 2 61671 88790
0 37966 5 1 1 37965
0 37967 7 1 2 77153 79732
0 37968 5 1 1 37967
0 37969 7 1 2 82468 37968
0 37970 5 2 1 37969
0 37971 7 1 2 87534 91142
0 37972 7 1 2 93918 37971
0 37973 5 1 1 37972
0 37974 7 1 2 37966 37973
0 37975 5 1 1 37974
0 37976 7 1 2 76654 37975
0 37977 5 1 1 37976
0 37978 7 1 2 73468 88650
0 37979 5 1 1 37978
0 37980 7 1 2 64719 93910
0 37981 5 1 1 37980
0 37982 7 1 2 37979 37981
0 37983 5 1 1 37982
0 37984 7 1 2 57734 37983
0 37985 5 1 1 37984
0 37986 7 1 2 88655 19991
0 37987 5 2 1 37986
0 37988 7 1 2 59141 93920
0 37989 5 1 1 37988
0 37990 7 1 2 88742 37989
0 37991 5 1 1 37990
0 37992 7 1 2 65656 37991
0 37993 5 1 1 37992
0 37994 7 1 2 79517 93921
0 37995 5 1 1 37994
0 37996 7 1 2 65657 88669
0 37997 5 1 1 37996
0 37998 7 1 2 88743 37997
0 37999 5 1 1 37998
0 38000 7 1 2 68395 37999
0 38001 5 1 1 38000
0 38002 7 1 2 37995 38001
0 38003 5 1 1 38002
0 38004 7 1 2 77154 38003
0 38005 5 1 1 38004
0 38006 7 1 2 37993 38005
0 38007 7 1 2 37985 38006
0 38008 5 1 1 38007
0 38009 7 1 2 86567 38008
0 38010 5 1 1 38009
0 38011 7 1 2 87151 90033
0 38012 5 1 1 38011
0 38013 7 1 2 38010 38012
0 38014 5 1 1 38013
0 38015 7 1 2 64592 38014
0 38016 5 1 1 38015
0 38017 7 1 2 37977 38016
0 38018 5 1 1 38017
0 38019 7 1 2 75683 38018
0 38020 5 1 1 38019
0 38021 7 1 2 37964 38020
0 38022 5 1 1 38021
0 38023 7 1 2 67931 38022
0 38024 5 1 1 38023
0 38025 7 4 2 91827 92222
0 38026 7 4 2 65658 86614
0 38027 7 1 2 90076 93926
0 38028 7 1 2 93922 38027
0 38029 7 1 2 80916 38028
0 38030 5 1 1 38029
0 38031 7 1 2 38024 38030
0 38032 5 1 1 38031
0 38033 7 1 2 68024 38032
0 38034 5 1 1 38033
0 38035 7 1 2 79366 87550
0 38036 5 1 1 38035
0 38037 7 1 2 72766 82233
0 38038 5 1 1 38037
0 38039 7 1 2 68025 87535
0 38040 7 1 2 38038 38039
0 38041 5 1 1 38040
0 38042 7 1 2 38036 38041
0 38043 5 1 1 38042
0 38044 7 1 2 89268 38043
0 38045 5 1 1 38044
0 38046 7 2 2 60025 60635
0 38047 7 1 2 59876 93930
0 38048 7 1 2 90195 38047
0 38049 5 1 1 38048
0 38050 7 1 2 38045 38049
0 38051 5 1 1 38050
0 38052 7 1 2 61382 38051
0 38053 5 1 1 38052
0 38054 7 1 2 86881 89657
0 38055 5 1 1 38054
0 38056 7 1 2 89632 93902
0 38057 5 1 1 38056
0 38058 7 1 2 38055 38057
0 38059 5 1 1 38058
0 38060 7 1 2 64720 38059
0 38061 5 1 1 38060
0 38062 7 1 2 31539 38061
0 38063 5 1 1 38062
0 38064 7 1 2 59877 38063
0 38065 5 1 1 38064
0 38066 7 1 2 70331 88791
0 38067 7 2 2 87559 87543
0 38068 5 1 1 93932
0 38069 7 2 2 79271 86681
0 38070 7 1 2 93933 93934
0 38071 7 1 2 38066 38070
0 38072 5 1 1 38071
0 38073 7 1 2 38065 38072
0 38074 5 1 1 38073
0 38075 7 1 2 68026 38074
0 38076 5 1 1 38075
0 38077 7 1 2 38053 38076
0 38078 5 1 1 38077
0 38079 7 1 2 58767 38078
0 38080 5 1 1 38079
0 38081 7 3 2 64593 87137
0 38082 5 3 1 93936
0 38083 7 3 2 73562 91546
0 38084 5 1 1 93942
0 38085 7 1 2 73794 93943
0 38086 5 1 1 38085
0 38087 7 1 2 93939 38086
0 38088 5 1 1 38087
0 38089 7 1 2 75786 38088
0 38090 5 1 1 38089
0 38091 7 3 2 64594 73634
0 38092 7 1 2 60026 93945
0 38093 5 1 1 38092
0 38094 7 2 2 84005 86107
0 38095 5 1 1 93948
0 38096 7 3 2 59142 59878
0 38097 7 3 2 57735 93950
0 38098 7 1 2 72479 87577
0 38099 7 2 2 93953 38098
0 38100 5 1 1 93956
0 38101 7 1 2 38095 38100
0 38102 5 1 1 38101
0 38103 7 1 2 68625 38102
0 38104 5 1 1 38103
0 38105 7 1 2 38093 38104
0 38106 7 1 2 38090 38105
0 38107 5 1 1 38106
0 38108 7 1 2 66510 38107
0 38109 5 1 1 38108
0 38110 7 1 2 73469 78207
0 38111 5 2 1 38110
0 38112 7 1 2 73436 93958
0 38113 5 1 1 38112
0 38114 7 1 2 57456 38113
0 38115 5 2 1 38114
0 38116 7 1 2 7109 93960
0 38117 5 1 1 38116
0 38118 7 1 2 87501 88651
0 38119 7 1 2 38117 38118
0 38120 5 1 1 38119
0 38121 7 1 2 38109 38120
0 38122 5 1 1 38121
0 38123 7 1 2 66293 38122
0 38124 5 1 1 38123
0 38125 7 1 2 70352 86840
0 38126 7 1 2 80605 74849
0 38127 7 1 2 38125 38126
0 38128 5 1 1 38127
0 38129 7 1 2 87560 38128
0 38130 5 1 1 38129
0 38131 7 1 2 66511 38130
0 38132 5 1 1 38131
0 38133 7 1 2 87608 91249
0 38134 7 1 2 78366 38133
0 38135 5 1 1 38134
0 38136 7 1 2 38132 38135
0 38137 5 1 1 38136
0 38138 7 1 2 59879 38137
0 38139 5 1 1 38138
0 38140 7 1 2 90258 92060
0 38141 5 1 1 38140
0 38142 7 1 2 38139 38141
0 38143 5 1 1 38142
0 38144 7 1 2 71903 38143
0 38145 5 1 1 38144
0 38146 7 1 2 79057 84244
0 38147 5 1 1 38146
0 38148 7 1 2 87551 89428
0 38149 7 1 2 38147 38148
0 38150 5 1 1 38149
0 38151 7 1 2 38145 38150
0 38152 7 1 2 38124 38151
0 38153 5 1 1 38152
0 38154 7 1 2 76014 38153
0 38155 5 1 1 38154
0 38156 7 1 2 38080 38155
0 38157 5 1 1 38156
0 38158 7 1 2 58616 38157
0 38159 5 1 1 38158
0 38160 7 1 2 75239 88823
0 38161 5 1 1 38160
0 38162 7 1 2 80495 92265
0 38163 5 1 1 38162
0 38164 7 1 2 38161 38163
0 38165 5 1 1 38164
0 38166 7 1 2 59143 38165
0 38167 5 1 1 38166
0 38168 7 1 2 79078 92266
0 38169 5 1 1 38168
0 38170 7 1 2 38167 38169
0 38171 5 1 1 38170
0 38172 7 1 2 57736 38171
0 38173 5 1 1 38172
0 38174 7 1 2 79132 92267
0 38175 5 1 1 38174
0 38176 7 1 2 38173 38175
0 38177 5 1 1 38176
0 38178 7 1 2 65659 38177
0 38179 5 1 1 38178
0 38180 7 2 2 74007 74895
0 38181 7 1 2 75423 88734
0 38182 7 1 2 93962 38181
0 38183 5 1 1 38182
0 38184 7 1 2 38179 38183
0 38185 5 1 1 38184
0 38186 7 1 2 86568 38185
0 38187 5 1 1 38186
0 38188 7 1 2 66854 93898
0 38189 5 1 1 38188
0 38190 7 1 2 38187 38189
0 38191 5 1 1 38190
0 38192 7 1 2 88415 38191
0 38193 5 1 1 38192
0 38194 7 1 2 38159 38193
0 38195 5 1 1 38194
0 38196 7 1 2 66603 38195
0 38197 5 1 1 38196
0 38198 7 1 2 83006 92577
0 38199 7 1 2 93906 38198
0 38200 5 1 1 38199
0 38201 7 1 2 38197 38200
0 38202 5 1 1 38201
0 38203 7 1 2 70525 38202
0 38204 5 1 1 38203
0 38205 7 6 2 66604 80433
0 38206 7 1 2 76934 89288
0 38207 7 1 2 93964 38206
0 38208 7 1 2 91275 38207
0 38209 5 1 1 38208
0 38210 7 1 2 38204 38209
0 38211 7 1 2 38034 38210
0 38212 5 1 1 38211
0 38213 7 1 2 66713 38212
0 38214 5 1 1 38213
0 38215 7 1 2 86890 81644
0 38216 5 1 1 38215
0 38217 7 3 2 76608 90311
0 38218 7 1 2 81188 93379
0 38219 7 1 2 89319 38218
0 38220 7 1 2 93970 38219
0 38221 7 1 2 38216 38220
0 38222 5 1 1 38221
0 38223 7 1 2 76762 81402
0 38224 5 1 1 38223
0 38225 7 1 2 89392 38224
0 38226 5 1 1 38225
0 38227 7 1 2 64721 38226
0 38228 5 1 1 38227
0 38229 7 6 2 84006 86803
0 38230 5 1 1 93973
0 38231 7 1 2 38228 38230
0 38232 5 1 1 38231
0 38233 7 1 2 66004 38232
0 38234 5 1 1 38233
0 38235 7 1 2 75205 82567
0 38236 5 1 1 38235
0 38237 7 1 2 17752 38236
0 38238 5 1 1 38237
0 38239 7 1 2 70970 38238
0 38240 5 1 1 38239
0 38241 7 1 2 83297 93565
0 38242 5 1 1 38241
0 38243 7 1 2 68781 87455
0 38244 5 1 1 38243
0 38245 7 1 2 91874 38244
0 38246 5 1 1 38245
0 38247 7 1 2 75874 38246
0 38248 5 1 1 38247
0 38249 7 1 2 38242 38248
0 38250 7 1 2 38240 38249
0 38251 5 1 1 38250
0 38252 7 1 2 82641 38251
0 38253 5 1 1 38252
0 38254 7 1 2 38234 38253
0 38255 5 1 1 38254
0 38256 7 1 2 58768 38255
0 38257 5 1 1 38256
0 38258 7 1 2 87456 79733
0 38259 5 1 1 38258
0 38260 7 2 2 61672 73383
0 38261 5 2 1 93979
0 38262 7 1 2 38259 93981
0 38263 5 1 1 38262
0 38264 7 1 2 65067 38263
0 38265 5 1 1 38264
0 38266 7 1 2 75875 82568
0 38267 5 1 1 38266
0 38268 7 1 2 38265 38267
0 38269 5 1 1 38268
0 38270 7 1 2 91841 38269
0 38271 5 1 1 38270
0 38272 7 1 2 57737 86651
0 38273 7 2 2 59144 84007
0 38274 7 4 2 58769 69398
0 38275 5 1 1 93985
0 38276 7 1 2 93983 93986
0 38277 7 1 2 38272 38276
0 38278 5 1 1 38277
0 38279 7 1 2 38271 38278
0 38280 5 1 1 38279
0 38281 7 1 2 68626 38280
0 38282 5 1 1 38281
0 38283 7 2 2 58617 73365
0 38284 5 1 1 93989
0 38285 7 1 2 61024 83086
0 38286 5 2 1 38285
0 38287 7 1 2 71904 93991
0 38288 5 1 1 38287
0 38289 7 1 2 65660 75787
0 38290 5 2 1 38289
0 38291 7 2 2 70782 75788
0 38292 5 1 1 93995
0 38293 7 1 2 93993 38292
0 38294 7 1 2 38288 38293
0 38295 5 1 1 38294
0 38296 7 1 2 93990 38295
0 38297 5 1 1 38296
0 38298 7 1 2 77884 73263
0 38299 5 1 1 38298
0 38300 7 1 2 38297 38299
0 38301 5 1 1 38300
0 38302 7 1 2 66294 38301
0 38303 5 1 1 38302
0 38304 7 2 2 61383 70008
0 38305 5 1 1 93997
0 38306 7 1 2 73283 82760
0 38307 5 1 1 38306
0 38308 7 1 2 77541 38307
0 38309 7 1 2 93998 38308
0 38310 7 1 2 93827 38309
0 38311 5 1 1 38310
0 38312 7 1 2 89354 38311
0 38313 5 1 1 38312
0 38314 7 1 2 38303 38313
0 38315 5 1 1 38314
0 38316 7 1 2 79862 38315
0 38317 5 1 1 38316
0 38318 7 1 2 38282 38317
0 38319 7 1 2 38257 38318
0 38320 5 1 1 38319
0 38321 7 1 2 70526 38320
0 38322 5 1 1 38321
0 38323 7 1 2 68627 80333
0 38324 7 1 2 83155 38323
0 38325 7 1 2 91679 38324
0 38326 5 1 1 38325
0 38327 7 1 2 86490 89341
0 38328 5 1 1 38327
0 38329 7 1 2 66512 38328
0 38330 7 1 2 38326 38329
0 38331 7 1 2 38322 38330
0 38332 5 1 1 38331
0 38333 7 1 2 63372 34425
0 38334 5 1 1 38333
0 38335 7 1 2 66005 38334
0 38336 5 1 1 38335
0 38337 7 1 2 65296 11082
0 38338 5 1 1 38337
0 38339 7 1 2 61025 38338
0 38340 5 1 1 38339
0 38341 7 2 2 58618 85960
0 38342 5 1 1 93999
0 38343 7 1 2 38340 94000
0 38344 5 1 1 38343
0 38345 7 1 2 38336 38344
0 38346 5 2 1 38345
0 38347 7 1 2 82211 94001
0 38348 5 1 1 38347
0 38349 7 1 2 79737 89355
0 38350 5 1 1 38349
0 38351 7 1 2 38348 38350
0 38352 5 1 1 38351
0 38353 7 1 2 79974 38352
0 38354 5 1 1 38353
0 38355 7 1 2 58865 82688
0 38356 7 1 2 73366 81026
0 38357 7 1 2 38355 38356
0 38358 5 1 1 38357
0 38359 7 3 2 73563 82529
0 38360 7 1 2 70527 92683
0 38361 7 1 2 94003 38360
0 38362 5 1 1 38361
0 38363 7 1 2 38358 38362
0 38364 5 1 1 38363
0 38365 7 1 2 57738 38364
0 38366 5 1 1 38365
0 38367 7 1 2 71905 79200
0 38368 7 1 2 89568 38367
0 38369 7 1 2 87879 38368
0 38370 5 1 1 38369
0 38371 7 1 2 38366 38370
0 38372 5 1 1 38371
0 38373 7 1 2 58994 38372
0 38374 5 1 1 38373
0 38375 7 2 2 67932 87713
0 38376 7 1 2 76077 87262
0 38377 7 1 2 94006 38376
0 38378 5 1 1 38377
0 38379 7 1 2 38374 38378
0 38380 5 1 1 38379
0 38381 7 1 2 57457 38380
0 38382 5 1 1 38381
0 38383 7 1 2 90339 92233
0 38384 7 1 2 83817 38383
0 38385 5 1 1 38384
0 38386 7 1 2 38382 38385
0 38387 5 1 1 38386
0 38388 7 1 2 66921 38387
0 38389 5 1 1 38388
0 38390 7 1 2 61864 38389
0 38391 7 1 2 38354 38390
0 38392 5 1 1 38391
0 38393 7 1 2 38332 38392
0 38394 5 1 1 38393
0 38395 7 1 2 66605 38394
0 38396 5 1 1 38395
0 38397 7 2 2 67674 94004
0 38398 7 1 2 92179 94008
0 38399 5 1 1 38398
0 38400 7 2 2 79903 89387
0 38401 5 2 1 94010
0 38402 7 1 2 38399 94012
0 38403 7 1 2 88288 93957
0 38404 5 1 1 38403
0 38405 7 3 2 60027 80434
0 38406 7 2 2 79555 94014
0 38407 5 1 1 94017
0 38408 7 3 2 61673 94018
0 38409 5 2 1 94019
0 38410 7 1 2 38404 94022
0 38411 7 1 2 38402 38410
0 38412 5 1 1 38411
0 38413 7 1 2 66513 38412
0 38414 5 1 1 38413
0 38415 7 1 2 75876 89682
0 38416 7 1 2 93890 38415
0 38417 5 1 1 38416
0 38418 7 1 2 38414 38417
0 38419 5 1 1 38418
0 38420 7 1 2 60139 38419
0 38421 5 1 1 38420
0 38422 7 1 2 79724 79810
0 38423 7 3 2 66006 89907
0 38424 7 3 2 57739 91828
0 38425 7 1 2 94024 94027
0 38426 7 1 2 38422 38425
0 38427 5 1 1 38426
0 38428 7 1 2 38421 38427
0 38429 5 1 1 38428
0 38430 7 1 2 58866 38429
0 38431 5 1 1 38430
0 38432 7 2 2 92559 94028
0 38433 7 2 2 70461 94030
0 38434 7 1 2 70783 79266
0 38435 7 1 2 94032 38434
0 38436 5 1 1 38435
0 38437 7 1 2 38431 38436
0 38438 5 1 1 38437
0 38439 7 1 2 57458 38438
0 38440 5 1 1 38439
0 38441 7 1 2 81260 92985
0 38442 7 1 2 93971 38441
0 38443 5 1 1 38442
0 38444 7 1 2 38440 38443
0 38445 5 1 1 38444
0 38446 7 1 2 71743 38445
0 38447 5 1 1 38446
0 38448 7 1 2 93721 94009
0 38449 5 1 1 38448
0 38450 7 1 2 61674 92578
0 38451 5 1 1 38450
0 38452 7 1 2 38449 38451
0 38453 5 1 1 38452
0 38454 7 1 2 58995 38453
0 38455 5 1 1 38454
0 38456 7 1 2 86997 87514
0 38457 5 1 1 38456
0 38458 7 1 2 38455 38457
0 38459 5 1 1 38458
0 38460 7 1 2 65068 38459
0 38461 5 1 1 38460
0 38462 7 1 2 70971 82569
0 38463 5 1 1 38462
0 38464 7 1 2 61026 38463
0 38465 5 1 1 38464
0 38466 7 1 2 86998 87339
0 38467 7 1 2 38465 38466
0 38468 5 1 1 38467
0 38469 7 1 2 63513 38468
0 38470 7 1 2 38461 38469
0 38471 5 1 1 38470
0 38472 7 1 2 74494 94005
0 38473 5 1 1 38472
0 38474 7 1 2 26977 38473
0 38475 5 1 1 38474
0 38476 7 1 2 57740 38475
0 38477 5 1 1 38476
0 38478 7 1 2 81602 91664
0 38479 5 1 1 38478
0 38480 7 1 2 58619 87536
0 38481 7 1 2 83253 38480
0 38482 5 1 1 38481
0 38483 7 1 2 38479 38482
0 38484 7 1 2 38477 38483
0 38485 5 1 1 38484
0 38486 7 1 2 64595 38485
0 38487 5 1 1 38486
0 38488 7 1 2 84245 81595
0 38489 5 1 1 38488
0 38490 7 1 2 82642 82570
0 38491 7 1 2 38489 38490
0 38492 5 1 1 38491
0 38493 7 1 2 58770 38492
0 38494 7 1 2 38487 38493
0 38495 5 1 1 38494
0 38496 7 1 2 38471 38495
0 38497 5 1 1 38496
0 38498 7 1 2 66514 38497
0 38499 5 1 1 38498
0 38500 7 1 2 73284 87047
0 38501 5 1 1 38500
0 38502 7 2 2 59145 73564
0 38503 7 1 2 78321 94034
0 38504 5 1 1 38503
0 38505 7 1 2 38501 38504
0 38506 5 1 1 38505
0 38507 7 1 2 93891 38506
0 38508 5 1 1 38507
0 38509 7 1 2 93893 38508
0 38510 5 1 1 38509
0 38511 7 1 2 82530 38510
0 38512 5 1 1 38511
0 38513 7 1 2 77962 93895
0 38514 5 1 1 38513
0 38515 7 4 2 58771 59880
0 38516 5 2 1 94036
0 38517 7 2 2 61675 94037
0 38518 7 1 2 70935 86999
0 38519 7 1 2 94042 38518
0 38520 5 1 1 38519
0 38521 7 1 2 61865 38520
0 38522 7 1 2 38514 38521
0 38523 7 1 2 38512 38522
0 38524 5 1 1 38523
0 38525 7 1 2 60140 38524
0 38526 7 1 2 38499 38525
0 38527 5 1 1 38526
0 38528 7 1 2 80040 79811
0 38529 7 1 2 94031 38528
0 38530 5 1 1 38529
0 38531 7 1 2 38527 38530
0 38532 5 1 1 38531
0 38533 7 1 2 58867 38532
0 38534 5 1 1 38533
0 38535 7 2 2 69878 89296
0 38536 7 1 2 74896 94044
0 38537 7 1 2 94033 38536
0 38538 5 1 1 38537
0 38539 7 1 2 61959 38538
0 38540 7 1 2 38534 38539
0 38541 7 1 2 38447 38540
0 38542 5 1 1 38541
0 38543 7 1 2 66714 38542
0 38544 7 1 2 38396 38543
0 38545 5 1 1 38544
0 38546 7 1 2 38222 38545
0 38547 5 1 1 38546
0 38548 7 1 2 67357 38547
0 38549 5 1 1 38548
0 38550 7 1 2 57741 73442
0 38551 5 4 1 38550
0 38552 7 2 2 73957 94046
0 38553 5 1 1 94050
0 38554 7 1 2 65069 38553
0 38555 5 1 1 38554
0 38556 7 1 2 73333 38555
0 38557 5 1 1 38556
0 38558 7 1 2 68628 38557
0 38559 5 1 1 38558
0 38560 7 1 2 71830 72049
0 38561 5 1 1 38560
0 38562 7 1 2 91151 38561
0 38563 5 1 1 38562
0 38564 7 1 2 70830 38563
0 38565 5 1 1 38564
0 38566 7 1 2 66007 38565
0 38567 5 1 1 38566
0 38568 7 1 2 68782 73443
0 38569 5 1 1 38568
0 38570 7 1 2 86277 38569
0 38571 5 1 1 38570
0 38572 7 1 2 57742 38571
0 38573 5 1 1 38572
0 38574 7 1 2 38567 38573
0 38575 7 1 2 38559 38574
0 38576 5 1 1 38575
0 38577 7 2 2 83561 89320
0 38578 7 4 2 59377 86314
0 38579 7 1 2 82412 94054
0 38580 7 1 2 94052 38579
0 38581 7 1 2 38576 38580
0 38582 5 1 1 38581
0 38583 7 1 2 38549 38582
0 38584 7 1 2 38214 38583
0 38585 5 1 1 38584
0 38586 7 1 2 71509 38585
0 38587 5 1 1 38586
0 38588 7 1 2 67358 93588
0 38589 5 2 1 38588
0 38590 7 3 2 72031 94058
0 38591 5 1 1 94060
0 38592 7 1 2 80400 94061
0 38593 5 1 1 38592
0 38594 7 1 2 63075 93612
0 38595 7 1 2 13064 38594
0 38596 7 1 2 93050 38595
0 38597 5 1 1 38596
0 38598 7 1 2 63373 38597
0 38599 5 1 1 38598
0 38600 7 1 2 38593 38599
0 38601 5 1 1 38600
0 38602 7 1 2 59629 38601
0 38603 5 1 1 38602
0 38604 7 1 2 64382 94059
0 38605 5 1 1 38604
0 38606 7 2 2 67774 79087
0 38607 5 3 1 94063
0 38608 7 1 2 65661 84553
0 38609 5 1 1 38608
0 38610 7 1 2 92962 38609
0 38611 5 1 1 38610
0 38612 7 1 2 80496 85368
0 38613 7 1 2 92660 38612
0 38614 7 1 2 38611 38613
0 38615 7 2 2 94065 38614
0 38616 5 1 1 94068
0 38617 7 1 2 38605 94069
0 38618 5 1 1 38617
0 38619 7 1 2 91850 38618
0 38620 5 2 1 38619
0 38621 7 2 2 85046 72874
0 38622 5 1 1 94072
0 38623 7 1 2 83254 94073
0 38624 5 1 1 38623
0 38625 7 1 2 94070 38624
0 38626 7 1 2 38603 38625
0 38627 5 1 1 38626
0 38628 7 1 2 66515 38627
0 38629 5 1 1 38628
0 38630 7 1 2 71906 85747
0 38631 5 1 1 38630
0 38632 7 1 2 78322 80328
0 38633 5 1 1 38632
0 38634 7 1 2 38631 38633
0 38635 5 1 1 38634
0 38636 7 1 2 86293 89497
0 38637 7 1 2 38635 38636
0 38638 5 1 1 38637
0 38639 7 1 2 38629 38638
0 38640 5 1 1 38639
0 38641 7 1 2 66295 38640
0 38642 5 1 1 38641
0 38643 7 1 2 68027 80057
0 38644 5 1 1 38643
0 38645 7 1 2 63374 38644
0 38646 5 1 1 38645
0 38647 7 1 2 71195 89658
0 38648 7 1 2 38646 38647
0 38649 5 1 1 38648
0 38650 7 1 2 38642 38649
0 38651 5 1 1 38650
0 38652 7 1 2 59881 38651
0 38653 5 1 1 38652
0 38654 7 1 2 64596 83255
0 38655 5 1 1 38654
0 38656 7 1 2 72394 91748
0 38657 5 2 1 38656
0 38658 7 1 2 38655 94074
0 38659 5 1 1 38658
0 38660 7 1 2 82444 38659
0 38661 5 1 1 38660
0 38662 7 1 2 77830 38661
0 38663 5 1 1 38662
0 38664 7 2 2 71196 38663
0 38665 5 1 1 94076
0 38666 7 1 2 89908 94077
0 38667 5 1 1 38666
0 38668 7 1 2 38653 38667
0 38669 5 1 1 38668
0 38670 7 1 2 63514 38669
0 38671 5 1 1 38670
0 38672 7 1 2 80566 72287
0 38673 7 1 2 86380 38672
0 38674 7 1 2 89751 38673
0 38675 7 1 2 80058 38674
0 38676 5 1 1 38675
0 38677 7 1 2 38671 38676
0 38678 5 1 1 38677
0 38679 7 1 2 60028 38678
0 38680 5 1 1 38679
0 38681 7 1 2 63515 83256
0 38682 5 2 1 38681
0 38683 7 1 2 94075 94078
0 38684 5 1 1 38683
0 38685 7 3 2 86960 89429
0 38686 5 1 1 94080
0 38687 7 2 2 83048 83349
0 38688 7 1 2 94081 94083
0 38689 7 1 2 38684 38688
0 38690 5 1 1 38689
0 38691 7 1 2 70216 92823
0 38692 5 1 1 38691
0 38693 7 1 2 80739 73130
0 38694 5 1 1 38693
0 38695 7 2 2 38692 38694
0 38696 5 1 1 94085
0 38697 7 1 2 64383 38696
0 38698 5 1 1 38697
0 38699 7 3 2 63912 78766
0 38700 5 2 1 94087
0 38701 7 1 2 81173 94090
0 38702 5 1 1 38701
0 38703 7 1 2 72942 38702
0 38704 5 1 1 38703
0 38705 7 1 2 63785 69399
0 38706 7 1 2 68200 38705
0 38707 7 1 2 81145 38706
0 38708 5 1 1 38707
0 38709 7 1 2 38704 38708
0 38710 5 1 1 38709
0 38711 7 1 2 62501 38710
0 38712 5 1 1 38711
0 38713 7 1 2 38698 38712
0 38714 5 1 1 38713
0 38715 7 1 2 62771 38714
0 38716 5 1 1 38715
0 38717 7 1 2 92831 38716
0 38718 5 1 1 38717
0 38719 7 1 2 63076 38718
0 38720 5 1 1 38719
0 38721 7 2 2 77993 83590
0 38722 7 1 2 78460 94092
0 38723 5 1 1 38722
0 38724 7 2 2 38720 38723
0 38725 5 1 1 94094
0 38726 7 1 2 64597 38725
0 38727 5 1 1 38726
0 38728 7 1 2 77482 92383
0 38729 5 1 1 38728
0 38730 7 2 2 71510 38729
0 38731 5 1 1 94096
0 38732 7 2 2 84928 75907
0 38733 7 1 2 38731 94098
0 38734 5 1 1 38733
0 38735 7 1 2 70831 78351
0 38736 7 1 2 84376 38735
0 38737 5 1 1 38736
0 38738 7 1 2 71438 5838
0 38739 5 1 1 38738
0 38740 7 1 2 71306 81860
0 38741 7 2 2 84285 38740
0 38742 7 1 2 78228 94100
0 38743 5 1 1 38742
0 38744 7 1 2 38739 38743
0 38745 7 3 2 38737 38744
0 38746 5 1 1 94102
0 38747 7 2 2 38734 94103
0 38748 7 1 2 68253 85697
0 38749 5 1 1 38748
0 38750 7 1 2 82846 38749
0 38751 5 3 1 38750
0 38752 7 1 2 78870 94107
0 38753 5 1 1 38752
0 38754 7 2 2 71307 67880
0 38755 5 1 1 94110
0 38756 7 4 2 84382 38755
0 38757 5 1 1 94112
0 38758 7 1 2 38753 94113
0 38759 5 1 1 38758
0 38760 7 1 2 60636 38759
0 38761 5 1 1 38760
0 38762 7 1 2 71511 25698
0 38763 5 1 1 38762
0 38764 7 1 2 71308 69892
0 38765 7 1 2 38763 38764
0 38766 5 1 1 38765
0 38767 7 1 2 71439 14505
0 38768 5 1 1 38767
0 38769 7 1 2 71309 93394
0 38770 5 1 1 38769
0 38771 7 1 2 38768 38770
0 38772 7 3 2 38766 38771
0 38773 5 1 1 94116
0 38774 7 1 2 38761 94117
0 38775 5 2 1 38774
0 38776 7 1 2 61027 94119
0 38777 5 1 1 38776
0 38778 7 1 2 94105 38777
0 38779 5 1 1 38778
0 38780 7 1 2 64598 38779
0 38781 5 1 1 38780
0 38782 7 2 2 78603 78451
0 38783 5 1 1 94121
0 38784 7 1 2 64384 87068
0 38785 7 1 2 94122 38784
0 38786 5 1 1 38785
0 38787 7 1 2 38781 38786
0 38788 5 1 1 38787
0 38789 7 1 2 61384 38788
0 38790 5 1 1 38789
0 38791 7 1 2 60029 38790
0 38792 7 1 2 38727 38791
0 38793 5 1 1 38792
0 38794 7 1 2 64385 83257
0 38795 5 1 1 38794
0 38796 7 1 2 65297 94062
0 38797 5 1 1 38796
0 38798 7 1 2 38795 38797
0 38799 5 1 1 38798
0 38800 7 1 2 64386 85041
0 38801 5 1 1 38800
0 38802 7 1 2 61385 38801
0 38803 7 1 2 38799 38802
0 38804 5 1 1 38803
0 38805 7 1 2 94071 38804
0 38806 5 1 1 38805
0 38807 7 1 2 59882 38806
0 38808 5 1 1 38807
0 38809 7 1 2 64722 38665
0 38810 7 1 2 38808 38809
0 38811 5 1 1 38810
0 38812 7 1 2 66516 38811
0 38813 7 1 2 38793 38812
0 38814 5 1 1 38813
0 38815 7 1 2 70832 82338
0 38816 5 1 1 38815
0 38817 7 1 2 8097 87061
0 38818 5 1 1 38817
0 38819 7 2 2 58063 38818
0 38820 5 1 1 94123
0 38821 7 1 2 38816 94124
0 38822 5 1 1 38821
0 38823 7 1 2 82632 73430
0 38824 5 1 1 38823
0 38825 7 1 2 38822 38824
0 38826 5 1 1 38825
0 38827 7 1 2 78323 38826
0 38828 5 1 1 38827
0 38829 7 1 2 82339 38820
0 38830 5 1 1 38829
0 38831 7 1 2 78208 38830
0 38832 5 1 1 38831
0 38833 7 1 2 13011 38832
0 38834 5 1 1 38833
0 38835 7 1 2 71907 38834
0 38836 5 1 1 38835
0 38837 7 1 2 38828 38836
0 38838 5 1 1 38837
0 38839 7 1 2 93305 38838
0 38840 5 1 1 38839
0 38841 7 1 2 78908 86169
0 38842 5 1 1 38841
0 38843 7 1 2 91851 38842
0 38844 5 1 1 38843
0 38845 7 1 2 64387 86784
0 38846 5 1 1 38845
0 38847 7 1 2 65298 38846
0 38848 5 1 1 38847
0 38849 7 1 2 58064 86182
0 38850 5 1 1 38849
0 38851 7 1 2 57743 69909
0 38852 5 1 1 38851
0 38853 7 2 2 60637 67214
0 38854 5 2 1 94125
0 38855 7 1 2 74026 94126
0 38856 5 1 1 38855
0 38857 7 1 2 58333 38856
0 38858 5 1 1 38857
0 38859 7 1 2 38852 38858
0 38860 7 1 2 38850 38859
0 38861 7 1 2 38848 38860
0 38862 5 1 1 38861
0 38863 7 3 2 65299 93601
0 38864 5 1 1 94129
0 38865 7 1 2 59630 38864
0 38866 5 1 1 38865
0 38867 7 1 2 73635 38866
0 38868 7 1 2 38862 38867
0 38869 5 1 1 38868
0 38870 7 1 2 38844 38869
0 38871 5 1 1 38870
0 38872 7 1 2 59883 38871
0 38873 5 1 1 38872
0 38874 7 1 2 73876 93356
0 38875 5 1 1 38874
0 38876 7 1 2 61028 93512
0 38877 5 1 1 38876
0 38878 7 1 2 38875 38877
0 38879 5 1 1 38878
0 38880 7 1 2 75877 37284
0 38881 7 1 2 38879 38880
0 38882 5 1 1 38881
0 38883 7 1 2 80064 83970
0 38884 5 1 1 38883
0 38885 7 2 2 71197 77827
0 38886 5 2 1 94132
0 38887 7 1 2 38884 94134
0 38888 7 1 2 38882 38887
0 38889 7 1 2 38873 38888
0 38890 5 1 1 38889
0 38891 7 1 2 60030 38890
0 38892 5 1 1 38891
0 38893 7 1 2 38840 38892
0 38894 5 1 1 38893
0 38895 7 1 2 61866 38894
0 38896 5 1 1 38895
0 38897 7 1 2 68396 29621
0 38898 5 1 1 38897
0 38899 7 1 2 67215 38898
0 38900 5 1 1 38899
0 38901 7 1 2 65662 38900
0 38902 5 1 1 38901
0 38903 7 1 2 63077 38902
0 38904 5 1 1 38903
0 38905 7 1 2 88792 38904
0 38906 5 1 1 38905
0 38907 7 1 2 69998 93727
0 38908 5 1 1 38907
0 38909 7 2 2 65070 75337
0 38910 5 1 1 94136
0 38911 7 1 2 70003 38910
0 38912 5 1 1 38911
0 38913 7 1 2 88803 38912
0 38914 5 1 1 38913
0 38915 7 1 2 38908 38914
0 38916 7 1 2 38906 38915
0 38917 5 1 1 38916
0 38918 7 1 2 73838 38917
0 38919 5 1 1 38918
0 38920 7 1 2 62772 35569
0 38921 5 1 1 38920
0 38922 7 1 2 77155 67872
0 38923 5 1 1 38922
0 38924 7 1 2 60638 70124
0 38925 7 1 2 38923 38924
0 38926 5 1 1 38925
0 38927 7 1 2 69796 2341
0 38928 5 1 1 38927
0 38929 7 1 2 68783 83935
0 38930 5 1 1 38929
0 38931 7 1 2 64097 38930
0 38932 7 1 2 38928 38931
0 38933 5 1 1 38932
0 38934 7 1 2 38926 38933
0 38935 7 1 2 38921 38934
0 38936 5 1 1 38935
0 38937 7 1 2 93139 38936
0 38938 5 1 1 38937
0 38939 7 2 2 78490 91993
0 38940 5 1 1 94138
0 38941 7 1 2 59884 38940
0 38942 5 1 1 38941
0 38943 7 1 2 69053 38942
0 38944 5 1 1 38943
0 38945 7 1 2 64599 87387
0 38946 5 1 1 38945
0 38947 7 1 2 66008 30191
0 38948 5 1 1 38947
0 38949 7 1 2 92796 38948
0 38950 5 1 1 38949
0 38951 7 1 2 38946 38950
0 38952 7 1 2 38944 38951
0 38953 5 1 1 38952
0 38954 7 1 2 67216 38953
0 38955 5 1 1 38954
0 38956 7 1 2 38938 38955
0 38957 5 1 1 38956
0 38958 7 1 2 61029 38957
0 38959 5 1 1 38958
0 38960 7 1 2 61030 93528
0 38961 5 1 1 38960
0 38962 7 1 2 59885 38961
0 38963 5 1 1 38962
0 38964 7 1 2 85670 38963
0 38965 5 1 1 38964
0 38966 7 1 2 76378 93140
0 38967 7 1 2 93856 38966
0 38968 5 1 1 38967
0 38969 7 1 2 58334 91484
0 38970 5 1 1 38969
0 38971 7 1 2 59886 72908
0 38972 5 7 1 38971
0 38973 7 1 2 85571 94140
0 38974 7 1 2 38970 38973
0 38975 5 1 1 38974
0 38976 7 1 2 38968 38975
0 38977 7 1 2 38965 38976
0 38978 7 1 2 62246 79125
0 38979 5 2 1 38978
0 38980 7 1 2 80049 94147
0 38981 5 1 1 38980
0 38982 7 1 2 62502 38981
0 38983 5 1 1 38982
0 38984 7 4 2 92820 38983
0 38985 5 7 1 94149
0 38986 7 1 2 84637 90928
0 38987 5 2 1 38986
0 38988 7 1 2 85426 94160
0 38989 5 1 1 38988
0 38990 7 3 2 62773 80672
0 38991 5 2 1 94162
0 38992 7 1 2 71310 94163
0 38993 5 1 1 38992
0 38994 7 1 2 85435 38993
0 38995 7 1 2 38989 38994
0 38996 5 1 1 38995
0 38997 7 1 2 94153 38996
0 38998 5 1 1 38997
0 38999 7 3 2 86909 30883
0 39000 5 2 1 94167
0 39001 7 1 2 85427 94168
0 39002 5 1 1 39001
0 39003 7 1 2 85432 78749
0 39004 5 1 1 39003
0 39005 7 1 2 39002 39004
0 39006 5 1 1 39005
0 39007 7 1 2 83954 39006
0 39008 5 1 1 39007
0 39009 7 1 2 38998 39008
0 39010 7 1 2 38977 39009
0 39011 7 1 2 38959 39010
0 39012 5 1 1 39011
0 39013 7 1 2 88675 39012
0 39014 5 1 1 39013
0 39015 7 1 2 38919 39014
0 39016 5 1 1 39015
0 39017 7 1 2 63375 39016
0 39018 5 1 1 39017
0 39019 7 1 2 66296 39018
0 39020 7 1 2 38896 39019
0 39021 7 1 2 38814 39020
0 39022 5 1 1 39021
0 39023 7 1 2 86584 81304
0 39024 5 1 1 39023
0 39025 7 1 2 76764 39024
0 39026 5 2 1 39025
0 39027 7 1 2 78593 94172
0 39028 5 1 1 39027
0 39029 7 2 2 61031 91564
0 39030 5 1 1 94174
0 39031 7 1 2 86585 94175
0 39032 5 1 1 39031
0 39033 7 1 2 39028 39032
0 39034 5 1 1 39033
0 39035 7 1 2 73692 39034
0 39036 5 1 1 39035
0 39037 7 1 2 84743 91371
0 39038 7 1 2 86350 39037
0 39039 5 1 1 39038
0 39040 7 1 2 39036 39039
0 39041 5 1 1 39040
0 39042 7 1 2 67775 39041
0 39043 5 1 1 39042
0 39044 7 1 2 78177 93432
0 39045 5 4 1 39044
0 39046 7 1 2 68397 94176
0 39047 5 1 1 39046
0 39048 7 1 2 33091 39047
0 39049 5 1 1 39048
0 39050 7 1 2 65663 39049
0 39051 5 1 1 39050
0 39052 7 1 2 86921 93703
0 39053 5 1 1 39052
0 39054 7 1 2 91852 39053
0 39055 5 1 1 39054
0 39056 7 1 2 64600 82911
0 39057 7 1 2 39055 39056
0 39058 7 1 2 39051 39057
0 39059 5 1 1 39058
0 39060 7 1 2 85665 85876
0 39061 5 3 1 39060
0 39062 7 1 2 93842 94180
0 39063 5 1 1 39062
0 39064 7 2 2 58620 93288
0 39065 5 1 1 94183
0 39066 7 1 2 85653 94184
0 39067 5 1 1 39066
0 39068 7 1 2 90013 39067
0 39069 5 1 1 39068
0 39070 7 1 2 39063 39069
0 39071 5 1 1 39070
0 39072 7 1 2 81951 39071
0 39073 5 1 1 39072
0 39074 7 2 2 76259 84638
0 39075 5 3 1 94185
0 39076 7 1 2 78594 94187
0 39077 5 1 1 39076
0 39078 7 1 2 39030 39077
0 39079 5 1 1 39078
0 39080 7 1 2 85879 39079
0 39081 5 1 1 39080
0 39082 7 1 2 85483 93093
0 39083 5 1 1 39082
0 39084 7 1 2 39081 39083
0 39085 5 1 1 39084
0 39086 7 1 2 67776 39085
0 39087 5 1 1 39086
0 39088 7 3 2 63078 73131
0 39089 5 1 1 94190
0 39090 7 1 2 58621 39089
0 39091 5 1 1 39090
0 39092 7 1 2 77677 39091
0 39093 5 1 1 39092
0 39094 7 1 2 70246 83466
0 39095 5 1 1 39094
0 39096 7 1 2 87076 39095
0 39097 7 1 2 39093 39096
0 39098 5 1 1 39097
0 39099 7 1 2 73693 39098
0 39100 5 1 1 39099
0 39101 7 1 2 76267 77678
0 39102 5 1 1 39101
0 39103 7 1 2 70217 83780
0 39104 5 1 1 39103
0 39105 7 1 2 39102 39104
0 39106 5 1 1 39105
0 39107 7 1 2 85880 39106
0 39108 5 1 1 39107
0 39109 7 1 2 59887 26983
0 39110 7 1 2 39108 39109
0 39111 7 1 2 39100 39110
0 39112 7 1 2 39087 39111
0 39113 7 1 2 39073 39112
0 39114 5 1 1 39113
0 39115 7 1 2 39059 39114
0 39116 5 1 1 39115
0 39117 7 1 2 39043 39116
0 39118 5 1 1 39117
0 39119 7 1 2 66517 39118
0 39120 5 1 1 39119
0 39121 7 1 2 86294 89239
0 39122 5 1 1 39121
0 39123 7 1 2 39120 39122
0 39124 5 1 1 39123
0 39125 7 1 2 60031 39124
0 39126 5 1 1 39125
0 39127 7 1 2 61676 38686
0 39128 7 1 2 39126 39127
0 39129 5 1 1 39128
0 39130 7 1 2 58772 39129
0 39131 7 1 2 39022 39130
0 39132 5 1 1 39131
0 39133 7 1 2 38690 39132
0 39134 7 1 2 38680 39133
0 39135 5 1 1 39134
0 39136 7 1 2 60141 39135
0 39137 5 1 1 39136
0 39138 7 1 2 71589 89909
0 39139 7 2 2 92582 39138
0 39140 5 1 1 94193
0 39141 7 3 2 57744 76857
0 39142 7 1 2 70175 94195
0 39143 7 1 2 94194 39142
0 39144 5 1 1 39143
0 39145 7 1 2 39137 39144
0 39146 5 1 1 39145
0 39147 7 1 2 58868 39146
0 39148 5 1 1 39147
0 39149 7 3 2 82275 77370
0 39150 7 1 2 80460 74761
0 39151 7 3 2 94198 39150
0 39152 7 1 2 73937 80059
0 39153 5 1 1 39152
0 39154 7 1 2 68028 79801
0 39155 5 1 1 39154
0 39156 7 1 2 39153 39155
0 39157 5 1 1 39156
0 39158 7 2 2 89910 39157
0 39159 7 1 2 94201 94204
0 39160 5 1 1 39159
0 39161 7 4 2 79812 80755
0 39162 5 1 1 94206
0 39163 7 1 2 94207 94205
0 39164 5 1 1 39163
0 39165 7 3 2 60032 78085
0 39166 7 1 2 86108 94210
0 39167 5 1 1 39166
0 39168 7 1 2 65071 79272
0 39169 5 1 1 39168
0 39170 7 1 2 78491 69324
0 39171 5 4 1 39170
0 39172 7 1 2 39169 94213
0 39173 5 1 1 39172
0 39174 7 3 2 64723 76690
0 39175 5 3 1 94217
0 39176 7 1 2 71198 94220
0 39177 7 1 2 39173 39176
0 39178 5 1 1 39177
0 39179 7 1 2 39167 39178
0 39180 5 1 1 39179
0 39181 7 1 2 68029 39180
0 39182 5 1 1 39181
0 39183 7 3 2 60033 72846
0 39184 7 1 2 92882 94223
0 39185 5 1 1 39184
0 39186 7 1 2 39182 39185
0 39187 5 1 1 39186
0 39188 7 1 2 58773 39187
0 39189 5 1 1 39188
0 39190 7 1 2 9697 94214
0 39191 5 1 1 39190
0 39192 7 2 2 60034 39191
0 39193 7 1 2 83828 94055
0 39194 7 1 2 94226 39193
0 39195 5 1 1 39194
0 39196 7 1 2 39189 39195
0 39197 5 1 1 39196
0 39198 7 1 2 66297 39197
0 39199 5 1 1 39198
0 39200 7 1 2 69461 89388
0 39201 5 1 1 39200
0 39202 7 1 2 77364 94215
0 39203 5 1 1 39202
0 39204 7 1 2 71199 39203
0 39205 5 1 1 39204
0 39206 7 6 2 75576 94141
0 39207 7 2 2 65072 94228
0 39208 5 1 1 94234
0 39209 7 1 2 39205 39208
0 39210 5 1 1 39209
0 39211 7 1 2 59146 66298
0 39212 7 1 2 39210 39211
0 39213 5 1 1 39212
0 39214 7 1 2 39201 39213
0 39215 5 1 1 39214
0 39216 7 1 2 57745 39215
0 39217 5 1 1 39216
0 39218 7 1 2 80050 89356
0 39219 5 1 1 39218
0 39220 7 1 2 39217 39219
0 39221 5 1 1 39220
0 39222 7 1 2 60035 39221
0 39223 5 1 1 39222
0 39224 7 1 2 2263 94216
0 39225 5 1 1 39224
0 39226 7 6 2 66299 73839
0 39227 7 2 2 92018 94236
0 39228 7 1 2 39225 94242
0 39229 5 1 1 39228
0 39230 7 1 2 39223 39229
0 39231 5 1 1 39230
0 39232 7 1 2 58774 39231
0 39233 5 1 1 39232
0 39234 7 1 2 94227 94243
0 39235 5 1 1 39234
0 39236 7 1 2 39233 39235
0 39237 5 1 1 39236
0 39238 7 1 2 67359 39237
0 39239 5 1 1 39238
0 39240 7 1 2 39199 39239
0 39241 5 1 1 39240
0 39242 7 1 2 65664 39241
0 39243 5 1 1 39242
0 39244 7 3 2 67675 90348
0 39245 7 2 2 81793 94244
0 39246 5 1 1 94247
0 39247 7 1 2 93484 94224
0 39248 7 1 2 94248 39247
0 39249 5 1 1 39248
0 39250 7 1 2 61867 39249
0 39251 7 1 2 39243 39250
0 39252 5 1 1 39251
0 39253 7 1 2 59147 79802
0 39254 5 1 1 39253
0 39255 7 1 2 79091 39254
0 39256 5 1 1 39255
0 39257 7 1 2 63516 39256
0 39258 5 1 1 39257
0 39259 7 2 2 75227 87060
0 39260 7 1 2 59148 94249
0 39261 5 1 1 39260
0 39262 7 1 2 39258 39261
0 39263 5 1 1 39262
0 39264 7 1 2 58065 39263
0 39265 5 1 1 39264
0 39266 7 1 2 75810 93181
0 39267 5 1 1 39266
0 39268 7 1 2 39265 39267
0 39269 5 1 1 39268
0 39270 7 1 2 92205 39269
0 39271 5 1 1 39270
0 39272 7 1 2 86381 94250
0 39273 5 1 1 39272
0 39274 7 3 2 80982 94142
0 39275 7 2 2 73877 94251
0 39276 5 1 1 94254
0 39277 7 1 2 69462 94255
0 39278 5 1 1 39277
0 39279 7 1 2 39273 39278
0 39280 5 1 1 39279
0 39281 7 1 2 59149 39280
0 39282 5 1 1 39281
0 39283 7 2 2 34411 93874
0 39284 5 2 1 94256
0 39285 7 1 2 39276 94257
0 39286 5 1 1 39285
0 39287 7 2 2 76351 39286
0 39288 5 1 1 94260
0 39289 7 1 2 39282 39288
0 39290 5 1 1 39289
0 39291 7 1 2 66922 39290
0 39292 5 1 1 39291
0 39293 7 1 2 39271 39292
0 39294 5 1 1 39293
0 39295 7 1 2 57746 39294
0 39296 5 1 1 39295
0 39297 7 1 2 69006 73490
0 39298 5 1 1 39297
0 39299 7 1 2 2976 39298
0 39300 5 1 1 39299
0 39301 7 1 2 58066 39300
0 39302 5 1 1 39301
0 39303 7 1 2 82004 71344
0 39304 5 1 1 39303
0 39305 7 1 2 39302 39304
0 39306 5 1 1 39305
0 39307 7 1 2 81058 39306
0 39308 5 1 1 39307
0 39309 7 1 2 79803 94258
0 39310 5 1 1 39309
0 39311 7 1 2 59150 94261
0 39312 5 1 1 39311
0 39313 7 1 2 39310 39312
0 39314 5 1 1 39313
0 39315 7 1 2 66923 39314
0 39316 5 1 1 39315
0 39317 7 1 2 39308 39316
0 39318 7 1 2 39296 39317
0 39319 5 1 1 39318
0 39320 7 1 2 66300 39319
0 39321 5 1 1 39320
0 39322 7 1 2 79456 93937
0 39323 5 1 1 39322
0 39324 7 1 2 88039 39323
0 39325 5 1 1 39324
0 39326 7 1 2 85356 87412
0 39327 7 1 2 39325 39326
0 39328 5 1 1 39327
0 39329 7 1 2 78098 82813
0 39330 5 1 1 39329
0 39331 7 2 2 79571 93430
0 39332 5 1 1 94262
0 39333 7 1 2 39330 39332
0 39334 7 1 2 39328 39333
0 39335 5 1 1 39334
0 39336 7 1 2 76568 81507
0 39337 7 1 2 39335 39336
0 39338 5 1 1 39337
0 39339 7 1 2 66518 39338
0 39340 7 1 2 39321 39339
0 39341 5 1 1 39340
0 39342 7 1 2 60142 39341
0 39343 7 1 2 39252 39342
0 39344 5 1 1 39343
0 39345 7 1 2 39164 39344
0 39346 5 1 1 39345
0 39347 7 1 2 58869 39346
0 39348 5 1 1 39347
0 39349 7 1 2 39160 39348
0 39350 5 1 1 39349
0 39351 7 1 2 57459 39350
0 39352 5 1 1 39351
0 39353 7 1 2 74524 81563
0 39354 5 2 1 39353
0 39355 7 1 2 87544 94264
0 39356 5 1 1 39355
0 39357 7 1 2 58067 39356
0 39358 5 1 1 39357
0 39359 7 2 2 66301 92809
0 39360 7 1 2 64724 94266
0 39361 5 1 1 39360
0 39362 7 1 2 39358 39361
0 39363 5 1 1 39362
0 39364 7 1 2 57747 39363
0 39365 5 1 1 39364
0 39366 7 1 2 65665 590
0 39367 5 1 1 39366
0 39368 7 1 2 78258 93503
0 39369 7 1 2 39367 39368
0 39370 5 1 1 39369
0 39371 7 2 2 66302 39370
0 39372 7 1 2 64725 94268
0 39373 5 1 1 39372
0 39374 7 1 2 39365 39373
0 39375 5 1 1 39374
0 39376 7 1 2 93306 39375
0 39377 5 1 1 39376
0 39378 7 1 2 58068 69463
0 39379 5 2 1 39378
0 39380 7 1 2 67360 87799
0 39381 5 1 1 39380
0 39382 7 1 2 94270 39381
0 39383 7 1 2 86185 39382
0 39384 5 1 1 39383
0 39385 7 1 2 82957 39384
0 39386 5 1 1 39385
0 39387 7 1 2 93377 39386
0 39388 5 1 1 39387
0 39389 7 1 2 85698 93602
0 39390 5 1 1 39389
0 39391 7 1 2 60405 93584
0 39392 5 1 1 39391
0 39393 7 1 2 39390 39392
0 39394 5 1 1 39393
0 39395 7 1 2 65300 39394
0 39396 5 1 1 39395
0 39397 7 1 2 58996 83585
0 39398 5 1 1 39397
0 39399 7 1 2 83687 39398
0 39400 5 1 1 39399
0 39401 7 1 2 57460 39400
0 39402 5 1 1 39401
0 39403 7 1 2 63376 88422
0 39404 5 1 1 39403
0 39405 7 1 2 65666 39404
0 39406 7 1 2 39402 39405
0 39407 7 1 2 39396 39406
0 39408 5 1 1 39407
0 39409 7 2 2 68136 93292
0 39410 5 1 1 94272
0 39411 7 1 2 85125 93055
0 39412 7 1 2 39410 39411
0 39413 5 2 1 39412
0 39414 7 1 2 59631 94274
0 39415 5 1 1 39414
0 39416 7 1 2 67217 78215
0 39417 5 3 1 39416
0 39418 7 1 2 71908 94276
0 39419 5 1 1 39418
0 39420 7 1 2 72514 37232
0 39421 7 1 2 39419 39420
0 39422 5 1 1 39421
0 39423 7 1 2 71311 39422
0 39424 5 1 1 39423
0 39425 7 1 2 61032 39424
0 39426 7 1 2 39415 39425
0 39427 5 1 1 39426
0 39428 7 1 2 39408 39427
0 39429 5 1 1 39428
0 39430 7 1 2 68137 89076
0 39431 5 2 1 39430
0 39432 7 1 2 70428 93813
0 39433 7 1 2 94279 39432
0 39434 5 1 1 39433
0 39435 7 1 2 59632 93072
0 39436 7 1 2 39434 39435
0 39437 5 1 1 39436
0 39438 7 1 2 59888 77786
0 39439 7 1 2 39437 39438
0 39440 7 1 2 39429 39439
0 39441 5 1 1 39440
0 39442 7 1 2 39388 39441
0 39443 5 1 1 39442
0 39444 7 1 2 66303 39443
0 39445 5 1 1 39444
0 39446 7 1 2 57748 69477
0 39447 5 1 1 39446
0 39448 7 1 2 73886 78625
0 39449 7 1 2 79108 39448
0 39450 7 1 2 39447 39449
0 39451 5 1 1 39450
0 39452 7 1 2 76655 39451
0 39453 5 1 1 39452
0 39454 7 2 2 71200 73744
0 39455 7 1 2 86180 82370
0 39456 7 1 2 94281 39455
0 39457 5 1 1 39456
0 39458 7 1 2 61677 39457
0 39459 7 1 2 39453 39458
0 39460 5 1 1 39459
0 39461 7 1 2 60036 39460
0 39462 7 1 2 39445 39461
0 39463 5 1 1 39462
0 39464 7 1 2 39377 39463
0 39465 5 1 1 39464
0 39466 7 1 2 58775 39465
0 39467 5 1 1 39466
0 39468 7 5 2 63517 66304
0 39469 5 1 1 94283
0 39470 7 1 2 94265 39469
0 39471 5 1 1 39470
0 39472 7 1 2 58069 39471
0 39473 5 1 1 39472
0 39474 7 1 2 63518 94267
0 39475 5 1 1 39474
0 39476 7 1 2 39473 39475
0 39477 5 1 1 39476
0 39478 7 1 2 57749 39477
0 39479 5 1 1 39478
0 39480 7 1 2 63519 94269
0 39481 5 1 1 39480
0 39482 7 1 2 39479 39481
0 39483 5 1 1 39482
0 39484 7 1 2 87000 83829
0 39485 7 1 2 39483 39484
0 39486 5 1 1 39485
0 39487 7 1 2 39467 39486
0 39488 5 1 1 39487
0 39489 7 1 2 90115 39488
0 39490 5 1 1 39489
0 39491 7 2 2 57461 89659
0 39492 5 1 1 94288
0 39493 7 1 2 22385 39492
0 39494 5 1 1 39493
0 39495 7 1 2 93638 39494
0 39496 5 1 1 39495
0 39497 7 1 2 76352 91762
0 39498 5 1 1 39497
0 39499 7 1 2 39496 39498
0 39500 5 1 1 39499
0 39501 7 1 2 59889 39500
0 39502 5 1 1 39501
0 39503 7 1 2 86382 91612
0 39504 5 1 1 39503
0 39505 7 1 2 39502 39504
0 39506 5 1 1 39505
0 39507 7 1 2 66924 39506
0 39508 5 1 1 39507
0 39509 7 1 2 76097 94082
0 39510 5 1 1 39509
0 39511 7 3 2 58776 82958
0 39512 5 1 1 94290
0 39513 7 1 2 61868 84008
0 39514 7 1 2 69464 39513
0 39515 7 1 2 94291 39514
0 39516 5 1 1 39515
0 39517 7 1 2 39510 39516
0 39518 5 1 1 39517
0 39519 7 1 2 66305 39518
0 39520 5 1 1 39519
0 39521 7 1 2 60143 39520
0 39522 7 1 2 39508 39521
0 39523 5 1 1 39522
0 39524 7 1 2 64824 39140
0 39525 5 1 1 39524
0 39526 7 1 2 58870 39525
0 39527 7 1 2 39523 39526
0 39528 5 1 1 39527
0 39529 7 2 2 59633 77371
0 39530 7 4 2 90259 94293
0 39531 7 3 2 58622 76110
0 39532 7 2 2 71590 94299
0 39533 7 1 2 66519 94302
0 39534 7 1 2 94295 39533
0 39535 5 1 1 39534
0 39536 7 1 2 39528 39535
0 39537 5 1 1 39536
0 39538 7 1 2 74717 39537
0 39539 5 1 1 39538
0 39540 7 1 2 76060 81054
0 39541 5 1 1 39540
0 39542 7 1 2 39162 39541
0 39543 5 1 1 39542
0 39544 7 1 2 93493 39543
0 39545 5 1 1 39544
0 39546 7 1 2 93302 93363
0 39547 5 1 1 39546
0 39548 7 1 2 76301 93357
0 39549 5 1 1 39548
0 39550 7 1 2 67361 77807
0 39551 5 1 1 39550
0 39552 7 1 2 39549 39551
0 39553 7 1 2 39547 39552
0 39554 5 1 1 39553
0 39555 7 1 2 85313 39554
0 39556 5 1 1 39555
0 39557 7 1 2 39545 39556
0 39558 5 1 1 39557
0 39559 7 1 2 58871 39558
0 39560 5 1 1 39559
0 39561 7 1 2 93494 94202
0 39562 5 1 1 39561
0 39563 7 1 2 39560 39562
0 39564 5 1 1 39563
0 39565 7 1 2 65667 39564
0 39566 5 1 1 39565
0 39567 7 1 2 78374 92777
0 39568 5 3 1 39567
0 39569 7 1 2 63079 94304
0 39570 5 1 1 39569
0 39571 7 1 2 68138 94154
0 39572 5 1 1 39571
0 39573 7 1 2 67362 85961
0 39574 5 1 1 39573
0 39575 7 1 2 86910 39574
0 39576 5 1 1 39575
0 39577 7 2 2 39572 39576
0 39578 5 2 1 94307
0 39579 7 1 2 39570 94308
0 39580 5 1 1 39579
0 39581 7 2 2 61033 39580
0 39582 5 1 1 94311
0 39583 7 1 2 76219 94155
0 39584 5 1 1 39583
0 39585 7 1 2 80880 86916
0 39586 5 1 1 39585
0 39587 7 1 2 68139 39586
0 39588 5 1 1 39587
0 39589 7 1 2 39584 39588
0 39590 7 1 2 39582 39589
0 39591 5 1 1 39590
0 39592 7 1 2 59634 39591
0 39593 5 1 1 39592
0 39594 7 1 2 85349 4067
0 39595 5 1 1 39594
0 39596 7 3 2 58997 74993
0 39597 7 1 2 64388 94313
0 39598 5 1 1 39597
0 39599 7 1 2 83688 39598
0 39600 5 1 1 39599
0 39601 7 1 2 39595 39600
0 39602 5 1 1 39601
0 39603 7 1 2 77994 35304
0 39604 5 1 1 39603
0 39605 7 1 2 63080 93695
0 39606 5 1 1 39605
0 39607 7 1 2 63377 39606
0 39608 5 1 1 39607
0 39609 7 1 2 39604 39608
0 39610 7 1 2 39602 39609
0 39611 7 1 2 39593 39610
0 39612 5 1 1 39611
0 39613 7 1 2 85314 90312
0 39614 7 1 2 39612 39613
0 39615 5 1 1 39614
0 39616 7 1 2 39566 39615
0 39617 5 1 1 39616
0 39618 7 1 2 66306 39617
0 39619 5 1 1 39618
0 39620 7 2 2 72657 83061
0 39621 5 1 1 94316
0 39622 7 1 2 87638 94317
0 39623 5 1 1 39622
0 39624 7 3 2 66307 77234
0 39625 7 1 2 59635 94318
0 39626 5 1 1 39625
0 39627 7 1 2 92725 39626
0 39628 5 1 1 39627
0 39629 7 1 2 66925 39628
0 39630 5 1 1 39629
0 39631 7 1 2 39623 39630
0 39632 5 1 1 39631
0 39633 7 1 2 59378 39632
0 39634 5 1 1 39633
0 39635 7 1 2 58070 87340
0 39636 7 1 2 91842 39635
0 39637 5 1 1 39636
0 39638 7 1 2 39634 39637
0 39639 5 1 1 39638
0 39640 7 1 2 60144 39639
0 39641 5 1 1 39640
0 39642 7 2 2 81876 79813
0 39643 7 1 2 80637 74762
0 39644 7 1 2 94321 39643
0 39645 5 1 1 39644
0 39646 7 1 2 39641 39645
0 39647 5 1 1 39646
0 39648 7 1 2 58872 39647
0 39649 5 1 1 39648
0 39650 7 2 2 81041 83400
0 39651 7 1 2 94296 94323
0 39652 5 1 1 39651
0 39653 7 1 2 39649 39652
0 39654 5 1 1 39653
0 39655 7 1 2 79518 39654
0 39656 5 1 1 39655
0 39657 7 1 2 76155 90559
0 39658 5 2 1 39657
0 39659 7 1 2 60639 94325
0 39660 5 1 1 39659
0 39661 7 1 2 68140 82469
0 39662 5 1 1 39661
0 39663 7 1 2 39660 39662
0 39664 5 1 1 39663
0 39665 7 1 2 78871 39664
0 39666 5 1 1 39665
0 39667 7 1 2 78135 93519
0 39668 5 1 1 39667
0 39669 7 1 2 76220 39668
0 39670 5 1 1 39669
0 39671 7 1 2 68141 79731
0 39672 5 1 1 39671
0 39673 7 1 2 70429 39672
0 39674 7 1 2 39670 39673
0 39675 7 1 2 39666 39674
0 39676 5 1 1 39675
0 39677 7 1 2 59636 39676
0 39678 5 1 1 39677
0 39679 7 1 2 77995 75338
0 39680 5 2 1 39679
0 39681 7 1 2 74202 94327
0 39682 5 1 1 39681
0 39683 7 1 2 69465 39682
0 39684 5 1 1 39683
0 39685 7 1 2 79575 83881
0 39686 5 1 1 39685
0 39687 7 1 2 39684 39686
0 39688 5 1 1 39687
0 39689 7 1 2 57462 39688
0 39690 5 1 1 39689
0 39691 7 1 2 85708 80358
0 39692 5 2 1 39691
0 39693 7 1 2 20661 94329
0 39694 5 1 1 39693
0 39695 7 1 2 65301 39694
0 39696 5 1 1 39695
0 39697 7 1 2 6733 39696
0 39698 5 1 1 39697
0 39699 7 1 2 65668 39698
0 39700 5 1 1 39699
0 39701 7 1 2 61034 3564
0 39702 5 1 1 39701
0 39703 7 1 2 67363 80593
0 39704 7 1 2 39702 39703
0 39705 5 1 1 39704
0 39706 7 1 2 64389 93666
0 39707 5 1 1 39706
0 39708 7 1 2 77787 39707
0 39709 7 1 2 39705 39708
0 39710 7 1 2 39700 39709
0 39711 7 1 2 39690 39710
0 39712 7 1 2 39678 39711
0 39713 5 1 1 39712
0 39714 7 1 2 64601 39713
0 39715 5 1 1 39714
0 39716 7 2 2 67777 91180
0 39717 7 1 2 88588 87966
0 39718 7 1 2 94331 39717
0 39719 5 1 1 39718
0 39720 7 1 2 39715 39719
0 39721 5 1 1 39720
0 39722 7 1 2 66855 39721
0 39723 5 1 1 39722
0 39724 7 1 2 73800 78767
0 39725 5 1 1 39724
0 39726 7 1 2 57750 39725
0 39727 5 1 1 39726
0 39728 7 1 2 80042 94271
0 39729 5 1 1 39728
0 39730 7 1 2 57463 39729
0 39731 5 1 1 39730
0 39732 7 1 2 39727 39731
0 39733 5 1 1 39732
0 39734 7 1 2 92166 39733
0 39735 5 1 1 39734
0 39736 7 1 2 39723 39735
0 39737 5 1 1 39736
0 39738 7 1 2 84536 39737
0 39739 5 1 1 39738
0 39740 7 1 2 39656 39739
0 39741 7 1 2 39619 39740
0 39742 5 1 1 39741
0 39743 7 1 2 66520 39742
0 39744 5 1 1 39743
0 39745 7 1 2 39539 39744
0 39746 7 1 2 39490 39745
0 39747 5 1 1 39746
0 39748 7 1 2 66009 39747
0 39749 5 1 1 39748
0 39750 7 1 2 83955 93129
0 39751 5 1 1 39750
0 39752 7 1 2 57751 39751
0 39753 5 1 1 39752
0 39754 7 1 2 14382 39753
0 39755 5 2 1 39754
0 39756 7 2 2 89911 94333
0 39757 5 1 1 94335
0 39758 7 3 2 81585 94025
0 39759 7 1 2 67364 94337
0 39760 5 1 1 39759
0 39761 7 1 2 39757 39760
0 39762 5 1 1 39761
0 39763 7 1 2 94203 39762
0 39764 5 1 1 39763
0 39765 7 1 2 86947 88652
0 39766 5 1 1 39765
0 39767 7 1 2 66308 94177
0 39768 5 1 1 39767
0 39769 7 1 2 93414 39768
0 39770 5 1 1 39769
0 39771 7 3 2 66521 68398
0 39772 7 1 2 64726 94340
0 39773 7 1 2 39770 39772
0 39774 5 1 1 39773
0 39775 7 1 2 39766 39774
0 39776 5 1 1 39775
0 39777 7 1 2 65669 39776
0 39778 5 1 1 39777
0 39779 7 2 2 57752 92966
0 39780 7 1 2 87609 89884
0 39781 7 1 2 94343 39780
0 39782 5 1 1 39781
0 39783 7 1 2 39778 39782
0 39784 5 1 1 39783
0 39785 7 1 2 58777 39784
0 39786 5 1 1 39785
0 39787 7 1 2 16468 17048
0 39788 5 1 1 39787
0 39789 7 1 2 68030 39788
0 39790 5 1 1 39789
0 39791 7 1 2 36760 39790
0 39792 5 1 1 39791
0 39793 7 1 2 66309 39792
0 39794 5 1 1 39793
0 39795 7 1 2 60037 86948
0 39796 5 1 1 39795
0 39797 7 1 2 39794 39796
0 39798 5 1 1 39797
0 39799 7 1 2 78136 39798
0 39800 5 1 1 39799
0 39801 7 4 2 65073 86569
0 39802 7 2 2 77508 94345
0 39803 5 1 1 94349
0 39804 7 1 2 92020 94350
0 39805 5 1 1 39804
0 39806 7 1 2 39800 39805
0 39807 5 1 1 39806
0 39808 7 1 2 92955 39807
0 39809 5 1 1 39808
0 39810 7 1 2 39786 39809
0 39811 5 1 1 39810
0 39812 7 1 2 59890 39811
0 39813 5 1 1 39812
0 39814 7 1 2 71201 94334
0 39815 5 1 1 39814
0 39816 7 1 2 85778 93710
0 39817 5 1 1 39816
0 39818 7 1 2 39815 39817
0 39819 5 1 1 39818
0 39820 7 1 2 86303 39819
0 39821 5 1 1 39820
0 39822 7 1 2 81704 93100
0 39823 5 1 1 39822
0 39824 7 1 2 81508 90107
0 39825 7 1 2 39823 39824
0 39826 5 1 1 39825
0 39827 7 1 2 39821 39826
0 39828 5 1 1 39827
0 39829 7 1 2 89269 39828
0 39830 5 1 1 39829
0 39831 7 1 2 39813 39830
0 39832 5 1 1 39831
0 39833 7 1 2 60145 39832
0 39834 5 1 1 39833
0 39835 7 1 2 73968 83000
0 39836 5 1 1 39835
0 39837 7 1 2 29299 39836
0 39838 5 1 1 39837
0 39839 7 1 2 94338 39838
0 39840 5 1 1 39839
0 39841 7 1 2 79904 94341
0 39842 5 1 1 39841
0 39843 7 1 2 29635 39842
0 39844 5 1 1 39843
0 39845 7 1 2 66010 39844
0 39846 5 1 1 39845
0 39847 7 1 2 61869 82363
0 39848 7 1 2 83696 39847
0 39849 5 1 1 39848
0 39850 7 1 2 39846 39849
0 39851 5 1 1 39850
0 39852 7 1 2 82571 39851
0 39853 5 1 1 39852
0 39854 7 1 2 39840 39853
0 39855 5 1 1 39854
0 39856 7 1 2 58623 39855
0 39857 5 1 1 39856
0 39858 7 1 2 68399 93375
0 39859 5 1 1 39858
0 39860 7 2 2 71202 92306
0 39861 5 1 1 94351
0 39862 7 1 2 65074 94352
0 39863 5 1 1 39862
0 39864 7 1 2 39859 39863
0 39865 5 1 1 39864
0 39866 7 1 2 86304 39865
0 39867 5 1 1 39866
0 39868 7 2 2 79457 92609
0 39869 5 1 1 94353
0 39870 7 1 2 81348 94354
0 39871 5 1 1 39870
0 39872 7 1 2 39867 39871
0 39873 5 1 1 39872
0 39874 7 1 2 90077 39873
0 39875 5 1 1 39874
0 39876 7 1 2 39857 39875
0 39877 5 1 1 39876
0 39878 7 1 2 60146 39877
0 39879 5 1 1 39878
0 39880 7 1 2 94208 94339
0 39881 5 1 1 39880
0 39882 7 1 2 39879 39881
0 39883 5 1 1 39882
0 39884 7 1 2 67365 39883
0 39885 5 1 1 39884
0 39886 7 1 2 94209 94336
0 39887 5 1 1 39886
0 39888 7 1 2 39885 39887
0 39889 7 1 2 39834 39888
0 39890 5 1 1 39889
0 39891 7 1 2 58873 39890
0 39892 5 1 1 39891
0 39893 7 1 2 39764 39892
0 39894 5 1 1 39893
0 39895 7 1 2 72356 39894
0 39896 5 1 1 39895
0 39897 7 2 2 71591 92518
0 39898 7 2 2 72437 89912
0 39899 7 1 2 80116 73536
0 39900 7 1 2 94357 39899
0 39901 7 1 2 94355 39900
0 39902 5 1 1 39901
0 39903 7 1 2 39896 39902
0 39904 7 1 2 39749 39903
0 39905 7 1 2 39352 39904
0 39906 7 1 2 39148 39905
0 39907 5 1 1 39906
0 39908 7 1 2 67529 39907
0 39909 5 1 1 39908
0 39910 7 1 2 71909 25171
0 39911 5 1 1 39910
0 39912 7 1 2 78367 73470
0 39913 5 1 1 39912
0 39914 7 1 2 5087 39913
0 39915 7 1 2 39911 39914
0 39916 5 1 1 39915
0 39917 7 2 2 86491 39916
0 39918 5 1 1 94359
0 39919 7 1 2 74380 87202
0 39920 5 1 1 39919
0 39921 7 1 2 39918 39920
0 39922 5 1 1 39921
0 39923 7 1 2 71512 39922
0 39924 5 1 1 39923
0 39925 7 2 2 68254 84329
0 39926 5 2 1 94361
0 39927 7 1 2 65670 94363
0 39928 5 1 1 39927
0 39929 7 1 2 61386 39928
0 39930 5 1 1 39929
0 39931 7 1 2 84063 39930
0 39932 5 1 1 39931
0 39933 7 1 2 39924 39932
0 39934 5 1 1 39933
0 39935 7 1 2 68031 39934
0 39936 5 1 1 39935
0 39937 7 1 2 71203 94360
0 39938 5 1 1 39937
0 39939 7 1 2 39936 39938
0 39940 5 1 1 39939
0 39941 7 1 2 79905 39940
0 39942 5 1 1 39941
0 39943 7 1 2 86922 92142
0 39944 7 1 2 84427 39943
0 39945 5 1 1 39944
0 39946 7 1 2 39942 39945
0 39947 5 1 1 39946
0 39948 7 1 2 66522 39947
0 39949 5 1 1 39948
0 39950 7 1 2 71910 24547
0 39951 5 1 1 39950
0 39952 7 1 2 73471 78194
0 39953 5 1 1 39952
0 39954 7 1 2 39951 39953
0 39955 5 1 1 39954
0 39956 7 1 2 66011 39955
0 39957 5 1 1 39956
0 39958 7 1 2 61035 93496
0 39959 5 1 1 39958
0 39960 7 1 2 57464 93499
0 39961 7 1 2 39959 39960
0 39962 5 1 1 39961
0 39963 7 1 2 39957 39962
0 39964 5 1 1 39963
0 39965 7 2 2 61678 39964
0 39966 5 1 1 94365
0 39967 7 1 2 87213 39966
0 39968 5 1 1 39967
0 39969 7 1 2 71513 39968
0 39970 5 1 1 39969
0 39971 7 1 2 65671 80946
0 39972 5 1 1 39971
0 39973 7 1 2 61387 39972
0 39974 7 1 2 81630 39973
0 39975 5 1 1 39974
0 39976 7 1 2 84064 39975
0 39977 5 1 1 39976
0 39978 7 1 2 39970 39977
0 39979 5 1 1 39978
0 39980 7 1 2 68032 39979
0 39981 5 1 1 39980
0 39982 7 1 2 71204 94366
0 39983 5 1 1 39982
0 39984 7 1 2 39981 39983
0 39985 5 1 1 39984
0 39986 7 1 2 92268 39985
0 39987 5 1 1 39986
0 39988 7 1 2 92584 93963
0 39989 5 1 1 39988
0 39990 7 1 2 69847 88670
0 39991 5 1 1 39990
0 39992 7 2 2 36748 39991
0 39993 5 1 1 94367
0 39994 7 1 2 58998 2288
0 39995 7 1 2 7537 39994
0 39996 7 1 2 88793 39995
0 39997 5 1 1 39996
0 39998 7 1 2 94368 39997
0 39999 5 1 1 39998
0 40000 7 1 2 67676 39999
0 40001 5 1 1 40000
0 40002 7 1 2 68400 81754
0 40003 7 1 2 92292 40002
0 40004 5 1 1 40003
0 40005 7 1 2 40001 40004
0 40006 5 1 1 40005
0 40007 7 1 2 61036 40006
0 40008 5 1 1 40007
0 40009 7 1 2 83750 89498
0 40010 7 1 2 92296 40009
0 40011 5 1 1 40010
0 40012 7 1 2 40008 40011
0 40013 5 1 1 40012
0 40014 7 1 2 57465 40013
0 40015 5 1 1 40014
0 40016 7 1 2 59151 39993
0 40017 5 1 1 40016
0 40018 7 1 2 65075 88737
0 40019 5 1 1 40018
0 40020 7 1 2 40017 40019
0 40021 5 1 1 40020
0 40022 7 1 2 58999 40021
0 40023 5 1 1 40022
0 40024 7 1 2 59152 88738
0 40025 5 1 1 40024
0 40026 7 1 2 40023 40025
0 40027 5 1 1 40026
0 40028 7 1 2 57753 40027
0 40029 5 1 1 40028
0 40030 7 1 2 80735 93728
0 40031 5 1 1 40030
0 40032 7 1 2 40029 40031
0 40033 5 1 1 40032
0 40034 7 1 2 61037 40033
0 40035 5 1 1 40034
0 40036 7 1 2 40015 40035
0 40037 5 1 1 40036
0 40038 7 1 2 84670 40037
0 40039 5 1 1 40038
0 40040 7 1 2 39989 40039
0 40041 5 1 1 40040
0 40042 7 1 2 58778 40041
0 40043 5 1 1 40042
0 40044 7 1 2 81403 77217
0 40045 7 1 2 81806 89509
0 40046 7 1 2 40044 40045
0 40047 7 1 2 75240 40046
0 40048 5 1 1 40047
0 40049 7 1 2 40043 40048
0 40050 5 1 1 40049
0 40051 7 1 2 78271 40050
0 40052 5 1 1 40051
0 40053 7 1 2 39987 40052
0 40054 7 1 2 39949 40053
0 40055 5 1 1 40054
0 40056 7 1 2 61960 40055
0 40057 5 1 1 40056
0 40058 7 1 2 86882 89770
0 40059 5 1 1 40058
0 40060 7 1 2 86492 78901
0 40061 5 1 1 40060
0 40062 7 1 2 40059 40061
0 40063 5 2 1 40062
0 40064 7 1 2 82858 94369
0 40065 5 1 1 40064
0 40066 7 2 2 78909 82386
0 40067 7 1 2 65672 87370
0 40068 5 1 1 40067
0 40069 7 1 2 82476 78638
0 40070 5 1 1 40069
0 40071 7 1 2 61388 40070
0 40072 7 1 2 40068 40071
0 40073 5 1 1 40072
0 40074 7 1 2 94371 40073
0 40075 5 1 1 40074
0 40076 7 1 2 40065 40075
0 40077 5 1 1 40076
0 40078 7 1 2 88713 40077
0 40079 5 1 1 40078
0 40080 7 1 2 40057 40079
0 40081 5 1 1 40080
0 40082 7 1 2 67933 40081
0 40083 5 1 1 40082
0 40084 7 1 2 86223 84588
0 40085 5 1 1 40084
0 40086 7 1 2 80917 89695
0 40087 5 1 1 40086
0 40088 7 1 2 40085 40087
0 40089 5 1 1 40088
0 40090 7 1 2 71514 40089
0 40091 5 1 1 40090
0 40092 7 1 2 61389 85054
0 40093 5 1 1 40092
0 40094 7 3 2 80497 40093
0 40095 7 1 2 68401 94373
0 40096 5 1 1 40095
0 40097 7 1 2 85783 76282
0 40098 5 1 1 40097
0 40099 7 1 2 68784 40098
0 40100 5 1 1 40099
0 40101 7 1 2 85898 93575
0 40102 5 1 1 40101
0 40103 7 1 2 66012 79519
0 40104 5 1 1 40103
0 40105 7 1 2 40102 40104
0 40106 7 1 2 40100 40105
0 40107 7 1 2 40096 40106
0 40108 5 1 1 40107
0 40109 7 1 2 84065 40108
0 40110 5 1 1 40109
0 40111 7 1 2 40091 40110
0 40112 5 1 1 40111
0 40113 7 1 2 67056 40112
0 40114 5 1 1 40113
0 40115 7 2 2 87680 93919
0 40116 7 1 2 59637 84117
0 40117 7 1 2 94376 40116
0 40118 5 1 1 40117
0 40119 7 1 2 40114 40118
0 40120 5 1 1 40119
0 40121 7 1 2 58874 40120
0 40122 5 1 1 40121
0 40123 7 1 2 84493 94377
0 40124 5 1 1 40123
0 40125 7 1 2 40122 40124
0 40126 5 1 1 40125
0 40127 7 1 2 88824 40126
0 40128 5 1 1 40127
0 40129 7 3 2 73694 85971
0 40130 5 5 1 94378
0 40131 7 2 2 67934 72452
0 40132 5 1 1 94386
0 40133 7 1 2 1275 40132
0 40134 5 1 1 40133
0 40135 7 1 2 68785 40134
0 40136 5 1 1 40135
0 40137 7 1 2 13387 72598
0 40138 5 1 1 40137
0 40139 7 1 2 40136 40138
0 40140 5 1 1 40139
0 40141 7 1 2 57754 40140
0 40142 5 1 1 40141
0 40143 7 1 2 68906 75160
0 40144 5 1 1 40143
0 40145 7 1 2 94387 40144
0 40146 5 1 1 40145
0 40147 7 1 2 40142 40146
0 40148 5 1 1 40147
0 40149 7 1 2 65673 40148
0 40150 5 1 1 40149
0 40151 7 1 2 72380 69166
0 40152 7 1 2 76849 40151
0 40153 5 1 1 40152
0 40154 7 1 2 40150 40153
0 40155 5 1 1 40154
0 40156 7 1 2 66856 40155
0 40157 5 1 1 40156
0 40158 7 1 2 72638 82255
0 40159 7 1 2 71127 40158
0 40160 5 1 1 40159
0 40161 7 1 2 40157 40160
0 40162 5 1 1 40161
0 40163 7 1 2 94381 40162
0 40164 5 1 1 40163
0 40165 7 1 2 7450 9877
0 40166 5 1 1 40165
0 40167 7 2 2 67436 40166
0 40168 5 1 1 94388
0 40169 7 1 2 87367 92420
0 40170 5 1 1 40169
0 40171 7 1 2 94389 40170
0 40172 5 1 1 40171
0 40173 7 2 2 58875 66857
0 40174 7 1 2 64825 91149
0 40175 5 1 1 40174
0 40176 7 1 2 71964 93260
0 40177 7 1 2 40175 40176
0 40178 5 1 1 40177
0 40179 7 1 2 75878 66975
0 40180 5 1 1 40179
0 40181 7 1 2 72505 40180
0 40182 7 1 2 40178 40181
0 40183 5 1 1 40182
0 40184 7 1 2 94390 40183
0 40185 5 1 1 40184
0 40186 7 1 2 40172 40185
0 40187 5 1 1 40186
0 40188 7 1 2 79049 40187
0 40189 5 1 1 40188
0 40190 7 1 2 40164 40189
0 40191 5 1 1 40190
0 40192 7 1 2 61679 40191
0 40193 5 1 1 40192
0 40194 7 1 2 66976 89771
0 40195 5 1 1 40194
0 40196 7 2 2 67057 89696
0 40197 5 1 1 94392
0 40198 7 1 2 40195 40197
0 40199 5 1 1 40198
0 40200 7 1 2 58876 40199
0 40201 5 1 1 40200
0 40202 7 1 2 63638 81027
0 40203 7 2 2 86524 40202
0 40204 5 1 1 94394
0 40205 7 1 2 60640 94395
0 40206 5 1 1 40205
0 40207 7 1 2 40201 40206
0 40208 5 1 1 40207
0 40209 7 1 2 59153 40208
0 40210 5 1 1 40209
0 40211 7 1 2 87230 72599
0 40212 5 1 1 40211
0 40213 7 1 2 40210 40212
0 40214 5 1 1 40213
0 40215 7 1 2 57755 40214
0 40216 5 1 1 40215
0 40217 7 1 2 86493 79725
0 40218 5 2 1 40217
0 40219 7 1 2 78688 84671
0 40220 5 2 1 40219
0 40221 7 1 2 94396 94398
0 40222 5 1 1 40221
0 40223 7 1 2 72600 40222
0 40224 5 1 1 40223
0 40225 7 1 2 40216 40224
0 40226 5 1 1 40225
0 40227 7 1 2 66858 40226
0 40228 5 1 1 40227
0 40229 7 1 2 66310 82771
0 40230 7 1 2 94007 40229
0 40231 5 1 1 40230
0 40232 7 1 2 40228 40231
0 40233 5 1 1 40232
0 40234 7 1 2 71515 40233
0 40235 5 1 1 40234
0 40236 7 1 2 72705 88462
0 40237 5 1 1 40236
0 40238 7 1 2 89043 40237
0 40239 5 1 1 40238
0 40240 7 1 2 73444 40239
0 40241 5 1 1 40240
0 40242 7 3 2 60147 66013
0 40243 7 2 2 71361 94400
0 40244 5 1 1 94403
0 40245 7 1 2 81890 94404
0 40246 5 1 1 40245
0 40247 7 1 2 71362 89477
0 40248 5 1 1 40247
0 40249 7 4 2 57756 60148
0 40250 7 2 2 74295 94405
0 40251 5 1 1 94409
0 40252 7 1 2 58877 40251
0 40253 7 1 2 40248 40252
0 40254 5 1 1 40253
0 40255 7 1 2 63639 40244
0 40256 5 1 1 40255
0 40257 7 1 2 66859 40256
0 40258 7 1 2 40254 40257
0 40259 5 1 1 40258
0 40260 7 1 2 40246 40259
0 40261 5 1 1 40260
0 40262 7 1 2 71911 40261
0 40263 5 1 1 40262
0 40264 7 1 2 40241 40263
0 40265 5 1 1 40264
0 40266 7 1 2 84066 40265
0 40267 5 1 1 40266
0 40268 7 1 2 40235 40267
0 40269 5 1 1 40268
0 40270 7 1 2 68629 40269
0 40271 5 1 1 40270
0 40272 7 1 2 72534 88463
0 40273 5 1 1 40272
0 40274 7 1 2 89044 40273
0 40275 5 1 1 40274
0 40276 7 1 2 68402 40275
0 40277 5 1 1 40276
0 40278 7 1 2 71625 67618
0 40279 5 1 1 40278
0 40280 7 1 2 60641 83717
0 40281 7 1 2 70572 40280
0 40282 5 1 1 40281
0 40283 7 1 2 40279 40282
0 40284 5 1 1 40283
0 40285 7 1 2 66860 40284
0 40286 5 1 1 40285
0 40287 7 1 2 82179 83705
0 40288 7 1 2 89334 40287
0 40289 5 1 1 40288
0 40290 7 1 2 40286 40289
0 40291 7 1 2 40277 40290
0 40292 5 1 1 40291
0 40293 7 1 2 71516 40292
0 40294 5 1 1 40293
0 40295 7 1 2 77940 88464
0 40296 5 1 1 40295
0 40297 7 1 2 40294 40296
0 40298 5 1 1 40297
0 40299 7 1 2 61038 40298
0 40300 5 1 1 40299
0 40301 7 1 2 58878 83366
0 40302 7 1 2 80334 40301
0 40303 7 1 2 83450 40302
0 40304 5 1 1 40303
0 40305 7 1 2 40300 40304
0 40306 5 1 1 40305
0 40307 7 1 2 84672 40306
0 40308 5 1 1 40307
0 40309 7 1 2 40271 40308
0 40310 7 1 2 40193 40309
0 40311 5 1 1 40310
0 40312 7 1 2 61870 40311
0 40313 5 1 1 40312
0 40314 7 1 2 40128 40313
0 40315 5 1 1 40314
0 40316 7 1 2 67366 40315
0 40317 5 1 1 40316
0 40318 7 2 2 61390 81235
0 40319 5 1 1 94411
0 40320 7 1 2 77156 40319
0 40321 5 1 1 40320
0 40322 7 1 2 57757 80742
0 40323 5 1 1 40322
0 40324 7 1 2 71974 86278
0 40325 7 1 2 40323 40324
0 40326 7 1 2 40321 40325
0 40327 5 2 1 40326
0 40328 7 1 2 88825 94413
0 40329 5 1 1 40328
0 40330 7 1 2 93904 94412
0 40331 5 1 1 40330
0 40332 7 1 2 92269 40331
0 40333 5 1 1 40332
0 40334 7 1 2 40329 40333
0 40335 5 1 1 40334
0 40336 7 1 2 94372 40335
0 40337 5 1 1 40336
0 40338 7 1 2 92270 94370
0 40339 5 1 1 40338
0 40340 7 1 2 66523 92102
0 40341 7 1 2 80732 40340
0 40342 5 1 1 40341
0 40343 7 1 2 40339 40342
0 40344 5 1 1 40343
0 40345 7 1 2 82859 40344
0 40346 5 1 1 40345
0 40347 7 1 2 40337 40346
0 40348 5 1 1 40347
0 40349 7 1 2 70573 40348
0 40350 5 1 1 40349
0 40351 7 1 2 40317 40350
0 40352 7 1 2 40083 40351
0 40353 5 1 1 40352
0 40354 7 1 2 66715 40353
0 40355 5 1 1 40354
0 40356 7 1 2 82005 76595
0 40357 7 2 2 73537 40356
0 40358 7 1 2 58335 74897
0 40359 7 1 2 91203 40358
0 40360 7 1 2 90702 40359
0 40361 7 1 2 94415 40360
0 40362 5 1 1 40361
0 40363 7 1 2 40355 40362
0 40364 5 1 1 40363
0 40365 7 1 2 75577 40364
0 40366 5 1 1 40365
0 40367 7 1 2 68255 72404
0 40368 7 1 2 83270 40367
0 40369 5 1 1 40368
0 40370 7 1 2 77885 40369
0 40371 5 1 1 40370
0 40372 7 2 2 58624 78099
0 40373 5 2 1 94417
0 40374 7 1 2 65076 94418
0 40375 5 1 1 40374
0 40376 7 1 2 40371 40375
0 40377 5 1 1 40376
0 40378 7 1 2 73264 40377
0 40379 5 1 1 40378
0 40380 7 1 2 58625 93946
0 40381 7 1 2 80728 40380
0 40382 5 1 1 40381
0 40383 7 1 2 40379 40382
0 40384 5 1 1 40383
0 40385 7 1 2 66311 40384
0 40386 5 1 1 40385
0 40387 7 1 2 89357 94414
0 40388 5 1 1 40387
0 40389 7 1 2 40386 40388
0 40390 5 1 1 40389
0 40391 7 1 2 70574 40390
0 40392 5 1 1 40391
0 40393 7 1 2 64602 82531
0 40394 5 5 1 40393
0 40395 7 1 2 91961 94421
0 40396 5 1 1 40395
0 40397 7 1 2 67677 40396
0 40398 5 1 1 40397
0 40399 7 1 2 65674 85899
0 40400 5 2 1 40399
0 40401 7 1 2 61391 94426
0 40402 5 1 1 40401
0 40403 7 1 2 87341 40402
0 40404 5 1 1 40403
0 40405 7 1 2 68403 83596
0 40406 5 1 1 40405
0 40407 7 1 2 83295 40406
0 40408 5 1 1 40407
0 40409 7 1 2 82607 40408
0 40410 5 1 1 40409
0 40411 7 1 2 72847 90349
0 40412 5 3 1 40411
0 40413 7 1 2 94422 94428
0 40414 5 1 1 40413
0 40415 7 1 2 68630 40414
0 40416 5 1 1 40415
0 40417 7 2 2 73548 87237
0 40418 5 1 1 94431
0 40419 7 1 2 40416 40418
0 40420 5 1 1 40419
0 40421 7 1 2 68404 40420
0 40422 5 1 1 40421
0 40423 7 1 2 40410 40422
0 40424 7 1 2 40404 40423
0 40425 7 1 2 40398 40424
0 40426 5 1 1 40425
0 40427 7 1 2 82697 40426
0 40428 5 1 1 40427
0 40429 7 1 2 40392 40428
0 40430 5 1 1 40429
0 40431 7 1 2 66524 40430
0 40432 5 1 1 40431
0 40433 7 1 2 79201 94406
0 40434 7 1 2 82159 40433
0 40435 7 1 2 82304 89988
0 40436 7 1 2 40434 40435
0 40437 5 1 1 40436
0 40438 7 1 2 40432 40437
0 40439 5 1 1 40438
0 40440 7 1 2 66926 40439
0 40441 5 1 1 40440
0 40442 7 1 2 61039 78341
0 40443 5 1 1 40442
0 40444 7 1 2 82572 40443
0 40445 5 1 1 40444
0 40446 7 1 2 94423 40445
0 40447 5 1 1 40446
0 40448 7 1 2 89039 40447
0 40449 5 1 1 40448
0 40450 7 3 2 81115 81739
0 40451 7 1 2 93972 94433
0 40452 5 1 1 40451
0 40453 7 1 2 57758 82212
0 40454 5 2 1 40453
0 40455 7 1 2 92720 94436
0 40456 5 1 1 40455
0 40457 7 1 2 72579 40456
0 40458 7 1 2 79975 40457
0 40459 5 1 1 40458
0 40460 7 1 2 40452 40459
0 40461 5 1 1 40460
0 40462 7 1 2 71744 40461
0 40463 5 1 1 40462
0 40464 7 2 2 65675 78324
0 40465 7 1 2 92710 94438
0 40466 5 1 1 40465
0 40467 7 1 2 17353 40466
0 40468 5 1 1 40467
0 40469 7 1 2 88465 40468
0 40470 5 1 1 40469
0 40471 7 1 2 40463 40470
0 40472 7 1 2 40449 40471
0 40473 5 1 1 40472
0 40474 7 1 2 89449 40473
0 40475 5 1 1 40474
0 40476 7 1 2 66525 75253
0 40477 7 1 2 84022 94434
0 40478 7 1 2 40476 40477
0 40479 5 1 1 40478
0 40480 7 1 2 72259 89574
0 40481 7 1 2 89195 40480
0 40482 5 1 1 40481
0 40483 7 1 2 40479 40482
0 40484 5 1 1 40483
0 40485 7 1 2 80435 40484
0 40486 5 1 1 40485
0 40487 7 1 2 40475 40486
0 40488 5 1 1 40487
0 40489 7 1 2 71912 40488
0 40490 5 1 1 40489
0 40491 7 1 2 86728 70575
0 40492 5 1 1 40491
0 40493 7 1 2 58879 72152
0 40494 7 1 2 72971 84101
0 40495 7 1 2 40493 40494
0 40496 5 1 1 40495
0 40497 7 1 2 40492 40496
0 40498 5 1 1 40497
0 40499 7 1 2 89660 40498
0 40500 5 1 1 40499
0 40501 7 3 2 65676 82658
0 40502 7 1 2 58626 90116
0 40503 7 1 2 94440 40502
0 40504 5 1 1 40503
0 40505 7 1 2 40500 40504
0 40506 5 1 1 40505
0 40507 7 1 2 66861 40506
0 40508 5 1 1 40507
0 40509 7 1 2 89338 91734
0 40510 5 1 1 40509
0 40511 7 1 2 40508 40510
0 40512 5 1 1 40511
0 40513 7 1 2 78325 40512
0 40514 5 1 1 40513
0 40515 7 2 2 65077 78969
0 40516 5 1 1 94443
0 40517 7 1 2 61392 40516
0 40518 5 1 1 40517
0 40519 7 1 2 89040 40518
0 40520 5 1 1 40519
0 40521 7 1 2 66014 93647
0 40522 5 2 1 40521
0 40523 7 1 2 94047 94445
0 40524 7 1 2 93961 40523
0 40525 5 1 1 40524
0 40526 7 1 2 88466 40525
0 40527 5 1 1 40526
0 40528 7 1 2 40520 40527
0 40529 5 1 1 40528
0 40530 7 1 2 91718 40529
0 40531 5 1 1 40530
0 40532 7 1 2 63913 70882
0 40533 5 1 1 40532
0 40534 7 2 2 61680 86729
0 40535 7 1 2 89313 94447
0 40536 7 1 2 40533 40535
0 40537 7 1 2 79976 40536
0 40538 5 1 1 40537
0 40539 7 1 2 40531 40538
0 40540 7 1 2 40514 40539
0 40541 5 1 1 40540
0 40542 7 1 2 64603 40541
0 40543 5 1 1 40542
0 40544 7 1 2 82213 73445
0 40545 5 1 1 40544
0 40546 7 1 2 76244 92718
0 40547 5 1 1 40546
0 40548 7 1 2 40545 40547
0 40549 5 1 1 40548
0 40550 7 1 2 88467 40549
0 40551 5 1 1 40550
0 40552 7 2 2 73472 82573
0 40553 5 1 1 94449
0 40554 7 1 2 89041 94450
0 40555 5 1 1 40554
0 40556 7 1 2 40551 40555
0 40557 5 1 1 40556
0 40558 7 1 2 89450 40557
0 40559 5 1 1 40558
0 40560 7 2 2 57466 66526
0 40561 7 1 2 81807 94451
0 40562 7 1 2 85757 40561
0 40563 7 2 2 58779 87263
0 40564 5 2 1 94453
0 40565 7 1 2 67619 94454
0 40566 7 1 2 40562 40565
0 40567 5 1 1 40566
0 40568 7 1 2 40559 40567
0 40569 5 1 1 40568
0 40570 7 1 2 71745 40569
0 40571 5 1 1 40570
0 40572 7 1 2 66977 94391
0 40573 5 1 1 40572
0 40574 7 1 2 40168 40573
0 40575 5 1 1 40574
0 40576 7 2 2 61393 93959
0 40577 5 1 1 94457
0 40578 7 1 2 73437 94458
0 40579 5 2 1 40578
0 40580 7 1 2 40575 94459
0 40581 5 1 1 40580
0 40582 7 2 2 66862 67620
0 40583 7 1 2 61394 84929
0 40584 7 1 2 76251 40583
0 40585 7 1 2 73992 40584
0 40586 5 1 1 40585
0 40587 7 1 2 94461 40586
0 40588 5 1 1 40587
0 40589 7 1 2 40581 40588
0 40590 5 1 1 40589
0 40591 7 1 2 90004 40590
0 40592 5 1 1 40591
0 40593 7 1 2 40571 40592
0 40594 7 1 2 40543 40593
0 40595 7 1 2 40490 40594
0 40596 7 1 2 40441 40595
0 40597 5 1 1 40596
0 40598 7 1 2 66716 40597
0 40599 5 1 1 40598
0 40600 7 1 2 79267 83697
0 40601 7 1 2 89013 40600
0 40602 7 1 2 79625 90703
0 40603 7 1 2 40601 40602
0 40604 5 1 1 40603
0 40605 7 1 2 40599 40604
0 40606 5 1 1 40605
0 40607 7 1 2 78272 40606
0 40608 5 1 1 40607
0 40609 7 1 2 70353 89063
0 40610 5 1 1 40609
0 40611 7 1 2 86730 89270
0 40612 5 1 1 40611
0 40613 7 1 2 40610 40612
0 40614 5 1 1 40613
0 40615 7 1 2 57467 40614
0 40616 5 1 1 40615
0 40617 7 1 2 89271 92883
0 40618 5 1 1 40617
0 40619 7 1 2 40616 40618
0 40620 5 2 1 40619
0 40621 7 1 2 61681 94463
0 40622 5 1 1 40621
0 40623 7 1 2 89597 93878
0 40624 5 1 1 40623
0 40625 7 1 2 40622 40624
0 40626 5 1 1 40625
0 40627 7 1 2 66606 40626
0 40628 5 1 1 40627
0 40629 7 3 2 71205 92014
0 40630 7 1 2 73384 89612
0 40631 7 1 2 94465 40630
0 40632 5 1 1 40631
0 40633 7 1 2 40628 40632
0 40634 5 1 1 40633
0 40635 7 1 2 59154 40634
0 40636 5 1 1 40635
0 40637 7 1 2 82659 93307
0 40638 5 1 1 40637
0 40639 7 2 2 63378 89179
0 40640 7 1 2 82103 94468
0 40641 5 1 1 40640
0 40642 7 1 2 40638 40641
0 40643 5 1 1 40642
0 40644 7 1 2 87465 40643
0 40645 5 1 1 40644
0 40646 7 1 2 87264 83036
0 40647 7 1 2 92884 40646
0 40648 5 1 1 40647
0 40649 7 1 2 40645 40648
0 40650 5 1 1 40649
0 40651 7 1 2 66527 40650
0 40652 5 1 1 40651
0 40653 7 3 2 85654 85881
0 40654 7 1 2 83037 90899
0 40655 7 1 2 94470 40654
0 40656 5 1 1 40655
0 40657 7 2 2 40652 40656
0 40658 5 1 1 94473
0 40659 7 1 2 40636 94474
0 40660 5 1 1 40659
0 40661 7 1 2 60149 40660
0 40662 5 1 1 40661
0 40663 7 3 2 81042 74056
0 40664 7 1 2 73670 76858
0 40665 7 1 2 91739 40664
0 40666 7 1 2 94475 40665
0 40667 5 1 1 40666
0 40668 7 1 2 40662 40667
0 40669 5 1 1 40668
0 40670 7 1 2 66863 40669
0 40671 5 1 1 40670
0 40672 7 1 2 73671 84102
0 40673 7 1 2 92956 40672
0 40674 7 2 2 66312 75738
0 40675 7 1 2 94476 94478
0 40676 7 1 2 40673 40675
0 40677 5 1 1 40676
0 40678 7 1 2 40671 40677
0 40679 5 1 1 40678
0 40680 7 1 2 67367 40679
0 40681 5 1 1 40680
0 40682 7 1 2 84575 94407
0 40683 5 1 1 40682
0 40684 7 1 2 83946 66978
0 40685 5 1 1 40684
0 40686 7 1 2 40683 40685
0 40687 5 1 1 40686
0 40688 7 1 2 57468 40687
0 40689 5 1 1 40688
0 40690 7 1 2 69193 82794
0 40691 5 1 1 40690
0 40692 7 1 2 40689 40691
0 40693 5 1 1 40692
0 40694 7 1 2 59155 40693
0 40695 5 1 1 40694
0 40696 7 1 2 66015 68194
0 40697 5 1 1 40696
0 40698 7 1 2 40695 40697
0 40699 5 1 1 40698
0 40700 7 1 2 66864 40699
0 40701 5 1 1 40700
0 40702 7 1 2 57469 73795
0 40703 5 1 1 40702
0 40704 7 1 2 61395 40703
0 40705 5 1 1 40704
0 40706 7 1 2 72328 82046
0 40707 7 1 2 40705 40706
0 40708 5 1 1 40707
0 40709 7 1 2 40701 40708
0 40710 5 1 1 40709
0 40711 7 1 2 89009 40710
0 40712 5 1 1 40711
0 40713 7 1 2 70176 88708
0 40714 7 1 2 93912 40713
0 40715 7 1 2 82042 40714
0 40716 5 1 1 40715
0 40717 7 1 2 40712 40716
0 40718 5 1 1 40717
0 40719 7 1 2 71206 40718
0 40720 5 1 1 40719
0 40721 7 1 2 68033 88709
0 40722 7 1 2 93951 40721
0 40723 7 2 2 61396 79458
0 40724 5 1 1 94480
0 40725 7 2 2 60038 72438
0 40726 7 1 2 94481 94482
0 40727 7 1 2 40722 40726
0 40728 5 1 1 40727
0 40729 7 1 2 40720 40728
0 40730 5 1 1 40729
0 40731 7 1 2 66313 40730
0 40732 5 1 1 40731
0 40733 7 1 2 82104 74827
0 40734 7 1 2 79696 40733
0 40735 7 4 2 57470 89510
0 40736 7 1 2 94483 94484
0 40737 7 1 2 40734 40736
0 40738 5 1 1 40737
0 40739 7 1 2 63640 40738
0 40740 7 1 2 40732 40739
0 40741 7 1 2 40681 40740
0 40742 5 1 1 40741
0 40743 7 2 2 73056 72288
0 40744 7 1 2 73969 94488
0 40745 5 1 1 40744
0 40746 7 1 2 60039 73549
0 40747 5 1 1 40746
0 40748 7 1 2 40745 40747
0 40749 5 1 1 40748
0 40750 7 1 2 58627 40749
0 40751 5 1 1 40750
0 40752 7 1 2 1395 87062
0 40753 5 1 1 40752
0 40754 7 1 2 71207 40753
0 40755 5 1 1 40754
0 40756 7 1 2 85602 40755
0 40757 5 1 1 40756
0 40758 7 1 2 60040 40757
0 40759 5 1 1 40758
0 40760 7 1 2 40751 40759
0 40761 5 1 1 40760
0 40762 7 1 2 58780 40761
0 40763 5 1 1 40762
0 40764 7 1 2 93850 94489
0 40765 5 1 1 40764
0 40766 7 1 2 40763 40765
0 40767 5 1 1 40766
0 40768 7 1 2 81719 40767
0 40769 5 1 1 40768
0 40770 7 1 2 85882 90940
0 40771 5 1 1 40770
0 40772 7 1 2 59891 40771
0 40773 5 1 1 40772
0 40774 7 1 2 64604 10514
0 40775 7 1 2 90801 40774
0 40776 5 1 1 40775
0 40777 7 1 2 77273 40776
0 40778 7 1 2 40773 40777
0 40779 5 1 1 40778
0 40780 7 1 2 40769 40779
0 40781 5 1 1 40780
0 40782 7 1 2 58071 40781
0 40783 5 1 1 40782
0 40784 7 1 2 78970 75661
0 40785 5 1 1 40784
0 40786 7 1 2 66016 75767
0 40787 5 1 1 40786
0 40788 7 1 2 40785 40787
0 40789 5 1 1 40788
0 40790 7 1 2 93358 40789
0 40791 5 1 1 40790
0 40792 7 1 2 75768 94471
0 40793 5 1 1 40792
0 40794 7 2 2 72972 82364
0 40795 7 1 2 57471 79459
0 40796 7 1 2 94490 40795
0 40797 5 1 1 40796
0 40798 7 1 2 40793 40797
0 40799 5 1 1 40798
0 40800 7 1 2 59892 40799
0 40801 5 1 1 40800
0 40802 7 1 2 40791 40801
0 40803 5 1 1 40802
0 40804 7 1 2 59379 40803
0 40805 5 1 1 40804
0 40806 7 1 2 60150 40805
0 40807 7 1 2 40783 40806
0 40808 5 1 1 40807
0 40809 7 1 2 67368 93879
0 40810 5 1 1 40809
0 40811 7 1 2 81070 93872
0 40812 5 1 1 40811
0 40813 7 1 2 40810 40812
0 40814 5 1 1 40813
0 40815 7 1 2 74487 40814
0 40816 5 1 1 40815
0 40817 7 1 2 64826 40816
0 40818 5 1 1 40817
0 40819 7 1 2 61871 40818
0 40820 7 1 2 40808 40819
0 40821 5 1 1 40820
0 40822 7 1 2 73887 87468
0 40823 5 1 1 40822
0 40824 7 1 2 85463 40823
0 40825 5 1 1 40824
0 40826 7 1 2 8915 40825
0 40827 5 1 1 40826
0 40828 7 1 2 61961 40827
0 40829 5 1 1 40828
0 40830 7 2 2 66607 67369
0 40831 7 1 2 64827 87686
0 40832 7 1 2 94492 40831
0 40833 5 1 1 40832
0 40834 7 1 2 40829 40833
0 40835 5 1 1 40834
0 40836 7 1 2 57759 40835
0 40837 5 1 1 40836
0 40838 7 3 2 57472 66979
0 40839 7 1 2 76331 74238
0 40840 7 1 2 94494 40839
0 40841 5 1 1 40840
0 40842 7 1 2 40837 40841
0 40843 5 1 1 40842
0 40844 7 1 2 93507 40843
0 40845 5 1 1 40844
0 40846 7 1 2 66314 40845
0 40847 7 1 2 40821 40846
0 40848 5 1 1 40847
0 40849 7 2 2 64390 81740
0 40850 7 1 2 93947 94497
0 40851 5 1 1 40850
0 40852 7 1 2 64605 37624
0 40853 5 1 1 40852
0 40854 7 1 2 94040 94282
0 40855 7 1 2 40853 40854
0 40856 5 1 1 40855
0 40857 7 1 2 40851 40856
0 40858 5 1 1 40857
0 40859 7 1 2 66528 40858
0 40860 5 1 1 40859
0 40861 7 1 2 91006 92986
0 40862 5 1 1 40861
0 40863 7 1 2 40860 40862
0 40864 5 1 1 40863
0 40865 7 1 2 58072 40864
0 40866 5 1 1 40865
0 40867 7 1 2 89511 91999
0 40868 5 1 1 40867
0 40869 7 1 2 89065 40868
0 40870 5 1 1 40869
0 40871 7 1 2 65677 76052
0 40872 7 1 2 40870 40871
0 40873 5 1 1 40872
0 40874 7 1 2 40866 40873
0 40875 5 1 1 40874
0 40876 7 1 2 77017 40875
0 40877 5 1 1 40876
0 40878 7 5 2 66608 85464
0 40879 7 1 2 67370 94464
0 40880 5 1 1 40879
0 40881 7 1 2 69746 88416
0 40882 7 1 2 94485 40881
0 40883 5 1 1 40882
0 40884 7 1 2 40880 40883
0 40885 5 1 1 40884
0 40886 7 1 2 94499 40885
0 40887 5 1 1 40886
0 40888 7 1 2 61682 40887
0 40889 7 1 2 40877 40888
0 40890 5 1 1 40889
0 40891 7 1 2 59156 40890
0 40892 7 1 2 40848 40891
0 40893 5 1 1 40892
0 40894 7 1 2 85465 40658
0 40895 5 1 1 40894
0 40896 7 3 2 57760 67117
0 40897 7 1 2 75662 91250
0 40898 7 1 2 94504 40897
0 40899 7 1 2 94252 40898
0 40900 5 1 1 40899
0 40901 7 1 2 40895 40900
0 40902 5 1 1 40901
0 40903 7 1 2 67371 40902
0 40904 5 1 1 40903
0 40905 7 1 2 81116 72439
0 40906 7 1 2 94263 40905
0 40907 5 1 1 40906
0 40908 7 1 2 68034 86637
0 40909 7 1 2 81055 40908
0 40910 5 1 1 40909
0 40911 7 1 2 40907 40910
0 40912 5 1 1 40911
0 40913 7 1 2 66529 40912
0 40914 5 1 1 40913
0 40915 7 1 2 58880 40914
0 40916 7 1 2 40904 40915
0 40917 7 1 2 40893 40916
0 40918 5 1 1 40917
0 40919 7 1 2 65302 40918
0 40920 7 1 2 40742 40919
0 40921 5 1 1 40920
0 40922 7 1 2 93881 94500
0 40923 5 1 1 40922
0 40924 7 2 2 77771 74052
0 40925 5 1 1 94507
0 40926 7 1 2 94221 94508
0 40927 5 1 1 40926
0 40928 7 3 2 66017 84009
0 40929 5 1 1 94509
0 40930 7 1 2 40927 40929
0 40931 5 1 1 40930
0 40932 7 1 2 71208 40931
0 40933 5 1 1 40932
0 40934 7 1 2 77831 22176
0 40935 5 4 1 40934
0 40936 7 1 2 87610 94512
0 40937 5 1 1 40936
0 40938 7 1 2 40933 40937
0 40939 5 1 1 40938
0 40940 7 1 2 58781 40939
0 40941 5 1 1 40940
0 40942 7 6 2 58073 81043
0 40943 7 4 2 72991 94516
0 40944 7 3 2 59893 94522
0 40945 7 1 2 94015 94526
0 40946 5 1 1 40945
0 40947 7 1 2 40941 40946
0 40948 5 1 1 40947
0 40949 7 1 2 67125 40948
0 40950 5 1 1 40949
0 40951 7 1 2 40923 40950
0 40952 5 1 1 40951
0 40953 7 1 2 66315 40952
0 40954 5 1 1 40953
0 40955 7 1 2 91518 93896
0 40956 5 1 1 40955
0 40957 7 1 2 93510 94501
0 40958 5 1 1 40957
0 40959 7 1 2 40956 40958
0 40960 5 1 1 40959
0 40961 7 1 2 67372 40960
0 40962 5 1 1 40961
0 40963 7 1 2 81117 94401
0 40964 7 1 2 92519 40963
0 40965 5 1 1 40964
0 40966 7 1 2 40962 40965
0 40967 7 1 2 40954 40966
0 40968 5 1 1 40967
0 40969 7 1 2 61872 40968
0 40970 5 1 1 40969
0 40971 7 2 2 64606 76609
0 40972 7 2 2 72973 88245
0 40973 7 1 2 94529 94531
0 40974 5 1 1 40973
0 40975 7 2 2 82712 72580
0 40976 7 1 2 92440 94533
0 40977 5 1 1 40976
0 40978 7 1 2 40974 40977
0 40979 5 1 1 40978
0 40980 7 1 2 58628 40979
0 40981 5 1 1 40980
0 40982 7 5 2 60151 81118
0 40983 7 1 2 92352 94535
0 40984 5 1 1 40983
0 40985 7 1 2 40981 40984
0 40986 5 1 1 40985
0 40987 7 1 2 71209 40986
0 40988 5 1 1 40987
0 40989 7 1 2 85741 87265
0 40990 7 1 2 94502 40989
0 40991 5 1 1 40990
0 40992 7 1 2 40988 40991
0 40993 5 1 1 40992
0 40994 7 1 2 68035 40993
0 40995 5 1 1 40994
0 40996 7 1 2 87266 72581
0 40997 7 1 2 85466 40996
0 40998 7 1 2 94472 40997
0 40999 5 1 1 40998
0 41000 7 1 2 40995 40999
0 41001 5 1 1 41000
0 41002 7 1 2 94452 41001
0 41003 5 1 1 41002
0 41004 7 1 2 40970 41003
0 41005 5 1 1 41004
0 41006 7 1 2 58881 41005
0 41007 5 1 1 41006
0 41008 7 4 2 63641 66609
0 41009 7 1 2 91322 93883
0 41010 5 1 1 41009
0 41011 7 1 2 72822 84118
0 41012 7 1 2 91124 41011
0 41013 7 1 2 72672 41012
0 41014 5 1 1 41013
0 41015 7 1 2 41010 41014
0 41016 5 1 1 41015
0 41017 7 1 2 66316 41016
0 41018 5 1 1 41017
0 41019 7 1 2 86989 93433
0 41020 5 2 1 41019
0 41021 7 3 2 57473 64607
0 41022 7 2 2 89661 94546
0 41023 5 1 1 94549
0 41024 7 1 2 72440 94550
0 41025 7 1 2 94544 41024
0 41026 5 1 1 41025
0 41027 7 1 2 41018 41026
0 41028 5 1 1 41027
0 41029 7 1 2 66865 41028
0 41030 5 1 1 41029
0 41031 7 1 2 72992 87884
0 41032 7 3 2 58336 72823
0 41033 7 1 2 94358 94551
0 41034 7 1 2 41031 41033
0 41035 5 1 1 41034
0 41036 7 1 2 41030 41035
0 41037 5 1 1 41036
0 41038 7 1 2 94540 41037
0 41039 5 1 1 41038
0 41040 7 1 2 41007 41039
0 41041 5 1 1 41040
0 41042 7 1 2 57761 41041
0 41043 5 1 1 41042
0 41044 7 1 2 73840 89996
0 41045 7 2 2 86607 41044
0 41046 7 1 2 83159 94554
0 41047 5 1 1 41046
0 41048 7 1 2 82786 92594
0 41049 5 1 1 41048
0 41050 7 1 2 89997 91168
0 41051 5 1 1 41050
0 41052 7 1 2 41049 41051
0 41053 5 1 1 41052
0 41054 7 1 2 70528 41053
0 41055 5 1 1 41054
0 41056 7 1 2 66786 84299
0 41057 7 1 2 90117 41056
0 41058 5 1 1 41057
0 41059 7 1 2 59638 71062
0 41060 7 1 2 85194 41059
0 41061 7 1 2 89998 41060
0 41062 5 1 1 41061
0 41063 7 1 2 41058 41062
0 41064 7 1 2 41055 41063
0 41065 5 1 1 41064
0 41066 7 1 2 89286 41065
0 41067 5 1 1 41066
0 41068 7 2 2 64391 84010
0 41069 7 1 2 81028 83555
0 41070 7 1 2 92294 41069
0 41071 7 1 2 94556 41070
0 41072 5 1 1 41071
0 41073 7 1 2 41067 41072
0 41074 5 1 1 41073
0 41075 7 1 2 67373 41074
0 41076 5 1 1 41075
0 41077 7 1 2 82993 94555
0 41078 5 1 1 41077
0 41079 7 1 2 41076 41078
0 41080 5 1 1 41079
0 41081 7 1 2 66018 41080
0 41082 5 1 1 41081
0 41083 7 1 2 41047 41082
0 41084 7 1 2 41043 41083
0 41085 5 1 1 41084
0 41086 7 1 2 71913 41085
0 41087 5 1 1 41086
0 41088 7 1 2 59894 93443
0 41089 5 1 1 41088
0 41090 7 1 2 94135 41089
0 41091 5 1 1 41090
0 41092 7 1 2 78950 41091
0 41093 5 1 1 41092
0 41094 7 1 2 73265 78100
0 41095 7 1 2 83644 41094
0 41096 5 1 1 41095
0 41097 7 1 2 41093 41096
0 41098 5 1 1 41097
0 41099 7 1 2 66530 41098
0 41100 5 1 1 41099
0 41101 7 1 2 83160 92121
0 41102 5 1 1 41101
0 41103 7 1 2 41100 41102
0 41104 5 1 1 41103
0 41105 7 1 2 66317 41104
0 41106 5 1 1 41105
0 41107 7 1 2 86295 89731
0 41108 5 1 1 41107
0 41109 7 1 2 64392 94486
0 41110 5 1 1 41109
0 41111 7 1 2 21782 41110
0 41112 5 1 1 41111
0 41113 7 1 2 68036 41112
0 41114 5 1 1 41113
0 41115 7 1 2 85909 94487
0 41116 5 1 1 41115
0 41117 7 1 2 89451 90009
0 41118 5 1 1 41117
0 41119 7 2 2 41116 41118
0 41120 5 1 1 94558
0 41121 7 1 2 41114 94559
0 41122 5 1 1 41121
0 41123 7 1 2 66318 41122
0 41124 5 1 1 41123
0 41125 7 1 2 85549 94289
0 41126 5 2 1 41125
0 41127 7 1 2 41124 94560
0 41128 5 1 1 41127
0 41129 7 1 2 59895 41128
0 41130 5 1 1 41129
0 41131 7 1 2 82543 92107
0 41132 7 1 2 94552 41131
0 41133 5 1 1 41132
0 41134 7 1 2 41130 41133
0 41135 5 1 1 41134
0 41136 7 1 2 81232 41135
0 41137 5 1 1 41136
0 41138 7 1 2 41108 41137
0 41139 7 1 2 41106 41138
0 41140 5 1 1 41139
0 41141 7 1 2 70529 41140
0 41142 5 1 1 41141
0 41143 7 1 2 68405 94545
0 41144 5 1 1 41143
0 41145 7 1 2 65303 94178
0 41146 5 1 1 41145
0 41147 7 1 2 41144 41146
0 41148 5 1 1 41147
0 41149 7 1 2 65678 41148
0 41150 5 1 1 41149
0 41151 7 1 2 84339 86731
0 41152 5 1 1 41151
0 41153 7 1 2 41150 41152
0 41154 5 1 1 41153
0 41155 7 2 2 79202 67118
0 41156 7 1 2 89885 94562
0 41157 7 1 2 41154 41156
0 41158 5 1 1 41157
0 41159 7 1 2 41142 41158
0 41160 5 1 1 41159
0 41161 7 1 2 66610 41160
0 41162 5 1 1 41161
0 41163 7 1 2 66319 41120
0 41164 5 1 1 41163
0 41165 7 1 2 94561 41164
0 41166 5 2 1 41165
0 41167 7 1 2 70576 94564
0 41168 5 1 1 41167
0 41169 7 2 2 60152 71210
0 41170 7 1 2 77025 81720
0 41171 7 1 2 91251 41170
0 41172 7 1 2 94566 41171
0 41173 5 1 1 41172
0 41174 7 1 2 41168 41173
0 41175 5 1 1 41174
0 41176 7 1 2 65304 41175
0 41177 5 1 1 41176
0 41178 7 1 2 66531 89014
0 41179 7 1 2 91836 41178
0 41180 5 1 1 41179
0 41181 7 1 2 41177 41180
0 41182 5 1 1 41181
0 41183 7 1 2 59896 41182
0 41184 5 1 1 41183
0 41185 7 1 2 82959 90771
0 41186 5 1 1 41185
0 41187 7 1 2 88710 88246
0 41188 7 1 2 87064 41187
0 41189 5 1 1 41188
0 41190 7 1 2 41186 41189
0 41191 5 1 1 41190
0 41192 7 1 2 67935 73513
0 41193 7 1 2 41191 41192
0 41194 5 1 1 41193
0 41195 7 1 2 41184 41194
0 41196 5 1 1 41195
0 41197 7 1 2 68406 41196
0 41198 5 1 1 41197
0 41199 7 1 2 79520 94565
0 41200 5 1 1 41199
0 41201 7 3 2 81404 90078
0 41202 7 1 2 84821 94568
0 41203 5 1 1 41202
0 41204 7 1 2 41200 41203
0 41205 5 1 1 41204
0 41206 7 1 2 87970 41205
0 41207 5 1 1 41206
0 41208 7 1 2 64828 94569
0 41209 7 1 2 85919 41208
0 41210 5 1 1 41209
0 41211 7 1 2 73072 85557
0 41212 7 1 2 67119 89886
0 41213 7 1 2 41211 41212
0 41214 7 1 2 93576 41213
0 41215 5 1 1 41214
0 41216 7 1 2 41210 41215
0 41217 5 1 1 41216
0 41218 7 1 2 58882 41217
0 41219 5 1 1 41218
0 41220 7 1 2 70462 94570
0 41221 7 1 2 85920 41220
0 41222 5 1 1 41221
0 41223 7 1 2 41219 41222
0 41224 5 1 1 41223
0 41225 7 1 2 78101 41224
0 41226 5 1 1 41225
0 41227 7 1 2 41207 41226
0 41228 5 1 1 41227
0 41229 7 1 2 66611 41228
0 41230 5 1 1 41229
0 41231 7 1 2 87469 76283
0 41232 5 1 1 41231
0 41233 7 1 2 93359 41232
0 41234 5 1 1 41233
0 41235 7 1 2 86225 73501
0 41236 5 1 1 41235
0 41237 7 1 2 41234 41236
0 41238 5 1 1 41237
0 41239 7 1 2 66320 41238
0 41240 5 1 1 41239
0 41241 7 1 2 89358 93577
0 41242 5 1 1 41241
0 41243 7 1 2 41240 41242
0 41244 5 1 1 41243
0 41245 7 1 2 88800 41244
0 41246 5 1 1 41245
0 41247 7 1 2 87466 93490
0 41248 5 1 1 41247
0 41249 7 1 2 41246 41248
0 41250 5 1 1 41249
0 41251 7 1 2 72601 41250
0 41252 5 1 1 41251
0 41253 7 1 2 41230 41252
0 41254 7 1 2 41198 41253
0 41255 5 1 1 41254
0 41256 7 1 2 67374 41255
0 41257 5 1 1 41256
0 41258 7 1 2 77813 79423
0 41259 5 1 1 41258
0 41260 7 1 2 86841 41259
0 41261 5 1 1 41260
0 41262 7 1 2 32556 41261
0 41263 5 1 1 41262
0 41264 7 1 2 82463 41263
0 41265 5 1 1 41264
0 41266 7 1 2 82960 87436
0 41267 5 1 1 41266
0 41268 7 1 2 89393 41267
0 41269 5 1 1 41268
0 41270 7 1 2 70099 41269
0 41271 5 1 1 41270
0 41272 7 1 2 41265 41271
0 41273 5 1 1 41272
0 41274 7 1 2 66532 41273
0 41275 5 1 1 41274
0 41276 7 1 2 57474 79734
0 41277 7 1 2 93491 41276
0 41278 5 1 1 41277
0 41279 7 1 2 41275 41278
0 41280 5 1 1 41279
0 41281 7 1 2 66019 41280
0 41282 5 1 1 41281
0 41283 7 1 2 80481 93875
0 41284 5 1 1 41283
0 41285 7 1 2 65305 41284
0 41286 5 1 1 41285
0 41287 7 1 2 68256 41286
0 41288 5 1 1 41287
0 41289 7 1 2 89999 94259
0 41290 7 1 2 41288 41289
0 41291 5 1 1 41290
0 41292 7 1 2 41282 41291
0 41293 5 1 1 41292
0 41294 7 1 2 72602 41293
0 41295 5 1 1 41294
0 41296 7 1 2 41257 41295
0 41297 7 1 2 41162 41296
0 41298 5 1 1 41297
0 41299 7 1 2 66927 41298
0 41300 5 1 1 41299
0 41301 7 1 2 90450 92000
0 41302 5 1 1 41301
0 41303 7 1 2 89250 41302
0 41304 5 1 1 41303
0 41305 7 1 2 67058 41304
0 41306 5 1 1 41305
0 41307 7 1 2 25203 92694
0 41308 5 2 1 41307
0 41309 7 1 2 94495 94571
0 41310 5 1 1 41309
0 41311 7 1 2 41306 41310
0 41312 5 1 1 41311
0 41313 7 1 2 61683 41312
0 41314 5 1 1 41313
0 41315 7 1 2 67090 1122
0 41316 5 1 1 41315
0 41317 7 1 2 93360 41316
0 41318 5 1 1 41317
0 41319 7 1 2 68941 83282
0 41320 5 1 1 41319
0 41321 7 1 2 63379 72632
0 41322 5 1 1 41321
0 41323 7 1 2 41320 41322
0 41324 5 1 1 41323
0 41325 7 1 2 59897 41324
0 41326 5 1 1 41325
0 41327 7 1 2 41318 41326
0 41328 5 1 1 41327
0 41329 7 1 2 89598 41328
0 41330 5 1 1 41329
0 41331 7 1 2 41314 41330
0 41332 5 1 1 41331
0 41333 7 1 2 58883 41332
0 41334 5 1 1 41333
0 41335 7 1 2 84300 94572
0 41336 5 1 1 41335
0 41337 7 1 2 91402 93364
0 41338 5 1 1 41337
0 41339 7 1 2 41336 41338
0 41340 5 1 1 41339
0 41341 7 1 2 60153 41340
0 41342 5 1 1 41341
0 41343 7 1 2 79181 90000
0 41344 7 1 2 94466 41343
0 41345 5 1 1 41344
0 41346 7 1 2 41342 41345
0 41347 5 2 1 41346
0 41348 7 1 2 94541 94573
0 41349 5 1 1 41348
0 41350 7 1 2 41334 41349
0 41351 5 1 1 41350
0 41352 7 1 2 66020 41351
0 41353 5 1 1 41352
0 41354 7 1 2 89748 41023
0 41355 5 1 1 41354
0 41356 7 2 2 92885 41355
0 41357 7 1 2 72588 94575
0 41358 5 1 1 41357
0 41359 7 1 2 41353 41358
0 41360 5 1 1 41359
0 41361 7 1 2 66866 41360
0 41362 5 1 1 41361
0 41363 7 1 2 66021 94574
0 41364 5 1 1 41363
0 41365 7 1 2 72441 94576
0 41366 5 1 1 41365
0 41367 7 1 2 41364 41366
0 41368 5 1 1 41367
0 41369 7 1 2 58884 41368
0 41370 5 1 1 41369
0 41371 7 1 2 72442 82289
0 41372 7 1 2 94026 41371
0 41373 7 1 2 94477 41372
0 41374 5 1 1 41373
0 41375 7 1 2 41370 41374
0 41376 5 1 1 41375
0 41377 7 1 2 77274 41376
0 41378 5 1 1 41377
0 41379 7 1 2 41362 41378
0 41380 5 1 1 41379
0 41381 7 1 2 73905 41380
0 41382 5 1 1 41381
0 41383 7 2 2 66612 75551
0 41384 7 2 2 72875 94577
0 41385 5 1 1 94579
0 41386 7 1 2 73385 84576
0 41387 7 1 2 94467 41386
0 41388 5 1 1 41387
0 41389 7 1 2 41385 41388
0 41390 5 1 1 41389
0 41391 7 1 2 57475 41390
0 41392 5 1 1 41391
0 41393 7 1 2 68407 85405
0 41394 5 1 1 41393
0 41395 7 1 2 76346 41394
0 41396 5 1 1 41395
0 41397 7 1 2 71211 84447
0 41398 7 1 2 41396 41397
0 41399 5 1 1 41398
0 41400 7 1 2 41392 41399
0 41401 5 1 1 41400
0 41402 7 1 2 66533 41401
0 41403 5 1 1 41402
0 41404 7 1 2 68037 87672
0 41405 7 1 2 89003 41404
0 41406 5 1 1 41405
0 41407 7 1 2 41403 41406
0 41408 5 1 1 41407
0 41409 7 1 2 66321 41408
0 41410 5 1 1 41409
0 41411 7 1 2 86494 88711
0 41412 7 1 2 71648 41411
0 41413 7 1 2 91007 41412
0 41414 5 1 1 41413
0 41415 7 1 2 41410 41414
0 41416 5 1 1 41415
0 41417 7 1 2 79977 41416
0 41418 5 1 1 41417
0 41419 7 1 2 86804 94342
0 41420 5 1 1 41419
0 41421 7 1 2 57476 89599
0 41422 7 1 2 82961 41421
0 41423 5 1 1 41422
0 41424 7 1 2 41420 41423
0 41425 5 1 1 41424
0 41426 7 1 2 64608 41425
0 41427 5 1 1 41426
0 41428 7 1 2 90006 41427
0 41429 5 1 1 41428
0 41430 7 1 2 73318 94462
0 41431 7 1 2 41429 41430
0 41432 5 1 1 41431
0 41433 7 1 2 41418 41432
0 41434 7 1 2 41382 41433
0 41435 7 1 2 41300 41434
0 41436 7 1 2 41087 41435
0 41437 7 1 2 40921 41436
0 41438 5 1 1 41437
0 41439 7 1 2 66717 41438
0 41440 5 1 1 41439
0 41441 7 1 2 84910 74072
0 41442 5 1 1 41441
0 41443 7 1 2 61397 84902
0 41444 5 1 1 41443
0 41445 7 1 2 57762 41444
0 41446 5 1 1 41445
0 41447 7 1 2 71914 73938
0 41448 5 1 1 41447
0 41449 7 1 2 73958 41448
0 41450 7 1 2 41446 41449
0 41451 5 1 1 41450
0 41452 7 1 2 66322 41451
0 41453 5 1 1 41452
0 41454 7 1 2 41442 41453
0 41455 5 1 1 41454
0 41456 7 1 2 57477 41455
0 41457 5 1 1 41456
0 41458 7 1 2 17729 41457
0 41459 5 1 1 41458
0 41460 7 1 2 93308 94053
0 41461 7 1 2 41459 41460
0 41462 5 1 1 41461
0 41463 7 1 2 41440 41462
0 41464 5 1 1 41463
0 41465 7 1 2 71746 41464
0 41466 5 1 1 41465
0 41467 7 1 2 40608 41466
0 41468 7 1 2 40366 41467
0 41469 7 1 2 39909 41468
0 41470 7 1 2 38587 41469
0 41471 7 1 2 37880 41470
0 41472 5 1 1 41471
0 41473 7 1 2 88344 41472
0 41474 5 1 1 41473
0 41475 7 1 2 59000 73988
0 41476 5 1 1 41475
0 41477 7 2 2 72493 41476
0 41478 5 1 1 94581
0 41479 7 1 2 61398 94582
0 41480 5 1 1 41479
0 41481 7 2 2 57763 86200
0 41482 7 1 2 41480 94583
0 41483 5 1 1 41482
0 41484 7 1 2 92277 41483
0 41485 5 1 1 41484
0 41486 7 1 2 83161 41485
0 41487 5 1 1 41486
0 41488 7 1 2 92792 32749
0 41489 5 1 1 41488
0 41490 7 1 2 69054 41489
0 41491 5 1 1 41490
0 41492 7 2 2 62503 81621
0 41493 5 1 1 94585
0 41494 7 1 2 87997 93020
0 41495 5 1 1 41494
0 41496 7 1 2 78254 86419
0 41497 7 1 2 41495 41496
0 41498 7 1 2 41493 41497
0 41499 7 2 2 41491 41498
0 41500 7 1 2 72658 76428
0 41501 7 1 2 94587 41500
0 41502 5 1 1 41501
0 41503 7 1 2 85020 86296
0 41504 5 1 1 41503
0 41505 7 1 2 28017 41504
0 41506 5 1 1 41505
0 41507 7 1 2 61040 41506
0 41508 5 1 1 41507
0 41509 7 1 2 66022 41508
0 41510 7 1 2 41502 41509
0 41511 5 1 1 41510
0 41512 7 1 2 80825 74994
0 41513 5 1 1 41512
0 41514 7 1 2 57764 41478
0 41515 5 1 1 41514
0 41516 7 1 2 63380 73438
0 41517 7 1 2 41515 41516
0 41518 5 1 1 41517
0 41519 7 1 2 61399 41518
0 41520 5 1 1 41519
0 41521 7 1 2 41513 41520
0 41522 7 1 2 41511 41521
0 41523 5 1 1 41522
0 41524 7 1 2 58782 41523
0 41525 5 1 1 41524
0 41526 7 1 2 41487 41525
0 41527 5 1 1 41526
0 41528 7 1 2 61962 41527
0 41529 5 1 1 41528
0 41530 7 1 2 71831 72195
0 41531 5 1 1 41530
0 41532 7 1 2 71643 82490
0 41533 5 1 1 41532
0 41534 7 1 2 41531 41533
0 41535 5 1 1 41534
0 41536 7 1 2 62247 41535
0 41537 5 1 1 41536
0 41538 7 1 2 87410 82491
0 41539 5 1 1 41538
0 41540 7 1 2 67218 84930
0 41541 5 1 1 41540
0 41542 7 1 2 41539 41541
0 41543 7 1 2 41537 41542
0 41544 5 1 1 41543
0 41545 7 1 2 71312 41544
0 41546 5 1 1 41545
0 41547 7 1 2 71832 91549
0 41548 5 1 1 41547
0 41549 7 1 2 57478 93482
0 41550 5 1 1 41549
0 41551 7 1 2 71440 41550
0 41552 5 1 1 41551
0 41553 7 1 2 41548 41552
0 41554 7 1 2 41546 41553
0 41555 5 1 1 41554
0 41556 7 1 2 63381 41555
0 41557 5 1 1 41556
0 41558 7 2 2 68142 77107
0 41559 5 1 1 94589
0 41560 7 1 2 67375 71517
0 41561 7 1 2 41559 41560
0 41562 5 1 1 41561
0 41563 7 1 2 82928 41562
0 41564 5 1 1 41563
0 41565 7 1 2 61041 77735
0 41566 7 1 2 91181 41565
0 41567 5 1 1 41566
0 41568 7 1 2 41564 41567
0 41569 5 1 1 41568
0 41570 7 1 2 70833 41569
0 41571 5 1 1 41570
0 41572 7 1 2 76342 77108
0 41573 5 2 1 41572
0 41574 7 1 2 83575 75942
0 41575 7 1 2 94591 41574
0 41576 5 1 1 41575
0 41577 7 1 2 80203 85164
0 41578 5 1 1 41577
0 41579 7 1 2 82962 41578
0 41580 5 2 1 41579
0 41581 7 3 2 57765 75943
0 41582 5 2 1 94595
0 41583 7 1 2 94593 94598
0 41584 7 1 2 41576 41583
0 41585 5 1 1 41584
0 41586 7 2 2 86018 78461
0 41587 5 1 1 94600
0 41588 7 1 2 60642 94601
0 41589 5 1 1 41588
0 41590 7 1 2 41585 41589
0 41591 7 1 2 41571 41590
0 41592 7 1 2 41557 41591
0 41593 5 1 1 41592
0 41594 7 1 2 61400 41593
0 41595 5 1 1 41594
0 41596 7 1 2 85497 38746
0 41597 5 1 1 41596
0 41598 7 2 2 61401 75275
0 41599 7 1 2 84803 94602
0 41600 5 1 1 41599
0 41601 7 1 2 76452 90058
0 41602 5 1 1 41601
0 41603 7 1 2 71518 41602
0 41604 5 1 1 41603
0 41605 7 1 2 63382 41604
0 41606 5 1 1 41605
0 41607 7 1 2 41600 41606
0 41608 5 1 1 41607
0 41609 7 1 2 62504 41608
0 41610 5 1 1 41609
0 41611 7 3 2 71695 77475
0 41612 5 1 1 94604
0 41613 7 2 2 59639 41612
0 41614 5 1 1 94607
0 41615 7 1 2 66023 77401
0 41616 5 1 1 41615
0 41617 7 1 2 41614 41616
0 41618 5 1 1 41617
0 41619 7 1 2 87703 28266
0 41620 5 1 1 41619
0 41621 7 1 2 91634 41620
0 41622 5 1 1 41621
0 41623 7 1 2 41618 41622
0 41624 5 1 1 41623
0 41625 7 1 2 63383 41624
0 41626 5 1 1 41625
0 41627 7 1 2 41610 41626
0 41628 5 1 1 41627
0 41629 7 1 2 61042 41628
0 41630 5 1 1 41629
0 41631 7 1 2 85803 84458
0 41632 7 1 2 87279 41631
0 41633 5 1 1 41632
0 41634 7 1 2 41630 41633
0 41635 5 1 1 41634
0 41636 7 1 2 75908 41635
0 41637 5 1 1 41636
0 41638 7 1 2 41597 41637
0 41639 7 1 2 41595 41638
0 41640 5 1 1 41639
0 41641 7 1 2 82619 41640
0 41642 5 1 1 41641
0 41643 7 1 2 41529 41642
0 41644 5 1 1 41643
0 41645 7 1 2 60041 41644
0 41646 5 1 1 41645
0 41647 7 1 2 66024 86433
0 41648 5 1 1 41647
0 41649 7 1 2 79588 41648
0 41650 5 1 1 41649
0 41651 7 1 2 67778 91150
0 41652 5 1 1 41651
0 41653 7 1 2 93774 41652
0 41654 5 1 1 41653
0 41655 7 1 2 62774 41654
0 41656 5 1 1 41655
0 41657 7 1 2 61402 83304
0 41658 5 1 1 41657
0 41659 7 1 2 41656 41658
0 41660 5 1 1 41659
0 41661 7 1 2 64098 41660
0 41662 5 1 1 41661
0 41663 7 1 2 41650 41662
0 41664 5 1 1 41663
0 41665 7 1 2 60643 41664
0 41666 5 1 1 41665
0 41667 7 1 2 91433 94592
0 41668 5 1 1 41667
0 41669 7 1 2 60644 41668
0 41670 5 1 1 41669
0 41671 7 1 2 76343 75488
0 41672 5 1 1 41671
0 41673 7 1 2 67376 41672
0 41674 5 1 1 41673
0 41675 7 1 2 68877 41674
0 41676 5 1 1 41675
0 41677 7 1 2 62505 93314
0 41678 5 1 1 41677
0 41679 7 1 2 62775 86429
0 41680 5 1 1 41679
0 41681 7 1 2 41678 41680
0 41682 7 1 2 41676 41681
0 41683 7 1 2 41670 41682
0 41684 5 1 1 41683
0 41685 7 1 2 61403 41684
0 41686 5 1 1 41685
0 41687 7 1 2 84568 31324
0 41688 5 1 1 41687
0 41689 7 1 2 69055 41688
0 41690 5 1 1 41689
0 41691 7 1 2 66025 26130
0 41692 5 1 1 41691
0 41693 7 1 2 78297 41692
0 41694 5 1 1 41693
0 41695 7 1 2 41690 41694
0 41696 5 1 1 41695
0 41697 7 1 2 61043 41696
0 41698 5 1 1 41697
0 41699 7 2 2 68143 70095
0 41700 5 3 1 94609
0 41701 7 1 2 88025 94610
0 41702 5 1 1 41701
0 41703 7 1 2 67377 41702
0 41704 5 1 1 41703
0 41705 7 1 2 61404 41704
0 41706 5 1 1 41705
0 41707 7 1 2 41698 41706
0 41708 5 1 1 41707
0 41709 7 1 2 63914 41708
0 41710 5 1 1 41709
0 41711 7 1 2 62776 83571
0 41712 5 1 1 41711
0 41713 7 1 2 25346 41712
0 41714 5 1 1 41713
0 41715 7 1 2 75489 41714
0 41716 5 1 1 41715
0 41717 7 1 2 80449 41716
0 41718 5 1 1 41717
0 41719 7 1 2 75909 41718
0 41720 5 1 1 41719
0 41721 7 1 2 41710 41720
0 41722 7 1 2 41686 41721
0 41723 7 2 2 41666 41722
0 41724 5 1 1 94614
0 41725 7 1 2 58783 41724
0 41726 5 1 1 41725
0 41727 7 1 2 74484 77195
0 41728 7 1 2 78462 41727
0 41729 5 1 1 41728
0 41730 7 1 2 41726 41729
0 41731 5 1 1 41730
0 41732 7 1 2 71313 41731
0 41733 5 1 1 41732
0 41734 7 2 2 89032 94150
0 41735 5 1 1 94616
0 41736 7 1 2 61044 41735
0 41737 5 1 1 41736
0 41738 7 2 2 78733 93697
0 41739 5 1 1 94618
0 41740 7 1 2 87037 94619
0 41741 5 1 1 41740
0 41742 7 1 2 93797 41741
0 41743 5 1 1 41742
0 41744 7 1 2 41737 41743
0 41745 5 1 1 41744
0 41746 7 1 2 58784 41745
0 41747 5 1 1 41746
0 41748 7 1 2 73319 94309
0 41749 5 1 1 41748
0 41750 7 1 2 41747 41749
0 41751 5 1 1 41750
0 41752 7 1 2 71441 41751
0 41753 5 1 1 41752
0 41754 7 1 2 41733 41753
0 41755 5 1 1 41754
0 41756 7 1 2 63384 41755
0 41757 5 1 1 41756
0 41758 7 1 2 87694 94066
0 41759 5 1 1 41758
0 41760 7 1 2 68144 41759
0 41761 5 1 1 41760
0 41762 7 2 2 68145 83884
0 41763 5 1 1 94620
0 41764 7 1 2 59380 83342
0 41765 5 1 1 41764
0 41766 7 1 2 68257 41765
0 41767 5 1 1 41766
0 41768 7 1 2 41763 41767
0 41769 5 1 1 41768
0 41770 7 1 2 62248 41769
0 41771 5 1 1 41770
0 41772 7 1 2 71212 13511
0 41773 5 2 1 41772
0 41774 7 1 2 74381 94622
0 41775 5 1 1 41774
0 41776 7 1 2 67219 83448
0 41777 5 1 1 41776
0 41778 7 1 2 63081 83359
0 41779 5 1 1 41778
0 41780 7 1 2 41777 41779
0 41781 7 1 2 41775 41780
0 41782 7 1 2 41771 41781
0 41783 7 1 2 41761 41782
0 41784 5 1 1 41783
0 41785 7 1 2 66026 41784
0 41786 5 1 1 41785
0 41787 7 1 2 79599 87741
0 41788 5 1 1 41787
0 41789 7 1 2 65679 86990
0 41790 7 1 2 41788 41789
0 41791 7 1 2 41786 41790
0 41792 5 1 1 41791
0 41793 7 1 2 62777 41739
0 41794 5 1 1 41793
0 41795 7 2 2 94617 41794
0 41796 5 1 1 94624
0 41797 7 2 2 58337 94625
0 41798 5 1 1 94626
0 41799 7 1 2 66027 94627
0 41800 5 1 1 41799
0 41801 7 1 2 59640 14191
0 41802 7 1 2 41800 41801
0 41803 5 1 1 41802
0 41804 7 1 2 69828 74078
0 41805 5 1 1 41804
0 41806 7 2 2 73695 41805
0 41807 7 1 2 68786 94628
0 41808 5 1 1 41807
0 41809 7 1 2 61045 27728
0 41810 7 1 2 41808 41809
0 41811 7 1 2 41803 41810
0 41812 5 1 1 41811
0 41813 7 1 2 41792 41812
0 41814 5 1 1 41813
0 41815 7 1 2 73473 93546
0 41816 5 1 1 41815
0 41817 7 1 2 69724 41816
0 41818 5 1 1 41817
0 41819 7 1 2 73096 41818
0 41820 5 1 1 41819
0 41821 7 1 2 85770 17803
0 41822 7 1 2 41820 41821
0 41823 7 1 2 41814 41822
0 41824 5 1 1 41823
0 41825 7 1 2 63520 41824
0 41826 5 1 1 41825
0 41827 7 6 2 58785 61405
0 41828 5 4 1 94630
0 41829 7 1 2 85165 94631
0 41830 7 1 2 93677 41829
0 41831 5 1 1 41830
0 41832 7 1 2 41826 41831
0 41833 7 1 2 41757 41832
0 41834 5 1 1 41833
0 41835 7 1 2 64727 41834
0 41836 5 1 1 41835
0 41837 7 1 2 92369 92844
0 41838 5 1 1 41837
0 41839 7 1 2 93322 41838
0 41840 5 1 1 41839
0 41841 7 1 2 63915 41840
0 41842 5 1 1 41841
0 41843 7 1 2 71442 87398
0 41844 5 1 1 41843
0 41845 7 1 2 41842 41844
0 41846 5 1 1 41845
0 41847 7 1 2 62506 41846
0 41848 5 1 1 41847
0 41849 7 1 2 70834 87393
0 41850 5 1 1 41849
0 41851 7 1 2 75910 75188
0 41852 5 1 1 41851
0 41853 7 1 2 41850 41852
0 41854 5 1 1 41853
0 41855 7 1 2 71443 41854
0 41856 5 1 1 41855
0 41857 7 1 2 41848 41856
0 41858 5 1 1 41857
0 41859 7 1 2 62778 41858
0 41860 5 1 1 41859
0 41861 7 1 2 81800 93693
0 41862 5 1 1 41861
0 41863 7 1 2 59157 89215
0 41864 5 1 1 41863
0 41865 7 1 2 59381 81617
0 41866 5 3 1 41865
0 41867 7 1 2 62249 94640
0 41868 7 1 2 41864 41867
0 41869 5 1 1 41868
0 41870 7 1 2 41862 41869
0 41871 5 1 1 41870
0 41872 7 1 2 62507 41871
0 41873 5 1 1 41872
0 41874 7 1 2 64099 92824
0 41875 5 1 1 41874
0 41876 7 3 2 41873 41875
0 41877 5 2 1 94643
0 41878 7 1 2 71444 94646
0 41879 5 1 1 41878
0 41880 7 1 2 41860 41879
0 41881 5 1 1 41880
0 41882 7 1 2 86042 74195
0 41883 7 1 2 41881 41882
0 41884 5 1 1 41883
0 41885 7 1 2 41836 41884
0 41886 5 1 1 41885
0 41887 7 1 2 66613 41886
0 41888 5 1 1 41887
0 41889 7 1 2 41646 41888
0 41890 5 1 1 41889
0 41891 7 1 2 64609 41890
0 41892 5 1 1 41891
0 41893 7 1 2 73474 75684
0 41894 7 1 2 85278 41893
0 41895 5 1 1 41894
0 41896 7 2 2 79169 82620
0 41897 7 1 2 85508 18336
0 41898 7 1 2 94648 41897
0 41899 5 1 1 41898
0 41900 7 1 2 41895 41899
0 41901 5 1 1 41900
0 41902 7 1 2 64728 41901
0 41903 5 1 1 41902
0 41904 7 1 2 79032 38284
0 41905 5 1 1 41904
0 41906 7 1 2 86923 41905
0 41907 5 1 1 41906
0 41908 7 1 2 92030 32796
0 41909 7 1 2 41907 41908
0 41910 5 1 1 41909
0 41911 7 1 2 73475 75961
0 41912 7 1 2 41910 41911
0 41913 5 1 1 41912
0 41914 7 1 2 41903 41913
0 41915 5 1 1 41914
0 41916 7 1 2 57766 41915
0 41917 5 1 1 41916
0 41918 7 1 2 63521 83176
0 41919 5 9 1 41918
0 41920 7 1 2 93913 94491
0 41921 7 1 2 94650 41920
0 41922 5 1 1 41921
0 41923 7 1 2 41917 41922
0 41924 5 1 1 41923
0 41925 7 1 2 65078 41924
0 41926 5 1 1 41925
0 41927 7 1 2 73970 94056
0 41928 5 2 1 41927
0 41929 7 1 2 78923 75552
0 41930 5 3 1 41929
0 41931 7 1 2 58786 94661
0 41932 5 1 1 41931
0 41933 7 1 2 94659 41932
0 41934 5 2 1 41933
0 41935 7 1 2 64729 94664
0 41936 5 1 1 41935
0 41937 7 1 2 79863 94662
0 41938 5 1 1 41937
0 41939 7 1 2 41936 41938
0 41940 5 3 1 41939
0 41941 7 2 2 86759 87106
0 41942 7 1 2 94666 94669
0 41943 5 1 1 41942
0 41944 7 1 2 83162 91697
0 41945 5 1 1 41944
0 41946 7 3 2 59641 77218
0 41947 7 1 2 66614 74657
0 41948 7 1 2 94671 41947
0 41949 5 1 1 41948
0 41950 7 1 2 41945 41949
0 41951 5 1 1 41950
0 41952 7 1 2 79985 41951
0 41953 5 1 1 41952
0 41954 7 1 2 41943 41953
0 41955 7 1 2 41926 41954
0 41956 5 1 1 41955
0 41957 7 1 2 68631 41956
0 41958 5 1 1 41957
0 41959 7 1 2 68439 84082
0 41960 5 2 1 41959
0 41961 7 1 2 93767 94674
0 41962 5 2 1 41961
0 41963 7 1 2 65680 94676
0 41964 5 1 1 41963
0 41965 7 1 2 68038 78826
0 41966 5 1 1 41965
0 41967 7 1 2 61046 41966
0 41968 5 1 1 41967
0 41969 7 1 2 67678 41968
0 41970 5 1 1 41969
0 41971 7 1 2 81071 78412
0 41972 5 1 1 41971
0 41973 7 1 2 75011 41972
0 41974 7 1 2 41970 41973
0 41975 5 1 1 41974
0 41976 7 1 2 41964 41975
0 41977 5 1 1 41976
0 41978 7 1 2 85166 41977
0 41979 5 1 1 41978
0 41980 7 2 2 68146 88953
0 41981 5 1 1 94678
0 41982 7 1 2 12984 41981
0 41983 5 1 1 41982
0 41984 7 1 2 61047 41983
0 41985 5 1 1 41984
0 41986 7 2 2 78245 75189
0 41987 5 1 1 94680
0 41988 7 1 2 78803 94681
0 41989 5 1 1 41988
0 41990 7 1 2 41985 41989
0 41991 5 1 1 41990
0 41992 7 1 2 67779 41991
0 41993 5 1 1 41992
0 41994 7 1 2 62250 77074
0 41995 7 1 2 93847 41994
0 41996 5 2 1 41995
0 41997 7 1 2 69428 76362
0 41998 5 1 1 41997
0 41999 7 1 2 94682 41998
0 42000 5 1 1 41999
0 42001 7 1 2 68147 42000
0 42002 5 1 1 42001
0 42003 7 1 2 75033 84083
0 42004 5 1 1 42003
0 42005 7 1 2 42002 42004
0 42006 5 1 1 42005
0 42007 7 1 2 68258 42006
0 42008 5 1 1 42007
0 42009 7 1 2 65079 72615
0 42010 5 1 1 42009
0 42011 7 1 2 94683 42010
0 42012 5 1 1 42011
0 42013 7 1 2 67220 42012
0 42014 5 1 1 42013
0 42015 7 1 2 42008 42014
0 42016 7 1 2 41993 42015
0 42017 5 1 1 42016
0 42018 7 1 2 71314 42017
0 42019 5 1 1 42018
0 42020 7 1 2 41979 42019
0 42021 5 1 1 42020
0 42022 7 1 2 66867 42021
0 42023 5 1 1 42022
0 42024 7 1 2 71315 90108
0 42025 5 1 1 42024
0 42026 7 1 2 83163 66928
0 42027 5 1 1 42026
0 42028 7 1 2 42025 42027
0 42029 5 1 1 42028
0 42030 7 1 2 75012 42029
0 42031 5 1 1 42030
0 42032 7 1 2 85254 92353
0 42033 5 1 1 42032
0 42034 7 2 2 64730 94651
0 42035 7 4 2 78910 91829
0 42036 5 2 1 94686
0 42037 7 1 2 73431 73841
0 42038 5 1 1 42037
0 42039 7 1 2 94690 42038
0 42040 5 1 1 42039
0 42041 7 1 2 94684 42040
0 42042 5 1 1 42041
0 42043 7 1 2 42033 42042
0 42044 5 1 1 42043
0 42045 7 1 2 57767 42044
0 42046 5 1 1 42045
0 42047 7 1 2 42031 42046
0 42048 7 1 2 42023 42047
0 42049 5 1 1 42048
0 42050 7 1 2 66028 42049
0 42051 5 1 1 42050
0 42052 7 1 2 84639 78657
0 42053 5 1 1 42052
0 42054 7 1 2 94064 42053
0 42055 5 1 1 42054
0 42056 7 1 2 76493 92925
0 42057 5 1 1 42056
0 42058 7 1 2 85710 82847
0 42059 7 1 2 42057 42058
0 42060 5 1 1 42059
0 42061 7 1 2 61048 42060
0 42062 5 1 1 42061
0 42063 7 1 2 85034 94623
0 42064 5 1 1 42063
0 42065 7 1 2 42062 42064
0 42066 7 1 2 42055 42065
0 42067 5 1 1 42066
0 42068 7 1 2 61406 42067
0 42069 5 1 1 42068
0 42070 7 1 2 61407 76357
0 42071 5 2 1 42070
0 42072 7 1 2 57479 94692
0 42073 5 1 1 42072
0 42074 7 1 2 88067 94108
0 42075 7 1 2 42073 42074
0 42076 5 1 1 42075
0 42077 7 1 2 88075 94111
0 42078 5 1 1 42077
0 42079 7 1 2 85484 86201
0 42080 5 1 1 42079
0 42081 7 1 2 42078 42080
0 42082 7 1 2 42076 42081
0 42083 7 1 2 42069 42082
0 42084 5 1 1 42083
0 42085 7 1 2 79268 42084
0 42086 5 1 1 42085
0 42087 7 3 2 86315 83924
0 42088 7 1 2 69879 82337
0 42089 7 1 2 94694 42088
0 42090 5 1 1 42089
0 42091 7 1 2 42086 42090
0 42092 5 1 1 42091
0 42093 7 1 2 58787 42092
0 42094 5 1 1 42093
0 42095 7 1 2 67595 92902
0 42096 5 1 1 42095
0 42097 7 1 2 73439 42096
0 42098 5 1 1 42097
0 42099 7 4 2 85291 79906
0 42100 5 2 1 94697
0 42101 7 1 2 92355 94701
0 42102 5 1 1 42101
0 42103 7 1 2 85829 42102
0 42104 5 1 1 42103
0 42105 7 1 2 85292 92154
0 42106 5 2 1 42105
0 42107 7 1 2 69821 87502
0 42108 5 1 1 42107
0 42109 7 1 2 94691 42108
0 42110 5 1 1 42109
0 42111 7 1 2 94685 42110
0 42112 5 1 1 42111
0 42113 7 1 2 94703 42112
0 42114 7 1 2 42104 42113
0 42115 5 1 1 42114
0 42116 7 1 2 42098 42115
0 42117 5 1 1 42116
0 42118 7 1 2 59898 23965
0 42119 5 1 1 42118
0 42120 7 1 2 82480 42119
0 42121 5 1 1 42120
0 42122 7 1 2 66029 42121
0 42123 5 1 1 42122
0 42124 7 3 2 59001 72032
0 42125 5 1 1 94705
0 42126 7 1 2 93952 94706
0 42127 5 1 1 42126
0 42128 7 1 2 42123 42127
0 42129 5 1 1 42128
0 42130 7 1 2 94698 42129
0 42131 5 1 1 42130
0 42132 7 1 2 61963 42131
0 42133 7 1 2 42117 42132
0 42134 7 1 2 42094 42133
0 42135 7 1 2 42051 42134
0 42136 5 1 1 42135
0 42137 7 1 2 66880 86682
0 42138 7 1 2 85077 42137
0 42139 5 1 1 42138
0 42140 7 1 2 4520 42139
0 42141 5 2 1 42140
0 42142 7 1 2 84416 94708
0 42143 5 1 1 42142
0 42144 7 1 2 71316 79038
0 42145 5 2 1 42144
0 42146 7 1 2 42143 94710
0 42147 5 1 1 42146
0 42148 7 1 2 78872 42147
0 42149 5 1 1 42148
0 42150 7 1 2 81168 79039
0 42151 5 1 1 42150
0 42152 7 1 2 42149 42151
0 42153 5 1 1 42152
0 42154 7 1 2 60645 42153
0 42155 5 1 1 42154
0 42156 7 1 2 85132 93324
0 42157 5 1 1 42156
0 42158 7 1 2 79040 42157
0 42159 5 1 1 42158
0 42160 7 1 2 42155 42159
0 42161 5 1 1 42160
0 42162 7 1 2 70218 42161
0 42163 5 1 1 42162
0 42164 7 4 2 84565 87787
0 42165 7 2 2 79852 94712
0 42166 7 1 2 61049 94716
0 42167 5 1 1 42166
0 42168 7 1 2 68148 34435
0 42169 5 1 1 42168
0 42170 7 1 2 81673 90166
0 42171 5 1 1 42170
0 42172 7 1 2 88775 42171
0 42173 5 1 1 42172
0 42174 7 1 2 58629 90560
0 42175 7 1 2 93788 42174
0 42176 7 1 2 42173 42175
0 42177 7 1 2 42169 42176
0 42178 5 1 1 42177
0 42179 7 1 2 71317 42178
0 42180 5 1 1 42179
0 42181 7 1 2 85167 93655
0 42182 5 1 1 42181
0 42183 7 1 2 93289 42182
0 42184 7 1 2 42180 42183
0 42185 5 1 1 42184
0 42186 7 1 2 79828 42185
0 42187 5 1 1 42186
0 42188 7 1 2 42167 42187
0 42189 5 1 1 42188
0 42190 7 1 2 63522 42189
0 42191 5 1 1 42190
0 42192 7 1 2 75375 79027
0 42193 7 1 2 90748 42192
0 42194 5 1 1 42193
0 42195 7 2 2 73132 94709
0 42196 5 1 1 94718
0 42197 7 1 2 77698 94719
0 42198 5 1 1 42197
0 42199 7 1 2 42194 42198
0 42200 5 1 1 42199
0 42201 7 1 2 62251 42200
0 42202 5 1 1 42201
0 42203 7 1 2 85133 34503
0 42204 5 1 1 42203
0 42205 7 1 2 79041 42204
0 42206 5 1 1 42205
0 42207 7 1 2 42202 42206
0 42208 5 1 1 42207
0 42209 7 1 2 69056 42208
0 42210 5 1 1 42209
0 42211 7 2 2 78086 94713
0 42212 7 1 2 74467 94720
0 42213 5 1 1 42212
0 42214 7 1 2 62779 88001
0 42215 5 1 1 42214
0 42216 7 1 2 92755 42215
0 42217 5 1 1 42216
0 42218 7 1 2 42196 94711
0 42219 5 1 1 42218
0 42220 7 1 2 42217 42219
0 42221 5 1 1 42220
0 42222 7 1 2 42213 42221
0 42223 7 1 2 42210 42222
0 42224 7 1 2 42191 42223
0 42225 7 1 2 42163 42224
0 42226 5 1 1 42225
0 42227 7 1 2 61408 42226
0 42228 5 1 1 42227
0 42229 7 1 2 79340 85485
0 42230 5 1 1 42229
0 42231 7 2 2 68149 85168
0 42232 5 1 1 94722
0 42233 7 1 2 73320 94723
0 42234 5 1 1 42233
0 42235 7 1 2 42230 42234
0 42236 5 1 1 42235
0 42237 7 1 2 94156 42236
0 42238 5 1 1 42237
0 42239 7 1 2 74729 74196
0 42240 5 1 1 42239
0 42241 7 1 2 25850 93735
0 42242 5 1 1 42241
0 42243 7 1 2 62252 93464
0 42244 5 2 1 42243
0 42245 7 1 2 76312 94724
0 42246 5 1 1 42245
0 42247 7 1 2 42242 42246
0 42248 5 1 1 42247
0 42249 7 1 2 42240 42248
0 42250 7 1 2 63082 92797
0 42251 5 1 1 42250
0 42252 7 1 2 58630 42251
0 42253 5 1 1 42252
0 42254 7 1 2 73341 79351
0 42255 5 1 1 42254
0 42256 7 1 2 63385 76310
0 42257 5 1 1 42256
0 42258 7 1 2 57480 42257
0 42259 5 1 1 42258
0 42260 7 1 2 42255 42259
0 42261 7 1 2 42253 42260
0 42262 5 1 1 42261
0 42263 7 2 2 62780 85169
0 42264 5 1 1 94726
0 42265 7 1 2 78750 94727
0 42266 5 1 1 42265
0 42267 7 1 2 92384 93501
0 42268 5 1 1 42267
0 42269 7 1 2 82963 42268
0 42270 7 1 2 42266 42269
0 42271 5 1 1 42270
0 42272 7 1 2 70219 73638
0 42273 7 1 2 79991 42272
0 42274 7 1 2 42271 42273
0 42275 5 1 1 42274
0 42276 7 1 2 42262 42275
0 42277 7 1 2 42249 42276
0 42278 7 1 2 42238 42277
0 42279 5 1 1 42278
0 42280 7 1 2 66787 42279
0 42281 5 1 1 42280
0 42282 7 1 2 66615 42281
0 42283 7 1 2 42228 42282
0 42284 5 1 1 42283
0 42285 7 1 2 42136 42284
0 42286 5 1 1 42285
0 42287 7 1 2 41958 42286
0 42288 7 1 2 41892 42287
0 42289 5 1 1 42288
0 42290 7 1 2 82184 88296
0 42291 7 1 2 42289 42290
0 42292 5 1 1 42291
0 42293 7 3 2 67959 88297
0 42294 7 1 2 19526 93825
0 42295 5 3 1 42294
0 42296 7 1 2 59158 78102
0 42297 7 1 2 94731 42296
0 42298 5 1 1 42297
0 42299 7 2 2 70305 75578
0 42300 5 1 1 94734
0 42301 7 1 2 66030 42300
0 42302 7 1 2 42298 42301
0 42303 5 1 1 42302
0 42304 7 1 2 61409 80775
0 42305 5 1 1 42304
0 42306 7 1 2 79907 42305
0 42307 7 1 2 42303 42306
0 42308 5 1 1 42307
0 42309 7 1 2 70784 87578
0 42310 7 1 2 94041 42309
0 42311 7 1 2 85279 42310
0 42312 7 1 2 94732 42311
0 42313 5 1 1 42312
0 42314 7 1 2 42308 42313
0 42315 5 1 1 42314
0 42316 7 1 2 94728 42315
0 42317 5 1 1 42316
0 42318 7 2 2 91106 91205
0 42319 7 2 2 94517 94736
0 42320 7 2 2 66031 94038
0 42321 7 1 2 92287 94740
0 42322 7 1 2 94738 42321
0 42323 5 1 1 42322
0 42324 7 1 2 61410 94729
0 42325 7 1 2 94667 42324
0 42326 5 1 1 42325
0 42327 7 1 2 42323 42326
0 42328 5 1 1 42327
0 42329 7 1 2 90561 42328
0 42330 5 1 1 42329
0 42331 7 1 2 42317 42330
0 42332 5 1 1 42331
0 42333 7 1 2 59642 42332
0 42334 5 1 1 42333
0 42335 7 1 2 76691 81146
0 42336 5 1 1 42335
0 42337 7 1 2 58338 42336
0 42338 5 1 1 42337
0 42339 7 1 2 59899 90854
0 42340 5 1 1 42339
0 42341 7 2 2 42338 42340
0 42342 7 1 2 62781 94742
0 42343 5 1 1 42342
0 42344 7 1 2 71519 76656
0 42345 5 6 1 42344
0 42346 7 1 2 81088 94744
0 42347 7 1 2 85572 42346
0 42348 5 1 1 42347
0 42349 7 1 2 42343 42348
0 42350 5 1 1 42349
0 42351 7 1 2 78873 42350
0 42352 5 1 1 42351
0 42353 7 1 2 65681 75891
0 42354 5 1 1 42353
0 42355 7 1 2 78874 42354
0 42356 5 1 1 42355
0 42357 7 1 2 62508 12936
0 42358 5 1 1 42357
0 42359 7 1 2 73923 34592
0 42360 7 1 2 42358 42359
0 42361 7 1 2 42356 42360
0 42362 5 1 1 42361
0 42363 7 1 2 85216 42362
0 42364 5 1 1 42363
0 42365 7 1 2 93674 94745
0 42366 5 1 1 42365
0 42367 7 1 2 42364 42366
0 42368 7 1 2 42352 42367
0 42369 5 1 1 42368
0 42370 7 1 2 66868 42369
0 42371 5 1 1 42370
0 42372 7 1 2 93900 94427
0 42373 5 1 1 42372
0 42374 7 1 2 57768 42373
0 42375 5 2 1 42374
0 42376 7 1 2 72480 88887
0 42377 5 1 1 42376
0 42378 7 1 2 94750 42377
0 42379 5 2 1 42378
0 42380 7 1 2 92155 94752
0 42381 5 1 1 42380
0 42382 7 1 2 61411 42381
0 42383 7 1 2 42371 42382
0 42384 5 1 1 42383
0 42385 7 1 2 80274 75024
0 42386 5 1 1 42385
0 42387 7 1 2 91605 42386
0 42388 5 1 1 42387
0 42389 7 1 2 62782 42388
0 42390 5 1 1 42389
0 42391 7 1 2 61050 88636
0 42392 5 1 1 42391
0 42393 7 1 2 42390 42392
0 42394 5 1 1 42393
0 42395 7 1 2 71318 42394
0 42396 5 1 1 42395
0 42397 7 1 2 80275 78671
0 42398 5 1 1 42397
0 42399 7 1 2 42396 42398
0 42400 5 1 1 42399
0 42401 7 1 2 62509 42400
0 42402 5 1 1 42401
0 42403 7 1 2 36813 42402
0 42404 5 1 1 42403
0 42405 7 1 2 70835 42404
0 42406 5 1 1 42405
0 42407 7 1 2 76771 78048
0 42408 5 1 1 42407
0 42409 7 1 2 78673 42408
0 42410 5 1 1 42409
0 42411 7 1 2 63786 42410
0 42412 5 1 1 42411
0 42413 7 1 2 60406 79705
0 42414 5 1 1 42413
0 42415 7 1 2 42412 42414
0 42416 5 1 1 42415
0 42417 7 1 2 62253 42416
0 42418 5 1 1 42417
0 42419 7 1 2 78298 79706
0 42420 5 1 1 42419
0 42421 7 1 2 42418 42420
0 42422 5 1 1 42421
0 42423 7 1 2 75911 42422
0 42424 5 1 1 42423
0 42425 7 1 2 85350 94590
0 42426 5 1 1 42425
0 42427 7 1 2 75339 42426
0 42428 5 1 1 42427
0 42429 7 1 2 71319 42428
0 42430 5 1 1 42429
0 42431 7 1 2 71445 93189
0 42432 5 1 1 42431
0 42433 7 1 2 42430 42432
0 42434 5 1 1 42433
0 42435 7 1 2 72153 42434
0 42436 5 1 1 42435
0 42437 7 1 2 93172 94101
0 42438 5 1 1 42437
0 42439 7 1 2 93221 42438
0 42440 7 1 2 42436 42439
0 42441 7 1 2 42424 42440
0 42442 7 1 2 42406 42441
0 42443 5 1 1 42442
0 42444 7 1 2 85095 42443
0 42445 5 1 1 42444
0 42446 7 2 2 86316 83062
0 42447 7 1 2 70332 82633
0 42448 7 1 2 94754 42447
0 42449 5 1 1 42448
0 42450 7 1 2 42445 42449
0 42451 5 1 1 42450
0 42452 7 1 2 59900 42451
0 42453 5 1 1 42452
0 42454 7 1 2 59901 76817
0 42455 5 1 1 42454
0 42456 7 1 2 80776 42455
0 42457 5 1 1 42456
0 42458 7 1 2 61051 42457
0 42459 5 1 1 42458
0 42460 7 1 2 68039 77182
0 42461 5 1 1 42460
0 42462 7 1 2 73386 42461
0 42463 5 1 1 42462
0 42464 7 1 2 42459 42463
0 42465 5 1 1 42464
0 42466 7 1 2 60646 42465
0 42467 5 1 1 42466
0 42468 7 2 2 64610 85293
0 42469 5 1 1 94756
0 42470 7 1 2 59902 84487
0 42471 5 1 1 42470
0 42472 7 1 2 42469 42471
0 42473 5 1 1 42472
0 42474 7 1 2 70333 42473
0 42475 5 1 1 42474
0 42476 7 2 2 59382 79112
0 42477 7 1 2 69194 94758
0 42478 5 1 1 42477
0 42479 7 1 2 65306 42478
0 42480 5 1 1 42479
0 42481 7 2 2 93162 42480
0 42482 7 1 2 61052 94760
0 42483 5 1 1 42482
0 42484 7 1 2 78649 93586
0 42485 5 1 1 42484
0 42486 7 1 2 83413 42485
0 42487 5 1 1 42486
0 42488 7 1 2 59903 42487
0 42489 7 1 2 42483 42488
0 42490 5 1 1 42489
0 42491 7 1 2 42475 42490
0 42492 7 1 2 42467 42491
0 42493 5 1 1 42492
0 42494 7 1 2 66929 42493
0 42495 5 1 1 42494
0 42496 7 1 2 66032 42495
0 42497 7 1 2 42453 42496
0 42498 5 1 1 42497
0 42499 7 1 2 42384 42498
0 42500 5 1 1 42499
0 42501 7 1 2 61412 94753
0 42502 5 1 1 42501
0 42503 7 1 2 86883 73532
0 42504 5 1 1 42503
0 42505 7 1 2 42502 42504
0 42506 5 1 1 42505
0 42507 7 1 2 78911 87164
0 42508 5 1 1 42507
0 42509 7 1 2 94702 42508
0 42510 5 1 1 42509
0 42511 7 1 2 42506 42510
0 42512 5 1 1 42511
0 42513 7 1 2 78875 81236
0 42514 5 2 1 42513
0 42515 7 1 2 67780 82465
0 42516 5 1 1 42515
0 42517 7 1 2 94762 42516
0 42518 5 1 1 42517
0 42519 7 1 2 85486 42518
0 42520 5 1 1 42519
0 42521 7 1 2 91177 42520
0 42522 5 1 1 42521
0 42523 7 1 2 64611 42522
0 42524 5 1 1 42523
0 42525 7 2 2 64612 85170
0 42526 5 1 1 94764
0 42527 7 1 2 59904 89931
0 42528 5 1 1 42527
0 42529 7 1 2 77037 81160
0 42530 7 1 2 42528 42529
0 42531 5 1 1 42530
0 42532 7 1 2 42526 42531
0 42533 5 1 1 42532
0 42534 7 1 2 84084 42533
0 42535 5 1 1 42534
0 42536 7 1 2 60407 91399
0 42537 5 1 1 42536
0 42538 7 1 2 25653 42537
0 42539 5 1 1 42538
0 42540 7 1 2 75838 78049
0 42541 7 1 2 42539 42540
0 42542 5 1 1 42541
0 42543 7 1 2 76284 94765
0 42544 5 1 1 42543
0 42545 7 1 2 42542 42544
0 42546 7 1 2 42535 42545
0 42547 5 1 1 42546
0 42548 7 1 2 68150 42547
0 42549 5 1 1 42548
0 42550 7 1 2 42524 42549
0 42551 5 1 1 42550
0 42552 7 1 2 66869 42551
0 42553 5 1 1 42552
0 42554 7 1 2 78668 6337
0 42555 5 1 1 42554
0 42556 7 1 2 76692 66870
0 42557 7 1 2 42555 42556
0 42558 5 1 1 42557
0 42559 7 1 2 88040 42558
0 42560 5 1 1 42559
0 42561 7 1 2 72961 42560
0 42562 5 1 1 42561
0 42563 7 1 2 61964 42562
0 42564 7 1 2 42553 42563
0 42565 7 1 2 42512 42564
0 42566 7 1 2 42500 42565
0 42567 5 1 1 42566
0 42568 7 3 2 62112 88298
0 42569 7 1 2 71213 93319
0 42570 7 1 2 92911 42569
0 42571 5 1 1 42570
0 42572 7 1 2 62254 42571
0 42573 5 1 1 42572
0 42574 7 1 2 61053 75839
0 42575 5 1 1 42574
0 42576 7 1 2 42573 42575
0 42577 5 1 1 42576
0 42578 7 1 2 69057 42577
0 42579 5 1 1 42578
0 42580 7 1 2 73888 93021
0 42581 5 1 1 42580
0 42582 7 1 2 71214 42581
0 42583 5 1 1 42582
0 42584 7 1 2 76332 86756
0 42585 5 1 1 42584
0 42586 7 1 2 63083 42585
0 42587 5 1 1 42586
0 42588 7 1 2 87988 42587
0 42589 5 1 1 42588
0 42590 7 1 2 42583 42589
0 42591 5 1 1 42590
0 42592 7 2 2 65682 69804
0 42593 5 1 1 94769
0 42594 7 1 2 67378 94770
0 42595 5 1 1 42594
0 42596 7 1 2 84549 42595
0 42597 5 1 1 42596
0 42598 7 1 2 64393 10600
0 42599 5 1 1 42598
0 42600 7 1 2 78612 42599
0 42601 7 1 2 42597 42600
0 42602 7 1 2 42591 42601
0 42603 7 1 2 83925 94416
0 42604 5 1 1 42603
0 42605 7 1 2 61413 42604
0 42606 5 1 1 42605
0 42607 7 1 2 83956 81622
0 42608 5 1 1 42607
0 42609 7 1 2 68151 76379
0 42610 5 1 1 42609
0 42611 7 1 2 42608 42610
0 42612 5 1 1 42611
0 42613 7 1 2 62510 42612
0 42614 5 1 1 42613
0 42615 7 1 2 42606 42614
0 42616 7 1 2 42602 42615
0 42617 7 1 2 42579 42616
0 42618 5 1 1 42617
0 42619 7 1 2 75553 42618
0 42620 5 1 1 42619
0 42621 7 1 2 85021 72481
0 42622 5 1 1 42621
0 42623 7 1 2 71446 42622
0 42624 5 1 1 42623
0 42625 7 1 2 83957 94157
0 42626 5 1 1 42625
0 42627 7 1 2 78751 81305
0 42628 5 1 1 42627
0 42629 7 1 2 78613 80947
0 42630 7 1 2 42628 42629
0 42631 7 1 2 42626 42630
0 42632 5 1 1 42631
0 42633 7 1 2 71320 42632
0 42634 5 1 1 42633
0 42635 7 1 2 42624 42634
0 42636 5 1 1 42635
0 42637 7 1 2 61414 42636
0 42638 5 1 1 42637
0 42639 7 1 2 68152 78595
0 42640 5 1 1 42639
0 42641 7 2 2 67379 42640
0 42642 5 1 1 94771
0 42643 7 1 2 71447 42642
0 42644 5 1 1 42643
0 42645 7 1 2 71520 83474
0 42646 5 1 1 42645
0 42647 7 1 2 92372 42646
0 42648 5 1 1 42647
0 42649 7 1 2 84323 42648
0 42650 5 1 1 42649
0 42651 7 1 2 75103 42650
0 42652 5 1 1 42651
0 42653 7 1 2 71521 83592
0 42654 5 1 1 42653
0 42655 7 1 2 71321 42654
0 42656 7 1 2 79589 42655
0 42657 5 1 1 42656
0 42658 7 1 2 20618 89784
0 42659 7 1 2 84377 42658
0 42660 5 1 1 42659
0 42661 7 1 2 42657 42660
0 42662 7 1 2 42652 42661
0 42663 7 1 2 42644 42662
0 42664 5 1 1 42663
0 42665 7 1 2 61054 42664
0 42666 5 2 1 42665
0 42667 7 1 2 77736 92769
0 42668 5 1 1 42667
0 42669 7 2 2 70836 80276
0 42670 5 1 1 94775
0 42671 7 1 2 90728 94776
0 42672 5 1 1 42671
0 42673 7 1 2 73906 42672
0 42674 7 1 2 42668 42673
0 42675 5 2 1 42674
0 42676 7 1 2 71448 94777
0 42677 5 1 1 42676
0 42678 7 1 2 94773 42677
0 42679 7 1 2 42638 42678
0 42680 5 1 1 42679
0 42681 7 1 2 76693 42680
0 42682 5 1 1 42681
0 42683 7 1 2 42620 42682
0 42684 5 1 1 42683
0 42685 7 1 2 66788 42684
0 42686 5 1 1 42685
0 42687 7 1 2 62783 92829
0 42688 5 1 1 42687
0 42689 7 1 2 92835 42688
0 42690 5 1 1 42689
0 42691 7 1 2 76694 66789
0 42692 5 1 1 42691
0 42693 7 1 2 66802 75579
0 42694 5 1 1 42693
0 42695 7 1 2 71449 66881
0 42696 7 1 2 42694 42695
0 42697 5 1 1 42696
0 42698 7 1 2 42692 42697
0 42699 5 1 1 42698
0 42700 7 1 2 61415 42699
0 42701 7 1 2 42690 42700
0 42702 5 1 1 42701
0 42703 7 1 2 66616 42702
0 42704 7 1 2 42686 42703
0 42705 5 1 1 42704
0 42706 7 1 2 94766 42705
0 42707 7 1 2 42567 42706
0 42708 5 1 1 42707
0 42709 7 1 2 42334 42708
0 42710 5 1 1 42709
0 42711 7 1 2 66323 42710
0 42712 5 1 1 42711
0 42713 7 1 2 61416 5079
0 42714 5 2 1 42713
0 42715 7 1 2 58788 87431
0 42716 7 1 2 89018 42715
0 42717 7 1 2 86757 42716
0 42718 7 1 2 94739 42717
0 42719 5 1 1 42718
0 42720 7 2 2 64731 94687
0 42721 5 1 1 94781
0 42722 7 1 2 94704 42721
0 42723 5 2 1 42722
0 42724 7 1 2 84301 94730
0 42725 7 1 2 94783 42724
0 42726 5 1 1 42725
0 42727 7 1 2 42719 42726
0 42728 5 1 1 42727
0 42729 7 1 2 94779 42728
0 42730 5 1 1 42729
0 42731 7 1 2 42712 42730
0 42732 7 1 2 42292 42731
0 42733 5 1 1 42732
0 42734 7 1 2 60154 42733
0 42735 5 1 1 42734
0 42736 7 1 2 60647 38757
0 42737 5 1 1 42736
0 42738 7 1 2 94118 42737
0 42739 5 1 1 42738
0 42740 7 1 2 61055 42739
0 42741 5 1 1 42740
0 42742 7 1 2 94106 42741
0 42743 5 1 1 42742
0 42744 7 1 2 61417 42743
0 42745 5 1 1 42744
0 42746 7 1 2 94095 42745
0 42747 5 1 1 42746
0 42748 7 1 2 63386 42747
0 42749 5 1 1 42748
0 42750 7 1 2 68259 91182
0 42751 5 1 1 42750
0 42752 7 1 2 68153 82929
0 42753 5 1 1 42752
0 42754 7 1 2 42751 42753
0 42755 5 1 1 42754
0 42756 7 1 2 86088 75276
0 42757 7 1 2 42755 42756
0 42758 5 1 1 42757
0 42759 7 1 2 42749 42758
0 42760 5 1 1 42759
0 42761 7 1 2 66324 42760
0 42762 5 1 1 42761
0 42763 7 1 2 78452 93283
0 42764 5 1 1 42763
0 42765 7 1 2 76268 81610
0 42766 5 1 1 42765
0 42767 7 1 2 70257 42766
0 42768 5 1 1 42767
0 42769 7 1 2 62784 42768
0 42770 5 1 1 42769
0 42771 7 1 2 63084 92815
0 42772 5 1 1 42771
0 42773 7 1 2 42770 42772
0 42774 5 1 1 42773
0 42775 7 1 2 68260 42774
0 42776 5 1 1 42775
0 42777 7 1 2 62785 92816
0 42778 5 1 1 42777
0 42779 7 1 2 73133 76380
0 42780 5 1 1 42779
0 42781 7 1 2 42778 42780
0 42782 5 1 1 42781
0 42783 7 1 2 63085 42782
0 42784 5 1 1 42783
0 42785 7 1 2 42776 42784
0 42786 5 1 1 42785
0 42787 7 1 2 62255 42786
0 42788 5 1 1 42787
0 42789 7 1 2 42764 42788
0 42790 5 1 1 42789
0 42791 7 1 2 66325 42790
0 42792 5 1 1 42791
0 42793 7 1 2 86924 93524
0 42794 5 1 1 42793
0 42795 7 1 2 81261 42794
0 42796 5 2 1 42795
0 42797 7 1 2 83976 86495
0 42798 5 1 1 42797
0 42799 7 1 2 94785 42798
0 42800 7 1 2 42792 42799
0 42801 5 1 1 42800
0 42802 7 1 2 64394 42801
0 42803 5 1 1 42802
0 42804 7 1 2 78255 67877
0 42805 5 1 1 42804
0 42806 7 1 2 61056 42805
0 42807 5 1 1 42806
0 42808 7 1 2 28131 42807
0 42809 5 1 1 42808
0 42810 7 1 2 73672 42809
0 42811 5 1 1 42810
0 42812 7 1 2 16332 42811
0 42813 5 1 1 42812
0 42814 7 1 2 91472 42813
0 42815 5 1 1 42814
0 42816 7 1 2 84804 92654
0 42817 5 1 1 42816
0 42818 7 1 2 86496 84744
0 42819 7 1 2 77679 42818
0 42820 5 1 1 42819
0 42821 7 1 2 42817 42820
0 42822 5 1 1 42821
0 42823 7 1 2 60648 42822
0 42824 5 1 1 42823
0 42825 7 1 2 83467 84130
0 42826 5 1 1 42825
0 42827 7 1 2 42824 42826
0 42828 5 1 1 42827
0 42829 7 1 2 70220 42828
0 42830 5 1 1 42829
0 42831 7 1 2 81342 94191
0 42832 7 1 2 77685 42831
0 42833 5 1 1 42832
0 42834 7 1 2 42830 42833
0 42835 7 1 2 42815 42834
0 42836 5 1 1 42835
0 42837 7 1 2 69058 42836
0 42838 5 1 1 42837
0 42839 7 1 2 75457 33115
0 42840 5 1 1 42839
0 42841 7 1 2 78596 42840
0 42842 5 1 1 42841
0 42843 7 1 2 68154 73673
0 42844 7 1 2 80529 42843
0 42845 5 1 1 42844
0 42846 7 1 2 42842 42845
0 42847 5 1 1 42846
0 42848 7 1 2 61684 42847
0 42849 5 1 1 42848
0 42850 7 2 2 62256 80518
0 42851 7 1 2 85573 94787
0 42852 5 1 1 42851
0 42853 7 1 2 78614 42852
0 42854 5 1 1 42853
0 42855 7 1 2 81560 42854
0 42856 5 1 1 42855
0 42857 7 1 2 42849 42856
0 42858 5 1 1 42857
0 42859 7 1 2 67781 42858
0 42860 5 1 1 42859
0 42861 7 1 2 62786 92811
0 42862 5 1 1 42861
0 42863 7 1 2 76269 83345
0 42864 5 1 1 42863
0 42865 7 1 2 70258 42864
0 42866 7 1 2 42862 42865
0 42867 5 1 1 42866
0 42868 7 1 2 87477 42867
0 42869 5 1 1 42868
0 42870 7 1 2 83958 81611
0 42871 5 1 1 42870
0 42872 7 1 2 73939 42871
0 42873 5 1 1 42872
0 42874 7 1 2 87478 42873
0 42875 5 1 1 42874
0 42876 7 1 2 58339 42875
0 42877 5 1 1 42876
0 42878 7 1 2 79679 90520
0 42879 5 1 1 42878
0 42880 7 1 2 86700 42879
0 42881 5 1 1 42880
0 42882 7 1 2 68261 42881
0 42883 7 1 2 42877 42882
0 42884 5 1 1 42883
0 42885 7 1 2 42869 42884
0 42886 7 1 2 42860 42885
0 42887 7 1 2 42838 42886
0 42888 7 1 2 42803 42887
0 42889 7 1 2 71696 81098
0 42890 5 1 1 42889
0 42891 7 1 2 73482 42890
0 42892 5 1 1 42891
0 42893 7 1 2 62257 42892
0 42894 5 1 1 42893
0 42895 7 1 2 93239 42894
0 42896 5 1 1 42895
0 42897 7 1 2 62511 42896
0 42898 5 1 1 42897
0 42899 7 1 2 94086 42898
0 42900 5 1 1 42899
0 42901 7 1 2 62787 42900
0 42902 5 1 1 42901
0 42903 7 1 2 83959 78752
0 42904 5 1 1 42903
0 42905 7 1 2 73940 42904
0 42906 7 1 2 94151 42905
0 42907 5 1 1 42906
0 42908 7 1 2 18090 42907
0 42909 5 1 1 42908
0 42910 7 2 2 66326 85667
0 42911 7 1 2 92827 94789
0 42912 7 1 2 42909 42911
0 42913 7 1 2 42902 42912
0 42914 5 1 1 42913
0 42915 7 2 2 61685 85972
0 42916 7 1 2 64395 85784
0 42917 5 1 1 42916
0 42918 7 2 2 68787 42917
0 42919 5 1 1 94793
0 42920 7 1 2 65683 94794
0 42921 5 1 1 42920
0 42922 7 1 2 94791 42921
0 42923 5 1 1 42922
0 42924 7 1 2 63387 42923
0 42925 7 1 2 42914 42924
0 42926 5 1 1 42925
0 42927 7 2 2 66327 94120
0 42928 5 1 1 94795
0 42929 7 2 2 68040 87372
0 42930 5 1 1 94797
0 42931 7 1 2 42928 42930
0 42932 5 1 1 42931
0 42933 7 1 2 61057 42932
0 42934 5 1 1 42933
0 42935 7 1 2 83885 88812
0 42936 5 1 1 42935
0 42937 7 1 2 67221 76381
0 42938 5 1 1 42937
0 42939 7 1 2 42936 42938
0 42940 5 1 1 42939
0 42941 7 1 2 62258 42940
0 42942 5 1 1 42941
0 42943 7 4 2 63916 93750
0 42944 5 3 1 94799
0 42945 7 1 2 42942 94803
0 42946 5 1 1 42945
0 42947 7 1 2 71322 42946
0 42948 5 1 1 42947
0 42949 7 1 2 68440 74231
0 42950 5 1 1 42949
0 42951 7 1 2 93768 42950
0 42952 5 1 1 42951
0 42953 7 1 2 71450 42952
0 42954 5 1 1 42953
0 42955 7 1 2 42948 42954
0 42956 5 1 1 42955
0 42957 7 1 2 66328 42956
0 42958 5 1 1 42957
0 42959 7 1 2 78836 84378
0 42960 5 1 1 42959
0 42961 7 1 2 78273 42960
0 42962 5 1 1 42961
0 42963 7 1 2 66329 42962
0 42964 5 1 1 42963
0 42965 7 1 2 84314 89459
0 42966 5 2 1 42965
0 42967 7 1 2 42964 94806
0 42968 5 1 1 42967
0 42969 7 1 2 69059 42968
0 42970 5 1 1 42969
0 42971 7 1 2 80519 86827
0 42972 7 1 2 84379 42971
0 42973 5 1 1 42972
0 42974 7 1 2 80520 81262
0 42975 5 2 1 42974
0 42976 7 1 2 68155 81561
0 42977 5 1 1 42976
0 42978 7 1 2 85091 91473
0 42979 5 1 1 42978
0 42980 7 1 2 42977 42979
0 42981 7 1 2 94808 42980
0 42982 7 1 2 42973 42981
0 42983 5 1 1 42982
0 42984 7 1 2 67782 42983
0 42985 5 1 1 42984
0 42986 7 1 2 94786 42985
0 42987 7 1 2 42970 42986
0 42988 7 1 2 42958 42987
0 42989 7 1 2 42934 42988
0 42990 5 1 1 42989
0 42991 7 1 2 61418 42990
0 42992 5 1 1 42991
0 42993 7 1 2 42926 42992
0 42994 7 1 2 42888 42993
0 42995 5 1 1 42994
0 42996 7 1 2 64613 42995
0 42997 5 1 1 42996
0 42998 7 1 2 42762 42997
0 42999 5 1 1 42998
0 43000 7 1 2 64732 42999
0 43001 5 1 1 43000
0 43002 7 2 2 72909 85847
0 43003 5 1 1 94810
0 43004 7 1 2 72910 73878
0 43005 5 1 1 43004
0 43006 7 2 2 43003 43005
0 43007 5 1 1 94812
0 43008 7 1 2 60649 94813
0 43009 5 1 1 43008
0 43010 7 1 2 77911 77109
0 43011 5 1 1 43010
0 43012 7 1 2 43009 43011
0 43013 5 1 1 43012
0 43014 7 1 2 63086 43013
0 43015 5 1 1 43014
0 43016 7 2 2 80628 72928
0 43017 5 1 1 94814
0 43018 7 1 2 84193 94815
0 43019 5 1 1 43018
0 43020 7 1 2 43015 43019
0 43021 5 1 1 43020
0 43022 7 1 2 67783 43021
0 43023 5 1 1 43022
0 43024 7 1 2 85646 93342
0 43025 5 1 1 43024
0 43026 7 1 2 85671 93284
0 43027 5 1 1 43026
0 43028 7 1 2 43025 43027
0 43029 7 1 2 43023 43028
0 43030 5 2 1 43029
0 43031 7 1 2 93974 94816
0 43032 5 1 1 43031
0 43033 7 1 2 61686 70221
0 43034 7 2 2 12922 43033
0 43035 7 1 2 84011 94818
0 43036 5 1 1 43035
0 43037 7 1 2 71215 11413
0 43038 5 1 1 43037
0 43039 7 2 2 81099 43038
0 43040 7 1 2 87624 94820
0 43041 5 1 1 43040
0 43042 7 1 2 72783 15319
0 43043 7 1 2 82432 43042
0 43044 7 1 2 78022 43043
0 43045 5 1 1 43044
0 43046 7 1 2 43041 43045
0 43047 5 1 1 43046
0 43048 7 1 2 62512 43047
0 43049 5 1 1 43048
0 43050 7 1 2 43036 43049
0 43051 5 1 1 43050
0 43052 7 1 2 62788 43051
0 43053 5 1 1 43052
0 43054 7 1 2 71323 93670
0 43055 5 1 1 43054
0 43056 7 1 2 64396 81280
0 43057 5 1 1 43056
0 43058 7 1 2 43055 43057
0 43059 5 2 1 43058
0 43060 7 1 2 87625 94822
0 43061 5 1 1 43060
0 43062 7 1 2 43053 43061
0 43063 5 1 1 43062
0 43064 7 1 2 61419 43063
0 43065 5 1 1 43064
0 43066 7 1 2 68156 70115
0 43067 5 1 1 43066
0 43068 7 1 2 79675 43067
0 43069 5 1 1 43068
0 43070 7 1 2 64397 43069
0 43071 5 1 1 43070
0 43072 7 1 2 94804 43071
0 43073 5 1 1 43072
0 43074 7 1 2 63087 43073
0 43075 5 1 1 43074
0 43076 7 1 2 70951 75059
0 43077 5 1 1 43076
0 43078 7 1 2 43075 43077
0 43079 5 1 1 43078
0 43080 7 1 2 61058 43079
0 43081 5 1 1 43080
0 43082 7 1 2 85361 78572
0 43083 5 1 1 43082
0 43084 7 1 2 43081 43083
0 43085 5 2 1 43084
0 43086 7 1 2 87626 94824
0 43087 5 1 1 43086
0 43088 7 1 2 43065 43087
0 43089 5 1 1 43088
0 43090 7 1 2 63388 43089
0 43091 5 1 1 43090
0 43092 7 1 2 78246 79853
0 43093 7 1 2 80662 43092
0 43094 7 1 2 84798 92249
0 43095 7 1 2 43093 43094
0 43096 5 1 1 43095
0 43097 7 1 2 43091 43096
0 43098 5 1 1 43097
0 43099 7 1 2 78876 43098
0 43100 5 1 1 43099
0 43101 7 1 2 43032 43100
0 43102 7 1 2 43001 43101
0 43103 5 1 1 43102
0 43104 7 1 2 63523 43103
0 43105 5 1 1 43104
0 43106 7 4 2 63389 88264
0 43107 5 1 1 94826
0 43108 7 1 2 94817 94827
0 43109 5 1 1 43108
0 43110 7 1 2 88265 94821
0 43111 5 1 1 43110
0 43112 7 2 2 78247 81658
0 43113 7 1 2 81368 94830
0 43114 5 1 1 43113
0 43115 7 1 2 43111 43114
0 43116 5 1 1 43115
0 43117 7 1 2 63390 43116
0 43118 5 1 1 43117
0 43119 7 1 2 77592 88266
0 43120 7 1 2 86426 43119
0 43121 5 1 1 43120
0 43122 7 1 2 43118 43121
0 43123 5 1 1 43122
0 43124 7 1 2 62513 43123
0 43125 5 1 1 43124
0 43126 7 1 2 82808 94819
0 43127 5 1 1 43126
0 43128 7 1 2 43125 43127
0 43129 5 1 1 43128
0 43130 7 1 2 62789 43129
0 43131 5 1 1 43130
0 43132 7 1 2 94823 94828
0 43133 5 1 1 43132
0 43134 7 1 2 43131 43133
0 43135 5 1 1 43134
0 43136 7 1 2 61420 43135
0 43137 5 1 1 43136
0 43138 7 1 2 94825 94829
0 43139 5 1 1 43138
0 43140 7 1 2 43137 43139
0 43141 5 1 1 43140
0 43142 7 1 2 78877 43141
0 43143 5 1 1 43142
0 43144 7 1 2 43109 43143
0 43145 5 1 1 43144
0 43146 7 1 2 86671 43145
0 43147 5 1 1 43146
0 43148 7 1 2 43105 43147
0 43149 5 1 1 43148
0 43150 7 1 2 66718 43149
0 43151 5 1 1 43150
0 43152 7 2 2 67784 80359
0 43153 7 1 2 85945 94832
0 43154 5 1 1 43153
0 43155 7 1 2 63391 68632
0 43156 7 1 2 93829 43155
0 43157 5 1 1 43156
0 43158 7 1 2 43154 43157
0 43159 5 1 1 43158
0 43160 7 1 2 64614 43159
0 43161 5 1 1 43160
0 43162 7 1 2 66033 80160
0 43163 7 1 2 94332 43162
0 43164 5 1 1 43163
0 43165 7 1 2 43161 43164
0 43166 5 1 1 43165
0 43167 7 1 2 64733 43166
0 43168 5 1 1 43167
0 43169 7 2 2 84613 94833
0 43170 7 1 2 80682 94834
0 43171 5 1 1 43170
0 43172 7 1 2 43168 43171
0 43173 5 1 1 43172
0 43174 7 1 2 63524 43173
0 43175 5 1 1 43174
0 43176 7 1 2 86672 80763
0 43177 7 1 2 94835 43176
0 43178 5 1 1 43177
0 43179 7 1 2 43175 43178
0 43180 5 1 1 43179
0 43181 7 1 2 88923 43180
0 43182 5 1 1 43181
0 43183 7 2 2 59002 72669
0 43184 7 2 2 90260 94836
0 43185 7 1 2 74890 86323
0 43186 7 1 2 94838 43185
0 43187 5 1 1 43186
0 43188 7 1 2 43182 43187
0 43189 5 1 1 43188
0 43190 7 1 2 65684 43189
0 43191 5 1 1 43190
0 43192 7 1 2 73387 72201
0 43193 5 1 1 43192
0 43194 7 1 2 84917 87275
0 43195 5 1 1 43194
0 43196 7 1 2 43193 43195
0 43197 5 1 1 43196
0 43198 7 1 2 73674 43197
0 43199 5 1 1 43198
0 43200 7 1 2 83076 82611
0 43201 5 1 1 43200
0 43202 7 1 2 43199 43201
0 43203 5 1 1 43202
0 43204 7 1 2 58631 43203
0 43205 5 1 1 43204
0 43206 7 1 2 87467 83049
0 43207 7 1 2 92698 43206
0 43208 5 1 1 43207
0 43209 7 1 2 43205 43208
0 43210 5 1 1 43209
0 43211 7 1 2 86925 43210
0 43212 5 1 1 43211
0 43213 7 3 2 58632 82413
0 43214 7 1 2 85830 75716
0 43215 7 1 2 94840 43214
0 43216 5 1 1 43215
0 43217 7 1 2 43212 43216
0 43218 5 1 1 43217
0 43219 7 1 2 74250 43218
0 43220 5 1 1 43219
0 43221 7 2 2 73321 88924
0 43222 7 2 2 91654 94843
0 43223 5 1 1 94845
0 43224 7 2 2 62514 70883
0 43225 5 9 1 94847
0 43226 7 1 2 66790 91288
0 43227 5 1 1 43226
0 43228 7 2 2 73322 74251
0 43229 7 1 2 66330 94858
0 43230 7 1 2 85280 43229
0 43231 5 1 1 43230
0 43232 7 1 2 43227 43231
0 43233 5 1 1 43232
0 43234 7 1 2 59643 43233
0 43235 5 1 1 43234
0 43236 7 2 2 74468 91594
0 43237 7 1 2 69777 87913
0 43238 7 1 2 94860 43237
0 43239 5 1 1 43238
0 43240 7 1 2 43235 43239
0 43241 5 1 1 43240
0 43242 7 1 2 94849 43241
0 43243 5 1 1 43242
0 43244 7 1 2 43223 43243
0 43245 7 1 2 43220 43244
0 43246 5 1 1 43245
0 43247 7 1 2 59159 43246
0 43248 5 1 1 43247
0 43249 7 1 2 43191 43248
0 43250 5 1 1 43249
0 43251 7 1 2 65307 43250
0 43252 5 1 1 43251
0 43253 7 1 2 61687 73696
0 43254 5 1 1 43253
0 43255 7 2 2 65685 43254
0 43256 7 1 2 84918 94862
0 43257 5 1 1 43256
0 43258 7 2 2 66331 84249
0 43259 5 1 1 94864
0 43260 7 1 2 72911 94865
0 43261 5 1 1 43260
0 43262 7 1 2 43257 43261
0 43263 5 1 1 43262
0 43264 7 3 2 86317 74763
0 43265 7 3 2 74416 94866
0 43266 7 1 2 62113 94869
0 43267 7 1 2 43263 43266
0 43268 5 1 1 43267
0 43269 7 1 2 73917 94181
0 43270 5 1 1 43269
0 43271 7 2 2 32946 43270
0 43272 5 1 1 94872
0 43273 7 1 2 67785 43272
0 43274 5 1 1 43273
0 43275 7 1 2 62790 84436
0 43276 5 1 1 43275
0 43277 7 1 2 72950 43276
0 43278 5 1 1 43277
0 43279 7 1 2 68262 43278
0 43280 5 1 1 43279
0 43281 7 1 2 43280 43007
0 43282 5 1 1 43281
0 43283 7 1 2 63088 43282
0 43284 5 1 1 43283
0 43285 7 1 2 73697 39065
0 43286 5 1 1 43285
0 43287 7 1 2 85883 93843
0 43288 5 1 1 43287
0 43289 7 1 2 43286 43288
0 43290 7 1 2 43284 43289
0 43291 5 1 1 43290
0 43292 7 1 2 60650 43291
0 43293 5 1 1 43292
0 43294 7 1 2 43274 43293
0 43295 5 1 1 43294
0 43296 7 1 2 63525 43295
0 43297 5 1 1 43296
0 43298 7 2 2 68263 90059
0 43299 5 1 1 94874
0 43300 7 1 2 86441 94875
0 43301 5 1 1 43300
0 43302 7 1 2 58789 43301
0 43303 5 1 1 43302
0 43304 7 1 2 60651 80819
0 43305 7 1 2 43303 43304
0 43306 5 1 1 43305
0 43307 7 1 2 43297 43306
0 43308 5 1 1 43307
0 43309 7 1 2 78878 43308
0 43310 5 1 1 43309
0 43311 7 1 2 67820 32825
0 43312 5 1 1 43311
0 43313 7 1 2 77686 90932
0 43314 5 1 1 43313
0 43315 7 1 2 70222 91928
0 43316 5 1 1 43315
0 43317 7 1 2 43314 43316
0 43318 7 1 2 43312 43317
0 43319 5 1 1 43318
0 43320 7 1 2 85171 43319
0 43321 5 1 1 43320
0 43322 7 1 2 63392 78597
0 43323 5 1 1 43322
0 43324 7 1 2 78492 81306
0 43325 5 1 1 43324
0 43326 7 1 2 43323 43325
0 43327 5 1 1 43326
0 43328 7 1 2 67786 43327
0 43329 5 1 1 43328
0 43330 7 1 2 58633 43299
0 43331 5 1 1 43330
0 43332 7 1 2 70223 43331
0 43333 5 1 1 43332
0 43334 7 1 2 85989 77653
0 43335 5 1 1 43334
0 43336 7 1 2 87039 43335
0 43337 5 1 1 43336
0 43338 7 1 2 85079 43337
0 43339 7 1 2 43333 43338
0 43340 7 1 2 43329 43339
0 43341 5 1 1 43340
0 43342 7 1 2 71324 43341
0 43343 5 1 1 43342
0 43344 7 2 2 43321 43343
0 43345 5 1 1 94876
0 43346 7 1 2 63526 43345
0 43347 5 1 1 43346
0 43348 7 1 2 43310 43347
0 43349 5 1 1 43348
0 43350 7 4 2 64734 66719
0 43351 7 1 2 61688 94878
0 43352 7 1 2 43349 43351
0 43353 5 1 1 43352
0 43354 7 1 2 43268 43353
0 43355 5 1 1 43354
0 43356 7 1 2 59905 43355
0 43357 5 1 1 43356
0 43358 7 1 2 82695 94688
0 43359 5 1 1 43358
0 43360 7 1 2 69987 87914
0 43361 7 1 2 94861 43360
0 43362 5 1 1 43361
0 43363 7 1 2 43359 43362
0 43364 5 1 1 43363
0 43365 7 1 2 57769 43364
0 43366 5 1 1 43365
0 43367 7 1 2 85281 87432
0 43368 5 1 1 43367
0 43369 7 1 2 94660 43368
0 43370 5 2 1 43369
0 43371 7 1 2 94859 94882
0 43372 5 1 1 43371
0 43373 7 1 2 74431 91289
0 43374 5 1 1 43373
0 43375 7 1 2 43372 43374
0 43376 5 1 1 43375
0 43377 7 1 2 73228 43376
0 43378 5 1 1 43377
0 43379 7 1 2 43366 43378
0 43380 5 1 1 43379
0 43381 7 1 2 65308 43380
0 43382 5 1 1 43381
0 43383 7 1 2 57770 94846
0 43384 5 1 1 43383
0 43385 7 1 2 43382 43384
0 43386 5 1 1 43385
0 43387 7 1 2 76460 43386
0 43388 5 1 1 43387
0 43389 7 3 2 60042 83023
0 43390 7 1 2 73842 94884
0 43391 7 1 2 94689 43390
0 43392 5 1 1 43391
0 43393 7 1 2 72033 91595
0 43394 7 1 2 91655 43393
0 43395 5 1 1 43394
0 43396 7 1 2 43392 43395
0 43397 5 1 1 43396
0 43398 7 1 2 59160 43397
0 43399 5 1 1 43398
0 43400 7 1 2 43388 43399
0 43401 7 1 2 43357 43400
0 43402 7 1 2 43252 43401
0 43403 7 1 2 43151 43402
0 43404 5 1 1 43403
0 43405 7 1 2 61965 43404
0 43406 5 1 1 43405
0 43407 7 1 2 58074 94091
0 43408 7 1 2 79079 43407
0 43409 5 1 1 43408
0 43410 7 1 2 62515 43409
0 43411 5 1 1 43410
0 43412 7 1 2 74875 75190
0 43413 5 1 1 43412
0 43414 7 1 2 70837 80704
0 43415 5 1 1 43414
0 43416 7 1 2 43413 43415
0 43417 7 2 2 43411 43416
0 43418 7 1 2 71522 94887
0 43419 5 1 1 43418
0 43420 7 1 2 85217 43419
0 43421 5 1 1 43420
0 43422 7 1 2 76382 81021
0 43423 7 1 2 94746 43422
0 43424 7 1 2 94088 43423
0 43425 5 1 1 43424
0 43426 7 1 2 43421 43425
0 43427 5 1 1 43426
0 43428 7 1 2 70224 43427
0 43429 5 1 1 43428
0 43430 7 1 2 62259 93651
0 43431 5 1 1 43430
0 43432 7 1 2 83337 81801
0 43433 5 1 1 43432
0 43434 7 1 2 43431 43433
0 43435 5 1 1 43434
0 43436 7 1 2 62516 43435
0 43437 5 1 1 43436
0 43438 7 1 2 62791 92825
0 43439 5 1 1 43438
0 43440 7 1 2 43437 43439
0 43441 5 2 1 43440
0 43442 7 1 2 94743 94889
0 43443 5 1 1 43442
0 43444 7 1 2 76695 91590
0 43445 7 1 2 81773 43444
0 43446 5 1 1 43445
0 43447 7 1 2 69822 80184
0 43448 7 1 2 72838 43447
0 43449 5 1 1 43448
0 43450 7 1 2 75554 43449
0 43451 5 1 1 43450
0 43452 7 1 2 43446 43451
0 43453 7 1 2 43443 43452
0 43454 7 1 2 43429 43453
0 43455 5 1 1 43454
0 43456 7 1 2 61421 43455
0 43457 5 1 1 43456
0 43458 7 1 2 12088 21625
0 43459 5 1 1 43458
0 43460 7 1 2 62260 43459
0 43461 5 1 1 43460
0 43462 7 1 2 59003 70049
0 43463 5 1 1 43462
0 43464 7 1 2 93530 43463
0 43465 5 1 1 43464
0 43466 7 1 2 81603 43465
0 43467 7 1 2 43461 43466
0 43468 5 1 1 43467
0 43469 7 1 2 61059 43468
0 43470 5 1 1 43469
0 43471 7 1 2 71216 34306
0 43472 7 1 2 94763 43471
0 43473 5 1 1 43472
0 43474 7 1 2 68157 43473
0 43475 5 1 1 43474
0 43476 7 1 2 71523 72482
0 43477 5 1 1 43476
0 43478 7 1 2 85699 43477
0 43479 5 1 1 43478
0 43480 7 1 2 43475 43479
0 43481 7 1 2 43470 43480
0 43482 5 1 1 43481
0 43483 7 1 2 63393 43482
0 43484 5 1 1 43483
0 43485 7 1 2 84194 77407
0 43486 5 1 1 43485
0 43487 7 1 2 85499 43486
0 43488 5 1 1 43487
0 43489 7 1 2 67787 43488
0 43490 5 1 1 43489
0 43491 7 1 2 80277 90384
0 43492 5 1 1 43491
0 43493 7 1 2 43490 43492
0 43494 5 1 1 43493
0 43495 7 1 2 68158 43494
0 43496 5 1 1 43495
0 43497 7 1 2 83305 91183
0 43498 5 1 1 43497
0 43499 7 1 2 43496 43498
0 43500 7 1 2 43484 43499
0 43501 5 1 1 43500
0 43502 7 1 2 64615 43501
0 43503 5 1 1 43502
0 43504 7 1 2 67380 34137
0 43505 5 1 1 43504
0 43506 7 1 2 78573 43505
0 43507 5 1 1 43506
0 43508 7 1 2 94774 43507
0 43509 5 1 1 43508
0 43510 7 1 2 76696 43509
0 43511 5 1 1 43510
0 43512 7 1 2 43503 43511
0 43513 7 1 2 43457 43512
0 43514 5 1 1 43513
0 43515 7 1 2 58790 43514
0 43516 5 1 1 43515
0 43517 7 1 2 76927 90096
0 43518 5 1 1 43517
0 43519 7 1 2 58634 74148
0 43520 5 1 1 43519
0 43521 7 2 2 69829 93208
0 43522 5 1 1 94891
0 43523 7 1 2 67679 94892
0 43524 5 1 1 43523
0 43525 7 1 2 43520 43524
0 43526 5 1 1 43525
0 43527 7 1 2 61422 79028
0 43528 7 1 2 43526 43527
0 43529 5 1 1 43528
0 43530 7 1 2 43518 43529
0 43531 7 1 2 43516 43530
0 43532 5 1 1 43531
0 43533 7 1 2 66332 43532
0 43534 5 1 1 43533
0 43535 7 1 2 63394 73334
0 43536 5 1 1 43535
0 43537 7 1 2 94615 43536
0 43538 5 1 1 43537
0 43539 7 1 2 71325 43538
0 43540 5 1 1 43539
0 43541 7 2 2 62517 75265
0 43542 5 1 1 94893
0 43543 7 1 2 90060 94894
0 43544 5 1 1 43543
0 43545 7 1 2 85134 43544
0 43546 5 1 1 43545
0 43547 7 1 2 69060 43546
0 43548 5 1 1 43547
0 43549 7 1 2 91340 93659
0 43550 7 1 2 43548 43549
0 43551 5 1 1 43550
0 43552 7 1 2 75912 43551
0 43553 5 1 1 43552
0 43554 7 1 2 62261 94164
0 43555 5 1 1 43554
0 43556 7 1 2 91341 43555
0 43557 5 1 1 43556
0 43558 7 1 2 70838 43557
0 43559 5 1 1 43558
0 43560 7 1 2 64100 94139
0 43561 5 1 1 43560
0 43562 7 1 2 42264 43561
0 43563 7 1 2 43559 43562
0 43564 5 1 1 43563
0 43565 7 1 2 69061 43564
0 43566 5 1 1 43565
0 43567 7 1 2 93660 94165
0 43568 5 1 1 43567
0 43569 7 1 2 78299 43568
0 43570 5 1 1 43569
0 43571 7 1 2 42232 43570
0 43572 5 1 1 43571
0 43573 7 1 2 70839 43572
0 43574 5 1 1 43573
0 43575 7 1 2 61423 80204
0 43576 5 1 1 43575
0 43577 7 1 2 93661 43576
0 43578 5 1 1 43577
0 43579 7 1 2 78200 43578
0 43580 5 1 1 43579
0 43581 7 1 2 62792 67103
0 43582 5 1 1 43581
0 43583 7 1 2 66034 43582
0 43584 5 1 1 43583
0 43585 7 1 2 85172 43584
0 43586 5 1 1 43585
0 43587 7 1 2 43580 43586
0 43588 7 1 2 43574 43587
0 43589 7 1 2 43566 43588
0 43590 7 1 2 43553 43589
0 43591 5 1 1 43590
0 43592 7 1 2 61060 43591
0 43593 5 1 1 43592
0 43594 7 1 2 80205 77483
0 43595 5 1 1 43594
0 43596 7 1 2 85135 43595
0 43597 5 1 1 43596
0 43598 7 1 2 69062 43597
0 43599 5 1 1 43598
0 43600 7 1 2 60652 84423
0 43601 5 2 1 43600
0 43602 7 1 2 68041 87384
0 43603 5 1 1 43602
0 43604 7 1 2 85173 43603
0 43605 5 1 1 43604
0 43606 7 1 2 94895 43605
0 43607 7 1 2 43599 43606
0 43608 5 1 1 43607
0 43609 7 1 2 61424 43608
0 43610 5 1 1 43609
0 43611 7 1 2 43593 43610
0 43612 7 1 2 43540 43611
0 43613 5 1 1 43612
0 43614 7 1 2 94043 43613
0 43615 5 1 1 43614
0 43616 7 2 2 78912 81263
0 43617 5 1 1 94897
0 43618 7 1 2 83077 94898
0 43619 5 1 1 43618
0 43620 7 2 2 70840 92410
0 43621 5 1 1 94899
0 43622 7 1 2 59906 82508
0 43623 7 1 2 43621 43622
0 43624 5 1 1 43623
0 43625 7 1 2 43619 43624
0 43626 5 1 1 43625
0 43627 7 1 2 63527 43626
0 43628 5 1 1 43627
0 43629 7 1 2 72729 76697
0 43630 5 1 1 43629
0 43631 7 1 2 76494 94800
0 43632 5 2 1 43631
0 43633 7 1 2 43630 94901
0 43634 5 1 1 43633
0 43635 7 1 2 88267 43634
0 43636 5 1 1 43635
0 43637 7 2 2 59907 87238
0 43638 7 1 2 84875 94903
0 43639 5 2 1 43638
0 43640 7 1 2 71833 88268
0 43641 5 1 1 43640
0 43642 7 1 2 94905 43641
0 43643 5 1 1 43642
0 43644 7 1 2 62518 43643
0 43645 5 1 1 43644
0 43646 7 1 2 61689 93987
0 43647 5 1 1 43646
0 43648 7 1 2 94906 43647
0 43649 5 1 1 43648
0 43650 7 1 2 63917 43649
0 43651 5 1 1 43650
0 43652 7 1 2 43645 43651
0 43653 5 1 1 43652
0 43654 7 1 2 64101 43653
0 43655 5 1 1 43654
0 43656 7 2 2 76698 88269
0 43657 5 1 1 94907
0 43658 7 1 2 85252 82078
0 43659 5 1 1 43658
0 43660 7 1 2 77242 90883
0 43661 5 1 1 43660
0 43662 7 1 2 43659 43661
0 43663 5 1 1 43662
0 43664 7 1 2 68527 43663
0 43665 5 1 1 43664
0 43666 7 1 2 43657 43665
0 43667 7 1 2 43655 43666
0 43668 5 1 1 43667
0 43669 7 1 2 64398 43668
0 43670 5 1 1 43669
0 43671 7 1 2 43636 43670
0 43672 5 1 1 43671
0 43673 7 1 2 63089 43672
0 43674 5 1 1 43673
0 43675 7 2 2 88270 94747
0 43676 7 1 2 78352 94909
0 43677 5 1 1 43676
0 43678 7 2 2 84266 82612
0 43679 7 1 2 92607 94911
0 43680 5 1 1 43679
0 43681 7 1 2 43677 43680
0 43682 5 1 1 43681
0 43683 7 1 2 68159 43682
0 43684 5 1 1 43683
0 43685 7 1 2 67222 94748
0 43686 5 1 1 43685
0 43687 7 1 2 85215 43686
0 43688 5 2 1 43687
0 43689 7 1 2 88271 94913
0 43690 5 1 1 43689
0 43691 7 1 2 43684 43690
0 43692 5 1 1 43691
0 43693 7 1 2 70841 43692
0 43694 5 1 1 43693
0 43695 7 1 2 78229 94910
0 43696 5 1 1 43695
0 43697 7 1 2 86659 94912
0 43698 5 1 1 43697
0 43699 7 1 2 43696 43698
0 43700 5 1 1 43699
0 43701 7 1 2 75913 43700
0 43702 5 1 1 43701
0 43703 7 1 2 76657 93683
0 43704 5 1 1 43703
0 43705 7 1 2 2337 28897
0 43706 5 1 1 43705
0 43707 7 1 2 43704 43706
0 43708 5 1 1 43707
0 43709 7 1 2 84931 76699
0 43710 7 1 2 84286 43709
0 43711 5 1 1 43710
0 43712 7 1 2 75580 43711
0 43713 7 1 2 43708 43712
0 43714 5 1 1 43713
0 43715 7 1 2 88272 43714
0 43716 5 1 1 43715
0 43717 7 1 2 71326 94908
0 43718 5 1 1 43717
0 43719 7 1 2 68264 69848
0 43720 7 1 2 89864 43719
0 43721 7 1 2 91462 43720
0 43722 5 1 1 43721
0 43723 7 1 2 43718 43722
0 43724 5 1 1 43723
0 43725 7 1 2 68160 43724
0 43726 5 1 1 43725
0 43727 7 1 2 68878 80820
0 43728 7 1 2 79508 43727
0 43729 7 1 2 94904 43728
0 43730 5 1 1 43729
0 43731 7 1 2 43726 43730
0 43732 7 1 2 43716 43731
0 43733 7 1 2 43702 43732
0 43734 7 1 2 43694 43733
0 43735 7 1 2 43674 43734
0 43736 5 1 1 43735
0 43737 7 1 2 65686 43736
0 43738 5 1 1 43737
0 43739 7 1 2 43628 43738
0 43740 5 1 1 43739
0 43741 7 1 2 66035 43740
0 43742 5 1 1 43741
0 43743 7 1 2 43615 43742
0 43744 7 1 2 43534 43743
0 43745 5 1 1 43744
0 43746 7 1 2 60043 43745
0 43747 5 1 1 43746
0 43748 7 3 2 61690 85294
0 43749 7 2 2 83194 88021
0 43750 7 1 2 86760 94918
0 43751 5 1 1 43750
0 43752 7 1 2 64616 83177
0 43753 5 1 1 43752
0 43754 7 1 2 73455 94749
0 43755 5 1 1 43754
0 43756 7 1 2 43753 43755
0 43757 5 1 1 43756
0 43758 7 1 2 43751 43757
0 43759 5 1 1 43758
0 43760 7 1 2 94915 43759
0 43761 5 1 1 43760
0 43762 7 1 2 91921 94759
0 43763 5 1 1 43762
0 43764 7 1 2 65309 43763
0 43765 5 1 1 43764
0 43766 7 2 2 93163 43765
0 43767 7 1 2 2544 94920
0 43768 5 1 1 43767
0 43769 7 1 2 65687 43768
0 43770 5 1 1 43769
0 43771 7 1 2 68633 72494
0 43772 7 1 2 86411 43771
0 43773 5 1 1 43772
0 43774 7 1 2 64399 77718
0 43775 7 1 2 43773 43774
0 43776 7 1 2 43770 43775
0 43777 5 1 1 43776
0 43778 7 1 2 68161 75840
0 43779 5 1 1 43778
0 43780 7 1 2 93320 43779
0 43781 5 1 1 43780
0 43782 7 1 2 77110 43781
0 43783 5 1 1 43782
0 43784 7 1 2 68528 93316
0 43785 5 1 1 43784
0 43786 7 1 2 59644 43785
0 43787 7 1 2 43783 43786
0 43788 5 1 1 43787
0 43789 7 1 2 43777 43788
0 43790 5 1 1 43789
0 43791 7 1 2 65688 92049
0 43792 5 1 1 43791
0 43793 7 1 2 78536 43792
0 43794 5 1 1 43793
0 43795 7 1 2 93042 43794
0 43796 5 1 1 43795
0 43797 7 1 2 67788 93156
0 43798 5 1 1 43797
0 43799 7 1 2 74786 43798
0 43800 5 1 1 43799
0 43801 7 1 2 68162 43800
0 43802 5 1 1 43801
0 43803 7 1 2 58635 90337
0 43804 5 1 1 43803
0 43805 7 1 2 65310 43804
0 43806 5 1 1 43805
0 43807 7 1 2 43802 43806
0 43808 5 1 1 43807
0 43809 7 1 2 65689 43808
0 43810 5 1 1 43809
0 43811 7 1 2 43796 43810
0 43812 7 1 2 43790 43811
0 43813 5 1 1 43812
0 43814 7 1 2 59908 43813
0 43815 5 1 1 43814
0 43816 7 1 2 57481 86412
0 43817 5 1 1 43816
0 43818 7 1 2 72050 81802
0 43819 7 2 2 43817 43818
0 43820 5 1 1 94922
0 43821 7 1 2 57771 91152
0 43822 5 1 1 43821
0 43823 7 1 2 85174 43822
0 43824 7 1 2 94923 43823
0 43825 5 1 1 43824
0 43826 7 1 2 94757 43825
0 43827 5 1 1 43826
0 43828 7 1 2 43815 43827
0 43829 5 1 1 43828
0 43830 7 1 2 66333 43829
0 43831 5 1 1 43830
0 43832 7 1 2 43761 43831
0 43833 5 1 1 43832
0 43834 7 1 2 66036 43833
0 43835 5 1 1 43834
0 43836 7 2 2 81405 78951
0 43837 5 3 1 94924
0 43838 7 1 2 69823 94925
0 43839 5 1 1 43838
0 43840 7 1 2 82574 79726
0 43841 5 1 1 43840
0 43842 7 1 2 24741 43841
0 43843 5 1 1 43842
0 43844 7 1 2 76461 43843
0 43845 5 1 1 43844
0 43846 7 7 2 66334 78952
0 43847 5 2 1 94929
0 43848 7 2 2 70785 72002
0 43849 5 1 1 94938
0 43850 7 1 2 94930 94939
0 43851 5 1 1 43850
0 43852 7 1 2 91809 43851
0 43853 7 1 2 43845 43852
0 43854 5 1 1 43853
0 43855 7 1 2 59004 43854
0 43856 5 1 1 43855
0 43857 7 1 2 43839 43856
0 43858 5 1 1 43857
0 43859 7 1 2 57772 43858
0 43860 5 1 1 43859
0 43861 7 1 2 8383 82399
0 43862 5 1 1 43861
0 43863 7 1 2 59909 43862
0 43864 5 1 1 43863
0 43865 7 1 2 61691 81072
0 43866 5 1 1 43865
0 43867 7 1 2 12362 43866
0 43868 5 1 1 43867
0 43869 7 1 2 71217 43868
0 43870 5 1 1 43869
0 43871 7 1 2 43864 43870
0 43872 5 1 1 43871
0 43873 7 1 2 58636 43872
0 43874 5 1 1 43873
0 43875 7 1 2 87214 82596
0 43876 5 3 1 43875
0 43877 7 1 2 70786 94940
0 43878 5 1 1 43877
0 43879 7 1 2 93982 43878
0 43880 5 1 1 43879
0 43881 7 1 2 59645 43880
0 43882 5 1 1 43881
0 43883 7 1 2 43874 43882
0 43884 7 1 2 43860 43883
0 43885 5 1 1 43884
0 43886 7 1 2 85295 43885
0 43887 5 1 1 43886
0 43888 7 1 2 43835 43887
0 43889 5 1 1 43888
0 43890 7 1 2 66930 43889
0 43891 5 1 1 43890
0 43892 7 1 2 68042 93598
0 43893 5 1 1 43892
0 43894 7 1 2 60653 43893
0 43895 5 1 1 43894
0 43896 7 2 2 67896 43895
0 43897 5 1 1 94943
0 43898 7 2 2 78989 94944
0 43899 5 1 1 94945
0 43900 7 1 2 61425 93547
0 43901 5 1 1 43900
0 43902 7 1 2 65690 43901
0 43903 5 1 1 43902
0 43904 7 1 2 43899 43903
0 43905 5 1 1 43904
0 43906 7 1 2 58637 43905
0 43907 5 1 1 43906
0 43908 7 2 2 73456 77737
0 43909 5 1 1 94947
0 43910 7 1 2 75468 94948
0 43911 5 1 1 43910
0 43912 7 1 2 66335 43911
0 43913 7 1 2 43907 43912
0 43914 5 1 1 43913
0 43915 7 1 2 70100 90494
0 43916 7 1 2 78848 43915
0 43917 5 1 1 43916
0 43918 7 1 2 43914 43917
0 43919 5 1 1 43918
0 43920 7 1 2 59910 43919
0 43921 5 1 1 43920
0 43922 7 1 2 72410 89182
0 43923 7 1 2 94346 43922
0 43924 5 1 1 43923
0 43925 7 1 2 43921 43924
0 43926 5 1 1 43925
0 43927 7 1 2 63528 43926
0 43928 5 1 1 43927
0 43929 7 1 2 83941 32522
0 43930 7 1 2 94611 43929
0 43931 5 1 1 43930
0 43932 7 1 2 79556 91498
0 43933 7 1 2 43931 43932
0 43934 5 1 1 43933
0 43935 7 1 2 60044 43934
0 43936 7 1 2 43928 43935
0 43937 5 1 1 43936
0 43938 7 2 2 68788 77219
0 43939 7 1 2 87486 94045
0 43940 7 1 2 94949 43939
0 43941 7 1 2 85296 43940
0 43942 5 1 1 43941
0 43943 7 1 2 70842 74818
0 43944 5 1 1 43943
0 43945 7 1 2 83164 88273
0 43946 7 1 2 43944 43945
0 43947 5 1 1 43946
0 43948 7 1 2 64735 43947
0 43949 7 1 2 43942 43948
0 43950 5 1 1 43949
0 43951 7 1 2 59646 43950
0 43952 7 1 2 43937 43951
0 43953 5 1 1 43952
0 43954 7 1 2 78166 80450
0 43955 5 1 1 43954
0 43956 7 1 2 59647 94946
0 43957 5 1 1 43956
0 43958 7 1 2 61426 93408
0 43959 5 1 1 43958
0 43960 7 1 2 65691 43959
0 43961 5 1 1 43960
0 43962 7 1 2 61427 79778
0 43963 5 1 1 43962
0 43964 7 1 2 64400 94900
0 43965 5 1 1 43964
0 43966 7 1 2 43963 43965
0 43967 5 1 1 43966
0 43968 7 1 2 63395 43967
0 43969 5 1 1 43968
0 43970 7 1 2 43961 43969
0 43971 7 1 2 43957 43970
0 43972 5 1 1 43971
0 43973 7 1 2 43955 43972
0 43974 5 1 1 43973
0 43975 7 1 2 58791 43974
0 43976 5 1 1 43975
0 43977 7 1 2 65692 88499
0 43978 5 1 1 43977
0 43979 7 2 2 78009 43978
0 43980 7 1 2 94652 94951
0 43981 5 1 1 43980
0 43982 7 1 2 68634 72034
0 43983 7 1 2 94498 43982
0 43984 5 1 1 43983
0 43985 7 1 2 43981 43984
0 43986 5 1 1 43985
0 43987 7 1 2 61428 70787
0 43988 7 1 2 43986 43987
0 43989 5 1 1 43988
0 43990 7 1 2 43976 43989
0 43991 5 1 1 43990
0 43992 7 1 2 87647 43991
0 43993 5 1 1 43992
0 43994 7 1 2 74469 94237
0 43995 5 1 1 43994
0 43996 7 1 2 74519 81509
0 43997 7 1 2 93984 43996
0 43998 5 1 1 43997
0 43999 7 1 2 43995 43998
0 44000 5 1 1 43999
0 44001 7 1 2 59005 44000
0 44002 5 1 1 44001
0 44003 7 1 2 65080 87639
0 44004 5 1 1 44003
0 44005 7 1 2 87633 44004
0 44006 5 3 1 44005
0 44007 7 1 2 74543 94953
0 44008 5 1 1 44007
0 44009 7 1 2 44002 44008
0 44010 5 1 1 44009
0 44011 7 1 2 61429 44010
0 44012 5 1 1 44011
0 44013 7 1 2 59006 82214
0 44014 5 1 1 44013
0 44015 7 1 2 82597 44014
0 44016 5 3 1 44015
0 44017 7 1 2 60408 20700
0 44018 5 1 1 44017
0 44019 7 1 2 64736 73675
0 44020 7 1 2 73432 44019
0 44021 7 1 2 44018 44020
0 44022 7 1 2 94956 44021
0 44023 5 1 1 44022
0 44024 7 1 2 44012 44023
0 44025 5 1 1 44024
0 44026 7 1 2 57482 44025
0 44027 5 1 1 44026
0 44028 7 1 2 87215 94397
0 44029 5 2 1 44028
0 44030 7 1 2 91547 94959
0 44031 5 1 1 44030
0 44032 7 2 2 84012 86652
0 44033 5 1 1 94961
0 44034 7 1 2 44031 44033
0 44035 5 1 1 44034
0 44036 7 1 2 59007 44035
0 44037 5 1 1 44036
0 44038 7 1 2 88247 93949
0 44039 5 1 1 44038
0 44040 7 1 2 44037 44039
0 44041 5 1 1 44040
0 44042 7 1 2 59648 44041
0 44043 5 1 1 44042
0 44044 7 1 2 44027 44043
0 44045 5 1 1 44044
0 44046 7 1 2 57773 44045
0 44047 5 1 1 44046
0 44048 7 3 2 73728 75694
0 44049 7 1 2 68789 84799
0 44050 7 1 2 94963 44049
0 44051 5 1 1 44050
0 44052 7 1 2 44047 44051
0 44053 5 1 1 44052
0 44054 7 1 2 94653 44053
0 44055 5 1 1 44054
0 44056 7 4 2 87503 94284
0 44057 5 1 1 94966
0 44058 7 1 2 39246 44057
0 44059 5 1 1 44058
0 44060 7 1 2 76462 44059
0 44061 5 1 1 44060
0 44062 7 3 2 59911 86570
0 44063 7 1 2 77220 94970
0 44064 5 1 1 44063
0 44065 7 1 2 44061 44064
0 44066 5 1 1 44065
0 44067 7 1 2 65693 44066
0 44068 5 1 1 44067
0 44069 7 1 2 74819 69893
0 44070 5 1 1 44069
0 44071 7 1 2 57483 44070
0 44072 5 1 1 44071
0 44073 7 1 2 81803 44072
0 44074 5 1 1 44073
0 44075 7 1 2 94967 44074
0 44076 5 1 1 44075
0 44077 7 1 2 44068 44076
0 44078 5 1 1 44077
0 44079 7 1 2 78913 82643
0 44080 7 1 2 44078 44079
0 44081 5 1 1 44080
0 44082 7 1 2 44055 44081
0 44083 7 1 2 43993 44082
0 44084 7 1 2 43953 44083
0 44085 7 1 2 43891 44084
0 44086 7 1 2 43747 44085
0 44087 5 1 1 44086
0 44088 7 1 2 67481 44087
0 44089 5 1 1 44088
0 44090 7 1 2 43406 44089
0 44091 5 1 1 44090
0 44092 7 1 2 64829 88299
0 44093 7 1 2 44091 44092
0 44094 5 1 1 44093
0 44095 7 1 2 42735 44094
0 44096 5 1 1 44095
0 44097 7 1 2 58885 44096
0 44098 5 1 1 44097
0 44099 7 1 2 86089 83821
0 44100 7 1 2 94238 44099
0 44101 5 1 1 44100
0 44102 7 1 2 74156 90350
0 44103 7 1 2 94518 44102
0 44104 7 1 2 94850 44103
0 44105 5 1 1 44104
0 44106 7 1 2 44101 44105
0 44107 5 1 1 44106
0 44108 7 1 2 69119 44107
0 44109 5 1 1 44108
0 44110 7 1 2 89753 94312
0 44111 5 1 1 44110
0 44112 7 1 2 44109 44111
0 44113 5 1 1 44112
0 44114 7 1 2 64830 44113
0 44115 5 1 1 44114
0 44116 7 2 2 61430 91235
0 44117 5 1 1 94973
0 44118 7 2 2 70306 94974
0 44119 7 1 2 69212 94714
0 44120 7 1 2 94975 44119
0 44121 5 1 1 44120
0 44122 7 1 2 44115 44121
0 44123 5 1 1 44122
0 44124 7 1 2 60045 44123
0 44125 5 1 1 44124
0 44126 7 1 2 75277 87220
0 44127 5 1 1 44126
0 44128 7 1 2 86238 91491
0 44129 5 1 1 44128
0 44130 7 1 2 44127 44129
0 44131 5 1 1 44130
0 44132 7 1 2 62519 44131
0 44133 5 1 1 44132
0 44134 7 1 2 89483 91492
0 44135 5 1 1 44134
0 44136 7 1 2 44133 44135
0 44137 5 2 1 44136
0 44138 7 1 2 84876 89957
0 44139 7 1 2 94977 44138
0 44140 5 1 1 44139
0 44141 7 1 2 44125 44140
0 44142 5 1 1 44141
0 44143 7 1 2 61966 44142
0 44144 5 1 1 44143
0 44145 7 1 2 82964 93290
0 44146 5 1 1 44145
0 44147 7 1 2 90802 44146
0 44148 5 1 1 44147
0 44149 7 1 2 84274 37815
0 44150 5 1 1 44149
0 44151 7 1 2 85175 83960
0 44152 7 1 2 85351 44151
0 44153 5 1 1 44152
0 44154 7 1 2 44150 44153
0 44155 7 1 2 44148 44154
0 44156 5 1 1 44155
0 44157 7 1 2 60654 44156
0 44158 5 1 1 44157
0 44159 7 1 2 94873 44158
0 44160 5 1 1 44159
0 44161 7 1 2 93552 44160
0 44162 5 1 1 44161
0 44163 7 1 2 94877 44162
0 44164 5 1 1 44163
0 44165 7 1 2 94536 44164
0 44166 5 1 1 44165
0 44167 7 5 2 60655 84673
0 44168 7 1 2 84886 94979
0 44169 5 1 1 44168
0 44170 7 2 2 66037 92803
0 44171 5 1 1 94984
0 44172 7 1 2 87781 94985
0 44173 5 1 1 44172
0 44174 7 1 2 44169 44173
0 44175 5 1 1 44174
0 44176 7 1 2 87998 44175
0 44177 5 1 1 44176
0 44178 7 1 2 65081 81202
0 44179 5 2 1 44178
0 44180 7 1 2 60409 76973
0 44181 5 1 1 44180
0 44182 7 2 2 94986 44181
0 44183 5 1 1 94988
0 44184 7 1 2 61431 44183
0 44185 5 1 1 44184
0 44186 7 1 2 78738 73018
0 44187 7 1 2 73219 44186
0 44188 5 1 1 44187
0 44189 7 1 2 44185 44188
0 44190 5 1 1 44189
0 44191 7 1 2 84993 44190
0 44192 5 1 1 44191
0 44193 7 1 2 75472 77575
0 44194 5 1 1 44193
0 44195 7 1 2 44192 44194
0 44196 5 1 1 44195
0 44197 7 1 2 61692 44196
0 44198 5 1 1 44197
0 44199 7 1 2 44177 44198
0 44200 5 1 1 44199
0 44201 7 1 2 61061 44200
0 44202 5 1 1 44201
0 44203 7 1 2 80942 84589
0 44204 5 1 1 44203
0 44205 7 2 2 61693 84349
0 44206 7 1 2 66038 94990
0 44207 5 1 1 44206
0 44208 7 1 2 44204 44207
0 44209 5 1 1 44208
0 44210 7 1 2 77168 44209
0 44211 5 1 1 44210
0 44212 7 1 2 81237 86497
0 44213 5 1 1 44212
0 44214 7 1 2 44211 44213
0 44215 5 1 1 44214
0 44216 7 1 2 63396 44215
0 44217 5 1 1 44216
0 44218 7 3 2 72154 84781
0 44219 7 1 2 86877 94992
0 44220 5 1 1 44219
0 44221 7 1 2 80436 81447
0 44222 7 1 2 84827 44221
0 44223 5 1 1 44222
0 44224 7 1 2 44220 44223
0 44225 7 1 2 44217 44224
0 44226 5 1 1 44225
0 44227 7 1 2 71327 44226
0 44228 5 1 1 44227
0 44229 7 1 2 91685 92388
0 44230 5 2 1 44229
0 44231 7 1 2 92501 94995
0 44232 5 1 1 44231
0 44233 7 1 2 85176 78554
0 44234 7 1 2 75776 44233
0 44235 5 1 1 44234
0 44236 7 1 2 44232 44235
0 44237 5 1 1 44236
0 44238 7 1 2 60656 44237
0 44239 5 1 1 44238
0 44240 7 1 2 85177 84503
0 44241 7 1 2 84044 44240
0 44242 5 1 1 44241
0 44243 7 1 2 44239 44242
0 44244 5 1 1 44243
0 44245 7 1 2 61694 44244
0 44246 5 1 1 44245
0 44247 7 1 2 80821 84755
0 44248 5 1 1 44247
0 44249 7 1 2 44246 44248
0 44250 5 1 1 44249
0 44251 7 1 2 61062 44250
0 44252 5 1 1 44251
0 44253 7 1 2 44228 44252
0 44254 5 1 1 44253
0 44255 7 1 2 68163 44254
0 44256 5 1 1 44255
0 44257 7 2 2 61432 69508
0 44258 5 1 1 94997
0 44259 7 1 2 86742 44258
0 44260 5 3 1 44259
0 44261 7 1 2 67789 94999
0 44262 5 1 1 44261
0 44263 7 1 2 60410 92392
0 44264 5 1 1 44263
0 44265 7 1 2 44262 44264
0 44266 5 1 1 44265
0 44267 7 1 2 60657 44266
0 44268 5 1 1 44267
0 44269 7 1 2 68265 95000
0 44270 5 1 1 44269
0 44271 7 1 2 44268 44270
0 44272 5 1 1 44271
0 44273 7 1 2 61695 44272
0 44274 5 1 1 44273
0 44275 7 1 2 84195 84674
0 44276 5 2 1 44275
0 44277 7 1 2 91075 95002
0 44278 5 1 1 44277
0 44279 7 1 2 63397 44278
0 44280 5 1 1 44279
0 44281 7 2 2 65311 84782
0 44282 7 1 2 79497 95004
0 44283 5 1 1 44282
0 44284 7 1 2 44280 44283
0 44285 5 1 1 44284
0 44286 7 1 2 76966 44285
0 44287 5 1 1 44286
0 44288 7 1 2 94991 95001
0 44289 5 1 1 44288
0 44290 7 1 2 79498 90485
0 44291 5 1 1 44290
0 44292 7 1 2 44289 44291
0 44293 5 1 1 44292
0 44294 7 1 2 68879 44293
0 44295 5 1 1 44294
0 44296 7 1 2 44287 44295
0 44297 7 1 2 44274 44296
0 44298 5 1 1 44297
0 44299 7 1 2 61063 44298
0 44300 5 1 1 44299
0 44301 7 1 2 93630 94448
0 44302 5 1 1 44301
0 44303 7 1 2 44300 44302
0 44304 5 1 1 44303
0 44305 7 1 2 76221 44304
0 44306 5 1 1 44305
0 44307 7 1 2 86660 84600
0 44308 5 1 1 44307
0 44309 7 1 2 73019 87782
0 44310 7 1 2 93632 44309
0 44311 5 1 1 44310
0 44312 7 1 2 44308 44311
0 44313 5 1 1 44312
0 44314 7 1 2 69063 44313
0 44315 5 1 1 44314
0 44316 7 2 2 60658 84994
0 44317 7 1 2 78189 77898
0 44318 7 1 2 95006 44317
0 44319 5 1 1 44318
0 44320 7 1 2 12870 44319
0 44321 5 1 1 44320
0 44322 7 1 2 86498 44321
0 44323 5 1 1 44322
0 44324 7 1 2 44315 44323
0 44325 7 1 2 44306 44324
0 44326 7 1 2 44256 44325
0 44327 7 1 2 44202 44326
0 44328 5 1 1 44327
0 44329 7 1 2 66617 44328
0 44330 5 1 1 44329
0 44331 7 1 2 85178 94273
0 44332 5 1 1 44331
0 44333 7 1 2 93058 44332
0 44334 5 1 1 44333
0 44335 7 1 2 85487 44334
0 44336 5 1 1 44335
0 44337 7 1 2 91178 44336
0 44338 5 1 1 44337
0 44339 7 1 2 90634 44338
0 44340 5 1 1 44339
0 44341 7 1 2 73573 81705
0 44342 5 2 1 44341
0 44343 7 1 2 57774 95008
0 44344 5 1 1 44343
0 44345 7 1 2 74079 81706
0 44346 5 1 1 44345
0 44347 7 1 2 70873 44346
0 44348 5 1 1 44347
0 44349 7 1 2 93833 44348
0 44350 7 1 2 44344 44349
0 44351 5 1 1 44350
0 44352 7 1 2 83165 82660
0 44353 7 1 2 44351 44352
0 44354 5 1 1 44353
0 44355 7 1 2 44340 44354
0 44356 5 1 1 44355
0 44357 7 1 2 65694 44356
0 44358 5 1 1 44357
0 44359 7 3 2 66618 84783
0 44360 7 1 2 73918 85179
0 44361 5 1 1 44360
0 44362 7 1 2 82965 44361
0 44363 5 1 1 44362
0 44364 7 1 2 95010 44363
0 44365 5 1 1 44364
0 44366 7 2 2 67596 87660
0 44367 7 1 2 71345 94519
0 44368 7 1 2 95013 44367
0 44369 5 1 1 44368
0 44370 7 1 2 44365 44369
0 44371 5 1 1 44370
0 44372 7 1 2 69429 44371
0 44373 5 1 1 44372
0 44374 7 3 2 88248 91771
0 44375 7 1 2 93118 95015
0 44376 5 2 1 44375
0 44377 7 1 2 68043 84954
0 44378 7 3 2 65312 82661
0 44379 7 1 2 86855 95020
0 44380 7 1 2 44377 44379
0 44381 5 1 1 44380
0 44382 7 1 2 95018 44381
0 44383 5 1 1 44382
0 44384 7 1 2 68408 44383
0 44385 5 1 1 44384
0 44386 7 1 2 78734 86318
0 44387 7 1 2 83124 87661
0 44388 7 1 2 44386 44387
0 44389 5 1 1 44388
0 44390 7 1 2 95019 44389
0 44391 5 1 1 44390
0 44392 7 1 2 58340 44391
0 44393 5 1 1 44392
0 44394 7 1 2 44385 44393
0 44395 7 1 2 44373 44394
0 44396 7 1 2 44358 44395
0 44397 7 1 2 44330 44396
0 44398 5 1 1 44397
0 44399 7 1 2 64831 44398
0 44400 5 1 1 44399
0 44401 7 1 2 44166 44400
0 44402 5 1 1 44401
0 44403 7 1 2 59912 44402
0 44404 5 1 1 44403
0 44405 7 1 2 85762 84784
0 44406 5 2 1 44405
0 44407 7 4 2 66336 91184
0 44408 5 1 1 95025
0 44409 7 1 2 60411 95026
0 44410 5 1 1 44409
0 44411 7 1 2 91407 44410
0 44412 5 1 1 44411
0 44413 7 1 2 66039 44412
0 44414 5 1 1 44413
0 44415 7 1 2 95023 44414
0 44416 5 1 1 44415
0 44417 7 1 2 68880 44416
0 44418 5 1 1 44417
0 44419 7 1 2 84504 95027
0 44420 5 1 1 44419
0 44421 7 1 2 44418 44420
0 44422 5 1 1 44421
0 44423 7 1 2 84350 44422
0 44424 5 1 1 44423
0 44425 7 1 2 79050 33210
0 44426 5 1 1 44425
0 44427 7 1 2 58638 85593
0 44428 7 1 2 44426 44427
0 44429 5 1 1 44428
0 44430 7 1 2 66040 93037
0 44431 5 1 1 44430
0 44432 7 1 2 61696 44431
0 44433 7 1 2 44429 44432
0 44434 5 1 1 44433
0 44435 7 1 2 93626 94996
0 44436 5 1 1 44435
0 44437 7 1 2 66337 92394
0 44438 7 1 2 44436 44437
0 44439 5 1 1 44438
0 44440 7 1 2 68164 44439
0 44441 7 1 2 44434 44440
0 44442 5 1 1 44441
0 44443 7 2 2 84675 92804
0 44444 5 1 1 95029
0 44445 7 1 2 86701 44444
0 44446 5 1 1 44445
0 44447 7 1 2 76222 44446
0 44448 5 1 1 44447
0 44449 7 1 2 84676 93783
0 44450 5 1 1 44449
0 44451 7 1 2 44448 44450
0 44452 5 1 1 44451
0 44453 7 1 2 71785 44452
0 44454 5 1 1 44453
0 44455 7 1 2 84532 86499
0 44456 5 1 1 44455
0 44457 7 1 2 72807 86828
0 44458 7 1 2 92856 44457
0 44459 5 1 1 44458
0 44460 7 1 2 44456 44459
0 44461 5 1 1 44460
0 44462 7 1 2 60659 44461
0 44463 5 1 1 44462
0 44464 7 1 2 44454 44463
0 44465 5 1 1 44464
0 44466 7 1 2 69064 44465
0 44467 5 1 1 44466
0 44468 7 1 2 77047 74011
0 44469 5 1 1 44468
0 44470 7 1 2 60412 86023
0 44471 5 1 1 44470
0 44472 7 1 2 44469 44471
0 44473 5 1 1 44472
0 44474 7 1 2 58639 44473
0 44475 5 1 1 44474
0 44476 7 1 2 73862 84513
0 44477 7 1 2 89717 44476
0 44478 5 1 1 44477
0 44479 7 1 2 44475 44478
0 44480 5 1 1 44479
0 44481 7 1 2 61697 44480
0 44482 5 1 1 44481
0 44483 7 1 2 87808 44482
0 44484 5 1 1 44483
0 44485 7 1 2 66041 44484
0 44486 5 1 1 44485
0 44487 7 1 2 91408 44408
0 44488 5 1 1 44487
0 44489 7 1 2 66042 44488
0 44490 5 1 1 44489
0 44491 7 1 2 44490 95024
0 44492 5 1 1 44491
0 44493 7 1 2 81089 44492
0 44494 5 1 1 44493
0 44495 7 1 2 87226 84745
0 44496 5 1 1 44495
0 44497 7 1 2 67026 89932
0 44498 7 1 2 84756 44497
0 44499 5 1 1 44498
0 44500 7 1 2 44496 44499
0 44501 5 1 1 44500
0 44502 7 1 2 76223 44501
0 44503 5 1 1 44502
0 44504 7 1 2 84677 93792
0 44505 5 1 1 44504
0 44506 7 1 2 44503 44505
0 44507 5 1 1 44506
0 44508 7 1 2 79121 44507
0 44509 5 1 1 44508
0 44510 7 1 2 69849 77496
0 44511 5 2 1 44510
0 44512 7 1 2 58640 67569
0 44513 5 1 1 44512
0 44514 7 1 2 95031 44513
0 44515 5 1 1 44514
0 44516 7 1 2 85472 44515
0 44517 5 1 1 44516
0 44518 7 1 2 60660 83329
0 44519 5 1 1 44518
0 44520 7 1 2 95032 44519
0 44521 5 1 1 44520
0 44522 7 1 2 84995 44521
0 44523 5 1 1 44522
0 44524 7 1 2 44517 44523
0 44525 5 1 1 44524
0 44526 7 1 2 66338 44525
0 44527 5 1 1 44526
0 44528 7 1 2 78537 77719
0 44529 7 1 2 76975 44528
0 44530 5 1 1 44529
0 44531 7 1 2 86863 44530
0 44532 5 1 1 44531
0 44533 7 1 2 44527 44532
0 44534 5 1 1 44533
0 44535 7 1 2 61433 44534
0 44536 5 1 1 44535
0 44537 7 1 2 44509 44536
0 44538 7 1 2 44494 44537
0 44539 7 1 2 44486 44538
0 44540 7 1 2 44467 44539
0 44541 7 1 2 44442 44540
0 44542 7 1 2 44424 44541
0 44543 5 1 1 44542
0 44544 7 1 2 61064 44543
0 44545 5 1 1 44544
0 44546 7 1 2 74134 93634
0 44547 5 1 1 44546
0 44548 7 1 2 75449 93385
0 44549 5 1 1 44548
0 44550 7 1 2 44547 44549
0 44551 5 1 1 44550
0 44552 7 1 2 78879 44551
0 44553 5 1 1 44552
0 44554 7 1 2 89851 92912
0 44555 5 1 1 44554
0 44556 7 1 2 90993 44555
0 44557 5 1 1 44556
0 44558 7 1 2 44553 44557
0 44559 5 1 1 44558
0 44560 7 1 2 61698 44559
0 44561 5 1 1 44560
0 44562 7 2 2 80542 91465
0 44563 5 1 1 95033
0 44564 7 1 2 84196 78880
0 44565 7 1 2 95034 44564
0 44566 5 1 1 44565
0 44567 7 1 2 44561 44566
0 44568 5 1 1 44567
0 44569 7 1 2 66043 44568
0 44570 5 1 1 44569
0 44571 7 1 2 59649 69880
0 44572 5 1 1 44571
0 44573 7 1 2 73335 44572
0 44574 5 1 1 44573
0 44575 7 1 2 57775 44574
0 44576 5 1 1 44575
0 44577 7 1 2 59161 85824
0 44578 5 1 1 44577
0 44579 7 1 2 44576 44578
0 44580 5 1 1 44579
0 44581 7 1 2 68790 44580
0 44582 5 1 1 44581
0 44583 7 1 2 12184 44582
0 44584 5 1 1 44583
0 44585 7 1 2 65313 44584
0 44586 5 1 1 44585
0 44587 7 1 2 73676 81660
0 44588 5 1 1 44587
0 44589 7 1 2 44586 44588
0 44590 5 1 1 44589
0 44591 7 1 2 61699 44590
0 44592 5 1 1 44591
0 44593 7 1 2 66044 94796
0 44594 5 1 1 44593
0 44595 7 1 2 44592 44594
0 44596 5 1 1 44595
0 44597 7 1 2 63398 44596
0 44598 5 1 1 44597
0 44599 7 1 2 85180 93386
0 44600 5 1 1 44599
0 44601 7 1 2 80943 78666
0 44602 5 1 1 44601
0 44603 7 1 2 44600 44602
0 44604 5 1 1 44603
0 44605 7 1 2 78881 44604
0 44606 5 1 1 44605
0 44607 7 1 2 85181 33145
0 44608 5 1 1 44607
0 44609 7 1 2 44606 44608
0 44610 5 1 1 44609
0 44611 7 1 2 65695 44610
0 44612 5 1 1 44611
0 44613 7 1 2 68881 90385
0 44614 5 1 1 44613
0 44615 7 1 2 82930 44614
0 44616 5 1 1 44615
0 44617 7 1 2 66339 44616
0 44618 7 1 2 44612 44617
0 44619 5 1 1 44618
0 44620 7 1 2 80589 94275
0 44621 5 1 1 44620
0 44622 7 1 2 61700 93815
0 44623 7 1 2 44621 44622
0 44624 5 1 1 44623
0 44625 7 1 2 61434 44624
0 44626 7 1 2 44619 44625
0 44627 5 1 1 44626
0 44628 7 1 2 44598 44627
0 44629 7 1 2 44570 44628
0 44630 7 1 2 44545 44629
0 44631 5 1 1 44630
0 44632 7 1 2 66980 44631
0 44633 5 1 1 44632
0 44634 7 1 2 81961 94612
0 44635 5 1 1 44634
0 44636 7 1 2 63918 44635
0 44637 5 1 1 44636
0 44638 7 1 2 94772 44637
0 44639 5 1 1 44638
0 44640 7 1 2 62520 44639
0 44641 5 1 1 44640
0 44642 7 1 2 67223 80740
0 44643 5 1 1 44642
0 44644 7 1 2 83848 28970
0 44645 5 1 1 44644
0 44646 7 1 2 68165 44645
0 44647 5 1 1 44646
0 44648 7 1 2 44643 44647
0 44649 7 1 2 44641 44648
0 44650 5 1 1 44649
0 44651 7 1 2 61435 44650
0 44652 5 1 1 44651
0 44653 7 1 2 81840 91550
0 44654 5 1 1 44653
0 44655 7 1 2 44652 44654
0 44656 5 1 1 44655
0 44657 7 1 2 71328 44656
0 44658 5 1 1 44657
0 44659 7 1 2 85182 94310
0 44660 5 1 1 44659
0 44661 7 1 2 14413 94305
0 44662 5 1 1 44661
0 44663 7 1 2 94603 94801
0 44664 5 1 1 44663
0 44665 7 1 2 66340 44664
0 44666 7 1 2 44662 44665
0 44667 7 1 2 44660 44666
0 44668 7 1 2 44658 44667
0 44669 5 1 1 44668
0 44670 7 1 2 58341 93390
0 44671 5 1 1 44670
0 44672 7 1 2 73677 44671
0 44673 5 1 1 44672
0 44674 7 1 2 85790 93996
0 44675 5 1 1 44674
0 44676 7 2 2 68044 86267
0 44677 5 3 1 95035
0 44678 7 1 2 73698 95036
0 44679 5 1 1 44678
0 44680 7 1 2 44675 44679
0 44681 7 2 2 44673 44680
0 44682 7 1 2 61701 95040
0 44683 5 1 1 44682
0 44684 7 1 2 61065 44683
0 44685 7 1 2 44669 44684
0 44686 5 1 1 44685
0 44687 7 1 2 90014 41796
0 44688 5 1 1 44687
0 44689 7 1 2 80260 92845
0 44690 5 3 1 44689
0 44691 7 1 2 58075 95042
0 44692 5 2 1 44691
0 44693 7 1 2 94644 95043
0 44694 5 1 1 44693
0 44695 7 1 2 95045 44694
0 44696 5 2 1 44695
0 44697 7 1 2 94790 95047
0 44698 7 1 2 44688 44697
0 44699 5 1 1 44698
0 44700 7 2 2 78342 72730
0 44701 5 1 1 95049
0 44702 7 1 2 77498 70050
0 44703 5 1 1 44702
0 44704 7 1 2 95050 44703
0 44705 5 1 1 44704
0 44706 7 1 2 66045 44705
0 44707 5 1 1 44706
0 44708 7 1 2 81712 44707
0 44709 5 1 1 44708
0 44710 7 1 2 65696 44709
0 44711 5 1 1 44710
0 44712 7 1 2 94792 44711
0 44713 5 1 1 44712
0 44714 7 1 2 63399 44713
0 44715 7 1 2 44699 44714
0 44716 5 1 1 44715
0 44717 7 2 2 66341 80521
0 44718 7 1 2 80869 95051
0 44719 5 1 1 44718
0 44720 7 1 2 16294 44719
0 44721 5 1 1 44720
0 44722 7 1 2 62262 44721
0 44723 5 1 1 44722
0 44724 7 2 2 66342 69065
0 44725 7 1 2 85451 95053
0 44726 5 1 1 44725
0 44727 7 1 2 94809 44726
0 44728 7 1 2 44723 44727
0 44729 5 1 1 44728
0 44730 7 1 2 67790 44729
0 44731 5 1 1 44730
0 44732 7 1 2 94807 44563
0 44733 5 1 1 44732
0 44734 7 1 2 69066 44733
0 44735 5 1 1 44734
0 44736 7 2 2 79228 89890
0 44737 5 1 1 95055
0 44738 7 1 2 81270 44737
0 44739 5 1 1 44738
0 44740 7 1 2 94641 44739
0 44741 5 1 1 44740
0 44742 7 1 2 44735 44741
0 44743 7 1 2 75402 81474
0 44744 7 1 2 93623 44743
0 44745 5 1 1 44744
0 44746 7 1 2 81271 44745
0 44747 5 1 1 44746
0 44748 7 1 2 77680 44747
0 44749 5 1 1 44748
0 44750 7 1 2 66343 94805
0 44751 5 1 1 44750
0 44752 7 1 2 63090 86807
0 44753 7 1 2 44751 44752
0 44754 5 1 1 44753
0 44755 7 1 2 44749 44754
0 44756 7 1 2 44742 44755
0 44757 7 1 2 44731 44756
0 44758 5 1 1 44757
0 44759 7 1 2 73699 44758
0 44760 5 1 1 44759
0 44761 7 1 2 86966 31320
0 44762 5 1 1 44761
0 44763 7 1 2 68529 44762
0 44764 5 1 1 44763
0 44765 7 1 2 60661 91766
0 44766 5 1 1 44765
0 44767 7 1 2 22671 95003
0 44768 5 1 1 44767
0 44769 7 1 2 68882 44768
0 44770 5 1 1 44769
0 44771 7 1 2 44766 44770
0 44772 7 1 2 44764 44771
0 44773 5 1 1 44772
0 44774 7 1 2 76224 44773
0 44775 5 1 1 44774
0 44776 7 2 2 68166 85647
0 44777 5 1 1 95057
0 44778 7 1 2 66344 95058
0 44779 5 1 1 44778
0 44780 7 1 2 73097 80161
0 44781 7 1 2 92550 44780
0 44782 5 1 1 44781
0 44783 7 1 2 44779 44782
0 44784 7 1 2 44775 44783
0 44785 5 1 1 44784
0 44786 7 1 2 67791 44785
0 44787 5 1 1 44786
0 44788 7 2 2 77593 84678
0 44789 5 1 1 95059
0 44790 7 1 2 69400 87479
0 44791 5 1 1 44790
0 44792 7 1 2 44789 44791
0 44793 5 1 1 44792
0 44794 7 1 2 83781 44793
0 44795 5 1 1 44794
0 44796 7 1 2 77576 91689
0 44797 5 1 1 44796
0 44798 7 1 2 24587 44797
0 44799 5 1 1 44798
0 44800 7 1 2 77681 44799
0 44801 5 1 1 44800
0 44802 7 1 2 44795 44801
0 44803 5 1 1 44802
0 44804 7 1 2 68883 44803
0 44805 5 1 1 44804
0 44806 7 1 2 76890 34985
0 44807 5 1 1 44806
0 44808 7 1 2 84757 44807
0 44809 5 1 1 44808
0 44810 7 1 2 68167 86007
0 44811 5 1 1 44810
0 44812 7 1 2 76225 84962
0 44813 5 1 1 44812
0 44814 7 1 2 70430 44813
0 44815 7 1 2 44811 44814
0 44816 5 1 1 44815
0 44817 7 1 2 91767 44816
0 44818 5 1 1 44817
0 44819 7 1 2 44809 44818
0 44820 7 1 2 44805 44819
0 44821 7 1 2 44787 44820
0 44822 7 1 2 44760 44821
0 44823 7 1 2 44716 44822
0 44824 7 1 2 44686 44823
0 44825 5 1 1 44824
0 44826 7 1 2 67059 44825
0 44827 5 1 1 44826
0 44828 7 1 2 44633 44827
0 44829 5 1 1 44828
0 44830 7 1 2 64617 44829
0 44831 5 1 1 44830
0 44832 7 1 2 66981 93741
0 44833 5 1 1 44832
0 44834 7 1 2 69894 91050
0 44835 5 1 1 44834
0 44836 7 1 2 74820 93649
0 44837 5 1 1 44836
0 44838 7 1 2 93752 44837
0 44839 7 1 2 44835 44838
0 44840 5 1 1 44839
0 44841 7 1 2 61066 44840
0 44842 5 1 1 44841
0 44843 7 1 2 94645 44842
0 44844 5 1 1 44843
0 44845 7 1 2 62793 44844
0 44846 5 1 1 44845
0 44847 7 1 2 80081 89420
0 44848 5 1 1 44847
0 44849 7 1 2 60662 44848
0 44850 5 1 1 44849
0 44851 7 1 2 76082 79513
0 44852 5 1 1 44851
0 44853 7 1 2 44850 44852
0 44854 5 1 1 44853
0 44855 7 1 2 62263 44854
0 44856 5 1 1 44855
0 44857 7 1 2 60663 87999
0 44858 5 1 1 44857
0 44859 7 1 2 79122 78305
0 44860 5 1 1 44859
0 44861 7 1 2 74946 92896
0 44862 7 1 2 44860 44861
0 44863 7 1 2 44858 44862
0 44864 5 1 1 44863
0 44865 7 1 2 61067 44864
0 44866 5 1 1 44865
0 44867 7 1 2 44856 44866
0 44868 5 1 1 44867
0 44869 7 1 2 64102 44868
0 44870 5 1 1 44869
0 44871 7 1 2 44846 44870
0 44872 5 1 1 44871
0 44873 7 1 2 61436 44872
0 44874 5 1 1 44873
0 44875 7 1 2 77157 83407
0 44876 5 1 1 44875
0 44877 7 1 2 61437 44876
0 44878 5 1 1 44877
0 44879 7 1 2 64103 84999
0 44880 5 1 1 44879
0 44881 7 1 2 44878 44880
0 44882 5 1 1 44881
0 44883 7 1 2 60664 75934
0 44884 7 1 2 44882 44883
0 44885 5 1 1 44884
0 44886 7 1 2 44874 44885
0 44887 5 1 1 44886
0 44888 7 1 2 71329 44887
0 44889 5 1 1 44888
0 44890 7 1 2 94158 94161
0 44891 5 1 1 44890
0 44892 7 1 2 73134 78753
0 44893 5 1 1 44892
0 44894 7 1 2 72936 44893
0 44895 5 1 1 44894
0 44896 7 1 2 62794 44895
0 44897 5 1 1 44896
0 44898 7 1 2 83961 94169
0 44899 5 1 1 44898
0 44900 7 1 2 87028 44899
0 44901 7 1 2 44897 44900
0 44902 7 1 2 44891 44901
0 44903 5 1 1 44902
0 44904 7 1 2 71451 44903
0 44905 5 1 1 44904
0 44906 7 1 2 44889 44905
0 44907 5 1 1 44906
0 44908 7 1 2 67060 44907
0 44909 5 1 1 44908
0 44910 7 1 2 44833 44909
0 44911 5 1 1 44910
0 44912 7 1 2 82883 44911
0 44913 5 1 1 44912
0 44914 7 1 2 67061 91185
0 44915 7 1 2 94978 44914
0 44916 5 1 1 44915
0 44917 7 1 2 44913 44916
0 44918 7 1 2 44831 44917
0 44919 7 1 2 44404 44918
0 44920 5 1 1 44919
0 44921 7 1 2 64737 44920
0 44922 5 1 1 44921
0 44923 7 1 2 44144 44922
0 44924 5 1 1 44923
0 44925 7 1 2 63529 44924
0 44926 5 1 1 44925
0 44927 7 2 2 84679 74909
0 44928 5 1 1 95061
0 44929 7 1 2 94527 95062
0 44930 5 1 1 44929
0 44931 7 1 2 86500 91329
0 44932 5 1 1 44931
0 44933 7 1 2 44930 44932
0 44934 5 1 1 44933
0 44935 7 1 2 57776 44934
0 44936 5 1 1 44935
0 44937 7 2 2 84785 94654
0 44938 7 1 2 94964 95063
0 44939 5 1 1 44938
0 44940 7 1 2 44936 44939
0 44941 5 1 1 44940
0 44942 7 1 2 68934 44941
0 44943 5 1 1 44942
0 44944 7 1 2 73550 72912
0 44945 7 1 2 74850 44944
0 44946 7 1 2 91813 44945
0 44947 5 1 1 44946
0 44948 7 1 2 44943 44947
0 44949 5 1 1 44948
0 44950 7 1 2 64832 44949
0 44951 5 1 1 44950
0 44952 7 3 2 76061 87915
0 44953 7 2 2 81119 95065
0 44954 7 1 2 61068 94629
0 44955 7 1 2 95068 44954
0 44956 5 1 1 44955
0 44957 7 1 2 44951 44956
0 44958 5 1 1 44957
0 44959 7 1 2 59162 44958
0 44960 5 1 1 44959
0 44961 7 2 2 59650 67062
0 44962 5 1 1 95070
0 44963 7 1 2 72706 92228
0 44964 5 1 1 44963
0 44965 7 1 2 44962 44964
0 44966 5 1 1 44965
0 44967 7 1 2 66791 44966
0 44968 5 1 1 44967
0 44969 7 1 2 75685 82278
0 44970 5 1 1 44969
0 44971 7 1 2 44968 44970
0 44972 5 1 1 44971
0 44973 7 1 2 75555 81510
0 44974 7 1 2 44972 44973
0 44975 5 1 1 44974
0 44976 7 1 2 44960 44975
0 44977 5 1 1 44976
0 44978 7 1 2 65314 44977
0 44979 5 1 1 44978
0 44980 7 1 2 70307 89823
0 44981 5 1 1 44980
0 44982 7 1 2 32346 44981
0 44983 5 1 1 44982
0 44984 7 1 2 87846 91776
0 44985 7 1 2 44983 44984
0 44986 5 1 1 44985
0 44987 7 1 2 44979 44986
0 44988 5 1 1 44987
0 44989 7 1 2 68635 44988
0 44990 5 1 1 44989
0 44991 7 1 2 78882 82850
0 44992 5 1 1 44991
0 44993 7 1 2 94114 44992
0 44994 5 1 1 44993
0 44995 7 1 2 76700 44994
0 44996 5 1 1 44995
0 44997 7 1 2 87069 94914
0 44998 5 1 1 44997
0 44999 7 1 2 44996 44998
0 45000 5 1 1 44999
0 45001 7 1 2 60665 45000
0 45002 5 1 1 45001
0 45003 7 1 2 76701 38773
0 45004 5 1 1 45003
0 45005 7 1 2 45002 45004
0 45006 5 1 1 45005
0 45007 7 1 2 61069 45006
0 45008 5 1 1 45007
0 45009 7 1 2 75581 94097
0 45010 5 1 1 45009
0 45011 7 1 2 94099 45010
0 45012 5 1 1 45011
0 45013 7 1 2 94104 45012
0 45014 5 1 1 45013
0 45015 7 1 2 76702 45014
0 45016 5 1 1 45015
0 45017 7 1 2 70843 88488
0 45018 5 1 1 45017
0 45019 7 1 2 85931 77537
0 45020 5 1 1 45019
0 45021 7 1 2 61070 45020
0 45022 5 1 1 45021
0 45023 7 1 2 62264 78201
0 45024 5 2 1 45023
0 45025 7 1 2 64104 86387
0 45026 5 1 1 45025
0 45027 7 1 2 71218 78222
0 45028 7 1 2 45026 45027
0 45029 7 1 2 95072 45028
0 45030 7 1 2 45022 45029
0 45031 7 1 2 45018 45030
0 45032 5 1 1 45031
0 45033 7 1 2 75556 45032
0 45034 5 1 1 45033
0 45035 7 1 2 45016 45034
0 45036 7 1 2 45008 45035
0 45037 5 1 1 45036
0 45038 7 1 2 61438 45037
0 45039 5 1 1 45038
0 45040 7 1 2 58342 94888
0 45041 5 1 1 45040
0 45042 7 1 2 75557 45041
0 45043 5 1 1 45042
0 45044 7 2 2 77400 94605
0 45045 7 1 2 92413 94089
0 45046 7 1 2 95074 45045
0 45047 5 1 1 45046
0 45048 7 1 2 45043 45047
0 45049 5 1 1 45048
0 45050 7 1 2 81147 45049
0 45051 5 1 1 45050
0 45052 7 1 2 63091 92749
0 45053 5 2 1 45052
0 45054 7 1 2 93466 95076
0 45055 5 1 1 45054
0 45056 7 1 2 62265 45055
0 45057 5 1 1 45056
0 45058 7 1 2 78216 87088
0 45059 5 1 1 45058
0 45060 7 1 2 73901 45059
0 45061 5 1 1 45060
0 45062 7 1 2 63092 45061
0 45063 5 1 1 45062
0 45064 7 1 2 45057 45063
0 45065 5 1 1 45064
0 45066 7 1 2 93330 45065
0 45067 5 1 1 45066
0 45068 7 1 2 81774 90847
0 45069 5 1 1 45068
0 45070 7 1 2 86444 45069
0 45071 5 1 1 45070
0 45072 7 1 2 75558 45071
0 45073 5 1 1 45072
0 45074 7 1 2 70225 80792
0 45075 7 1 2 94890 45074
0 45076 5 1 1 45075
0 45077 7 1 2 45073 45076
0 45078 7 1 2 45067 45077
0 45079 7 1 2 45051 45078
0 45080 7 1 2 45039 45079
0 45081 5 1 1 45080
0 45082 7 1 2 90261 45081
0 45083 5 1 1 45082
0 45084 7 1 2 93858 94469
0 45085 5 1 1 45084
0 45086 7 1 2 81974 82301
0 45087 7 1 2 94695 45086
0 45088 5 1 1 45087
0 45089 7 1 2 45085 45088
0 45090 5 1 1 45089
0 45091 7 1 2 76463 45090
0 45092 5 1 1 45091
0 45093 7 1 2 64618 95041
0 45094 5 1 1 45093
0 45095 7 1 2 76226 85884
0 45096 5 1 1 45095
0 45097 7 1 2 93388 45096
0 45098 5 1 1 45097
0 45099 7 1 2 94182 45098
0 45100 5 1 1 45099
0 45101 7 1 2 78883 90015
0 45102 7 1 2 94802 45101
0 45103 5 1 1 45102
0 45104 7 1 2 84996 73700
0 45105 5 1 1 45104
0 45106 7 1 2 59913 45105
0 45107 7 1 2 45103 45106
0 45108 7 1 2 45100 45107
0 45109 5 1 1 45108
0 45110 7 1 2 61071 45109
0 45111 7 1 2 45094 45110
0 45112 5 1 1 45111
0 45113 7 1 2 85700 78598
0 45114 5 1 1 45113
0 45115 7 1 2 61439 84085
0 45116 5 1 1 45115
0 45117 7 1 2 45114 45116
0 45118 5 1 1 45117
0 45119 7 1 2 67792 45118
0 45120 5 1 1 45119
0 45121 7 2 2 73581 78990
0 45122 5 1 1 95078
0 45123 7 1 2 88818 95079
0 45124 5 1 1 45123
0 45125 7 1 2 81952 45124
0 45126 5 1 1 45125
0 45127 7 1 2 68409 90010
0 45128 5 1 1 45127
0 45129 7 1 2 68441 45122
0 45130 7 1 2 45128 45129
0 45131 5 1 1 45130
0 45132 7 1 2 85668 45131
0 45133 7 1 2 45126 45132
0 45134 7 1 2 45120 45133
0 45135 5 1 1 45134
0 45136 7 1 2 59914 45135
0 45137 5 1 1 45136
0 45138 7 1 2 77235 72913
0 45139 5 1 1 45138
0 45140 7 1 2 29903 94330
0 45141 5 1 1 45140
0 45142 7 1 2 73565 45141
0 45143 5 1 1 45142
0 45144 7 1 2 59163 78942
0 45145 5 1 1 45144
0 45146 7 1 2 42919 45145
0 45147 5 1 1 45146
0 45148 7 1 2 64619 45147
0 45149 5 1 1 45148
0 45150 7 1 2 45143 45149
0 45151 5 1 1 45150
0 45152 7 1 2 65697 45151
0 45153 5 1 1 45152
0 45154 7 1 2 45139 45153
0 45155 7 1 2 45137 45154
0 45156 5 1 1 45155
0 45157 7 1 2 63400 45156
0 45158 5 1 1 45157
0 45159 7 2 2 75582 85619
0 45160 7 1 2 73701 95080
0 45161 5 1 1 45160
0 45162 7 1 2 76227 90409
0 45163 5 1 1 45162
0 45164 7 1 2 45161 45163
0 45165 5 1 1 45164
0 45166 7 1 2 78599 45165
0 45167 5 1 1 45166
0 45168 7 1 2 85428 84614
0 45169 5 1 1 45168
0 45170 7 1 2 90651 45169
0 45171 5 1 1 45170
0 45172 7 1 2 86239 45171
0 45173 5 1 1 45172
0 45174 7 1 2 61440 90087
0 45175 5 1 1 45174
0 45176 7 1 2 90584 45175
0 45177 5 1 1 45176
0 45178 7 1 2 71330 45177
0 45179 5 1 1 45178
0 45180 7 1 2 23527 45179
0 45181 7 1 2 45173 45180
0 45182 5 1 1 45181
0 45183 7 1 2 68530 45182
0 45184 5 1 1 45183
0 45185 7 1 2 45167 45184
0 45186 5 1 1 45185
0 45187 7 1 2 67793 45186
0 45188 5 1 1 45187
0 45189 7 2 2 70375 85352
0 45190 5 1 1 95082
0 45191 7 1 2 59915 95083
0 45192 5 2 1 45191
0 45193 7 1 2 77832 95084
0 45194 5 1 1 45193
0 45195 7 1 2 81953 45194
0 45196 5 1 1 45195
0 45197 7 1 2 58641 93237
0 45198 5 1 1 45197
0 45199 7 1 2 68266 95081
0 45200 5 1 1 45199
0 45201 7 1 2 45198 45200
0 45202 7 1 2 45196 45201
0 45203 5 1 1 45202
0 45204 7 1 2 73702 45203
0 45205 5 1 1 45204
0 45206 7 1 2 81954 93043
0 45207 5 1 1 45206
0 45208 7 1 2 93399 45207
0 45209 5 1 1 45208
0 45210 7 1 2 90410 45209
0 45211 5 1 1 45210
0 45212 7 1 2 45205 45211
0 45213 7 1 2 45188 45212
0 45214 7 1 2 45158 45213
0 45215 7 1 2 45112 45214
0 45216 5 1 1 45215
0 45217 7 1 2 60046 45216
0 45218 5 1 1 45217
0 45219 7 1 2 45092 45218
0 45220 5 1 1 45219
0 45221 7 1 2 61702 45220
0 45222 5 1 1 45221
0 45223 7 1 2 45083 45222
0 45224 5 1 1 45223
0 45225 7 1 2 58792 45224
0 45226 5 1 1 45225
0 45227 7 2 2 84151 86319
0 45228 7 1 2 82544 94993
0 45229 7 1 2 95086 45228
0 45230 7 1 2 83108 45229
0 45231 5 1 1 45230
0 45232 7 1 2 64833 45231
0 45233 7 1 2 45226 45232
0 45234 5 1 1 45233
0 45235 7 1 2 91372 92541
0 45236 5 1 1 45235
0 45237 7 1 2 74027 86090
0 45238 7 1 2 92526 45237
0 45239 5 1 1 45238
0 45240 7 1 2 45236 45239
0 45241 5 1 1 45240
0 45242 7 1 2 88776 45241
0 45243 5 1 1 45242
0 45244 7 2 2 61072 87349
0 45245 7 1 2 92751 95088
0 45246 5 1 1 45245
0 45247 7 1 2 45243 45246
0 45248 5 1 1 45247
0 45249 7 1 2 84891 45248
0 45250 5 1 1 45249
0 45251 7 1 2 60155 45250
0 45252 5 1 1 45251
0 45253 7 1 2 61967 45252
0 45254 7 1 2 45234 45253
0 45255 5 1 1 45254
0 45256 7 1 2 44990 45255
0 45257 7 1 2 44926 45256
0 45258 5 1 1 45257
0 45259 7 1 2 66720 45258
0 45260 5 1 1 45259
0 45261 7 1 2 61073 41798
0 45262 5 1 1 45261
0 45263 7 1 2 58642 45262
0 45264 5 1 1 45263
0 45265 7 1 2 59651 45264
0 45266 5 1 1 45265
0 45267 7 2 2 81373 82454
0 45268 5 1 1 95090
0 45269 7 1 2 65698 95091
0 45270 5 1 1 45269
0 45271 7 1 2 64401 43909
0 45272 7 1 2 45270 45271
0 45273 5 1 1 45272
0 45274 7 1 2 45266 45273
0 45275 5 1 1 45274
0 45276 7 1 2 64620 45275
0 45277 5 1 1 45276
0 45278 7 1 2 63093 94647
0 45279 5 1 1 45278
0 45280 7 1 2 93468 95077
0 45281 5 1 1 45280
0 45282 7 1 2 62266 45281
0 45283 5 1 1 45282
0 45284 7 1 2 75895 87086
0 45285 5 1 1 45284
0 45286 7 1 2 78217 45285
0 45287 5 1 1 45286
0 45288 7 1 2 72247 45287
0 45289 5 1 1 45288
0 45290 7 1 2 63094 45289
0 45291 5 1 1 45290
0 45292 7 1 2 45283 45291
0 45293 5 1 1 45292
0 45294 7 1 2 62795 45293
0 45295 5 1 1 45294
0 45296 7 1 2 45279 45295
0 45297 5 1 1 45296
0 45298 7 1 2 64402 45297
0 45299 5 1 1 45298
0 45300 7 1 2 64403 45268
0 45301 5 1 1 45300
0 45302 7 1 2 63095 92779
0 45303 5 1 1 45302
0 45304 7 1 2 59916 45303
0 45305 7 1 2 45301 45304
0 45306 7 1 2 92772 45305
0 45307 5 1 1 45306
0 45308 7 1 2 63401 45307
0 45309 5 1 1 45308
0 45310 7 1 2 63402 92758
0 45311 5 1 1 45310
0 45312 7 1 2 58343 45311
0 45313 5 1 1 45312
0 45314 7 1 2 58643 94896
0 45315 5 1 1 45314
0 45316 7 1 2 62267 45315
0 45317 7 1 2 45313 45316
0 45318 5 1 1 45317
0 45319 7 1 2 45309 45318
0 45320 7 1 2 45299 45319
0 45321 5 1 1 45320
0 45322 7 1 2 65699 45321
0 45323 5 1 1 45322
0 45324 7 1 2 45277 45323
0 45325 5 1 1 45324
0 45326 7 1 2 88274 45325
0 45327 5 1 1 45326
0 45328 7 1 2 68168 93158
0 45329 5 1 1 45328
0 45330 7 1 2 67224 93165
0 45331 5 1 1 45330
0 45332 7 1 2 45329 45331
0 45333 5 1 1 45332
0 45334 7 1 2 82532 89865
0 45335 7 1 2 45333 45334
0 45336 5 1 1 45335
0 45337 7 1 2 45327 45336
0 45338 5 1 1 45337
0 45339 7 1 2 66046 45338
0 45340 5 1 1 45339
0 45341 7 1 2 85701 94159
0 45342 5 1 1 45341
0 45343 7 1 2 71331 82087
0 45344 5 1 1 45343
0 45345 7 1 2 62268 93521
0 45346 5 1 1 45345
0 45347 7 1 2 45344 45346
0 45348 5 1 1 45347
0 45349 7 1 2 68169 45348
0 45350 5 1 1 45349
0 45351 7 1 2 85479 45350
0 45352 7 1 2 45342 45351
0 45353 5 1 1 45352
0 45354 7 1 2 64621 45353
0 45355 5 1 1 45354
0 45356 7 1 2 3588 95073
0 45357 5 1 1 45356
0 45358 7 1 2 94594 45357
0 45359 5 1 1 45358
0 45360 7 1 2 93658 94606
0 45361 5 1 1 45360
0 45362 7 1 2 82966 45361
0 45363 5 1 1 45362
0 45364 7 1 2 75914 67606
0 45365 7 1 2 45363 45364
0 45366 5 1 1 45365
0 45367 7 1 2 14002 45366
0 45368 7 1 2 45359 45367
0 45369 7 1 2 45355 45368
0 45370 5 1 1 45369
0 45371 7 1 2 66345 45370
0 45372 5 1 1 45371
0 45373 7 2 2 59917 90662
0 45374 5 1 1 95092
0 45375 7 1 2 62269 95028
0 45376 5 1 1 45375
0 45377 7 1 2 45374 45376
0 45378 5 1 1 45377
0 45379 7 1 2 78300 45378
0 45380 5 1 1 45379
0 45381 7 1 2 90133 93273
0 45382 5 2 1 45381
0 45383 7 1 2 45380 95094
0 45384 5 1 1 45383
0 45385 7 1 2 70844 45384
0 45386 5 1 1 45385
0 45387 7 2 2 73220 92655
0 45388 7 1 2 63403 95096
0 45389 5 1 1 45388
0 45390 7 4 2 62270 82575
0 45391 5 3 1 95098
0 45392 7 1 2 84351 95099
0 45393 5 1 1 45392
0 45394 7 1 2 45389 45393
0 45395 5 1 1 45394
0 45396 7 1 2 85702 45395
0 45397 5 1 1 45396
0 45398 7 1 2 79195 95097
0 45399 5 1 1 45398
0 45400 7 1 2 71834 82576
0 45401 7 1 2 93170 45400
0 45402 5 1 1 45401
0 45403 7 1 2 95095 45402
0 45404 7 1 2 45399 45403
0 45405 7 1 2 45397 45404
0 45406 5 1 1 45405
0 45407 7 1 2 69067 45406
0 45408 5 1 1 45407
0 45409 7 1 2 58344 94608
0 45410 5 1 1 45409
0 45411 7 1 2 75915 45410
0 45412 5 1 1 45411
0 45413 7 1 2 59652 81854
0 45414 5 1 1 45413
0 45415 7 1 2 78202 45414
0 45416 5 1 1 45415
0 45417 7 1 2 85136 45416
0 45418 7 1 2 45412 45417
0 45419 5 1 1 45418
0 45420 7 1 2 82577 45419
0 45421 5 1 1 45420
0 45422 7 1 2 45408 45421
0 45423 7 1 2 45386 45422
0 45424 7 1 2 45372 45423
0 45425 5 1 1 45424
0 45426 7 1 2 58793 45425
0 45427 5 1 1 45426
0 45428 7 1 2 75676 94655
0 45429 5 1 1 45428
0 45430 7 1 2 2217 45429
0 45431 5 1 1 45430
0 45432 7 1 2 59653 45431
0 45433 5 1 1 45432
0 45434 7 1 2 27651 45433
0 45435 5 1 1 45434
0 45436 7 1 2 87267 45435
0 45437 5 1 1 45436
0 45438 7 1 2 45427 45437
0 45439 5 1 1 45438
0 45440 7 1 2 61074 45439
0 45441 5 1 1 45440
0 45442 7 1 2 68201 95093
0 45443 5 1 1 45442
0 45444 7 1 2 90134 93264
0 45445 5 1 1 45444
0 45446 7 1 2 45443 45445
0 45447 5 1 1 45446
0 45448 7 1 2 62521 45447
0 45449 5 1 1 45448
0 45450 7 2 2 63919 76703
0 45451 7 2 2 66346 95105
0 45452 5 1 1 95107
0 45453 7 1 2 95102 45452
0 45454 5 1 1 45453
0 45455 7 1 2 82851 45454
0 45456 5 1 1 45455
0 45457 7 1 2 45449 45456
0 45458 5 1 1 45457
0 45459 7 1 2 69068 45458
0 45460 5 1 1 45459
0 45461 7 1 2 62271 90593
0 45462 5 1 1 45461
0 45463 7 1 2 82598 45462
0 45464 5 3 1 45463
0 45465 7 1 2 94109 95109
0 45466 5 1 1 45465
0 45467 7 1 2 77594 95056
0 45468 5 1 1 45467
0 45469 7 1 2 45466 45468
0 45470 5 1 1 45469
0 45471 7 1 2 71697 45470
0 45472 5 1 1 45471
0 45473 7 1 2 76704 88813
0 45474 5 1 1 45473
0 45475 7 1 2 85080 16522
0 45476 7 1 2 45474 45475
0 45477 5 1 1 45476
0 45478 7 1 2 90135 45477
0 45479 5 1 1 45478
0 45480 7 1 2 45472 45479
0 45481 7 1 2 45460 45480
0 45482 5 1 1 45481
0 45483 7 1 2 60666 45482
0 45484 5 1 1 45483
0 45485 7 1 2 75191 88814
0 45486 5 1 1 45485
0 45487 7 1 2 93810 45486
0 45488 5 1 1 45487
0 45489 7 1 2 82884 45488
0 45490 5 1 1 45489
0 45491 7 1 2 92933 95100
0 45492 5 1 1 45491
0 45493 7 1 2 45490 45492
0 45494 5 1 1 45493
0 45495 7 1 2 71332 45494
0 45496 5 1 1 45495
0 45497 7 1 2 75175 86148
0 45498 5 1 1 45497
0 45499 7 1 2 93247 45498
0 45500 5 1 1 45499
0 45501 7 1 2 71452 94306
0 45502 5 1 1 45501
0 45503 7 1 2 59654 74345
0 45504 5 1 1 45503
0 45505 7 1 2 63404 45504
0 45506 5 1 1 45505
0 45507 7 1 2 45502 45506
0 45508 7 1 2 45500 45507
0 45509 5 1 1 45508
0 45510 7 1 2 87342 45509
0 45511 5 1 1 45510
0 45512 7 1 2 85024 92675
0 45513 5 1 1 45512
0 45514 7 1 2 88615 45513
0 45515 5 1 1 45514
0 45516 7 1 2 64404 45515
0 45517 5 1 1 45516
0 45518 7 1 2 65700 87352
0 45519 5 1 1 45518
0 45520 7 1 2 88620 45519
0 45521 5 1 1 45520
0 45522 7 1 2 93548 45521
0 45523 5 1 1 45522
0 45524 7 2 2 67794 95110
0 45525 7 1 2 82852 80522
0 45526 7 1 2 95112 45525
0 45527 5 1 1 45526
0 45528 7 1 2 45523 45527
0 45529 7 1 2 45517 45528
0 45530 7 1 2 45511 45529
0 45531 7 1 2 45496 45530
0 45532 7 1 2 45484 45531
0 45533 5 1 1 45532
0 45534 7 1 2 58794 45533
0 45535 5 1 1 45534
0 45536 7 1 2 45441 45535
0 45537 5 1 1 45536
0 45538 7 1 2 61441 45537
0 45539 5 1 1 45538
0 45540 7 1 2 58644 95048
0 45541 5 1 1 45540
0 45542 7 1 2 82578 45541
0 45543 5 1 1 45542
0 45544 7 1 2 60667 87394
0 45545 5 1 1 45544
0 45546 7 1 2 16065 45545
0 45547 5 1 1 45546
0 45548 7 1 2 63920 45547
0 45549 5 1 1 45548
0 45550 7 1 2 41987 45549
0 45551 5 1 1 45550
0 45552 7 1 2 62522 45551
0 45553 5 1 1 45552
0 45554 7 1 2 78248 77534
0 45555 5 1 1 45554
0 45556 7 1 2 45553 45555
0 45557 5 1 1 45556
0 45558 7 1 2 62796 45557
0 45559 5 1 1 45558
0 45560 7 1 2 75583 95044
0 45561 7 1 2 45559 45560
0 45562 5 1 1 45561
0 45563 7 1 2 90594 45562
0 45564 5 1 1 45563
0 45565 7 1 2 45543 45564
0 45566 5 1 1 45565
0 45567 7 1 2 61075 45566
0 45568 5 1 1 45567
0 45569 7 2 2 70788 78849
0 45570 5 2 1 95114
0 45571 7 1 2 69204 95115
0 45572 5 1 1 45571
0 45573 7 1 2 88561 45572
0 45574 5 1 1 45573
0 45575 7 1 2 45568 45574
0 45576 5 1 1 45575
0 45577 7 1 2 71333 45576
0 45578 5 1 1 45577
0 45579 7 1 2 82215 94778
0 45580 5 1 1 45579
0 45581 7 1 2 87343 43897
0 45582 5 1 1 45581
0 45583 7 1 2 82579 83938
0 45584 5 1 1 45583
0 45585 7 1 2 69069 91470
0 45586 5 1 1 45585
0 45587 7 1 2 31255 95103
0 45588 7 1 2 45586 45587
0 45589 5 1 1 45588
0 45590 7 1 2 68442 45589
0 45591 5 1 1 45590
0 45592 7 1 2 45584 45591
0 45593 7 1 2 45582 45592
0 45594 5 1 1 45593
0 45595 7 1 2 61076 45594
0 45596 5 1 1 45595
0 45597 7 1 2 45580 45596
0 45598 5 1 1 45597
0 45599 7 1 2 85183 45598
0 45600 5 1 1 45599
0 45601 7 1 2 84133 25570
0 45602 5 1 1 45601
0 45603 7 1 2 63405 45602
0 45604 5 1 1 45603
0 45605 7 1 2 18455 45604
0 45606 5 1 1 45605
0 45607 7 1 2 64622 45606
0 45608 5 1 1 45607
0 45609 7 1 2 61077 94677
0 45610 5 1 1 45609
0 45611 7 1 2 68170 92478
0 45612 5 1 1 45611
0 45613 7 2 2 70308 75192
0 45614 5 1 1 95118
0 45615 7 1 2 45612 45614
0 45616 5 1 1 45615
0 45617 7 1 2 67795 45616
0 45618 5 1 1 45617
0 45619 7 3 2 85353 84550
0 45620 5 1 1 95120
0 45621 7 1 2 45618 45620
0 45622 7 1 2 45610 45621
0 45623 5 1 1 45622
0 45624 7 1 2 87805 45623
0 45625 5 1 1 45624
0 45626 7 1 2 45608 45625
0 45627 7 1 2 45600 45626
0 45628 7 1 2 45578 45627
0 45629 5 1 1 45628
0 45630 7 1 2 58795 45629
0 45631 5 1 1 45630
0 45632 7 1 2 45539 45631
0 45633 7 1 2 45340 45632
0 45634 5 1 1 45633
0 45635 7 1 2 60047 45634
0 45636 5 1 1 45635
0 45637 7 1 2 83166 94954
0 45638 5 1 1 45637
0 45639 7 1 2 58796 87627
0 45640 5 1 1 45639
0 45641 7 1 2 45638 45640
0 45642 5 1 1 45641
0 45643 7 1 2 74544 45642
0 45644 5 1 1 45643
0 45645 7 1 2 79170 87769
0 45646 7 1 2 82817 45645
0 45647 5 1 1 45646
0 45648 7 1 2 45644 45647
0 45649 5 1 1 45648
0 45650 7 1 2 68636 45649
0 45651 5 1 1 45650
0 45652 7 1 2 59655 78689
0 45653 5 1 1 45652
0 45654 7 1 2 65701 83758
0 45655 5 1 1 45654
0 45656 7 1 2 45653 45655
0 45657 5 1 1 45656
0 45658 7 1 2 87628 94656
0 45659 7 1 2 45657 45658
0 45660 5 1 1 45659
0 45661 7 1 2 74550 43849
0 45662 5 1 1 45661
0 45663 7 1 2 87640 76866
0 45664 7 1 2 94520 45663
0 45665 7 1 2 45662 45664
0 45666 5 1 1 45665
0 45667 7 1 2 45660 45666
0 45668 7 1 2 45651 45667
0 45669 5 1 1 45668
0 45670 7 1 2 61442 45669
0 45671 5 1 1 45670
0 45672 7 1 2 76464 73433
0 45673 5 1 1 45672
0 45674 7 1 2 64405 45673
0 45675 5 1 1 45674
0 45676 7 1 2 92731 94782
0 45677 7 1 2 45675 45676
0 45678 5 1 1 45677
0 45679 7 1 2 45671 45678
0 45680 5 1 1 45679
0 45681 7 1 2 57777 45680
0 45682 5 1 1 45681
0 45683 7 1 2 64406 88254
0 45684 5 1 1 45683
0 45685 7 2 2 74176 90297
0 45686 7 2 2 72035 87239
0 45687 7 2 2 58645 69120
0 45688 7 1 2 95125 95127
0 45689 7 1 2 95123 45688
0 45690 5 1 1 45689
0 45691 7 1 2 45684 45690
0 45692 5 1 1 45691
0 45693 7 1 2 64623 45692
0 45694 5 1 1 45693
0 45695 7 1 2 78653 94285
0 45696 5 1 1 45695
0 45697 7 1 2 74135 90351
0 45698 7 1 2 77725 45697
0 45699 5 1 1 45698
0 45700 7 1 2 45696 45699
0 45701 5 1 1 45700
0 45702 7 1 2 59164 45701
0 45703 5 1 1 45702
0 45704 7 1 2 37542 94286
0 45705 5 1 1 45704
0 45706 7 1 2 45703 45705
0 45707 5 1 1 45706
0 45708 7 1 2 79829 45707
0 45709 5 1 1 45708
0 45710 7 1 2 87552 94950
0 45711 5 1 1 45710
0 45712 7 1 2 45709 45711
0 45713 5 1 1 45712
0 45714 7 1 2 94057 45713
0 45715 5 1 1 45714
0 45716 7 1 2 45694 45715
0 45717 5 1 1 45716
0 45718 7 1 2 78991 45717
0 45719 5 1 1 45718
0 45720 7 2 2 81406 73502
0 45721 5 1 1 95129
0 45722 7 1 2 88277 45721
0 45723 5 1 1 45722
0 45724 7 1 2 82634 73761
0 45725 7 1 2 95087 45724
0 45726 7 1 2 45723 45725
0 45727 5 1 1 45726
0 45728 7 1 2 66619 45727
0 45729 7 1 2 45719 45728
0 45730 7 1 2 45682 45729
0 45731 7 1 2 45636 45730
0 45732 5 1 1 45731
0 45733 7 1 2 61443 94751
0 45734 5 1 1 45733
0 45735 7 1 2 84250 45734
0 45736 5 1 1 45735
0 45737 7 1 2 1293 45736
0 45738 5 1 1 45737
0 45739 7 1 2 82414 45738
0 45740 5 1 1 45739
0 45741 7 1 2 79617 74073
0 45742 5 1 1 45741
0 45743 7 1 2 43259 45742
0 45744 5 1 1 45743
0 45745 7 1 2 59918 45744
0 45746 5 1 1 45745
0 45747 7 2 2 66347 78850
0 45748 5 1 1 95131
0 45749 7 1 2 59919 76508
0 45750 5 1 1 45749
0 45751 7 1 2 45748 45750
0 45752 5 1 1 45751
0 45753 7 1 2 65702 45752
0 45754 5 1 1 45753
0 45755 7 1 2 87276 93823
0 45756 5 1 1 45755
0 45757 7 1 2 45754 45756
0 45758 5 1 1 45757
0 45759 7 1 2 94035 45758
0 45760 5 1 1 45759
0 45761 7 1 2 45746 45760
0 45762 5 1 1 45761
0 45763 7 1 2 59656 45762
0 45764 5 1 1 45763
0 45765 7 1 2 45740 45764
0 45766 5 1 1 45765
0 45767 7 1 2 94870 45766
0 45768 5 1 1 45767
0 45769 7 1 2 61968 45768
0 45770 5 1 1 45769
0 45771 7 1 2 60156 45770
0 45772 7 1 2 45732 45771
0 45773 5 1 1 45772
0 45774 7 1 2 66348 75176
0 45775 5 1 1 45774
0 45776 7 1 2 28154 45775
0 45777 5 1 1 45776
0 45778 7 1 2 85255 45777
0 45779 5 1 1 45778
0 45780 7 1 2 82415 92460
0 45781 5 1 1 45780
0 45782 7 1 2 45779 45781
0 45783 5 1 1 45782
0 45784 7 1 2 57778 45783
0 45785 5 1 1 45784
0 45786 7 1 2 82416 43820
0 45787 5 1 1 45786
0 45788 7 1 2 45785 45787
0 45789 5 1 1 45788
0 45790 7 1 2 66047 45789
0 45791 5 1 1 45790
0 45792 7 1 2 68410 94239
0 45793 7 1 2 42670 45792
0 45794 5 1 1 45793
0 45795 7 1 2 45791 45794
0 45796 5 1 1 45795
0 45797 7 1 2 66982 94871
0 45798 7 1 2 45796 45797
0 45799 5 1 1 45798
0 45800 7 1 2 45773 45799
0 45801 5 1 1 45800
0 45802 7 1 2 62114 45801
0 45803 5 1 1 45802
0 45804 7 1 2 85867 79600
0 45805 5 1 1 45804
0 45806 7 1 2 93029 45805
0 45807 5 1 1 45806
0 45808 7 1 2 61078 45807
0 45809 5 1 1 45808
0 45810 7 1 2 62797 13056
0 45811 5 1 1 45810
0 45812 7 1 2 37293 45811
0 45813 7 1 2 94152 45812
0 45814 5 1 1 45813
0 45815 7 1 2 58646 45814
0 45816 5 1 1 45815
0 45817 7 1 2 45809 45816
0 45818 5 1 1 45817
0 45819 7 1 2 71077 45818
0 45820 5 1 1 45819
0 45821 7 1 2 65703 76824
0 45822 7 1 2 94761 45821
0 45823 5 1 1 45822
0 45824 7 1 2 57484 18942
0 45825 5 1 1 45824
0 45826 7 1 2 80599 81804
0 45827 7 1 2 45825 45826
0 45828 5 1 1 45827
0 45829 7 1 2 45823 45828
0 45830 5 1 1 45829
0 45831 7 1 2 66048 45830
0 45832 5 1 1 45831
0 45833 7 1 2 72483 86152
0 45834 5 1 1 45833
0 45835 7 1 2 85984 45834
0 45836 5 1 1 45835
0 45837 7 1 2 82018 45836
0 45838 7 1 2 45832 45837
0 45839 5 1 1 45838
0 45840 7 2 2 67530 88981
0 45841 5 1 1 95133
0 45842 7 1 2 68171 95134
0 45843 5 1 1 45842
0 45844 7 1 2 87041 82019
0 45845 5 1 1 45844
0 45846 7 1 2 45843 45845
0 45847 5 1 1 45846
0 45848 7 1 2 72495 45847
0 45849 5 1 1 45848
0 45850 7 1 2 80545 82020
0 45851 5 1 1 45850
0 45852 7 1 2 45841 45851
0 45853 5 1 1 45852
0 45854 7 1 2 63096 45853
0 45855 5 1 1 45854
0 45856 7 1 2 45849 45855
0 45857 7 1 2 45839 45856
0 45858 7 1 2 45820 45857
0 45859 5 1 1 45858
0 45860 7 1 2 82417 45859
0 45861 5 1 1 45860
0 45862 7 2 2 64624 88925
0 45863 7 1 2 60157 80676
0 45864 7 2 2 91533 45863
0 45865 5 1 1 95137
0 45866 7 1 2 63097 95138
0 45867 5 1 1 45866
0 45868 7 4 2 64105 66983
0 45869 5 1 1 95139
0 45870 7 1 2 67085 45869
0 45871 5 2 1 45870
0 45872 7 1 2 63098 95143
0 45873 5 2 1 45872
0 45874 7 1 2 67063 90933
0 45875 5 1 1 45874
0 45876 7 1 2 95145 45875
0 45877 5 1 1 45876
0 45878 7 1 2 60413 45877
0 45879 5 1 1 45878
0 45880 7 1 2 61079 86532
0 45881 5 1 1 45880
0 45882 7 1 2 45879 45881
0 45883 5 1 1 45882
0 45884 7 1 2 71835 45883
0 45885 5 1 1 45884
0 45886 7 1 2 76270 79000
0 45887 7 5 2 90934 45886
0 45888 7 1 2 66984 95147
0 45889 5 1 1 45888
0 45890 7 1 2 45885 45889
0 45891 5 1 1 45890
0 45892 7 1 2 62798 45891
0 45893 5 1 1 45892
0 45894 7 1 2 84765 92172
0 45895 5 1 1 45894
0 45896 7 1 2 95148 45895
0 45897 5 1 1 45896
0 45898 7 1 2 45893 45897
0 45899 5 1 1 45898
0 45900 7 1 2 62523 45899
0 45901 5 1 1 45900
0 45902 7 2 2 62799 66985
0 45903 5 1 1 95152
0 45904 7 1 2 92173 45903
0 45905 5 2 1 45904
0 45906 7 1 2 70845 95154
0 45907 7 1 2 95149 45906
0 45908 5 1 1 45907
0 45909 7 1 2 45901 45908
0 45910 5 1 1 45909
0 45911 7 1 2 68884 45910
0 45912 5 1 1 45911
0 45913 7 2 2 3180 88880
0 45914 7 1 2 62524 95156
0 45915 5 1 1 45914
0 45916 7 1 2 86519 45915
0 45917 5 1 1 45916
0 45918 7 1 2 62800 45917
0 45919 5 1 1 45918
0 45920 7 1 2 60414 86533
0 45921 5 1 1 45920
0 45922 7 1 2 45919 45921
0 45923 5 1 1 45922
0 45924 7 1 2 72554 45923
0 45925 5 1 1 45924
0 45926 7 2 2 66620 72108
0 45927 7 2 2 68531 95158
0 45928 5 1 1 95160
0 45929 7 1 2 60668 95161
0 45930 5 1 1 45929
0 45931 7 1 2 86520 45930
0 45932 5 1 1 45931
0 45933 7 1 2 62525 45932
0 45934 5 1 1 45933
0 45935 7 1 2 76899 95157
0 45936 5 1 1 45935
0 45937 7 1 2 86534 45936
0 45938 7 1 2 45934 45937
0 45939 5 1 1 45938
0 45940 7 1 2 62801 45939
0 45941 5 1 1 45940
0 45942 7 2 2 68532 67064
0 45943 5 1 1 95162
0 45944 7 1 2 60669 95163
0 45945 5 1 1 45944
0 45946 7 1 2 86535 45945
0 45947 5 1 1 45946
0 45948 7 1 2 68267 45947
0 45949 5 1 1 45948
0 45950 7 1 2 86536 31995
0 45951 5 1 1 45950
0 45952 7 1 2 84352 45951
0 45953 5 1 1 45952
0 45954 7 1 2 70952 95155
0 45955 5 1 1 45954
0 45956 7 1 2 45953 45955
0 45957 5 1 1 45956
0 45958 7 1 2 68885 45957
0 45959 5 1 1 45958
0 45960 7 1 2 45949 45959
0 45961 7 1 2 45941 45960
0 45962 7 1 2 45925 45961
0 45963 5 1 1 45962
0 45964 7 1 2 61444 45963
0 45965 5 1 1 45964
0 45966 7 1 2 62802 93147
0 45967 5 1 1 45966
0 45968 7 1 2 66049 45967
0 45969 7 1 2 93328 45968
0 45970 5 1 1 45969
0 45971 7 1 2 61969 84114
0 45972 7 1 2 45970 45971
0 45973 5 1 1 45972
0 45974 7 1 2 45965 45973
0 45975 5 1 1 45974
0 45976 7 1 2 70226 45975
0 45977 5 1 1 45976
0 45978 7 1 2 67086 20301
0 45979 5 3 1 45978
0 45980 7 1 2 70907 95164
0 45981 5 1 1 45980
0 45982 7 1 2 71836 89470
0 45983 5 1 1 45982
0 45984 7 1 2 45981 45983
0 45985 5 1 1 45984
0 45986 7 1 2 68533 45985
0 45987 5 1 1 45986
0 45988 7 1 2 77542 95150
0 45989 5 1 1 45988
0 45990 7 1 2 85258 70908
0 45991 5 1 1 45990
0 45992 7 1 2 45989 45991
0 45993 5 1 1 45992
0 45994 7 1 2 66986 45993
0 45995 5 1 1 45994
0 45996 7 1 2 45987 45995
0 45997 5 1 1 45996
0 45998 7 1 2 62803 45997
0 45999 5 1 1 45998
0 46000 7 2 2 81029 68710
0 46001 5 1 1 95167
0 46002 7 1 2 60415 91777
0 46003 5 1 1 46002
0 46004 7 1 2 46001 46003
0 46005 5 1 1 46004
0 46006 7 1 2 64106 46005
0 46007 5 1 1 46006
0 46008 7 2 2 64834 93965
0 46009 7 1 2 60670 95169
0 46010 5 1 1 46009
0 46011 7 1 2 46007 46010
0 46012 5 1 1 46011
0 46013 7 1 2 63099 46012
0 46014 5 1 1 46013
0 46015 7 1 2 45999 46014
0 46016 5 1 1 46015
0 46017 7 1 2 62526 46016
0 46018 5 1 1 46017
0 46019 7 2 2 64107 67065
0 46020 5 1 1 95171
0 46021 7 1 2 27414 46020
0 46022 5 1 1 46021
0 46023 7 1 2 60671 46022
0 46024 5 1 1 46023
0 46025 7 1 2 83463 95165
0 46026 5 1 1 46025
0 46027 7 1 2 46024 46026
0 46028 5 1 1 46027
0 46029 7 1 2 61080 46028
0 46030 5 1 1 46029
0 46031 7 1 2 75403 91778
0 46032 5 1 1 46031
0 46033 7 1 2 46030 46032
0 46034 5 1 1 46033
0 46035 7 1 2 63921 46034
0 46036 5 1 1 46035
0 46037 7 1 2 80437 95140
0 46038 5 1 1 46037
0 46039 7 1 2 46036 46038
0 46040 5 1 1 46039
0 46041 7 1 2 63100 46040
0 46042 5 1 1 46041
0 46043 7 1 2 61081 95172
0 46044 5 1 1 46043
0 46045 7 1 2 95146 46044
0 46046 5 1 1 46045
0 46047 7 1 2 60672 46046
0 46048 5 1 1 46047
0 46049 7 1 2 66621 86527
0 46050 5 1 1 46049
0 46051 7 1 2 46048 46050
0 46052 5 1 1 46051
0 46053 7 1 2 86248 78465
0 46054 5 1 1 46053
0 46055 7 1 2 46052 46054
0 46056 5 1 1 46055
0 46057 7 1 2 70039 95166
0 46058 5 1 1 46057
0 46059 7 1 2 70024 95159
0 46060 5 1 1 46059
0 46061 7 1 2 46058 46060
0 46062 5 1 1 46061
0 46063 7 1 2 62527 46062
0 46064 5 1 1 46063
0 46065 7 1 2 60416 95153
0 46066 5 1 1 46065
0 46067 7 1 2 45943 46066
0 46068 5 1 1 46067
0 46069 7 1 2 70846 46068
0 46070 5 1 1 46069
0 46071 7 1 2 76509 84561
0 46072 5 1 1 46071
0 46073 7 1 2 74876 66987
0 46074 7 1 2 46072 46073
0 46075 5 1 1 46074
0 46076 7 1 2 31993 46075
0 46077 7 1 2 46070 46076
0 46078 7 1 2 46064 46077
0 46079 5 1 1 46078
0 46080 7 1 2 95151 46079
0 46081 5 1 1 46080
0 46082 7 1 2 46056 46081
0 46083 7 1 2 46042 46082
0 46084 7 1 2 46018 46083
0 46085 7 1 2 45977 46084
0 46086 7 1 2 45912 46085
0 46087 5 1 1 46086
0 46088 7 1 2 63406 46087
0 46089 5 1 1 46088
0 46090 7 1 2 45867 46089
0 46091 5 1 1 46090
0 46092 7 1 2 95135 46091
0 46093 5 1 1 46092
0 46094 7 1 2 45861 46093
0 46095 5 1 1 46094
0 46096 7 1 2 64407 46095
0 46097 5 1 1 46096
0 46098 7 1 2 16977 67066
0 46099 5 1 1 46098
0 46100 7 1 2 57779 46099
0 46101 5 1 1 46100
0 46102 7 1 2 67087 45928
0 46103 5 1 1 46102
0 46104 7 1 2 70847 46103
0 46105 7 1 2 46101 46104
0 46106 5 1 1 46105
0 46107 7 1 2 85928 84763
0 46108 5 1 1 46107
0 46109 7 1 2 62528 67067
0 46110 7 1 2 80278 46109
0 46111 5 1 1 46110
0 46112 7 1 2 46108 46111
0 46113 7 1 2 46106 46112
0 46114 5 1 1 46113
0 46115 7 1 2 85574 46114
0 46116 5 1 1 46115
0 46117 7 1 2 66622 93335
0 46118 5 1 1 46117
0 46119 7 1 2 73135 71965
0 46120 7 1 2 46118 46119
0 46121 5 1 1 46120
0 46122 7 1 2 80140 89488
0 46123 5 1 1 46122
0 46124 7 1 2 68268 92087
0 46125 5 1 1 46124
0 46126 7 1 2 46123 46125
0 46127 5 1 1 46126
0 46128 7 1 2 71698 46127
0 46129 5 1 1 46128
0 46130 7 1 2 71111 92088
0 46131 5 1 1 46130
0 46132 7 1 2 61082 95141
0 46133 5 1 1 46132
0 46134 7 1 2 46131 46133
0 46135 5 1 1 46134
0 46136 7 1 2 93806 46135
0 46137 5 1 1 46136
0 46138 7 1 2 46129 46137
0 46139 7 1 2 46121 46138
0 46140 5 1 1 46139
0 46141 7 1 2 62804 46140
0 46142 5 1 1 46141
0 46143 7 1 2 60158 68269
0 46144 7 1 2 75090 46143
0 46145 7 1 2 91418 46144
0 46146 5 1 1 46145
0 46147 7 1 2 46142 46146
0 46148 7 1 2 46116 46147
0 46149 5 1 1 46148
0 46150 7 1 2 61445 46149
0 46151 5 1 1 46150
0 46152 7 1 2 76935 93286
0 46153 7 1 2 91419 46152
0 46154 5 1 1 46153
0 46155 7 1 2 46151 46154
0 46156 5 1 1 46155
0 46157 7 1 2 63101 46156
0 46158 5 1 1 46157
0 46159 7 1 2 45865 46158
0 46160 5 1 1 46159
0 46161 7 1 2 91355 46160
0 46162 5 1 1 46161
0 46163 7 1 2 86003 71104
0 46164 5 1 1 46163
0 46165 7 1 2 67497 46164
0 46166 5 1 1 46165
0 46167 7 1 2 83167 46166
0 46168 5 1 1 46167
0 46169 7 1 2 76119 94696
0 46170 5 1 1 46169
0 46171 7 1 2 73762 82021
0 46172 7 1 2 93954 46171
0 46173 5 1 1 46172
0 46174 7 1 2 46170 46173
0 46175 5 1 1 46174
0 46176 7 1 2 70874 46175
0 46177 5 1 1 46176
0 46178 7 1 2 46168 46177
0 46179 5 1 1 46178
0 46180 7 1 2 66050 46179
0 46181 5 1 1 46180
0 46182 7 3 2 59008 64835
0 46183 7 1 2 72357 67531
0 46184 7 1 2 95173 46183
0 46185 5 1 1 46184
0 46186 7 1 2 67498 46185
0 46187 5 1 1 46186
0 46188 7 1 2 94523 46187
0 46189 5 1 1 46188
0 46190 7 1 2 46181 46189
0 46191 5 1 1 46190
0 46192 7 1 2 65704 46191
0 46193 5 1 1 46192
0 46194 7 2 2 67532 79182
0 46195 5 1 1 95176
0 46196 7 1 2 73954 84094
0 46197 5 1 1 46196
0 46198 7 1 2 46195 46197
0 46199 5 1 1 46198
0 46200 7 1 2 68045 46199
0 46201 5 1 1 46200
0 46202 7 2 2 72914 82022
0 46203 5 1 1 95178
0 46204 7 1 2 59920 95179
0 46205 5 1 1 46204
0 46206 7 1 2 46201 46205
0 46207 5 1 1 46206
0 46208 7 1 2 58345 46207
0 46209 5 1 1 46208
0 46210 7 1 2 90215 94294
0 46211 5 1 1 46210
0 46212 7 1 2 46209 46211
0 46213 5 1 1 46212
0 46214 7 1 2 58647 46213
0 46215 5 1 1 46214
0 46216 7 1 2 73476 83168
0 46217 7 1 2 67551 46216
0 46218 5 1 1 46217
0 46219 7 1 2 73388 84095
0 46220 7 1 2 93225 46219
0 46221 5 1 1 46220
0 46222 7 1 2 46218 46221
0 46223 5 1 1 46222
0 46224 7 1 2 74074 46223
0 46225 5 1 1 46224
0 46226 7 1 2 72644 94524
0 46227 5 1 1 46226
0 46228 7 1 2 46225 46227
0 46229 5 1 1 46228
0 46230 7 1 2 76465 46229
0 46231 5 1 1 46230
0 46232 7 1 2 46215 46231
0 46233 7 1 2 46193 46232
0 46234 7 1 2 46162 46233
0 46235 5 1 1 46234
0 46236 7 1 2 61703 46235
0 46237 5 1 1 46236
0 46238 7 1 2 76946 74995
0 46239 5 1 1 46238
0 46240 7 1 2 38591 46239
0 46241 5 1 1 46240
0 46242 7 1 2 61446 46241
0 46243 5 1 1 46242
0 46244 7 1 2 69007 71649
0 46245 5 1 1 46244
0 46246 7 1 2 73801 46245
0 46247 5 1 1 46246
0 46248 7 1 2 63407 46247
0 46249 5 1 1 46248
0 46250 7 1 2 46243 46249
0 46251 5 1 1 46250
0 46252 7 1 2 65315 46251
0 46253 5 1 1 46252
0 46254 7 1 2 67381 83442
0 46255 5 1 1 46254
0 46256 7 1 2 63102 46255
0 46257 5 1 1 46256
0 46258 7 1 2 94725 46257
0 46259 5 1 1 46258
0 46260 7 1 2 68172 46259
0 46261 5 1 1 46260
0 46262 7 1 2 62272 35532
0 46263 5 1 1 46262
0 46264 7 1 2 86004 46263
0 46265 7 1 2 94067 46264
0 46266 5 1 1 46265
0 46267 7 1 2 76228 46266
0 46268 5 1 1 46267
0 46269 7 1 2 46261 46268
0 46270 5 1 1 46269
0 46271 7 1 2 66051 46270
0 46272 5 1 1 46271
0 46273 7 1 2 69999 94851
0 46274 5 1 1 46273
0 46275 7 1 2 63103 46274
0 46276 5 1 1 46275
0 46277 7 1 2 63408 46276
0 46278 5 1 1 46277
0 46279 7 1 2 46272 46278
0 46280 7 1 2 46253 46279
0 46281 5 1 1 46280
0 46282 7 1 2 59657 46281
0 46283 5 1 1 46282
0 46284 7 1 2 66052 93401
0 46285 5 1 1 46284
0 46286 7 1 2 40925 46285
0 46287 5 1 1 46286
0 46288 7 1 2 59658 46287
0 46289 5 1 1 46288
0 46290 7 1 2 68046 80454
0 46291 5 1 1 46290
0 46292 7 1 2 46289 46291
0 46293 5 1 1 46292
0 46294 7 1 2 74382 46293
0 46295 5 1 1 46294
0 46296 7 1 2 57780 73989
0 46297 5 1 1 46296
0 46298 7 1 2 93613 46297
0 46299 5 1 1 46298
0 46300 7 1 2 65082 46299
0 46301 5 1 1 46300
0 46302 7 1 2 73440 46301
0 46303 5 1 1 46302
0 46304 7 1 2 86732 46303
0 46305 5 1 1 46304
0 46306 7 1 2 46295 46305
0 46307 7 1 2 46283 46306
0 46308 5 1 1 46307
0 46309 7 1 2 71078 46308
0 46310 5 1 1 46309
0 46311 7 1 2 78992 94588
0 46312 5 1 1 46311
0 46313 7 1 2 75469 77738
0 46314 5 1 1 46313
0 46315 7 1 2 61083 46314
0 46316 7 1 2 46312 46315
0 46317 5 1 1 46316
0 46318 7 1 2 73782 93148
0 46319 5 1 1 46318
0 46320 7 1 2 73639 46319
0 46321 5 1 1 46320
0 46322 7 1 2 68173 46321
0 46323 5 1 1 46322
0 46324 7 1 2 68791 84155
0 46325 5 1 1 46324
0 46326 7 1 2 61447 46325
0 46327 5 1 1 46326
0 46328 7 2 2 76229 73783
0 46329 5 1 1 95180
0 46330 7 1 2 58648 46329
0 46331 7 1 2 46327 46330
0 46332 5 1 1 46331
0 46333 7 1 2 80451 46332
0 46334 5 1 1 46333
0 46335 7 1 2 46323 46334
0 46336 7 1 2 46317 46335
0 46337 5 1 1 46336
0 46338 7 1 2 59659 46337
0 46339 5 1 1 46338
0 46340 7 1 2 58649 93176
0 46341 5 1 1 46340
0 46342 7 1 2 73323 46341
0 46343 5 1 1 46342
0 46344 7 1 2 59165 61448
0 46345 7 1 2 94952 46344
0 46346 5 1 1 46345
0 46347 7 1 2 46343 46346
0 46348 5 1 1 46347
0 46349 7 1 2 65316 46348
0 46350 5 1 1 46349
0 46351 7 1 2 72036 84505
0 46352 7 1 2 92914 46351
0 46353 5 1 1 46352
0 46354 7 1 2 46350 46353
0 46355 7 1 2 46339 46354
0 46356 5 1 1 46355
0 46357 7 1 2 82023 46356
0 46358 5 1 1 46357
0 46359 7 1 2 46310 46358
0 46360 5 1 1 46359
0 46361 7 1 2 59921 46360
0 46362 5 1 1 46361
0 46363 7 1 2 71079 38616
0 46364 5 1 1 46363
0 46365 7 1 2 7453 46364
0 46366 5 1 1 46365
0 46367 7 1 2 73503 46366
0 46368 5 1 1 46367
0 46369 7 1 2 71375 90216
0 46370 5 1 1 46369
0 46371 7 1 2 59383 72974
0 46372 7 1 2 80171 46371
0 46373 7 1 2 83891 46372
0 46374 5 1 1 46373
0 46375 7 1 2 46370 46374
0 46376 5 1 1 46375
0 46377 7 1 2 71524 46376
0 46378 5 1 1 46377
0 46379 7 2 2 67533 71348
0 46380 5 1 1 95182
0 46381 7 1 2 69338 93966
0 46382 5 1 1 46381
0 46383 7 1 2 46380 46382
0 46384 5 1 1 46383
0 46385 7 1 2 71219 46384
0 46386 5 1 1 46385
0 46387 7 1 2 46378 46386
0 46388 7 1 2 46368 46387
0 46389 5 1 1 46388
0 46390 7 1 2 58650 46389
0 46391 5 1 1 46390
0 46392 7 1 2 73678 93914
0 46393 7 1 2 75717 46392
0 46394 7 1 2 82031 46393
0 46395 5 1 1 46394
0 46396 7 1 2 46391 46395
0 46397 7 1 2 46362 46396
0 46398 5 1 1 46397
0 46399 7 1 2 66349 46398
0 46400 5 1 1 46399
0 46401 7 1 2 46237 46400
0 46402 7 1 2 46097 46401
0 46403 5 1 1 46402
0 46404 7 1 2 66931 46403
0 46405 5 1 1 46404
0 46406 7 1 2 90274 94530
0 46407 5 1 1 46406
0 46408 7 3 2 67534 79302
0 46409 7 1 2 74545 82418
0 46410 7 1 2 95184 46409
0 46411 5 1 1 46410
0 46412 7 1 2 46407 46411
0 46413 5 1 1 46412
0 46414 7 1 2 68174 69090
0 46415 5 1 1 46414
0 46416 7 1 2 57485 46415
0 46417 5 1 1 46416
0 46418 7 1 2 59384 86345
0 46419 5 1 1 46418
0 46420 7 2 2 46417 46419
0 46421 7 1 2 62529 95187
0 46422 5 1 1 46421
0 46423 7 1 2 86774 46422
0 46424 5 1 1 46423
0 46425 7 1 2 60673 46424
0 46426 5 1 1 46425
0 46427 7 1 2 63104 85025
0 46428 5 1 1 46427
0 46429 7 1 2 93811 46428
0 46430 7 1 2 94280 46429
0 46431 7 1 2 46426 46430
0 46432 5 1 1 46431
0 46433 7 1 2 93380 46432
0 46434 5 1 1 46433
0 46435 7 1 2 60674 86109
0 46436 7 1 2 79601 46435
0 46437 7 1 2 94657 46436
0 46438 5 1 1 46437
0 46439 7 1 2 46434 46438
0 46440 5 1 1 46439
0 46441 7 1 2 46413 46440
0 46442 5 1 1 46441
0 46443 7 1 2 82024 89764
0 46444 5 1 1 46443
0 46445 7 2 2 87203 67535
0 46446 7 1 2 72109 95189
0 46447 5 1 1 46446
0 46448 7 1 2 46444 46447
0 46449 5 1 1 46448
0 46450 7 1 2 59660 46449
0 46451 5 1 1 46450
0 46452 7 1 2 82327 93980
0 46453 5 1 1 46452
0 46454 7 1 2 46451 46453
0 46455 5 1 1 46454
0 46456 7 1 2 59009 46455
0 46457 5 1 1 46456
0 46458 7 1 2 59010 91485
0 46459 5 1 1 46458
0 46460 7 1 2 85832 46459
0 46461 5 1 1 46460
0 46462 7 1 2 69157 67437
0 46463 7 1 2 46461 46462
0 46464 5 1 1 46463
0 46465 7 1 2 87504 71080
0 46466 5 1 1 46465
0 46467 7 1 2 61704 46466
0 46468 7 1 2 46464 46467
0 46469 5 1 1 46468
0 46470 7 2 2 60159 85804
0 46471 7 1 2 83740 95191
0 46472 5 1 1 46471
0 46473 7 1 2 66053 95183
0 46474 5 1 1 46473
0 46475 7 1 2 46472 46474
0 46476 5 1 1 46475
0 46477 7 1 2 59011 46476
0 46478 5 1 1 46477
0 46479 7 1 2 59661 74996
0 46480 5 3 1 46479
0 46481 7 1 2 61449 95193
0 46482 5 1 1 46481
0 46483 7 1 2 66054 77365
0 46484 5 1 1 46483
0 46485 7 1 2 71081 46484
0 46486 7 1 2 46482 46485
0 46487 5 1 1 46486
0 46488 7 1 2 66350 46487
0 46489 7 1 2 46478 46488
0 46490 5 1 1 46489
0 46491 7 1 2 57486 46490
0 46492 7 1 2 46469 46491
0 46493 5 1 1 46492
0 46494 7 1 2 82309 91189
0 46495 5 1 1 46494
0 46496 7 1 2 46493 46495
0 46497 7 1 2 46457 46496
0 46498 5 1 1 46497
0 46499 7 1 2 57781 46498
0 46500 5 1 1 46499
0 46501 7 1 2 60417 11967
0 46502 5 1 1 46501
0 46503 7 1 2 59012 46502
0 46504 7 1 2 92711 46503
0 46505 5 1 1 46504
0 46506 7 1 2 94424 46505
0 46507 5 1 1 46506
0 46508 7 1 2 71082 46507
0 46509 5 1 1 46508
0 46510 7 1 2 82025 94941
0 46511 5 1 1 46510
0 46512 7 1 2 46509 46511
0 46513 5 1 1 46512
0 46514 7 1 2 59662 46513
0 46515 5 1 1 46514
0 46516 7 3 2 74296 69246
0 46517 5 1 1 95196
0 46518 7 1 2 7604 46517
0 46519 5 1 1 46518
0 46520 7 1 2 66055 87344
0 46521 7 1 2 46519 46520
0 46522 5 1 1 46521
0 46523 7 1 2 46515 46522
0 46524 7 1 2 46500 46523
0 46525 5 1 1 46524
0 46526 7 1 2 59166 46525
0 46527 5 1 1 46526
0 46528 7 1 2 76510 91427
0 46529 5 1 1 46528
0 46530 7 1 2 57487 87424
0 46531 5 1 1 46530
0 46532 7 1 2 46529 46531
0 46533 5 1 1 46532
0 46534 7 1 2 59663 46533
0 46535 5 1 1 46534
0 46536 7 1 2 72202 82580
0 46537 5 1 1 46536
0 46538 7 1 2 94437 46537
0 46539 5 1 1 46538
0 46540 7 1 2 73324 46539
0 46541 5 1 1 46540
0 46542 7 1 2 46535 46541
0 46543 5 1 1 46542
0 46544 7 1 2 71083 46543
0 46545 5 1 1 46544
0 46546 7 1 2 46527 46545
0 46547 5 1 1 46546
0 46548 7 1 2 65317 46547
0 46549 5 1 1 46548
0 46550 7 1 2 66056 44701
0 46551 5 1 1 46550
0 46552 7 1 2 81713 46551
0 46553 5 1 1 46552
0 46554 7 1 2 71084 46553
0 46555 5 1 1 46554
0 46556 7 1 2 46203 46555
0 46557 5 1 1 46556
0 46558 7 1 2 65705 46557
0 46559 5 1 1 46558
0 46560 7 1 2 57782 81696
0 46561 7 1 2 67494 46560
0 46562 5 1 1 46561
0 46563 7 1 2 46559 46562
0 46564 5 1 1 46563
0 46565 7 1 2 82581 46564
0 46566 5 1 1 46565
0 46567 7 1 2 86374 73522
0 46568 5 1 1 46567
0 46569 7 1 2 82026 46568
0 46570 5 1 1 46569
0 46571 7 1 2 12239 73523
0 46572 5 1 1 46571
0 46573 7 1 2 69881 67552
0 46574 7 1 2 46572 46573
0 46575 5 1 1 46574
0 46576 7 1 2 46570 46575
0 46577 5 1 1 46576
0 46578 7 1 2 59013 46577
0 46579 5 1 1 46578
0 46580 7 1 2 73514 95197
0 46581 5 1 1 46580
0 46582 7 1 2 86370 82027
0 46583 5 1 1 46582
0 46584 7 1 2 46581 46583
0 46585 5 1 1 46584
0 46586 7 1 2 65083 46585
0 46587 5 1 1 46586
0 46588 7 1 2 46579 46587
0 46589 5 1 1 46588
0 46590 7 1 2 57488 46589
0 46591 5 1 1 46590
0 46592 7 1 2 86110 81902
0 46593 5 1 1 46592
0 46594 7 1 2 73551 67553
0 46595 5 1 1 46594
0 46596 7 1 2 46593 46595
0 46597 5 1 1 46596
0 46598 7 1 2 81697 46597
0 46599 5 1 1 46598
0 46600 7 1 2 85588 71955
0 46601 5 1 1 46600
0 46602 7 1 2 46599 46601
0 46603 7 1 2 46591 46602
0 46604 5 1 1 46603
0 46605 7 1 2 57783 46604
0 46606 5 1 1 46605
0 46607 7 1 2 73426 94707
0 46608 5 1 1 46607
0 46609 7 1 2 60160 86413
0 46610 7 1 2 90217 46609
0 46611 5 1 1 46610
0 46612 7 1 2 46608 46611
0 46613 5 1 1 46612
0 46614 7 1 2 94547 46613
0 46615 5 1 1 46614
0 46616 7 1 2 71379 90545
0 46617 7 1 2 71980 46616
0 46618 5 1 1 46617
0 46619 7 1 2 46615 46618
0 46620 7 1 2 46606 46619
0 46621 5 1 1 46620
0 46622 7 1 2 66351 46621
0 46623 5 1 1 46622
0 46624 7 1 2 46566 46623
0 46625 7 1 2 46549 46624
0 46626 5 1 1 46625
0 46627 7 1 2 66932 46626
0 46628 5 1 1 46627
0 46629 7 2 2 79292 74915
0 46630 7 2 2 84786 69247
0 46631 7 1 2 95199 95201
0 46632 5 1 1 46631
0 46633 7 2 2 66057 83024
0 46634 7 1 2 69008 73763
0 46635 7 1 2 75215 46634
0 46636 7 1 2 95203 46635
0 46637 7 1 2 91700 46636
0 46638 5 1 1 46637
0 46639 7 1 2 46632 46638
0 46640 5 1 1 46639
0 46641 7 1 2 57489 46640
0 46642 5 1 1 46641
0 46643 7 1 2 69401 87916
0 46644 7 1 2 87695 46643
0 46645 7 1 2 79308 84800
0 46646 7 1 2 46644 46645
0 46647 5 1 1 46646
0 46648 7 1 2 46642 46647
0 46649 5 1 1 46648
0 46650 7 1 2 66623 46649
0 46651 5 1 1 46650
0 46652 7 1 2 79313 82832
0 46653 7 1 2 89754 46652
0 46654 7 1 2 94733 46653
0 46655 5 1 1 46654
0 46656 7 1 2 46651 46655
0 46657 7 1 2 46628 46656
0 46658 5 1 1 46657
0 46659 7 1 2 85297 46658
0 46660 5 1 1 46659
0 46661 7 1 2 46442 46660
0 46662 7 1 2 46405 46661
0 46663 7 1 2 45803 46662
0 46664 7 1 2 45260 46663
0 46665 5 1 1 46664
0 46666 7 1 2 60201 88090
0 46667 7 1 2 46665 46666
0 46668 5 1 1 46667
0 46669 7 3 2 58346 76658
0 46670 5 2 1 95205
0 46671 7 2 2 71525 75216
0 46672 5 1 1 95210
0 46673 7 1 2 71334 46672
0 46674 5 1 1 46673
0 46675 7 1 2 75584 80606
0 46676 7 1 2 46674 46675
0 46677 5 1 1 46676
0 46678 7 1 2 95208 46677
0 46679 5 1 1 46678
0 46680 7 1 2 75962 46679
0 46681 5 1 1 46680
0 46682 7 2 2 66624 86673
0 46683 7 1 2 72617 95212
0 46684 7 1 2 92886 46683
0 46685 5 1 1 46684
0 46686 7 1 2 46681 46685
0 46687 5 1 1 46686
0 46688 7 1 2 61705 46687
0 46689 5 1 1 46688
0 46690 7 1 2 93722 95211
0 46691 5 1 1 46690
0 46692 7 1 2 92207 46691
0 46693 5 1 1 46692
0 46694 7 1 2 73566 46693
0 46695 5 1 1 46694
0 46696 7 1 2 78087 72962
0 46697 5 1 1 46696
0 46698 7 1 2 34864 46697
0 46699 5 1 1 46698
0 46700 7 1 2 60048 46699
0 46701 5 1 1 46700
0 46702 7 1 2 92208 46701
0 46703 5 1 1 46702
0 46704 7 1 2 93578 46703
0 46705 5 1 1 46704
0 46706 7 1 2 60049 74736
0 46707 7 1 2 94735 46706
0 46708 5 1 1 46707
0 46709 7 1 2 46705 46708
0 46710 5 1 1 46709
0 46711 7 1 2 59014 46710
0 46712 5 1 1 46711
0 46713 7 1 2 46695 46712
0 46714 5 1 1 46713
0 46715 7 1 2 82662 46714
0 46716 5 1 1 46715
0 46717 7 1 2 46689 46716
0 46718 5 1 1 46717
0 46719 7 1 2 65084 46718
0 46720 5 1 1 46719
0 46721 7 1 2 59015 85221
0 46722 5 1 1 46721
0 46723 7 1 2 27901 46722
0 46724 5 1 1 46723
0 46725 7 1 2 61706 46724
0 46726 5 1 1 46725
0 46727 7 3 2 66352 94229
0 46728 7 1 2 65318 95214
0 46729 5 1 1 46728
0 46730 7 1 2 46726 46729
0 46731 5 1 1 46730
0 46732 7 1 2 67680 75963
0 46733 7 1 2 46731 46732
0 46734 5 1 1 46733
0 46735 7 1 2 78935 92307
0 46736 7 1 2 87616 46735
0 46737 5 1 1 46736
0 46738 7 1 2 46734 46737
0 46739 5 1 1 46738
0 46740 7 1 2 65706 46739
0 46741 5 1 1 46740
0 46742 7 1 2 69850 95130
0 46743 5 1 1 46742
0 46744 7 1 2 69851 87204
0 46745 5 1 1 46744
0 46746 7 1 2 59922 92732
0 46747 5 1 1 46746
0 46748 7 1 2 46745 46747
0 46749 5 1 1 46748
0 46750 7 1 2 58651 46749
0 46751 5 1 1 46750
0 46752 7 1 2 46743 46751
0 46753 5 1 1 46752
0 46754 7 1 2 75964 46753
0 46755 5 1 1 46754
0 46756 7 1 2 75376 79986
0 46757 7 1 2 81216 46756
0 46758 7 1 2 90635 46757
0 46759 5 1 1 46758
0 46760 7 1 2 46755 46759
0 46761 5 1 1 46760
0 46762 7 1 2 71526 46761
0 46763 5 1 1 46762
0 46764 7 3 2 59664 76287
0 46765 5 1 1 95217
0 46766 7 1 2 93723 95218
0 46767 5 1 1 46766
0 46768 7 1 2 77833 93373
0 46769 5 1 1 46768
0 46770 7 1 2 60050 46769
0 46771 5 1 1 46770
0 46772 7 1 2 46767 46771
0 46773 5 1 1 46772
0 46774 7 1 2 95021 46773
0 46775 5 1 1 46774
0 46776 7 2 2 83981 84315
0 46777 7 1 2 81971 92001
0 46778 7 1 2 95220 46777
0 46779 5 1 1 46778
0 46780 7 1 2 46775 46779
0 46781 5 1 1 46780
0 46782 7 1 2 59016 46781
0 46783 5 1 1 46782
0 46784 7 2 2 75585 76288
0 46785 7 1 2 59665 95222
0 46786 5 1 1 46785
0 46787 7 1 2 76705 46786
0 46788 5 1 1 46787
0 46789 7 2 2 81120 81755
0 46790 7 1 2 46788 95224
0 46791 5 1 1 46790
0 46792 7 1 2 46783 46791
0 46793 5 1 1 46792
0 46794 7 1 2 66058 46793
0 46795 5 1 1 46794
0 46796 7 1 2 46763 46795
0 46797 7 1 2 46741 46796
0 46798 7 1 2 46720 46797
0 46799 5 1 1 46798
0 46800 7 1 2 57490 46799
0 46801 5 1 1 46800
0 46802 7 5 2 66353 79830
0 46803 7 1 2 59017 95226
0 46804 5 1 1 46803
0 46805 7 1 2 87561 46804
0 46806 5 1 1 46805
0 46807 7 1 2 58652 46806
0 46808 5 2 1 46807
0 46809 7 1 2 60051 94957
0 46810 5 1 1 46809
0 46811 7 1 2 95231 46810
0 46812 5 1 1 46811
0 46813 7 1 2 73679 46812
0 46814 5 1 1 46813
0 46815 7 1 2 78088 84680
0 46816 5 3 1 46815
0 46817 7 1 2 92726 95233
0 46818 5 1 1 46817
0 46819 7 1 2 60052 46818
0 46820 5 1 1 46819
0 46821 7 1 2 46814 46820
0 46822 5 1 1 46821
0 46823 7 1 2 75217 46822
0 46824 5 1 1 46823
0 46825 7 1 2 86501 92579
0 46826 5 1 1 46825
0 46827 7 1 2 18039 95232
0 46828 5 1 1 46827
0 46829 7 1 2 73680 46828
0 46830 5 1 1 46829
0 46831 7 1 2 79269 84758
0 46832 5 1 1 46831
0 46833 7 1 2 46830 46832
0 46834 5 1 1 46833
0 46835 7 1 2 58347 46834
0 46836 5 1 1 46835
0 46837 7 1 2 46826 46836
0 46838 7 1 2 46824 46837
0 46839 5 1 1 46838
0 46840 7 1 2 69167 46839
0 46841 5 1 1 46840
0 46842 7 1 2 65319 92137
0 46843 5 1 1 46842
0 46844 7 1 2 65707 77635
0 46845 7 1 2 90636 46844
0 46846 5 1 1 46845
0 46847 7 1 2 46843 46846
0 46848 5 1 1 46847
0 46849 7 1 2 59018 46848
0 46850 5 1 1 46849
0 46851 7 1 2 87001 95022
0 46852 5 1 1 46851
0 46853 7 1 2 77438 87617
0 46854 5 1 1 46853
0 46855 7 1 2 46852 46854
0 46856 7 1 2 46850 46855
0 46857 5 1 1 46856
0 46858 7 1 2 77236 46857
0 46859 5 1 1 46858
0 46860 7 1 2 46841 46859
0 46861 5 1 1 46860
0 46862 7 1 2 65085 46861
0 46863 5 1 1 46862
0 46864 7 1 2 86158 94211
0 46865 5 1 1 46864
0 46866 7 1 2 60053 94230
0 46867 5 1 1 46866
0 46868 7 1 2 93868 46867
0 46869 5 1 1 46868
0 46870 7 1 2 72411 46869
0 46871 5 1 1 46870
0 46872 7 1 2 46865 46871
0 46873 5 1 1 46872
0 46874 7 1 2 67681 46873
0 46875 5 1 1 46874
0 46876 7 1 2 86192 94212
0 46877 5 1 1 46876
0 46878 7 1 2 46875 46877
0 46879 5 1 1 46878
0 46880 7 1 2 61970 46879
0 46881 5 1 1 46880
0 46882 7 1 2 64738 94580
0 46883 5 1 1 46882
0 46884 7 1 2 46881 46883
0 46885 5 1 1 46884
0 46886 7 1 2 66354 46885
0 46887 5 1 1 46886
0 46888 7 1 2 76659 75218
0 46889 5 1 1 46888
0 46890 7 1 2 73681 95223
0 46891 5 1 1 46890
0 46892 7 1 2 46889 46891
0 46893 5 1 1 46892
0 46894 7 1 2 59019 46893
0 46895 5 1 1 46894
0 46896 7 1 2 95209 46895
0 46897 5 1 1 46896
0 46898 7 1 2 95225 46897
0 46899 5 1 1 46898
0 46900 7 1 2 85610 82117
0 46901 5 1 1 46900
0 46902 7 1 2 85779 81756
0 46903 7 1 2 88459 46902
0 46904 5 1 1 46903
0 46905 7 1 2 46901 46904
0 46906 5 1 1 46905
0 46907 7 1 2 93365 46906
0 46908 5 1 1 46907
0 46909 7 1 2 85611 83443
0 46910 5 1 1 46909
0 46911 7 1 2 86743 46910
0 46912 5 1 1 46911
0 46913 7 1 2 95213 46912
0 46914 5 1 1 46913
0 46915 7 1 2 87002 91410
0 46916 7 1 2 80082 46915
0 46917 5 1 1 46916
0 46918 7 1 2 46914 46917
0 46919 5 1 1 46918
0 46920 7 1 2 61707 46919
0 46921 5 1 1 46920
0 46922 7 1 2 75586 83898
0 46923 7 1 2 91749 46922
0 46924 5 1 1 46923
0 46925 7 1 2 35618 46924
0 46926 5 1 1 46925
0 46927 7 1 2 61971 90262
0 46928 7 1 2 46926 46927
0 46929 5 1 1 46928
0 46930 7 1 2 46921 46929
0 46931 5 1 1 46930
0 46932 7 1 2 71527 46931
0 46933 5 1 1 46932
0 46934 7 1 2 46908 46933
0 46935 7 1 2 46899 46934
0 46936 7 1 2 46887 46935
0 46937 7 1 2 46863 46936
0 46938 7 1 2 46801 46937
0 46939 5 1 1 46938
0 46940 7 1 2 63530 46939
0 46941 5 1 1 46940
0 46942 7 2 2 69009 82967
0 46943 5 1 1 95236
0 46944 7 1 2 63409 46765
0 46945 5 1 1 46944
0 46946 7 1 2 71747 46945
0 46947 5 1 1 46946
0 46948 7 1 2 84156 72037
0 46949 5 1 1 46948
0 46950 7 1 2 46947 46949
0 46951 5 1 1 46950
0 46952 7 1 2 65320 46951
0 46953 5 1 1 46952
0 46954 7 1 2 46943 46953
0 46955 5 1 1 46954
0 46956 7 1 2 57491 46955
0 46957 5 1 1 46956
0 46958 7 1 2 76302 95219
0 46959 5 1 1 46958
0 46960 7 1 2 64625 46959
0 46961 7 1 2 46957 46960
0 46962 5 1 1 46961
0 46963 7 1 2 59020 77996
0 46964 7 1 2 77313 46963
0 46965 5 1 1 46964
0 46966 7 1 2 36136 46965
0 46967 5 1 1 46966
0 46968 7 1 2 57492 46967
0 46969 5 1 1 46968
0 46970 7 1 2 77997 81217
0 46971 5 1 1 46970
0 46972 7 1 2 59923 46971
0 46973 7 1 2 46969 46972
0 46974 5 1 1 46973
0 46975 7 1 2 66059 46974
0 46976 7 1 2 46962 46975
0 46977 5 1 1 46976
0 46978 7 1 2 70059 94235
0 46979 5 1 1 46978
0 46980 7 1 2 70889 94253
0 46981 5 1 1 46980
0 46982 7 2 2 65321 76466
0 46983 7 1 2 94231 95238
0 46984 5 1 1 46983
0 46985 7 1 2 46981 46984
0 46986 5 1 1 46985
0 46987 7 1 2 67682 46986
0 46988 5 1 1 46987
0 46989 7 1 2 80767 94143
0 46990 5 1 1 46989
0 46991 7 1 2 58653 73729
0 46992 5 1 1 46991
0 46993 7 1 2 46990 46992
0 46994 7 1 2 46988 46993
0 46995 5 1 1 46994
0 46996 7 1 2 65708 46995
0 46997 5 1 1 46996
0 46998 7 1 2 46979 46997
0 46999 7 1 2 46977 46998
0 47000 5 1 1 46999
0 47001 7 1 2 66355 47000
0 47002 5 1 1 47001
0 47003 7 1 2 85805 81407
0 47004 5 1 1 47003
0 47005 7 2 2 73325 81538
0 47006 5 1 1 95240
0 47007 7 1 2 47004 47006
0 47008 5 1 1 47007
0 47009 7 1 2 67683 47008
0 47010 5 1 1 47009
0 47011 7 1 2 75241 87205
0 47012 5 1 1 47011
0 47013 7 1 2 47010 47012
0 47014 5 1 1 47013
0 47015 7 1 2 71528 47014
0 47016 5 1 1 47015
0 47017 7 1 2 70364 88888
0 47018 5 1 1 47017
0 47019 7 1 2 85849 47018
0 47020 5 1 1 47019
0 47021 7 1 2 66060 47020
0 47022 5 1 1 47021
0 47023 7 2 2 57493 72831
0 47024 7 1 2 76123 95242
0 47025 5 1 1 47024
0 47026 7 1 2 47022 47025
0 47027 5 1 1 47026
0 47028 7 1 2 82387 47027
0 47029 5 1 1 47028
0 47030 7 1 2 47016 47029
0 47031 5 1 1 47030
0 47032 7 1 2 75587 47031
0 47033 5 1 1 47032
0 47034 7 1 2 78385 93580
0 47035 5 1 1 47034
0 47036 7 1 2 76467 47035
0 47037 5 1 1 47036
0 47038 7 1 2 72681 9455
0 47039 5 1 1 47038
0 47040 7 1 2 57494 47039
0 47041 5 1 1 47040
0 47042 7 1 2 64408 79741
0 47043 5 1 1 47042
0 47044 7 1 2 65709 47043
0 47045 5 1 1 47044
0 47046 7 1 2 78727 47045
0 47047 7 1 2 47041 47046
0 47048 7 1 2 47037 47047
0 47049 5 1 1 47048
0 47050 7 1 2 89359 47049
0 47051 5 1 1 47050
0 47052 7 1 2 47033 47051
0 47053 7 1 2 47002 47052
0 47054 5 1 1 47053
0 47055 7 1 2 64739 47054
0 47056 5 1 1 47055
0 47057 7 6 2 61708 84013
0 47058 5 1 1 95244
0 47059 7 1 2 61450 79387
0 47060 5 1 1 47059
0 47061 7 1 2 74920 47060
0 47062 5 1 1 47061
0 47063 7 1 2 61084 47062
0 47064 5 1 1 47063
0 47065 7 1 2 70101 85742
0 47066 5 1 1 47065
0 47067 7 1 2 47064 47066
0 47068 5 1 1 47067
0 47069 7 1 2 71748 47068
0 47070 5 1 1 47069
0 47071 7 1 2 69466 87078
0 47072 5 1 1 47071
0 47073 7 1 2 74721 47072
0 47074 5 1 1 47073
0 47075 7 1 2 61085 47074
0 47076 5 1 1 47075
0 47077 7 1 2 67597 87375
0 47078 5 1 1 47077
0 47079 7 1 2 63105 47078
0 47080 5 1 1 47079
0 47081 7 1 2 85743 47080
0 47082 5 1 1 47081
0 47083 7 1 2 47076 47082
0 47084 7 1 2 47070 47083
0 47085 5 2 1 47084
0 47086 7 1 2 95245 95250
0 47087 5 1 1 47086
0 47088 7 1 2 47056 47087
0 47089 5 1 1 47088
0 47090 7 1 2 75686 47089
0 47091 5 1 1 47090
0 47092 7 1 2 46941 47091
0 47093 5 1 1 47092
0 47094 7 1 2 64836 47093
0 47095 5 1 1 47094
0 47096 7 1 2 95251 95069
0 47097 5 1 1 47096
0 47098 7 1 2 66721 47097
0 47099 7 1 2 47095 47098
0 47100 5 1 1 47099
0 47101 7 1 2 63531 93569
0 47102 5 1 1 47101
0 47103 7 1 2 86029 81691
0 47104 5 1 1 47103
0 47105 7 1 2 47102 47104
0 47106 5 1 1 47105
0 47107 7 1 2 92206 47106
0 47108 5 1 1 47107
0 47109 7 1 2 83626 43522
0 47110 5 1 1 47109
0 47111 7 1 2 59924 47110
0 47112 5 1 1 47111
0 47113 7 1 2 58654 83623
0 47114 5 1 1 47113
0 47115 7 1 2 85937 81692
0 47116 5 1 1 47115
0 47117 7 1 2 47114 47116
0 47118 7 1 2 47112 47117
0 47119 5 1 1 47118
0 47120 7 1 2 61451 47119
0 47121 5 1 1 47120
0 47122 7 1 2 82968 93570
0 47123 5 1 1 47122
0 47124 7 1 2 86240 86848
0 47125 5 1 1 47124
0 47126 7 1 2 47123 47125
0 47127 5 1 1 47126
0 47128 7 1 2 64626 47127
0 47129 5 1 1 47128
0 47130 7 1 2 87505 87743
0 47131 5 1 1 47130
0 47132 7 1 2 47129 47131
0 47133 7 1 2 47121 47132
0 47134 5 1 1 47133
0 47135 7 1 2 66933 47134
0 47136 5 1 1 47135
0 47137 7 1 2 47108 47136
0 47138 5 1 1 47137
0 47139 7 1 2 66625 47138
0 47140 5 1 1 47139
0 47141 7 1 2 68792 83258
0 47142 5 1 1 47141
0 47143 7 1 2 63106 47142
0 47144 5 1 1 47143
0 47145 7 2 2 66061 47144
0 47146 5 1 1 95252
0 47147 7 1 2 75663 91745
0 47148 7 1 2 95253 47147
0 47149 5 1 1 47148
0 47150 7 1 2 47140 47149
0 47151 5 1 1 47150
0 47152 7 1 2 66356 47151
0 47153 5 1 1 47152
0 47154 7 3 2 58797 72876
0 47155 5 1 1 95254
0 47156 7 1 2 64627 95255
0 47157 5 1 1 47156
0 47158 7 1 2 39621 47157
0 47159 5 1 1 47158
0 47160 7 1 2 68637 47159
0 47161 5 1 1 47160
0 47162 7 1 2 80609 82708
0 47163 5 1 1 47162
0 47164 7 2 2 58348 47163
0 47165 7 1 2 79029 95257
0 47166 5 1 1 47165
0 47167 7 1 2 47161 47166
0 47168 5 2 1 47167
0 47169 7 1 2 65086 95259
0 47170 5 1 1 47169
0 47171 7 1 2 85806 79642
0 47172 5 1 1 47171
0 47173 7 1 2 79033 47172
0 47174 5 1 1 47173
0 47175 7 1 2 58655 47174
0 47176 5 1 1 47175
0 47177 7 1 2 85807 79557
0 47178 5 1 1 47177
0 47179 7 1 2 47176 47178
0 47180 5 1 1 47179
0 47181 7 1 2 68793 47180
0 47182 5 1 1 47181
0 47183 7 1 2 47170 47182
0 47184 5 1 1 47183
0 47185 7 1 2 65322 47184
0 47186 5 1 1 47185
0 47187 7 1 2 63532 84488
0 47188 5 7 1 47187
0 47189 7 2 2 70875 78493
0 47190 5 1 1 95268
0 47191 7 1 2 92308 95269
0 47192 7 1 2 95261 47191
0 47193 5 1 1 47192
0 47194 7 1 2 47186 47193
0 47195 5 1 1 47194
0 47196 7 1 2 65710 47195
0 47197 5 1 1 47196
0 47198 7 1 2 85717 79558
0 47199 5 1 1 47198
0 47200 7 1 2 80438 79559
0 47201 5 2 1 47200
0 47202 7 2 2 63533 75588
0 47203 7 1 2 92194 95272
0 47204 5 1 1 47203
0 47205 7 1 2 95270 47204
0 47206 5 1 1 47205
0 47207 7 1 2 58349 47206
0 47208 5 1 1 47207
0 47209 7 1 2 47199 47208
0 47210 7 1 2 47197 47209
0 47211 5 1 1 47210
0 47212 7 1 2 60054 47211
0 47213 5 1 1 47212
0 47214 7 3 2 59925 86849
0 47215 5 1 1 95274
0 47216 7 1 2 93611 95275
0 47217 5 1 1 47216
0 47218 7 1 2 74346 78971
0 47219 5 1 1 47218
0 47220 7 1 2 61452 47219
0 47221 5 1 1 47220
0 47222 7 1 2 59666 47221
0 47223 5 1 1 47222
0 47224 7 1 2 85780 72412
0 47225 5 1 1 47224
0 47226 7 1 2 76706 47225
0 47227 7 1 2 47223 47226
0 47228 5 1 1 47227
0 47229 7 1 2 80768 47228
0 47230 5 1 1 47229
0 47231 7 1 2 47217 47230
0 47232 5 1 1 47231
0 47233 7 1 2 79433 47232
0 47234 5 1 1 47233
0 47235 7 1 2 47213 47234
0 47236 5 1 1 47235
0 47237 7 1 2 82105 47236
0 47238 5 1 1 47237
0 47239 7 3 2 66871 84448
0 47240 5 1 1 95277
0 47241 7 1 2 76303 94863
0 47242 5 1 1 47241
0 47243 7 1 2 7447 47242
0 47244 5 1 1 47243
0 47245 7 1 2 58350 47244
0 47246 5 1 1 47245
0 47247 7 1 2 82540 93760
0 47248 5 1 1 47247
0 47249 7 1 2 47246 47248
0 47250 5 1 1 47249
0 47251 7 1 2 57495 47250
0 47252 5 1 1 47251
0 47253 7 1 2 69830 83928
0 47254 5 1 1 47253
0 47255 7 1 2 86571 47254
0 47256 5 1 1 47255
0 47257 7 1 2 47252 47256
0 47258 5 1 1 47257
0 47259 7 1 2 95278 47258
0 47260 5 1 1 47259
0 47261 7 1 2 68794 70060
0 47262 5 1 1 47261
0 47263 7 2 2 71529 80498
0 47264 7 1 2 65711 95280
0 47265 5 1 1 47264
0 47266 7 1 2 47262 47265
0 47267 5 1 1 47266
0 47268 7 1 2 95227 47267
0 47269 5 1 1 47268
0 47270 7 1 2 81434 82365
0 47271 5 1 1 47270
0 47272 7 1 2 47269 47271
0 47273 5 1 1 47272
0 47274 7 1 2 76928 47273
0 47275 5 1 1 47274
0 47276 7 2 2 75589 82388
0 47277 5 1 1 95282
0 47278 7 1 2 82216 95281
0 47279 5 1 1 47278
0 47280 7 1 2 47277 47279
0 47281 5 1 1 47280
0 47282 7 1 2 65712 47281
0 47283 5 1 1 47282
0 47284 7 1 2 87515 81374
0 47285 5 1 1 47284
0 47286 7 1 2 47283 47285
0 47287 5 1 1 47286
0 47288 7 1 2 66934 47287
0 47289 5 1 1 47288
0 47290 7 1 2 47275 47289
0 47291 5 1 1 47290
0 47292 7 1 2 66062 47291
0 47293 5 1 1 47292
0 47294 7 1 2 83259 94011
0 47295 5 1 1 47294
0 47296 7 1 2 77158 87641
0 47297 5 1 1 47296
0 47298 7 2 2 76511 87553
0 47299 7 1 2 64628 95284
0 47300 5 1 1 47299
0 47301 7 1 2 47297 47300
0 47302 5 1 1 47301
0 47303 7 1 2 65323 47302
0 47304 5 1 1 47303
0 47305 7 3 2 60055 81448
0 47306 5 1 1 95286
0 47307 7 1 2 92311 95287
0 47308 5 1 1 47307
0 47309 7 1 2 61086 47308
0 47310 7 1 2 47304 47309
0 47311 5 1 1 47310
0 47312 7 3 2 66357 75377
0 47313 5 1 1 95289
0 47314 7 1 2 59926 95290
0 47315 5 1 1 47314
0 47316 7 1 2 84014 82689
0 47317 5 2 1 47316
0 47318 7 1 2 65713 95292
0 47319 7 1 2 47315 47318
0 47320 5 1 1 47319
0 47321 7 1 2 95262 47320
0 47322 7 1 2 47311 47321
0 47323 5 1 1 47322
0 47324 7 3 2 82969 79908
0 47325 5 1 1 95294
0 47326 7 1 2 92356 47325
0 47327 5 1 1 47326
0 47328 7 1 2 66358 80074
0 47329 7 1 2 92461 47328
0 47330 7 1 2 47327 47329
0 47331 5 1 1 47330
0 47332 7 1 2 47323 47331
0 47333 5 1 1 47332
0 47334 7 1 2 61453 47333
0 47335 5 1 1 47334
0 47336 7 1 2 47295 47335
0 47337 7 1 2 47293 47336
0 47338 5 1 1 47337
0 47339 7 1 2 66626 47338
0 47340 5 1 1 47339
0 47341 7 1 2 47260 47340
0 47342 5 1 1 47341
0 47343 7 1 2 67684 47342
0 47344 5 1 1 47343
0 47345 7 1 2 47238 47344
0 47346 7 1 2 47153 47345
0 47347 5 1 1 47346
0 47348 7 1 2 60161 47347
0 47349 5 1 1 47348
0 47350 7 2 2 59667 74223
0 47351 5 1 1 95297
0 47352 7 2 2 72679 95298
0 47353 5 1 1 95299
0 47354 7 2 2 65324 76578
0 47355 5 1 1 95301
0 47356 7 1 2 74149 47355
0 47357 5 1 1 47356
0 47358 7 1 2 59021 47357
0 47359 5 1 1 47358
0 47360 7 1 2 60675 76453
0 47361 5 1 1 47360
0 47362 7 1 2 82292 47361
0 47363 5 1 1 47362
0 47364 7 1 2 47359 47363
0 47365 5 1 1 47364
0 47366 7 1 2 66063 47365
0 47367 5 1 1 47366
0 47368 7 1 2 47353 47367
0 47369 5 1 1 47368
0 47370 7 1 2 67685 47369
0 47371 5 1 1 47370
0 47372 7 1 2 90016 47371
0 47373 5 1 1 47372
0 47374 7 1 2 66627 82713
0 47375 7 1 2 92520 47374
0 47376 7 1 2 47373 47375
0 47377 5 1 1 47376
0 47378 7 1 2 62115 47377
0 47379 7 1 2 47349 47378
0 47380 5 1 1 47379
0 47381 7 1 2 63642 47380
0 47382 7 1 2 47100 47381
0 47383 5 1 1 47382
0 47384 7 2 2 58351 78895
0 47385 7 2 2 75590 79434
0 47386 5 1 1 95305
0 47387 7 1 2 92357 47386
0 47388 5 3 1 47387
0 47389 7 1 2 67482 95307
0 47390 7 2 2 95303 47389
0 47391 5 1 1 95310
0 47392 7 1 2 60162 95311
0 47393 5 1 1 47392
0 47394 7 1 2 67068 91656
0 47395 5 1 1 47394
0 47396 7 4 2 75591 79909
0 47397 7 2 2 80736 72832
0 47398 7 1 2 95312 95316
0 47399 5 1 1 47398
0 47400 7 1 2 85388 47399
0 47401 5 1 1 47400
0 47402 7 1 2 61972 47401
0 47403 5 1 1 47402
0 47404 7 1 2 74432 94578
0 47405 5 1 1 47404
0 47406 7 1 2 80769 84340
0 47407 7 1 2 88845 47406
0 47408 5 1 1 47407
0 47409 7 1 2 47405 47408
0 47410 5 1 1 47409
0 47411 7 1 2 76468 47410
0 47412 5 1 1 47411
0 47413 7 1 2 47403 47412
0 47414 5 1 1 47413
0 47415 7 1 2 64837 47414
0 47416 5 1 1 47415
0 47417 7 1 2 47395 47416
0 47418 5 1 1 47417
0 47419 7 1 2 66722 47418
0 47420 5 1 1 47419
0 47421 7 1 2 47393 47420
0 47422 5 1 1 47421
0 47423 7 1 2 63643 47422
0 47424 5 1 1 47423
0 47425 7 1 2 67536 91657
0 47426 5 1 1 47425
0 47427 7 1 2 47391 47426
0 47428 5 1 1 47427
0 47429 7 1 2 70458 47428
0 47430 5 1 1 47429
0 47431 7 1 2 47424 47430
0 47432 5 1 1 47431
0 47433 7 1 2 65714 47432
0 47434 5 1 1 47433
0 47435 7 1 2 70555 88036
0 47436 5 1 1 47435
0 47437 7 1 2 47434 47436
0 47438 5 1 1 47437
0 47439 7 1 2 61709 47438
0 47440 5 1 1 47439
0 47441 7 1 2 82333 83427
0 47442 5 1 1 47441
0 47443 7 1 2 60056 85763
0 47444 7 1 2 70547 47443
0 47445 7 1 2 95304 47444
0 47446 5 1 1 47445
0 47447 7 1 2 47442 47446
0 47448 5 1 1 47447
0 47449 7 1 2 58798 47448
0 47450 5 1 1 47449
0 47451 7 1 2 63410 76030
0 47452 7 1 2 72563 81984
0 47453 7 1 2 47451 47452
0 47454 5 1 1 47453
0 47455 7 1 2 47450 47454
0 47456 5 1 1 47455
0 47457 7 1 2 82461 47456
0 47458 5 1 1 47457
0 47459 7 1 2 47440 47458
0 47460 5 1 1 47459
0 47461 7 1 2 72915 47460
0 47462 5 1 1 47461
0 47463 7 2 2 74997 94510
0 47464 5 1 1 95318
0 47465 7 1 2 58656 95319
0 47466 5 1 1 47465
0 47467 7 1 2 79439 93940
0 47468 5 2 1 47467
0 47469 7 1 2 58657 95320
0 47470 5 1 1 47469
0 47471 7 1 2 92161 47470
0 47472 5 1 1 47471
0 47473 7 1 2 72413 47472
0 47474 5 1 1 47473
0 47475 7 1 2 47466 47474
0 47476 5 1 1 47475
0 47477 7 1 2 57496 47476
0 47478 5 1 1 47477
0 47479 7 1 2 87152 91455
0 47480 7 1 2 81944 47479
0 47481 5 1 1 47480
0 47482 7 1 2 47478 47481
0 47483 5 1 1 47482
0 47484 7 1 2 67686 47483
0 47485 5 1 1 47484
0 47486 7 1 2 79864 85550
0 47487 7 1 2 93714 47486
0 47488 5 1 1 47487
0 47489 7 1 2 47485 47488
0 47490 5 1 1 47489
0 47491 7 1 2 61973 47490
0 47492 5 1 1 47491
0 47493 7 1 2 91755 93967
0 47494 5 1 1 47493
0 47495 7 1 2 47492 47494
0 47496 5 1 1 47495
0 47497 7 1 2 60163 47496
0 47498 5 1 1 47497
0 47499 7 1 2 84439 76929
0 47500 5 1 1 47499
0 47501 7 1 2 47500 95271
0 47502 5 1 1 47501
0 47503 7 1 2 60057 66988
0 47504 7 1 2 47502 47503
0 47505 5 1 1 47504
0 47506 7 1 2 47498 47505
0 47507 5 1 1 47506
0 47508 7 1 2 71530 47507
0 47509 5 1 1 47508
0 47510 7 1 2 60058 95260
0 47511 5 1 1 47510
0 47512 7 1 2 95306 95258
0 47513 5 1 1 47512
0 47514 7 1 2 47511 47513
0 47515 5 1 1 47514
0 47516 7 1 2 74347 47515
0 47517 5 1 1 47516
0 47518 7 3 2 66064 95308
0 47519 7 1 2 73233 95322
0 47520 5 1 1 47519
0 47521 7 1 2 47517 47520
0 47522 5 1 1 47521
0 47523 7 1 2 64838 47522
0 47524 5 1 1 47523
0 47525 7 1 2 91756 95192
0 47526 5 1 1 47525
0 47527 7 1 2 64839 88037
0 47528 5 1 1 47527
0 47529 7 1 2 47526 47528
0 47530 5 1 1 47529
0 47531 7 1 2 78896 47530
0 47532 5 1 1 47531
0 47533 7 1 2 73770 86111
0 47534 7 1 2 95066 47533
0 47535 7 1 2 71633 47534
0 47536 5 1 1 47535
0 47537 7 1 2 47532 47536
0 47538 7 1 2 47524 47537
0 47539 5 1 1 47538
0 47540 7 1 2 65715 47539
0 47541 5 1 1 47540
0 47542 7 1 2 74348 89397
0 47543 5 1 1 47542
0 47544 7 1 2 80439 92364
0 47545 7 1 2 69478 47544
0 47546 5 1 1 47545
0 47547 7 1 2 47543 47546
0 47548 5 1 1 47547
0 47549 7 1 2 67687 47548
0 47550 5 1 1 47549
0 47551 7 2 2 80770 92195
0 47552 5 1 1 95325
0 47553 7 1 2 76031 95326
0 47554 5 1 1 47553
0 47555 7 1 2 90249 92365
0 47556 5 1 1 47555
0 47557 7 1 2 47554 47556
0 47558 7 1 2 47550 47557
0 47559 5 1 1 47558
0 47560 7 1 2 63534 47559
0 47561 5 1 1 47560
0 47562 7 1 2 65087 89297
0 47563 7 1 2 94344 47562
0 47564 5 1 1 47563
0 47565 7 1 2 47552 47564
0 47566 5 1 1 47565
0 47567 7 1 2 64740 47566
0 47568 5 1 1 47567
0 47569 7 1 2 84015 90250
0 47570 5 1 1 47569
0 47571 7 1 2 47568 47570
0 47572 5 1 1 47571
0 47573 7 1 2 82352 47572
0 47574 5 1 1 47573
0 47575 7 1 2 47561 47574
0 47576 7 1 2 47541 47575
0 47577 5 1 1 47576
0 47578 7 1 2 66628 47577
0 47579 5 1 1 47578
0 47580 7 1 2 78735 92403
0 47581 5 1 1 47580
0 47582 7 1 2 93941 47581
0 47583 5 1 1 47582
0 47584 7 1 2 76304 47583
0 47585 5 1 1 47584
0 47586 7 1 2 47464 47585
0 47587 5 1 1 47586
0 47588 7 1 2 67069 47587
0 47589 5 1 1 47588
0 47590 7 1 2 68795 77314
0 47591 5 1 1 47590
0 47592 7 1 2 65716 81220
0 47593 7 1 2 47591 47592
0 47594 5 1 1 47593
0 47595 7 1 2 84016 79521
0 47596 7 1 2 91779 47595
0 47597 7 1 2 80096 47596
0 47598 7 1 2 47594 47597
0 47599 5 1 1 47598
0 47600 7 1 2 47589 47599
0 47601 5 1 1 47600
0 47602 7 1 2 47601 95263
0 47603 5 1 1 47602
0 47604 7 1 2 59927 94693
0 47605 5 1 1 47604
0 47606 7 1 2 87526 92866
0 47607 5 1 1 47606
0 47608 7 1 2 47605 47607
0 47609 5 1 1 47608
0 47610 7 1 2 82970 47609
0 47611 5 1 1 47610
0 47612 7 1 2 63107 85785
0 47613 5 2 1 47612
0 47614 7 1 2 78827 73843
0 47615 7 1 2 95327 47614
0 47616 5 1 1 47615
0 47617 7 1 2 47611 47616
0 47618 5 1 1 47617
0 47619 7 1 2 66935 47618
0 47620 5 1 1 47619
0 47621 7 1 2 73737 77221
0 47622 7 1 2 68903 94225
0 47623 7 1 2 47621 47622
0 47624 5 1 1 47623
0 47625 7 1 2 76469 77402
0 47626 7 2 2 95328 47625
0 47627 5 1 1 95329
0 47628 7 1 2 72395 95330
0 47629 5 1 1 47628
0 47630 7 1 2 79001 47629
0 47631 5 1 1 47630
0 47632 7 1 2 82644 83638
0 47633 7 1 2 47631 47632
0 47634 5 1 1 47633
0 47635 7 1 2 47624 47634
0 47636 7 1 2 47620 47635
0 47637 5 1 1 47636
0 47638 7 1 2 67070 47637
0 47639 5 1 1 47638
0 47640 7 1 2 47603 47639
0 47641 7 1 2 47579 47640
0 47642 7 1 2 47509 47641
0 47643 5 1 1 47642
0 47644 7 1 2 62116 47643
0 47645 5 1 1 47644
0 47646 7 1 2 92512 95185
0 47647 7 1 2 93732 47646
0 47648 5 1 1 47647
0 47649 7 1 2 69467 73266
0 47650 5 1 1 47649
0 47651 7 5 2 57784 61454
0 47652 7 1 2 65717 95331
0 47653 7 1 2 87376 47652
0 47654 5 1 1 47653
0 47655 7 1 2 47650 47654
0 47656 5 1 1 47655
0 47657 7 1 2 57497 47656
0 47658 5 1 1 47657
0 47659 7 1 2 67688 73267
0 47660 5 1 1 47659
0 47661 7 1 2 86194 47660
0 47662 7 1 2 47658 47661
0 47663 5 1 1 47662
0 47664 7 1 2 79479 71085
0 47665 7 1 2 47663 47664
0 47666 5 1 1 47665
0 47667 7 1 2 47648 47666
0 47668 7 1 2 47645 47667
0 47669 5 1 1 47668
0 47670 7 1 2 61710 47669
0 47671 5 1 1 47670
0 47672 7 1 2 73552 82787
0 47673 5 1 1 47672
0 47674 7 1 2 63535 76707
0 47675 5 2 1 47674
0 47676 7 1 2 67689 70309
0 47677 7 1 2 95336 47676
0 47678 5 1 1 47677
0 47679 7 1 2 47673 47678
0 47680 5 1 1 47679
0 47681 7 2 2 71531 86572
0 47682 7 1 2 47680 95338
0 47683 5 1 1 47682
0 47684 7 1 2 57498 91830
0 47685 7 1 2 91900 47684
0 47686 5 1 1 47685
0 47687 7 1 2 47683 47686
0 47688 5 1 1 47687
0 47689 7 1 2 69339 47688
0 47690 5 1 1 47689
0 47691 7 1 2 79987 95202
0 47692 5 1 1 47691
0 47693 7 1 2 58658 69340
0 47694 7 1 2 87506 82533
0 47695 7 1 2 47693 47694
0 47696 5 1 1 47695
0 47697 7 1 2 47692 47696
0 47698 5 2 1 47697
0 47699 7 1 2 79388 95340
0 47700 5 1 1 47699
0 47701 7 1 2 74098 71349
0 47702 7 1 2 88926 47701
0 47703 7 1 2 85509 86249
0 47704 7 1 2 47702 47703
0 47705 5 1 1 47704
0 47706 7 1 2 47700 47705
0 47707 5 1 1 47706
0 47708 7 1 2 63536 47707
0 47709 5 1 1 47708
0 47710 7 1 2 47690 47709
0 47711 5 1 1 47710
0 47712 7 1 2 61974 47711
0 47713 5 1 1 47712
0 47714 7 1 2 79564 92031
0 47715 5 2 1 47714
0 47716 7 2 2 71532 73326
0 47717 5 1 1 95344
0 47718 7 1 2 95342 95345
0 47719 5 1 1 47718
0 47720 7 1 2 58799 80983
0 47721 5 1 1 47720
0 47722 7 1 2 93309 47721
0 47723 5 1 1 47722
0 47724 7 1 2 74224 80440
0 47725 7 1 2 47723 47724
0 47726 5 1 1 47725
0 47727 7 1 2 47719 47726
0 47728 5 1 1 47727
0 47729 7 1 2 82714 47728
0 47730 5 1 1 47729
0 47731 7 1 2 92024 94994
0 47732 5 1 1 47731
0 47733 7 1 2 47730 47732
0 47734 5 1 1 47733
0 47735 7 1 2 67690 67483
0 47736 7 1 2 47734 47735
0 47737 5 1 1 47736
0 47738 7 1 2 47713 47737
0 47739 5 1 1 47738
0 47740 7 1 2 64741 47739
0 47741 5 1 1 47740
0 47742 7 2 2 82582 67071
0 47743 5 2 1 95346
0 47744 7 2 2 87206 66989
0 47745 5 1 1 95350
0 47746 7 1 2 67691 95351
0 47747 5 1 1 47746
0 47748 7 1 2 95348 47747
0 47749 5 1 1 47748
0 47750 7 1 2 58659 47749
0 47751 5 1 1 47750
0 47752 7 2 2 61455 85436
0 47753 5 1 1 95352
0 47754 7 1 2 86631 94196
0 47755 7 1 2 95353 47754
0 47756 5 1 1 47755
0 47757 7 1 2 47751 47756
0 47758 5 1 1 47757
0 47759 7 1 2 74225 47758
0 47760 5 1 1 47759
0 47761 7 1 2 67692 87790
0 47762 5 1 1 47761
0 47763 7 1 2 22185 47762
0 47764 5 1 1 47763
0 47765 7 6 2 66065 71533
0 47766 5 1 1 95354
0 47767 7 1 2 67072 95355
0 47768 7 1 2 47764 47767
0 47769 5 1 1 47768
0 47770 7 1 2 47760 47769
0 47771 5 1 1 47770
0 47772 7 1 2 63537 47771
0 47773 5 1 1 47772
0 47774 7 3 2 76859 83038
0 47775 5 1 1 95360
0 47776 7 1 2 61087 95361
0 47777 5 1 1 47776
0 47778 7 1 2 82 47777
0 47779 5 1 1 47778
0 47780 7 1 2 95264 95005
0 47781 7 1 2 47779 47780
0 47782 5 1 1 47781
0 47783 7 1 2 67091 47775
0 47784 5 1 1 47783
0 47785 7 1 2 81985 95339
0 47786 7 1 2 47784 47785
0 47787 5 1 1 47786
0 47788 7 1 2 47782 47787
0 47789 5 1 1 47788
0 47790 7 1 2 64629 47789
0 47791 5 1 1 47790
0 47792 7 1 2 47773 47791
0 47793 5 1 1 47792
0 47794 7 1 2 74797 47793
0 47795 5 1 1 47794
0 47796 7 1 2 47741 47795
0 47797 5 1 1 47796
0 47798 7 1 2 71749 47797
0 47799 5 1 1 47798
0 47800 7 1 2 75219 66990
0 47801 5 1 1 47800
0 47802 7 2 2 59022 72502
0 47803 5 1 1 95363
0 47804 7 1 2 65325 95364
0 47805 5 1 1 47804
0 47806 7 1 2 47801 47805
0 47807 5 1 1 47806
0 47808 7 1 2 57499 47807
0 47809 5 1 1 47808
0 47810 7 1 2 70102 66991
0 47811 5 1 1 47810
0 47812 7 1 2 47803 47811
0 47813 5 1 1 47812
0 47814 7 1 2 65718 47813
0 47815 5 1 1 47814
0 47816 7 1 2 47809 47815
0 47817 5 1 1 47816
0 47818 7 1 2 87687 47817
0 47819 5 1 1 47818
0 47820 7 2 2 57785 88882
0 47821 7 1 2 69130 95365
0 47822 7 1 2 77326 47821
0 47823 5 1 1 47822
0 47824 7 1 2 47819 47823
0 47825 5 1 1 47824
0 47826 7 1 2 71534 47825
0 47827 5 1 1 47826
0 47828 7 1 2 82836 93571
0 47829 5 1 1 47828
0 47830 7 1 2 85786 3094
0 47831 5 1 1 47830
0 47832 7 1 2 67693 47831
0 47833 5 1 1 47832
0 47834 7 1 2 47146 47833
0 47835 5 1 1 47834
0 47836 7 1 2 75664 47835
0 47837 5 1 1 47836
0 47838 7 1 2 47829 47837
0 47839 5 1 1 47838
0 47840 7 1 2 59668 47839
0 47841 5 1 1 47840
0 47842 7 1 2 76004 7291
0 47843 5 1 1 47842
0 47844 7 1 2 78993 83444
0 47845 7 1 2 47843 47844
0 47846 5 1 1 47845
0 47847 7 1 2 47841 47846
0 47848 5 1 1 47847
0 47849 7 1 2 64840 47848
0 47850 5 1 1 47849
0 47851 7 1 2 47827 47850
0 47852 5 1 1 47851
0 47853 7 1 2 76660 47852
0 47854 5 1 1 47853
0 47855 7 1 2 66953 87169
0 47856 5 4 1 47855
0 47857 7 1 2 69010 86030
0 47858 5 1 1 47857
0 47859 7 1 2 15628 47858
0 47860 5 2 1 47859
0 47861 7 1 2 67694 95371
0 47862 5 1 1 47861
0 47863 7 1 2 84618 81698
0 47864 5 1 1 47863
0 47865 7 1 2 47862 47864
0 47866 5 1 1 47865
0 47867 7 1 2 57500 47866
0 47868 5 1 1 47867
0 47869 7 1 2 74923 47868
0 47870 5 1 1 47869
0 47871 7 1 2 67073 47870
0 47872 5 1 1 47871
0 47873 7 1 2 67695 80084
0 47874 5 1 1 47873
0 47875 7 1 2 85236 47874
0 47876 5 1 1 47875
0 47877 7 1 2 59669 91780
0 47878 7 1 2 47876 47877
0 47879 5 1 1 47878
0 47880 7 1 2 47872 47879
0 47881 5 1 1 47880
0 47882 7 1 2 58352 47881
0 47883 5 1 1 47882
0 47884 7 1 2 74008 95071
0 47885 7 1 2 95372 47884
0 47886 5 1 1 47885
0 47887 7 1 2 47883 47886
0 47888 5 1 1 47887
0 47889 7 1 2 95367 47888
0 47890 5 1 1 47889
0 47891 7 1 2 68638 94232
0 47892 5 1 1 47891
0 47893 7 1 2 39861 47892
0 47894 5 1 1 47893
0 47895 7 1 2 74349 47894
0 47896 5 1 1 47895
0 47897 7 1 2 72363 93915
0 47898 7 1 2 95356 47897
0 47899 5 1 1 47898
0 47900 7 1 2 47896 47899
0 47901 5 1 1 47900
0 47902 7 1 2 65719 47901
0 47903 5 1 1 47902
0 47904 7 1 2 64409 86891
0 47905 5 1 1 47904
0 47906 7 1 2 77237 47905
0 47907 5 1 1 47906
0 47908 7 1 2 59928 87744
0 47909 5 1 1 47908
0 47910 7 1 2 77834 47909
0 47911 7 1 2 47907 47910
0 47912 5 1 1 47911
0 47913 7 1 2 66066 47912
0 47914 5 1 1 47913
0 47915 7 1 2 47903 47914
0 47916 5 1 1 47915
0 47917 7 1 2 66992 47916
0 47918 5 1 1 47917
0 47919 7 1 2 72506 26164
0 47920 5 1 1 47919
0 47921 7 1 2 76541 47920
0 47922 5 1 1 47921
0 47923 7 1 2 80085 95362
0 47924 5 1 1 47923
0 47925 7 1 2 67088 21166
0 47926 5 1 1 47925
0 47927 7 1 2 71535 47926
0 47928 5 1 1 47927
0 47929 7 1 2 47924 47928
0 47930 7 1 2 47922 47929
0 47931 5 1 1 47930
0 47932 7 1 2 61456 47931
0 47933 5 1 1 47932
0 47934 7 1 2 73533 67074
0 47935 5 1 1 47934
0 47936 7 1 2 47933 47935
0 47937 5 1 1 47936
0 47938 7 1 2 75592 47937
0 47939 5 1 1 47938
0 47940 7 1 2 78381 73515
0 47941 7 1 2 72503 93712
0 47942 7 1 2 47940 47941
0 47943 5 1 1 47942
0 47944 7 1 2 47939 47943
0 47945 7 1 2 47918 47944
0 47946 5 1 1 47945
0 47947 7 1 2 66936 47946
0 47948 5 1 1 47947
0 47949 7 1 2 47890 47948
0 47950 7 1 2 47854 47949
0 47951 5 1 1 47950
0 47952 7 1 2 66359 47951
0 47953 5 1 1 47952
0 47954 7 2 2 72707 88883
0 47955 7 1 2 81794 93851
0 47956 7 1 2 95373 47955
0 47957 7 1 2 94670 47956
0 47958 5 1 1 47957
0 47959 7 1 2 47953 47958
0 47960 5 1 1 47959
0 47961 7 1 2 62117 47960
0 47962 5 1 1 47961
0 47963 7 1 2 47799 47962
0 47964 7 1 2 47671 47963
0 47965 5 1 1 47964
0 47966 7 1 2 58886 47965
0 47967 5 1 1 47966
0 47968 7 1 2 47462 47967
0 47969 7 1 2 47383 47968
0 47970 5 1 1 47969
0 47971 7 1 2 88300 47970
0 47972 5 1 1 47971
0 47973 7 1 2 64630 83889
0 47974 5 1 1 47973
0 47975 7 1 2 94079 47974
0 47976 5 1 1 47975
0 47977 7 1 2 67075 47976
0 47978 5 1 1 47977
0 47979 7 1 2 60676 75266
0 47980 5 2 1 47979
0 47981 7 1 2 66993 81986
0 47982 7 1 2 95375 47981
0 47983 5 1 1 47982
0 47984 7 1 2 47978 47983
0 47985 5 1 1 47984
0 47986 7 1 2 60059 47985
0 47987 5 1 1 47986
0 47988 7 1 2 71363 72426
0 47989 5 1 1 47988
0 47990 7 1 2 92652 47989
0 47991 5 1 1 47990
0 47992 7 1 2 57501 47991
0 47993 5 1 1 47992
0 47994 7 1 2 65720 67115
0 47995 5 1 1 47994
0 47996 7 1 2 83260 67076
0 47997 5 1 1 47996
0 47998 7 1 2 47995 47997
0 47999 7 1 2 47993 47998
0 48000 5 1 1 47999
0 48001 7 1 2 79435 48000
0 48002 5 1 1 48001
0 48003 7 1 2 47987 48002
0 48004 5 1 1 48003
0 48005 7 1 2 58887 48004
0 48006 5 1 1 48005
0 48007 7 2 2 68796 79865
0 48008 5 1 1 95377
0 48009 7 1 2 66937 70887
0 48010 5 1 1 48009
0 48011 7 1 2 48008 48010
0 48012 5 1 1 48011
0 48013 7 1 2 72613 48012
0 48014 5 1 1 48013
0 48015 7 1 2 48006 48014
0 48016 5 1 1 48015
0 48017 7 1 2 62118 48016
0 48018 5 1 1 48017
0 48019 7 2 2 79910 67537
0 48020 7 1 2 68797 69556
0 48021 7 1 2 86241 48020
0 48022 7 1 2 95379 48021
0 48023 5 1 1 48022
0 48024 7 1 2 48018 48023
0 48025 5 1 1 48024
0 48026 7 1 2 86502 48025
0 48027 5 1 1 48026
0 48028 7 2 2 74383 80499
0 48029 7 1 2 86092 95381
0 48030 7 1 2 95190 48029
0 48031 5 1 1 48030
0 48032 7 1 2 48027 48031
0 48033 5 1 1 48032
0 48034 7 1 2 71536 48033
0 48035 5 1 1 48034
0 48036 7 1 2 78944 93573
0 48037 5 1 1 48036
0 48038 7 2 2 58800 86333
0 48039 5 3 1 95383
0 48040 7 1 2 63538 22270
0 48041 7 1 2 38068 48040
0 48042 5 1 1 48041
0 48043 7 1 2 95385 48042
0 48044 5 1 1 48043
0 48045 7 1 2 48037 48044
0 48046 5 1 1 48045
0 48047 7 1 2 81699 92588
0 48048 5 1 1 48047
0 48049 7 1 2 87562 48048
0 48050 5 1 1 48049
0 48051 7 1 2 63539 48050
0 48052 5 1 1 48051
0 48053 7 1 2 95386 48052
0 48054 5 1 1 48053
0 48055 7 1 2 58353 48054
0 48056 5 1 1 48055
0 48057 7 1 2 48046 48056
0 48058 5 1 1 48057
0 48059 7 1 2 72568 48058
0 48060 5 1 1 48059
0 48061 7 1 2 72496 10256
0 48062 5 1 1 48061
0 48063 7 1 2 92103 48062
0 48064 5 1 1 48063
0 48065 7 1 2 66067 83418
0 48066 5 1 1 48065
0 48067 7 1 2 86627 48066
0 48068 5 1 1 48067
0 48069 7 1 2 58354 48068
0 48070 5 1 1 48069
0 48071 7 1 2 69824 86043
0 48072 5 1 1 48071
0 48073 7 1 2 48070 48072
0 48074 5 1 1 48073
0 48075 7 1 2 59023 48074
0 48076 5 1 1 48075
0 48077 7 1 2 73567 83063
0 48078 5 1 1 48077
0 48079 7 1 2 48076 48078
0 48080 5 1 1 48079
0 48081 7 1 2 57502 48080
0 48082 5 1 1 48081
0 48083 7 1 2 65326 83419
0 48084 7 1 2 95357 48083
0 48085 5 1 1 48084
0 48086 7 1 2 48082 48085
0 48087 5 1 1 48086
0 48088 7 1 2 91541 48087
0 48089 5 1 1 48088
0 48090 7 1 2 48064 48089
0 48091 5 1 1 48090
0 48092 7 1 2 66629 48091
0 48093 5 1 1 48092
0 48094 7 1 2 73764 92589
0 48095 5 1 1 48094
0 48096 7 1 2 87563 48095
0 48097 5 1 1 48096
0 48098 7 1 2 63540 48097
0 48099 5 1 1 48098
0 48100 7 1 2 84955 94980
0 48101 5 1 1 48100
0 48102 7 1 2 88278 48101
0 48103 5 1 1 48102
0 48104 7 1 2 64742 48103
0 48105 5 1 1 48104
0 48106 7 1 2 48099 48105
0 48107 5 1 1 48106
0 48108 7 1 2 72582 48107
0 48109 5 1 1 48108
0 48110 7 2 2 75687 90263
0 48111 7 2 2 94382 95388
0 48112 7 1 2 65327 95390
0 48113 5 1 1 48112
0 48114 7 1 2 48109 48113
0 48115 5 1 1 48114
0 48116 7 1 2 68639 48115
0 48117 5 1 1 48116
0 48118 7 1 2 85917 95391
0 48119 5 1 1 48118
0 48120 7 1 2 48117 48119
0 48121 7 1 2 48093 48120
0 48122 5 1 1 48121
0 48123 7 1 2 70530 48122
0 48124 5 1 1 48123
0 48125 7 2 2 66630 76470
0 48126 7 2 2 83519 95392
0 48127 7 1 2 72427 95394
0 48128 5 1 1 48127
0 48129 7 1 2 76512 82672
0 48130 5 1 1 48129
0 48131 7 1 2 48128 48130
0 48132 5 1 1 48131
0 48133 7 1 2 65328 48132
0 48134 5 1 1 48133
0 48135 7 2 2 67077 81881
0 48136 7 1 2 68798 86408
0 48137 5 1 1 48136
0 48138 7 1 2 7542 48137
0 48139 5 1 1 48138
0 48140 7 1 2 95396 48139
0 48141 5 1 1 48140
0 48142 7 1 2 48134 48141
0 48143 5 1 1 48142
0 48144 7 1 2 71537 48143
0 48145 5 1 1 48144
0 48146 7 1 2 59670 72583
0 48147 7 1 2 82069 48146
0 48148 7 1 2 70890 48147
0 48149 5 1 1 48148
0 48150 7 1 2 48145 48149
0 48151 5 1 1 48150
0 48152 7 1 2 66068 48151
0 48153 5 1 1 48152
0 48154 7 1 2 65329 92225
0 48155 5 1 1 48154
0 48156 7 1 2 76032 72584
0 48157 7 1 2 83610 48156
0 48158 5 1 1 48157
0 48159 7 1 2 48155 48158
0 48160 5 1 1 48159
0 48161 7 1 2 76471 48160
0 48162 5 1 1 48161
0 48163 7 1 2 61088 70892
0 48164 5 1 1 48163
0 48165 7 1 2 92226 48164
0 48166 5 1 1 48165
0 48167 7 1 2 48162 48166
0 48168 5 1 1 48167
0 48169 7 1 2 71220 48168
0 48170 5 1 1 48169
0 48171 7 1 2 48153 48170
0 48172 5 1 1 48171
0 48173 7 1 2 66360 48172
0 48174 5 1 1 48173
0 48175 7 1 2 81962 72603
0 48176 7 1 2 92104 48175
0 48177 5 1 1 48176
0 48178 7 1 2 48174 48177
0 48179 7 1 2 48124 48178
0 48180 5 1 1 48179
0 48181 7 1 2 62119 48180
0 48182 5 1 1 48181
0 48183 7 1 2 48060 48182
0 48184 5 1 1 48183
0 48185 7 1 2 59929 48184
0 48186 5 1 1 48185
0 48187 7 1 2 79440 24476
0 48188 5 2 1 48187
0 48189 7 1 2 58355 95398
0 48190 5 1 1 48189
0 48191 7 1 2 60418 82791
0 48192 5 2 1 48191
0 48193 7 1 2 87819 95400
0 48194 5 1 1 48193
0 48195 7 1 2 48190 48194
0 48196 5 1 1 48195
0 48197 7 1 2 82389 48196
0 48198 5 1 1 48197
0 48199 7 2 2 74384 76472
0 48200 7 1 2 79911 84681
0 48201 7 1 2 95402 48200
0 48202 5 1 1 48201
0 48203 7 1 2 48198 48202
0 48204 5 1 1 48203
0 48205 7 1 2 59024 48204
0 48206 5 1 1 48205
0 48207 7 1 2 3919 47190
0 48208 5 1 1 48207
0 48209 7 1 2 86305 48208
0 48210 5 1 1 48209
0 48211 7 1 2 65330 95399
0 48212 5 1 1 48211
0 48213 7 3 2 60419 78953
0 48214 7 1 2 84017 95404
0 48215 5 1 1 48214
0 48216 7 1 2 48212 48215
0 48217 5 1 1 48216
0 48218 7 1 2 84067 48217
0 48219 5 1 1 48218
0 48220 7 1 2 48210 48219
0 48221 7 1 2 48206 48220
0 48222 5 1 1 48221
0 48223 7 1 2 65721 48222
0 48224 5 1 1 48223
0 48225 7 1 2 61457 92610
0 48226 5 1 1 48225
0 48227 7 1 2 79441 48226
0 48228 5 1 1 48227
0 48229 7 2 2 61711 48228
0 48230 7 1 2 59025 95300
0 48231 7 1 2 95407 48230
0 48232 5 1 1 48231
0 48233 7 1 2 48224 48232
0 48234 5 1 1 48233
0 48235 7 1 2 70577 48234
0 48236 5 1 1 48235
0 48237 7 1 2 80534 86306
0 48238 5 1 1 48237
0 48239 7 1 2 71221 95246
0 48240 7 1 2 81963 48239
0 48241 5 1 1 48240
0 48242 7 1 2 48238 48241
0 48243 5 1 1 48242
0 48244 7 1 2 61458 48243
0 48245 5 1 1 48244
0 48246 7 1 2 73574 47627
0 48247 5 1 1 48246
0 48248 7 1 2 92143 92733
0 48249 7 1 2 48247 48248
0 48250 5 1 1 48249
0 48251 7 1 2 48245 48250
0 48252 5 1 1 48251
0 48253 7 1 2 72604 48252
0 48254 5 1 1 48253
0 48255 7 1 2 48236 48254
0 48256 5 1 1 48255
0 48257 7 1 2 62120 48256
0 48258 5 1 1 48257
0 48259 7 1 2 82222 82400
0 48260 5 1 1 48259
0 48261 7 1 2 86093 67538
0 48262 7 1 2 48260 48261
0 48263 7 1 2 94374 48262
0 48264 5 1 1 48263
0 48265 7 1 2 48258 48264
0 48266 7 1 2 48186 48265
0 48267 7 1 2 48035 48266
0 48268 5 1 1 48267
0 48269 7 1 2 58660 48268
0 48270 5 1 1 48269
0 48271 7 1 2 64410 74312
0 48272 5 1 1 48271
0 48273 7 1 2 61089 74282
0 48274 5 1 1 48273
0 48275 7 1 2 48272 48274
0 48276 5 1 1 48275
0 48277 7 1 2 78828 48276
0 48278 5 1 1 48277
0 48279 7 1 2 67484 79460
0 48280 7 1 2 82366 48279
0 48281 5 1 1 48280
0 48282 7 1 2 48278 48281
0 48283 5 1 1 48282
0 48284 7 1 2 65088 48283
0 48285 5 1 1 48284
0 48286 7 1 2 71538 88842
0 48287 5 1 1 48286
0 48288 7 1 2 48285 48287
0 48289 5 1 1 48288
0 48290 7 1 2 61459 48289
0 48291 5 1 1 48290
0 48292 7 1 2 73268 67539
0 48293 7 1 2 83015 48292
0 48294 5 1 1 48293
0 48295 7 1 2 76907 93105
0 48296 7 1 2 74283 48295
0 48297 5 1 1 48296
0 48298 7 1 2 48294 48297
0 48299 5 1 1 48298
0 48300 7 1 2 80500 48299
0 48301 5 1 1 48300
0 48302 7 1 2 48291 48301
0 48303 5 1 1 48302
0 48304 7 1 2 64631 48303
0 48305 5 1 1 48304
0 48306 7 1 2 59026 90197
0 48307 5 1 1 48306
0 48308 7 1 2 47717 48307
0 48309 5 1 1 48308
0 48310 7 1 2 70876 48309
0 48311 5 1 1 48310
0 48312 7 1 2 59027 76473
0 48313 5 1 1 48312
0 48314 7 1 2 60677 48313
0 48315 5 1 1 48314
0 48316 7 1 2 61460 70069
0 48317 5 2 1 48316
0 48318 7 1 2 74136 95409
0 48319 7 1 2 48315 48318
0 48320 5 1 1 48319
0 48321 7 1 2 48311 48320
0 48322 5 1 1 48321
0 48323 7 1 2 67485 92156
0 48324 7 1 2 48322 48323
0 48325 5 1 1 48324
0 48326 7 1 2 48305 48325
0 48327 5 1 1 48326
0 48328 7 1 2 70531 48327
0 48329 5 1 1 48328
0 48330 7 1 2 72155 69679
0 48331 5 1 1 48330
0 48332 7 1 2 78936 69274
0 48333 5 1 1 48332
0 48334 7 1 2 48331 48333
0 48335 5 1 1 48334
0 48336 7 1 2 68799 48335
0 48337 5 1 1 48336
0 48338 7 1 2 3068 72124
0 48339 5 1 1 48338
0 48340 7 1 2 64411 48339
0 48341 5 1 1 48340
0 48342 7 1 2 48337 48341
0 48343 5 1 1 48342
0 48344 7 1 2 77275 48343
0 48345 5 1 1 48344
0 48346 7 1 2 68640 69680
0 48347 5 1 1 48346
0 48348 7 1 2 83290 74099
0 48349 7 1 2 69579 48348
0 48350 5 1 1 48349
0 48351 7 1 2 48347 48350
0 48352 5 1 1 48351
0 48353 7 1 2 75665 48352
0 48354 5 1 1 48353
0 48355 7 1 2 48345 48354
0 48356 5 1 1 48355
0 48357 7 1 2 61461 48356
0 48358 5 1 1 48357
0 48359 7 2 2 66069 67540
0 48360 7 2 2 76111 79854
0 48361 5 1 1 95413
0 48362 7 1 2 71961 95414
0 48363 7 1 2 95411 48362
0 48364 5 1 1 48363
0 48365 7 1 2 64632 48364
0 48366 7 1 2 48358 48365
0 48367 5 1 1 48366
0 48368 7 5 2 67936 90546
0 48369 5 1 1 95415
0 48370 7 1 2 71626 95416
0 48371 5 1 1 48370
0 48372 7 1 2 85234 79002
0 48373 5 1 1 48372
0 48374 7 1 2 2665 69580
0 48375 7 1 2 48373 48374
0 48376 5 1 1 48375
0 48377 7 1 2 48371 48376
0 48378 5 1 1 48377
0 48379 7 1 2 59671 48378
0 48380 5 1 1 48379
0 48381 7 1 2 69248 80546
0 48382 7 1 2 92668 48381
0 48383 5 1 1 48382
0 48384 7 1 2 48380 48383
0 48385 5 1 1 48384
0 48386 7 1 2 88846 48385
0 48387 5 1 1 48386
0 48388 7 1 2 59930 48387
0 48389 5 1 1 48388
0 48390 7 1 2 65089 48389
0 48391 7 1 2 48367 48390
0 48392 5 1 1 48391
0 48393 7 1 2 75739 80885
0 48394 5 1 1 48393
0 48395 7 1 2 87611 77372
0 48396 7 1 2 82036 48395
0 48397 5 1 1 48396
0 48398 7 1 2 48394 48397
0 48399 5 1 1 48398
0 48400 7 1 2 63541 48399
0 48401 5 1 1 48400
0 48402 7 2 2 67960 94402
0 48403 7 1 2 81882 94039
0 48404 7 1 2 95420 48403
0 48405 5 1 1 48404
0 48406 7 1 2 48401 48405
0 48407 5 1 1 48406
0 48408 7 1 2 59672 48407
0 48409 5 1 1 48408
0 48410 7 2 2 75740 79943
0 48411 7 1 2 74690 79931
0 48412 7 1 2 80255 48411
0 48413 7 2 2 95422 48412
0 48414 5 1 1 95424
0 48415 7 1 2 48409 48414
0 48416 5 1 1 48415
0 48417 7 1 2 72618 48416
0 48418 5 1 1 48417
0 48419 7 1 2 67486 93106
0 48420 7 1 2 79207 48419
0 48421 5 1 1 48420
0 48422 7 1 2 71222 92157
0 48423 5 1 1 48422
0 48424 7 1 2 39869 48423
0 48425 5 1 1 48424
0 48426 7 1 2 69557 95412
0 48427 7 1 2 48425 48426
0 48428 5 1 1 48427
0 48429 7 1 2 48421 48428
0 48430 5 1 1 48429
0 48431 7 1 2 76908 48430
0 48432 5 1 1 48431
0 48433 7 1 2 71627 80034
0 48434 5 1 1 48433
0 48435 7 1 2 74737 76912
0 48436 5 1 1 48435
0 48437 7 1 2 48434 48436
0 48438 5 1 1 48437
0 48439 7 1 2 79572 48438
0 48440 5 1 1 48439
0 48441 7 1 2 76434 47351
0 48442 5 1 1 48441
0 48443 7 1 2 92158 95417
0 48444 7 1 2 48442 48443
0 48445 5 1 1 48444
0 48446 7 1 2 48440 48445
0 48447 5 1 1 48446
0 48448 7 1 2 61975 48447
0 48449 5 1 1 48448
0 48450 7 1 2 76474 72605
0 48451 5 1 1 48450
0 48452 7 1 2 72591 48451
0 48453 5 1 1 48452
0 48454 7 1 2 72419 92159
0 48455 7 1 2 48453 48454
0 48456 5 1 1 48455
0 48457 7 3 2 63542 79932
0 48458 7 1 2 73982 91107
0 48459 7 1 2 92045 48458
0 48460 7 1 2 95426 48459
0 48461 5 1 1 48460
0 48462 7 1 2 48456 48461
0 48463 5 1 1 48462
0 48464 7 1 2 95009 48463
0 48465 5 1 1 48464
0 48466 7 1 2 72877 95302
0 48467 5 1 1 48466
0 48468 7 1 2 93736 48467
0 48469 5 1 1 48468
0 48470 7 2 2 86674 82621
0 48471 7 1 2 69275 95429
0 48472 7 1 2 48469 48471
0 48473 5 1 1 48472
0 48474 7 1 2 48465 48473
0 48475 7 1 2 48449 48474
0 48476 7 1 2 48432 48475
0 48477 7 1 2 48418 48476
0 48478 7 1 2 48392 48477
0 48479 7 1 2 48329 48478
0 48480 5 1 1 48479
0 48481 7 1 2 61712 48480
0 48482 5 1 1 48481
0 48483 7 1 2 74738 95382
0 48484 5 1 1 48483
0 48485 7 1 2 76909 89791
0 48486 5 1 1 48485
0 48487 7 1 2 48484 48486
0 48488 5 1 1 48487
0 48489 7 1 2 61090 48488
0 48490 5 1 1 48489
0 48491 7 1 2 86031 79018
0 48492 5 1 1 48491
0 48493 7 1 2 86744 48492
0 48494 5 1 1 48493
0 48495 7 1 2 65090 48494
0 48496 5 1 1 48495
0 48497 7 1 2 48490 48496
0 48498 5 1 1 48497
0 48499 7 1 2 59931 48498
0 48500 5 1 1 48499
0 48501 7 1 2 79643 94375
0 48502 5 1 1 48501
0 48503 7 1 2 48500 48502
0 48504 5 1 1 48503
0 48505 7 1 2 69276 48504
0 48506 5 1 1 48505
0 48507 7 1 2 71539 90612
0 48508 5 1 1 48507
0 48509 7 2 2 71540 73516
0 48510 5 1 1 95431
0 48511 7 1 2 48508 48510
0 48512 7 1 2 47753 48511
0 48513 5 1 1 48512
0 48514 7 1 2 80535 68685
0 48515 7 1 2 48513 48514
0 48516 5 1 1 48515
0 48517 7 1 2 48506 48516
0 48518 5 1 1 48517
0 48519 7 1 2 61976 48518
0 48520 5 1 1 48519
0 48521 7 2 2 65331 78089
0 48522 5 1 1 95433
0 48523 7 1 2 85437 83222
0 48524 5 1 1 48523
0 48525 7 1 2 48522 48524
0 48526 5 1 1 48525
0 48527 7 1 2 61462 48526
0 48528 5 1 1 48527
0 48529 7 1 2 76454 81707
0 48530 5 1 1 48529
0 48531 7 1 2 95432 48530
0 48532 7 1 2 78413 48531
0 48533 5 1 1 48532
0 48534 7 1 2 48528 48533
0 48535 5 1 1 48534
0 48536 7 1 2 62121 72589
0 48537 7 1 2 48535 48536
0 48538 5 1 1 48537
0 48539 7 1 2 48520 48538
0 48540 5 1 1 48539
0 48541 7 1 2 86307 48540
0 48542 5 1 1 48541
0 48543 7 1 2 48482 48542
0 48544 7 1 2 48270 48543
0 48545 5 1 1 48544
0 48546 7 1 2 88301 48545
0 48547 5 1 1 48546
0 48548 7 2 2 84473 90716
0 48549 7 1 2 88519 95206
0 48550 7 2 2 95435 48549
0 48551 7 1 2 83657 95437
0 48552 7 1 2 85036 48551
0 48553 5 1 1 48552
0 48554 7 1 2 48547 48553
0 48555 5 1 1 48554
0 48556 7 1 2 68411 48555
0 48557 5 1 1 48556
0 48558 7 1 2 76513 92563
0 48559 5 1 1 48558
0 48560 7 1 2 79058 87634
0 48561 5 1 1 48560
0 48562 7 1 2 87648 95265
0 48563 7 1 2 48561 48562
0 48564 5 1 1 48563
0 48565 7 1 2 48559 48564
0 48566 5 1 1 48565
0 48567 7 1 2 61463 48566
0 48568 5 1 1 48567
0 48569 7 2 2 79391 81708
0 48570 5 1 1 95439
0 48571 7 1 2 780 95440
0 48572 5 1 1 48571
0 48573 7 1 2 95323 48572
0 48574 5 1 1 48573
0 48575 7 1 2 92168 48574
0 48576 5 1 1 48575
0 48577 7 1 2 61713 48576
0 48578 5 1 1 48577
0 48579 7 1 2 48568 48578
0 48580 5 1 1 48579
0 48581 7 1 2 60164 48580
0 48582 5 1 1 48581
0 48583 7 1 2 83926 91831
0 48584 7 1 2 94322 48583
0 48585 5 1 1 48584
0 48586 7 1 2 48582 48585
0 48587 5 1 1 48586
0 48588 7 1 2 58888 48587
0 48589 5 1 1 48588
0 48590 7 1 2 81044 83611
0 48591 7 1 2 94297 48590
0 48592 5 1 1 48591
0 48593 7 1 2 48589 48592
0 48594 5 1 1 48593
0 48595 7 1 2 62122 48594
0 48596 5 1 1 48595
0 48597 7 2 2 69558 90141
0 48598 5 1 1 95441
0 48599 7 1 2 87345 95442
0 48600 5 1 1 48599
0 48601 7 3 2 76514 84682
0 48602 5 1 1 95443
0 48603 7 1 2 69681 95444
0 48604 5 1 1 48603
0 48605 7 1 2 48600 48604
0 48606 5 1 1 48605
0 48607 7 1 2 95295 48606
0 48608 5 1 1 48607
0 48609 7 1 2 87564 87644
0 48610 5 1 1 48609
0 48611 7 2 2 63543 48610
0 48612 5 1 1 95446
0 48613 7 1 2 48612 95387
0 48614 5 1 1 48613
0 48615 7 2 2 92361 48614
0 48616 7 1 2 71223 80461
0 48617 7 1 2 95448 48616
0 48618 5 1 1 48617
0 48619 7 1 2 48608 48618
0 48620 7 1 2 48596 48619
0 48621 5 1 1 48620
0 48622 7 1 2 61977 48621
0 48623 5 1 1 48622
0 48624 7 1 2 95174 95395
0 48625 5 1 1 48624
0 48626 7 1 2 29475 48625
0 48627 5 1 1 48626
0 48628 7 1 2 91984 48627
0 48629 5 1 1 48628
0 48630 7 1 2 75688 94240
0 48631 5 1 1 48630
0 48632 7 1 2 83064 92734
0 48633 7 1 2 95393 48632
0 48634 5 1 1 48633
0 48635 7 1 2 48631 48634
0 48636 5 1 1 48635
0 48637 7 1 2 92041 48636
0 48638 5 1 1 48637
0 48639 7 3 2 63544 82419
0 48640 5 1 1 95450
0 48641 7 1 2 88279 48640
0 48642 5 1 1 48641
0 48643 7 1 2 71541 95397
0 48644 7 1 2 48642 48643
0 48645 5 1 1 48644
0 48646 7 1 2 48638 48645
0 48647 5 1 1 48646
0 48648 7 1 2 66070 48647
0 48649 5 1 1 48648
0 48650 7 1 2 48629 48649
0 48651 5 1 1 48650
0 48652 7 1 2 58661 48651
0 48653 5 1 1 48652
0 48654 7 1 2 82583 67621
0 48655 5 1 1 48654
0 48656 7 1 2 79203 88455
0 48657 5 1 1 48656
0 48658 7 1 2 48655 48657
0 48659 5 1 1 48658
0 48660 7 1 2 71542 48659
0 48661 5 1 1 48660
0 48662 7 1 2 65091 79389
0 48663 5 1 1 48662
0 48664 7 1 2 76475 81700
0 48665 5 1 1 48664
0 48666 7 1 2 48663 48665
0 48667 5 1 1 48666
0 48668 7 1 2 70578 91783
0 48669 7 1 2 48667 48668
0 48670 5 1 1 48669
0 48671 7 1 2 48661 48670
0 48672 5 1 1 48671
0 48673 7 1 2 66071 48672
0 48674 5 1 1 48673
0 48675 7 2 2 84683 72606
0 48676 5 1 1 95453
0 48677 7 1 2 80984 95454
0 48678 5 1 1 48677
0 48679 7 1 2 48674 48678
0 48680 5 1 1 48679
0 48681 7 1 2 66938 48680
0 48682 5 1 1 48681
0 48683 7 1 2 48653 48682
0 48684 5 1 1 48683
0 48685 7 1 2 62123 48684
0 48686 5 1 1 48685
0 48687 7 1 2 61714 95425
0 48688 5 1 1 48687
0 48689 7 4 2 61715 91108
0 48690 7 1 2 87925 95455
0 48691 5 1 1 48690
0 48692 7 2 2 75988 94841
0 48693 7 2 2 70532 72420
0 48694 7 1 2 95459 95461
0 48695 5 1 1 48694
0 48696 7 1 2 48691 48695
0 48697 5 1 1 48696
0 48698 7 1 2 72916 48697
0 48699 5 1 1 48698
0 48700 7 1 2 48688 48699
0 48701 7 1 2 48686 48700
0 48702 5 1 1 48701
0 48703 7 1 2 65332 48702
0 48704 5 1 1 48703
0 48705 7 1 2 83425 92349
0 48706 5 2 1 48705
0 48707 7 2 2 59028 70548
0 48708 7 1 2 81045 92144
0 48709 5 1 1 48708
0 48710 7 1 2 59932 95296
0 48711 5 1 1 48710
0 48712 7 1 2 48709 48711
0 48713 5 1 1 48712
0 48714 7 1 2 95465 48713
0 48715 5 1 1 48714
0 48716 7 1 2 95463 48715
0 48717 5 1 1 48716
0 48718 7 1 2 71364 84302
0 48719 7 1 2 48717 48718
0 48720 5 1 1 48719
0 48721 7 1 2 48704 48720
0 48722 7 1 2 48623 48721
0 48723 5 1 1 48722
0 48724 7 1 2 88302 48723
0 48725 5 1 1 48724
0 48726 7 1 2 87325 81701
0 48727 5 1 1 48726
0 48728 7 1 2 89394 48727
0 48729 5 1 1 48728
0 48730 7 1 2 57503 48729
0 48731 5 1 1 48730
0 48732 7 3 2 61716 82971
0 48733 5 2 1 95467
0 48734 7 1 2 89206 95468
0 48735 5 1 1 48734
0 48736 7 1 2 48731 48735
0 48737 5 1 1 48736
0 48738 7 1 2 79912 48737
0 48739 5 1 1 48738
0 48740 7 1 2 57504 94968
0 48741 5 1 1 48740
0 48742 7 1 2 61717 74764
0 48743 5 1 1 48742
0 48744 7 1 2 48741 48743
0 48745 5 1 1 48744
0 48746 7 1 2 82645 81702
0 48747 7 1 2 48745 48746
0 48748 5 1 1 48747
0 48749 7 1 2 48739 48748
0 48750 5 1 1 48749
0 48751 7 1 2 67110 48750
0 48752 5 1 1 48751
0 48753 7 1 2 86573 95279
0 48754 7 1 2 48570 48753
0 48755 5 1 1 48754
0 48756 7 1 2 48752 48755
0 48757 5 1 1 48756
0 48758 7 1 2 70533 48757
0 48759 5 1 1 48758
0 48760 7 2 2 87240 84474
0 48761 7 1 2 81711 95472
0 48762 7 1 2 93923 48761
0 48763 5 1 1 48762
0 48764 7 1 2 48759 48763
0 48765 5 1 1 48764
0 48766 7 1 2 94767 48765
0 48767 5 1 1 48766
0 48768 7 2 2 83562 92218
0 48769 7 1 2 68800 71224
0 48770 7 1 2 95436 48769
0 48771 7 1 2 95474 48770
0 48772 5 1 1 48771
0 48773 7 1 2 48767 48772
0 48774 5 1 1 48773
0 48775 7 1 2 83728 48774
0 48776 5 1 1 48775
0 48777 7 1 2 67937 83639
0 48778 7 1 2 79066 48777
0 48779 7 1 2 88380 93852
0 48780 7 1 2 95473 48779
0 48781 7 1 2 48778 48780
0 48782 5 1 1 48781
0 48783 7 1 2 48776 48782
0 48784 7 1 2 48725 48783
0 48785 5 1 1 48784
0 48786 7 1 2 79522 48785
0 48787 5 1 1 48786
0 48788 7 3 2 87487 91109
0 48789 7 1 2 67696 71225
0 48790 7 1 2 95476 48789
0 48791 7 1 2 95475 48790
0 48792 5 1 1 48791
0 48793 7 1 2 48787 48792
0 48794 7 1 2 48557 48793
0 48795 7 1 2 47972 48794
0 48796 5 1 1 48795
0 48797 7 1 2 67382 48796
0 48798 5 1 1 48797
0 48799 7 2 2 66792 94842
0 48800 5 2 1 95479
0 48801 7 1 2 82223 91789
0 48802 5 3 1 48801
0 48803 7 1 2 66939 95483
0 48804 5 1 1 48803
0 48805 7 1 2 95481 48804
0 48806 5 1 1 48805
0 48807 7 1 2 66072 48806
0 48808 5 1 1 48807
0 48809 7 1 2 95337 95405
0 48810 5 1 1 48809
0 48811 7 1 2 65092 95343
0 48812 5 1 1 48811
0 48813 7 1 2 48810 48812
0 48814 5 1 1 48813
0 48815 7 1 2 66361 48814
0 48816 5 1 1 48815
0 48817 7 1 2 75424 91784
0 48818 5 1 1 48817
0 48819 7 1 2 64743 48818
0 48820 7 1 2 48816 48819
0 48821 5 1 1 48820
0 48822 7 2 2 61718 77835
0 48823 5 1 1 95486
0 48824 7 3 2 58801 66362
0 48825 5 1 1 95488
0 48826 7 1 2 48825 95406
0 48827 7 1 2 48823 48826
0 48828 5 1 1 48827
0 48829 7 1 2 83420 95484
0 48830 5 1 1 48829
0 48831 7 1 2 60060 48830
0 48832 7 1 2 48828 48831
0 48833 5 1 1 48832
0 48834 7 1 2 59029 48833
0 48835 7 1 2 48821 48834
0 48836 5 1 1 48835
0 48837 7 1 2 58662 74503
0 48838 7 1 2 95288 48837
0 48839 5 1 1 48838
0 48840 7 1 2 48836 48839
0 48841 5 1 1 48840
0 48842 7 1 2 70354 48841
0 48843 5 1 1 48842
0 48844 7 1 2 48808 48843
0 48845 5 1 1 48844
0 48846 7 1 2 65333 48845
0 48847 5 1 1 48846
0 48848 7 1 2 63545 93718
0 48849 5 1 1 48848
0 48850 7 3 2 27113 48849
0 48851 7 1 2 68641 86574
0 48852 7 1 2 95491 48851
0 48853 5 1 1 48852
0 48854 7 1 2 84018 78494
0 48855 5 1 1 48854
0 48856 7 1 2 79442 48855
0 48857 5 1 1 48856
0 48858 7 1 2 58663 48857
0 48859 5 1 1 48858
0 48860 7 1 2 92162 48859
0 48861 5 1 1 48860
0 48862 7 5 2 57786 61719
0 48863 7 1 2 83291 95494
0 48864 7 1 2 48861 48863
0 48865 5 1 1 48864
0 48866 7 1 2 48853 48865
0 48867 5 1 1 48866
0 48868 7 1 2 65093 48867
0 48869 5 1 1 48868
0 48870 7 1 2 48847 48869
0 48871 5 1 1 48870
0 48872 7 1 2 59167 48871
0 48873 5 1 1 48872
0 48874 7 3 2 66073 80602
0 48875 7 2 2 66363 95492
0 48876 7 1 2 70936 95502
0 48877 5 1 1 48876
0 48878 7 2 2 79913 91785
0 48879 5 1 1 95504
0 48880 7 1 2 48877 48879
0 48881 5 1 1 48880
0 48882 7 1 2 95499 48881
0 48883 5 1 1 48882
0 48884 7 1 2 48873 48883
0 48885 5 1 1 48884
0 48886 7 1 2 66631 48885
0 48887 5 1 1 48886
0 48888 7 1 2 57505 40577
0 48889 5 1 1 48888
0 48890 7 1 2 61464 6290
0 48891 5 1 1 48890
0 48892 7 1 2 65722 48891
0 48893 5 1 1 48892
0 48894 7 1 2 94048 48893
0 48895 7 1 2 48889 48894
0 48896 5 1 1 48895
0 48897 7 1 2 95460 48896
0 48898 5 1 1 48897
0 48899 7 1 2 48887 48898
0 48900 5 1 1 48899
0 48901 7 1 2 70534 48900
0 48902 5 1 1 48901
0 48903 7 1 2 61465 93135
0 48904 5 1 1 48903
0 48905 7 1 2 94584 48904
0 48906 5 1 1 48905
0 48907 7 1 2 68642 86202
0 48908 7 1 2 94780 48907
0 48909 5 1 1 48908
0 48910 7 1 2 92278 48909
0 48911 7 1 2 48906 48910
0 48912 5 1 1 48911
0 48913 7 1 2 64633 48912
0 48914 5 1 1 48913
0 48915 7 1 2 63546 86197
0 48916 5 1 1 48915
0 48917 7 1 2 48914 48916
0 48918 5 1 1 48917
0 48919 7 1 2 60061 48918
0 48920 5 1 1 48919
0 48921 7 1 2 76476 92903
0 48922 5 1 1 48921
0 48923 7 1 2 61466 48922
0 48924 5 1 1 48923
0 48925 7 1 2 57787 48924
0 48926 5 1 1 48925
0 48927 7 1 2 71976 94446
0 48928 7 1 2 48926 48927
0 48929 5 2 1 48928
0 48930 7 1 2 79436 95506
0 48931 5 1 1 48930
0 48932 7 1 2 48920 48931
0 48933 5 1 1 48932
0 48934 7 1 2 58664 48933
0 48935 5 1 1 48934
0 48936 7 1 2 92160 95507
0 48937 5 1 1 48936
0 48938 7 1 2 48935 48937
0 48939 5 1 1 48938
0 48940 7 1 2 61720 48939
0 48941 5 1 1 48940
0 48942 7 1 2 57506 94460
0 48943 5 1 1 48942
0 48944 7 1 2 94051 48943
0 48945 5 1 1 48944
0 48946 7 1 2 66364 72963
0 48947 7 1 2 95368 48946
0 48948 7 1 2 48945 48947
0 48949 5 1 1 48948
0 48950 7 1 2 48941 48949
0 48951 5 1 1 48950
0 48952 7 1 2 72607 48951
0 48953 5 1 1 48952
0 48954 7 1 2 57788 72414
0 48955 5 1 1 48954
0 48956 7 1 2 85787 48955
0 48957 5 1 1 48956
0 48958 7 1 2 57507 48957
0 48959 5 1 1 48958
0 48960 7 1 2 61467 527
0 48961 5 2 1 48960
0 48962 7 1 2 69468 88072
0 48963 7 1 2 95508 48962
0 48964 5 1 1 48963
0 48965 7 1 2 48959 48964
0 48966 5 1 1 48965
0 48967 7 1 2 59168 48966
0 48968 5 1 1 48967
0 48969 7 1 2 70937 95500
0 48970 5 1 1 48969
0 48971 7 1 2 48968 48970
0 48972 5 1 1 48971
0 48973 7 1 2 86615 93924
0 48974 7 1 2 48972 48973
0 48975 5 1 1 48974
0 48976 7 1 2 48953 48975
0 48977 7 1 2 48902 48976
0 48978 5 1 1 48977
0 48979 7 1 2 62124 48978
0 48980 5 1 1 48979
0 48981 7 1 2 87667 80886
0 48982 5 1 1 48981
0 48983 7 1 2 69682 92148
0 48984 7 1 2 93724 48983
0 48985 5 1 1 48984
0 48986 7 1 2 48982 48985
0 48987 5 1 1 48986
0 48988 7 1 2 63547 48987
0 48989 5 1 1 48988
0 48990 7 1 2 64634 81883
0 48991 7 1 2 95489 48990
0 48992 7 1 2 95421 48991
0 48993 5 1 1 48992
0 48994 7 1 2 48989 48993
0 48995 5 1 1 48994
0 48996 7 1 2 70334 48995
0 48997 5 1 1 48996
0 48998 7 1 2 78209 72358
0 48999 5 1 1 48998
0 49000 7 1 2 72497 48999
0 49001 5 1 1 49000
0 49002 7 1 2 59169 49001
0 49003 5 1 1 49002
0 49004 7 1 2 6095 49003
0 49005 5 1 1 49004
0 49006 7 1 2 95503 49005
0 49007 5 1 1 49006
0 49008 7 1 2 73796 90352
0 49009 7 2 2 95313 49008
0 49010 5 1 1 95510
0 49011 7 1 2 49007 49010
0 49012 5 1 1 49011
0 49013 7 1 2 66074 49012
0 49014 5 1 1 49013
0 49015 7 1 2 94013 49014
0 49016 5 1 1 49015
0 49017 7 1 2 61978 49016
0 49018 5 1 1 49017
0 49019 7 1 2 76818 95011
0 49020 7 1 2 95200 49019
0 49021 5 1 1 49020
0 49022 7 1 2 49018 49021
0 49023 5 1 1 49022
0 49024 7 1 2 69277 49023
0 49025 5 1 1 49024
0 49026 7 1 2 48997 49025
0 49027 7 1 2 48980 49026
0 49028 5 1 1 49027
0 49029 7 1 2 59673 49028
0 49030 5 1 1 49029
0 49031 7 1 2 59170 67554
0 49032 7 1 2 75242 49031
0 49033 5 1 1 49032
0 49034 7 1 2 84148 49033
0 49035 5 1 1 49034
0 49036 7 1 2 63644 49035
0 49037 5 1 1 49036
0 49038 7 1 2 59030 70459
0 49039 7 1 2 91358 49038
0 49040 5 1 1 49039
0 49041 7 1 2 49037 49040
0 49042 5 1 1 49041
0 49043 7 1 2 57789 49042
0 49044 5 1 1 49043
0 49045 7 1 2 70789 70556
0 49046 5 1 1 49045
0 49047 7 1 2 49044 49046
0 49048 5 1 1 49047
0 49049 7 1 2 61091 49048
0 49050 5 1 1 49049
0 49051 7 1 2 2398 67966
0 49052 5 1 1 49051
0 49053 7 1 2 49050 49052
0 49054 5 1 1 49053
0 49055 7 1 2 84684 49054
0 49056 5 1 1 49055
0 49057 7 1 2 66632 69070
0 49058 5 1 1 49057
0 49059 7 1 2 58889 71966
0 49060 7 1 2 49058 49059
0 49061 5 1 1 49060
0 49062 7 1 2 249 49061
0 49063 5 1 1 49062
0 49064 7 1 2 57790 49063
0 49065 5 1 1 49064
0 49066 7 1 2 1656 49065
0 49067 5 1 1 49066
0 49068 7 2 2 81511 90547
0 49069 7 1 2 70790 95512
0 49070 7 1 2 49067 49069
0 49071 5 1 1 49070
0 49072 7 1 2 49056 49071
0 49073 5 1 1 49072
0 49074 7 1 2 75593 49073
0 49075 5 1 1 49074
0 49076 7 1 2 80121 95215
0 49077 5 1 1 49076
0 49078 7 1 2 92244 95513
0 49079 5 1 1 49078
0 49080 7 1 2 49077 49079
0 49081 5 1 1 49080
0 49082 7 1 2 74617 49081
0 49083 5 1 1 49082
0 49084 7 1 2 89180 95418
0 49085 5 1 1 49084
0 49086 7 1 2 69278 94233
0 49087 5 1 1 49086
0 49088 7 1 2 49085 49087
0 49089 5 1 1 49088
0 49090 7 1 2 86842 69121
0 49091 7 1 2 49089 49090
0 49092 5 1 1 49091
0 49093 7 1 2 49083 49092
0 49094 5 1 1 49093
0 49095 7 1 2 65094 49094
0 49096 5 1 1 49095
0 49097 7 1 2 59171 82217
0 49098 5 1 1 49097
0 49099 7 1 2 92721 49098
0 49100 5 1 1 49099
0 49101 7 1 2 58665 49100
0 49102 5 1 1 49101
0 49103 7 1 2 69988 91964
0 49104 5 1 1 49103
0 49105 7 1 2 49102 49104
0 49106 5 1 1 49105
0 49107 7 1 2 83568 49106
0 49108 5 1 1 49107
0 49109 7 1 2 49096 49108
0 49110 5 1 1 49109
0 49111 7 1 2 65334 49110
0 49112 5 1 1 49111
0 49113 7 1 2 27867 92727
0 49114 5 3 1 49113
0 49115 7 1 2 66075 95514
0 49116 5 1 1 49115
0 49117 7 1 2 88641 89360
0 49118 5 1 1 49117
0 49119 7 1 2 49116 49118
0 49120 5 1 1 49119
0 49121 7 1 2 69279 49120
0 49122 5 1 1 49121
0 49123 7 1 2 60165 82185
0 49124 7 1 2 90315 49123
0 49125 5 1 1 49124
0 49126 7 1 2 49122 49125
0 49127 7 1 2 49112 49126
0 49128 5 1 1 49127
0 49129 7 1 2 61979 49128
0 49130 5 1 1 49129
0 49131 7 1 2 40553 94425
0 49132 5 1 1 49131
0 49133 7 1 2 58666 49132
0 49134 5 1 1 49133
0 49135 7 1 2 73389 86688
0 49136 5 1 1 49135
0 49137 7 1 2 49134 49136
0 49138 5 1 1 49137
0 49139 7 1 2 70557 49138
0 49140 5 1 1 49139
0 49141 7 1 2 49130 49140
0 49142 7 1 2 49075 49141
0 49143 5 1 1 49142
0 49144 7 1 2 66940 49143
0 49145 5 1 1 49144
0 49146 7 1 2 68270 83271
0 49147 5 2 1 49146
0 49148 7 1 2 91519 95517
0 49149 5 1 1 49148
0 49150 7 1 2 71365 71099
0 49151 7 1 2 79602 49150
0 49152 5 1 1 49151
0 49153 7 1 2 49149 49152
0 49154 5 1 1 49153
0 49155 7 1 2 61468 49154
0 49156 5 1 1 49155
0 49157 7 1 2 86404 92670
0 49158 5 1 1 49157
0 49159 7 1 2 49156 49158
0 49160 5 1 1 49159
0 49161 7 1 2 64412 49160
0 49162 5 1 1 49161
0 49163 7 1 2 61092 94848
0 49164 5 1 1 49163
0 49165 7 1 2 86733 66994
0 49166 7 1 2 49164 49165
0 49167 5 1 1 49166
0 49168 7 1 2 49162 49167
0 49169 5 1 1 49168
0 49170 7 1 2 88451 49169
0 49171 5 1 1 49170
0 49172 7 1 2 64413 81891
0 49173 5 1 1 49172
0 49174 7 1 2 48361 49173
0 49175 5 1 1 49174
0 49176 7 1 2 72975 72428
0 49177 7 1 2 95518 49176
0 49178 7 1 2 49175 49177
0 49179 5 1 1 49178
0 49180 7 1 2 49171 49179
0 49181 5 1 1 49180
0 49182 7 1 2 66723 49181
0 49183 5 1 1 49182
0 49184 7 1 2 73477 74150
0 49185 7 1 2 88468 49184
0 49186 5 1 1 49185
0 49187 7 1 2 89045 49186
0 49188 5 1 1 49187
0 49189 7 1 2 80032 49188
0 49190 5 1 1 49189
0 49191 7 1 2 49183 49190
0 49192 5 1 1 49191
0 49193 7 1 2 64635 49192
0 49194 5 1 1 49193
0 49195 7 1 2 76245 79866
0 49196 5 1 1 49195
0 49197 7 2 2 72484 79437
0 49198 5 1 1 95519
0 49199 7 1 2 49196 49198
0 49200 5 1 1 49199
0 49201 7 1 2 68801 49200
0 49202 5 1 1 49201
0 49203 7 1 2 59172 95520
0 49204 5 1 1 49203
0 49205 7 1 2 49202 49204
0 49206 5 1 1 49205
0 49207 7 1 2 85551 92175
0 49208 7 1 2 49206 49207
0 49209 5 1 1 49208
0 49210 7 1 2 49194 49209
0 49211 5 1 1 49210
0 49212 7 1 2 61721 49211
0 49213 5 1 1 49212
0 49214 7 1 2 70877 92473
0 49215 5 1 1 49214
0 49216 7 1 2 70358 49215
0 49217 5 1 1 49216
0 49218 7 1 2 79954 49217
0 49219 5 1 1 49218
0 49220 7 1 2 58890 72708
0 49221 7 2 2 67120 49220
0 49222 7 1 2 74433 95521
0 49223 5 1 1 49222
0 49224 7 1 2 49219 49223
0 49225 5 1 1 49224
0 49226 7 1 2 70791 84577
0 49227 7 1 2 88470 49226
0 49228 7 1 2 49225 49227
0 49229 5 1 1 49228
0 49230 7 1 2 49213 49229
0 49231 7 1 2 49145 49230
0 49232 7 1 2 49030 49231
0 49233 5 1 1 49232
0 49234 7 1 2 88303 49233
0 49235 5 1 1 49234
0 49236 7 2 2 87579 82534
0 49237 7 3 2 81050 95523
0 49238 5 1 1 95525
0 49239 7 1 2 58667 95526
0 49240 5 1 1 49239
0 49241 7 1 2 57791 94020
0 49242 5 1 1 49241
0 49243 7 1 2 49240 49242
0 49244 5 1 1 49243
0 49245 7 1 2 57508 49244
0 49246 5 1 1 49245
0 49247 7 1 2 59933 86714
0 49248 5 1 1 49247
0 49249 7 1 2 86702 82224
0 49250 5 1 1 49249
0 49251 7 1 2 58668 49250
0 49252 5 1 1 49251
0 49253 7 1 2 49248 49252
0 49254 5 2 1 49253
0 49255 7 1 2 65723 95528
0 49256 5 1 1 49255
0 49257 7 2 2 76661 95495
0 49258 5 1 1 95530
0 49259 7 1 2 21645 49258
0 49260 5 1 1 49259
0 49261 7 1 2 57509 49260
0 49262 5 1 1 49261
0 49263 7 1 2 49256 49262
0 49264 5 1 1 49263
0 49265 7 1 2 66941 49264
0 49266 5 1 1 49265
0 49267 7 1 2 49246 49266
0 49268 5 1 1 49267
0 49269 7 1 2 64841 49268
0 49270 5 1 1 49269
0 49271 7 2 2 67598 84801
0 49272 7 1 2 95067 95532
0 49273 5 1 1 49272
0 49274 7 1 2 49270 49273
0 49275 5 1 1 49274
0 49276 7 1 2 61980 49275
0 49277 5 1 1 49276
0 49278 7 1 2 67599 72429
0 49279 7 1 2 79480 49278
0 49280 7 1 2 95012 49279
0 49281 5 1 1 49280
0 49282 7 1 2 49277 49281
0 49283 5 1 1 49282
0 49284 7 1 2 66724 49283
0 49285 5 1 1 49284
0 49286 7 4 2 57510 75594
0 49287 5 1 1 95534
0 49288 7 1 2 86703 87216
0 49289 5 3 1 49288
0 49290 7 1 2 95535 95538
0 49291 5 1 1 49290
0 49292 7 1 2 89395 49291
0 49293 5 1 1 49292
0 49294 7 1 2 66942 49293
0 49295 5 1 1 49294
0 49296 7 1 2 94023 49295
0 49297 5 1 1 49296
0 49298 7 1 2 82028 49297
0 49299 5 1 1 49298
0 49300 7 1 2 63645 49299
0 49301 7 1 2 49285 49300
0 49302 5 1 1 49301
0 49303 7 1 2 91757 95016
0 49304 5 1 1 49303
0 49305 7 1 2 57511 95228
0 49306 5 1 1 49305
0 49307 7 1 2 87565 49306
0 49308 5 1 1 49307
0 49309 7 1 2 86044 49308
0 49310 5 1 1 49309
0 49311 7 1 2 92131 49310
0 49312 5 1 1 49311
0 49313 7 1 2 74297 92015
0 49314 7 1 2 49312 49313
0 49315 5 1 1 49314
0 49316 7 1 2 49304 49315
0 49317 5 1 1 49316
0 49318 7 1 2 60166 49317
0 49319 5 1 1 49318
0 49320 7 1 2 76033 79560
0 49321 7 1 2 95017 49320
0 49322 5 1 1 49321
0 49323 7 1 2 57512 73517
0 49324 5 1 1 49323
0 49325 7 1 2 73073 49324
0 49326 5 1 1 49325
0 49327 7 1 2 94410 49326
0 49328 5 1 1 49327
0 49329 7 1 2 95536 95170
0 49330 5 1 1 49329
0 49331 7 1 2 49328 49330
0 49332 5 1 1 49331
0 49333 7 1 2 66365 49332
0 49334 5 1 1 49333
0 49335 7 1 2 76708 49287
0 49336 5 1 1 49335
0 49337 7 2 2 64842 82106
0 49338 7 1 2 92196 95541
0 49339 7 1 2 49336 49338
0 49340 5 1 1 49339
0 49341 7 1 2 49334 49340
0 49342 5 1 1 49341
0 49343 7 1 2 66943 49342
0 49344 5 1 1 49343
0 49345 7 1 2 49322 49344
0 49346 7 1 2 49319 49345
0 49347 5 1 1 49346
0 49348 7 1 2 62125 49347
0 49349 5 1 1 49348
0 49350 7 1 2 91758 95366
0 49351 7 1 2 86656 49350
0 49352 5 1 1 49351
0 49353 7 1 2 58891 49352
0 49354 7 1 2 49349 49353
0 49355 5 1 1 49354
0 49356 7 1 2 71750 49355
0 49357 7 1 2 49302 49356
0 49358 5 1 1 49357
0 49359 7 1 2 38305 95347
0 49360 5 1 1 49359
0 49361 7 2 2 71350 84475
0 49362 5 1 1 95543
0 49363 7 1 2 87836 83398
0 49364 5 1 1 49363
0 49365 7 1 2 49362 49364
0 49366 5 1 1 49365
0 49367 7 1 2 68802 49366
0 49368 5 1 1 49367
0 49369 7 1 2 84251 95544
0 49370 5 1 1 49369
0 49371 7 1 2 72443 81721
0 49372 7 1 2 95332 49371
0 49373 5 1 1 49372
0 49374 7 1 2 49370 49373
0 49375 7 1 2 49368 49374
0 49376 5 1 1 49375
0 49377 7 1 2 66366 49376
0 49378 5 1 1 49377
0 49379 7 1 2 49360 49378
0 49380 5 1 1 49379
0 49381 7 1 2 58892 49380
0 49382 5 1 1 49381
0 49383 7 2 2 73518 91156
0 49384 7 1 2 90306 94542
0 49385 7 1 2 95545 49384
0 49386 5 1 1 49385
0 49387 7 1 2 49382 49386
0 49388 5 1 1 49387
0 49389 7 1 2 62126 49388
0 49390 5 1 1 49389
0 49391 7 2 2 71351 72611
0 49392 7 1 2 86575 95547
0 49393 7 1 2 82061 49392
0 49394 5 1 1 49393
0 49395 7 1 2 49390 49394
0 49396 5 1 1 49395
0 49397 7 1 2 59674 49396
0 49398 5 1 1 49397
0 49399 7 3 2 77373 84027
0 49400 5 1 1 95549
0 49401 7 1 2 58669 95550
0 49402 5 1 1 49401
0 49403 7 1 2 95529 95198
0 49404 5 1 1 49403
0 49405 7 1 2 49402 49404
0 49406 5 1 1 49405
0 49407 7 1 2 63646 49406
0 49408 5 1 1 49407
0 49409 7 2 2 66995 82186
0 49410 7 1 2 90316 95552
0 49411 5 1 1 49410
0 49412 7 1 2 49408 49411
0 49413 5 1 1 49412
0 49414 7 1 2 70938 49413
0 49415 5 1 1 49414
0 49416 7 1 2 70558 95539
0 49417 5 1 1 49416
0 49418 7 1 2 69280 93761
0 49419 5 1 1 49418
0 49420 7 1 2 72125 49419
0 49421 5 1 1 49420
0 49422 7 1 2 84578 84303
0 49423 7 1 2 49421 49422
0 49424 5 1 1 49423
0 49425 7 1 2 49417 49424
0 49426 5 1 1 49425
0 49427 7 1 2 57792 49426
0 49428 5 1 1 49427
0 49429 7 1 2 69011 70579
0 49430 7 1 2 95540 49429
0 49431 5 1 1 49430
0 49432 7 1 2 48676 49431
0 49433 5 1 1 49432
0 49434 7 1 2 62127 49433
0 49435 5 1 1 49434
0 49436 7 1 2 49428 49435
0 49437 5 1 1 49436
0 49438 7 1 2 75595 49437
0 49439 5 1 1 49438
0 49440 7 3 2 80410 94958
0 49441 5 1 1 95554
0 49442 7 1 2 69147 88927
0 49443 7 1 2 85454 49442
0 49444 5 1 1 49443
0 49445 7 1 2 49441 49444
0 49446 5 1 1 49445
0 49447 7 1 2 61981 72709
0 49448 7 1 2 49446 49447
0 49449 5 1 1 49448
0 49450 7 1 2 49439 49449
0 49451 7 1 2 49415 49450
0 49452 7 1 2 49398 49451
0 49453 5 1 1 49452
0 49454 7 1 2 66944 49453
0 49455 5 1 1 49454
0 49456 7 2 2 70535 94852
0 49457 7 1 2 74900 95557
0 49458 5 1 1 49457
0 49459 7 1 2 78954 69683
0 49460 5 1 1 49459
0 49461 7 1 2 86045 69281
0 49462 5 1 1 49461
0 49463 7 1 2 49460 49462
0 49464 5 1 1 49463
0 49465 7 1 2 64744 78326
0 49466 7 1 2 49464 49465
0 49467 5 1 1 49466
0 49468 7 1 2 49458 49467
0 49469 5 1 1 49468
0 49470 7 1 2 61982 49469
0 49471 5 1 1 49470
0 49472 7 1 2 86071 90218
0 49473 5 1 1 49472
0 49474 7 1 2 49471 49473
0 49475 5 1 1 49474
0 49476 7 1 2 65724 49475
0 49477 5 1 1 49476
0 49478 7 2 2 66633 75789
0 49479 7 1 2 66793 95559
0 49480 5 1 1 49479
0 49481 7 1 2 76005 49480
0 49482 5 1 1 49481
0 49483 7 1 2 70536 49482
0 49484 5 1 1 49483
0 49485 7 1 2 82070 95560
0 49486 5 1 1 49485
0 49487 7 1 2 49484 49486
0 49488 5 1 1 49487
0 49489 7 1 2 90548 49488
0 49490 5 1 1 49489
0 49491 7 1 2 49477 49490
0 49492 5 1 1 49491
0 49493 7 1 2 82420 49492
0 49494 5 1 1 49493
0 49495 7 1 2 61093 92298
0 49496 5 1 1 49495
0 49497 7 1 2 79443 49496
0 49498 5 1 1 49497
0 49499 7 1 2 66076 49498
0 49500 5 1 1 49499
0 49501 7 1 2 68803 95321
0 49502 5 1 1 49501
0 49503 7 1 2 57793 93938
0 49504 5 1 1 49503
0 49505 7 1 2 49502 49504
0 49506 5 1 1 49505
0 49507 7 1 2 65725 49506
0 49508 5 1 1 49507
0 49509 7 1 2 49500 49508
0 49510 5 1 1 49509
0 49511 7 1 2 82037 89569
0 49512 7 1 2 49510 49511
0 49513 5 1 1 49512
0 49514 7 1 2 49494 49513
0 49515 5 1 1 49514
0 49516 7 1 2 59675 49515
0 49517 5 1 1 49516
0 49518 7 2 2 66367 74428
0 49519 5 1 1 95561
0 49520 7 1 2 59934 95562
0 49521 5 1 1 49520
0 49522 7 1 2 88280 49521
0 49523 5 1 1 49522
0 49524 7 1 2 76062 49523
0 49525 5 1 1 49524
0 49526 7 1 2 79183 82764
0 49527 7 1 2 95490 49526
0 49528 5 1 1 49527
0 49529 7 1 2 49525 49528
0 49530 5 1 1 49529
0 49531 7 1 2 57794 49530
0 49532 5 1 1 49531
0 49533 7 1 2 89570 95378
0 49534 5 1 1 49533
0 49535 7 1 2 49532 49534
0 49536 5 1 1 49535
0 49537 7 1 2 58893 49536
0 49538 5 1 1 49537
0 49539 7 2 2 77374 90264
0 49540 7 1 2 80117 82788
0 49541 7 1 2 95563 49540
0 49542 5 1 1 49541
0 49543 7 1 2 49538 49542
0 49544 5 1 1 49543
0 49545 7 1 2 67961 90819
0 49546 7 1 2 49544 49545
0 49547 5 1 1 49546
0 49548 7 1 2 49517 49547
0 49549 5 1 1 49548
0 49550 7 1 2 58670 49549
0 49551 5 1 1 49550
0 49552 7 1 2 67487 79955
0 49553 5 1 1 49552
0 49554 7 1 2 76141 49553
0 49555 5 1 1 49554
0 49556 7 1 2 70939 49555
0 49557 5 1 1 49556
0 49558 7 1 2 57795 76112
0 49559 7 1 2 74898 49558
0 49560 7 1 2 82310 49559
0 49561 5 1 1 49560
0 49562 7 1 2 69012 77222
0 49563 7 1 2 70537 49562
0 49564 7 1 2 74774 49563
0 49565 5 1 1 49564
0 49566 7 1 2 49561 49565
0 49567 7 1 2 49557 49566
0 49568 5 1 1 49567
0 49569 7 1 2 61094 49568
0 49570 5 1 1 49569
0 49571 7 1 2 69747 69559
0 49572 7 1 2 88258 49571
0 49573 7 1 2 95423 49572
0 49574 5 1 1 49573
0 49575 7 1 2 49570 49574
0 49576 5 1 1 49575
0 49577 7 1 2 61469 49576
0 49578 5 1 1 49577
0 49579 7 1 2 86734 79303
0 49580 7 1 2 79944 94543
0 49581 7 1 2 49579 49580
0 49582 5 1 1 49581
0 49583 7 1 2 49578 49582
0 49584 5 1 1 49583
0 49585 7 1 2 87268 49584
0 49586 5 1 1 49585
0 49587 7 1 2 49551 49586
0 49588 7 1 2 49455 49587
0 49589 7 1 2 49358 49588
0 49590 5 1 1 49589
0 49591 7 1 2 88304 49590
0 49592 5 1 1 49591
0 49593 7 1 2 75718 88866
0 49594 7 2 2 89150 91832
0 49595 7 1 2 94199 95565
0 49596 7 1 2 49593 49595
0 49597 7 1 2 95477 49596
0 49598 5 1 1 49597
0 49599 7 1 2 49592 49598
0 49600 5 1 1 49599
0 49601 7 1 2 71915 49600
0 49602 5 1 1 49601
0 49603 7 1 2 70580 89331
0 49604 5 1 1 49603
0 49605 7 2 2 72485 87662
0 49606 7 1 2 67938 93916
0 49607 7 1 2 95567 49606
0 49608 5 1 1 49607
0 49609 7 1 2 49604 49608
0 49610 5 1 1 49609
0 49611 7 1 2 62128 49610
0 49612 5 1 1 49611
0 49613 7 1 2 80750 95283
0 49614 5 1 1 49613
0 49615 7 1 2 65726 95216
0 49616 5 1 1 49615
0 49617 7 1 2 49614 49616
0 49618 5 1 1 49617
0 49619 7 1 2 57513 49618
0 49620 5 1 1 49619
0 49621 7 1 2 70792 89361
0 49622 5 1 1 49621
0 49623 7 1 2 49620 49622
0 49624 5 1 1 49623
0 49625 7 1 2 72569 49624
0 49626 5 1 1 49625
0 49627 7 1 2 49612 49626
0 49628 5 1 1 49627
0 49629 7 1 2 66945 49628
0 49630 5 1 1 49629
0 49631 7 1 2 58894 95341
0 49632 5 1 1 49631
0 49633 7 1 2 70463 91290
0 49634 5 1 1 49633
0 49635 7 1 2 49632 49634
0 49636 5 1 1 49635
0 49637 7 1 2 61983 49636
0 49638 5 1 1 49637
0 49639 7 1 2 85399 79935
0 49640 7 1 2 95456 49639
0 49641 5 1 1 49640
0 49642 7 1 2 49638 49641
0 49643 5 1 1 49642
0 49644 7 1 2 70793 49643
0 49645 5 1 1 49644
0 49646 7 1 2 80441 84167
0 49647 7 1 2 94563 49646
0 49648 5 1 1 49647
0 49649 7 1 2 49645 49648
0 49650 5 1 1 49649
0 49651 7 1 2 66794 49650
0 49652 5 1 1 49651
0 49653 7 1 2 57514 70559
0 49654 5 1 1 49653
0 49655 7 2 2 63647 76860
0 49656 7 1 2 74855 95569
0 49657 5 1 1 49656
0 49658 7 1 2 49654 49657
0 49659 5 1 1 49658
0 49660 7 1 2 94021 49659
0 49661 5 1 1 49660
0 49662 7 1 2 49652 49661
0 49663 7 1 2 49630 49662
0 49664 5 1 1 49663
0 49665 7 1 2 88305 49664
0 49666 5 1 1 49665
0 49667 7 1 2 72639 91206
0 49668 7 2 2 95478 49667
0 49669 7 1 2 73844 89151
0 49670 7 2 2 92967 49669
0 49671 7 1 2 82789 95573
0 49672 7 1 2 95571 49671
0 49673 5 1 1 49672
0 49674 7 1 2 49666 49673
0 49675 5 1 1 49674
0 49676 7 1 2 78327 49675
0 49677 5 1 1 49676
0 49678 7 1 2 94505 95505
0 49679 5 1 1 49678
0 49680 7 1 2 60167 92180
0 49681 5 1 1 49680
0 49682 7 1 2 37214 49681
0 49683 5 1 1 49682
0 49684 7 1 2 61095 67607
0 49685 5 2 1 49684
0 49686 7 1 2 66368 95575
0 49687 7 1 2 49683 49686
0 49688 5 1 1 49687
0 49689 7 1 2 49679 49688
0 49690 5 1 1 49689
0 49691 7 1 2 59676 49690
0 49692 5 1 1 49691
0 49693 7 1 2 94506 95511
0 49694 5 1 1 49693
0 49695 7 1 2 49692 49694
0 49696 5 1 1 49695
0 49697 7 1 2 66077 49696
0 49698 5 1 1 49697
0 49699 7 1 2 73229 87770
0 49700 5 1 1 49699
0 49701 7 1 2 87217 49700
0 49702 5 1 1 49701
0 49703 7 1 2 95309 49702
0 49704 5 1 1 49703
0 49705 7 1 2 88289 94016
0 49706 5 1 1 49705
0 49707 7 1 2 49704 49706
0 49708 5 1 1 49707
0 49709 7 1 2 57515 49708
0 49710 5 1 1 49709
0 49711 7 1 2 92169 38407
0 49712 5 1 1 49711
0 49713 7 1 2 61722 49712
0 49714 5 1 1 49713
0 49715 7 1 2 49710 49714
0 49716 5 1 1 49715
0 49717 7 1 2 94408 49716
0 49718 5 1 1 49717
0 49719 7 1 2 49698 49718
0 49720 5 1 1 49719
0 49721 7 1 2 66634 49720
0 49722 5 1 1 49721
0 49723 7 1 2 87663 91833
0 49724 7 1 2 94200 49723
0 49725 5 1 1 49724
0 49726 7 1 2 63648 49725
0 49727 7 1 2 49722 49726
0 49728 5 1 1 49727
0 49729 7 1 2 66635 95576
0 49730 7 1 2 95493 49729
0 49731 5 1 1 49730
0 49732 7 1 2 47240 49731
0 49733 5 1 1 49732
0 49734 7 1 2 64843 49733
0 49735 5 1 1 49734
0 49736 7 1 2 95369 95168
0 49737 5 1 1 49736
0 49738 7 1 2 49735 49737
0 49739 5 1 1 49738
0 49740 7 1 2 66078 49739
0 49741 5 1 1 49740
0 49742 7 1 2 79727 89471
0 49743 7 1 2 95370 49742
0 49744 5 1 1 49743
0 49745 7 1 2 66369 49744
0 49746 7 1 2 49741 49745
0 49747 5 1 1 49746
0 49748 7 1 2 87142 91843
0 49749 5 1 1 49748
0 49750 7 1 2 92163 49749
0 49751 5 1 1 49750
0 49752 7 1 2 66996 73446
0 49753 7 1 2 49751 49752
0 49754 5 1 1 49753
0 49755 7 1 2 76610 77828
0 49756 7 1 2 72976 49755
0 49757 7 1 2 73478 49756
0 49758 5 1 1 49757
0 49759 7 1 2 49754 49758
0 49760 5 1 1 49759
0 49761 7 1 2 67600 49760
0 49762 5 1 1 49761
0 49763 7 1 2 67078 95324
0 49764 5 1 1 49763
0 49765 7 1 2 61723 49764
0 49766 7 1 2 49762 49765
0 49767 5 1 1 49766
0 49768 7 1 2 59677 49767
0 49769 7 1 2 49747 49768
0 49770 5 1 1 49769
0 49771 7 1 2 72977 90307
0 49772 5 1 1 49771
0 49773 7 1 2 57796 94496
0 49774 7 1 2 94960 49773
0 49775 5 1 1 49774
0 49776 7 1 2 49772 49775
0 49777 5 1 1 49776
0 49778 7 1 2 75596 49777
0 49779 5 1 1 49778
0 49780 7 2 2 67121 93917
0 49781 7 1 2 95568 95577
0 49782 5 1 1 49781
0 49783 7 1 2 66997 95531
0 49784 5 1 1 49783
0 49785 7 1 2 49782 49784
0 49786 7 1 2 49779 49785
0 49787 5 1 1 49786
0 49788 7 1 2 66946 49787
0 49789 5 1 1 49788
0 49790 7 1 2 79988 95333
0 49791 7 1 2 94503 49790
0 49792 5 1 1 49791
0 49793 7 2 2 65335 92968
0 49794 7 1 2 63548 67079
0 49795 7 1 2 93859 49794
0 49796 7 1 2 95579 49795
0 49797 5 1 1 49796
0 49798 7 1 2 49792 49797
0 49799 5 1 1 49798
0 49800 7 1 2 61724 49799
0 49801 5 1 1 49800
0 49802 7 1 2 87885 67122
0 49803 7 1 2 79728 92149
0 49804 7 1 2 49802 49803
0 49805 5 1 1 49804
0 49806 7 1 2 58895 49805
0 49807 7 1 2 49801 49806
0 49808 7 1 2 49789 49807
0 49809 7 1 2 49770 49808
0 49810 5 1 1 49809
0 49811 7 1 2 49728 49810
0 49812 5 1 1 49811
0 49813 7 1 2 62129 49812
0 49814 5 1 1 49813
0 49815 7 1 2 80779 74075
0 49816 5 1 1 49815
0 49817 7 1 2 47215 49816
0 49818 5 1 1 49817
0 49819 7 1 2 59173 49818
0 49820 5 1 1 49819
0 49821 7 1 2 24389 49820
0 49822 5 1 1 49821
0 49823 7 1 2 86094 49822
0 49824 5 1 1 49823
0 49825 7 1 2 74151 73367
0 49826 7 1 2 73864 49825
0 49827 7 1 2 86072 49826
0 49828 5 1 1 49827
0 49829 7 1 2 49824 49828
0 49830 5 1 1 49829
0 49831 7 1 2 65336 49830
0 49832 5 1 1 49831
0 49833 7 1 2 80118 91104
0 49834 7 1 2 95314 49833
0 49835 5 1 1 49834
0 49836 7 1 2 49832 49835
0 49837 5 1 1 49836
0 49838 7 1 2 61725 49837
0 49839 5 1 1 49838
0 49840 7 1 2 73682 73990
0 49841 5 1 1 49840
0 49842 7 1 2 80594 49841
0 49843 5 1 1 49842
0 49844 7 1 2 64636 49843
0 49845 5 1 1 49844
0 49846 7 1 2 85603 49845
0 49847 5 1 1 49846
0 49848 7 1 2 79914 49847
0 49849 5 1 1 49848
0 49850 7 1 2 83001 95276
0 49851 7 1 2 80751 49850
0 49852 5 1 1 49851
0 49853 7 1 2 49849 49852
0 49854 5 1 1 49853
0 49855 7 1 2 69560 83050
0 49856 7 1 2 49854 49855
0 49857 5 1 1 49856
0 49858 7 1 2 49839 49857
0 49859 5 1 1 49858
0 49860 7 1 2 61984 49859
0 49861 5 1 1 49860
0 49862 7 1 2 78972 74658
0 49863 7 1 2 82995 49862
0 49864 7 1 2 88080 91919
0 49865 7 1 2 49863 49864
0 49866 5 1 1 49865
0 49867 7 1 2 66725 49866
0 49868 7 1 2 49861 49867
0 49869 5 1 1 49868
0 49870 7 1 2 88306 49869
0 49871 7 1 2 49814 49870
0 49872 5 1 1 49871
0 49873 7 1 2 81741 95574
0 49874 7 1 2 95572 49873
0 49875 5 1 1 49874
0 49876 7 1 2 49872 49875
0 49877 5 1 1 49876
0 49878 7 1 2 71751 49877
0 49879 5 1 1 49878
0 49880 7 1 2 49677 49879
0 49881 7 1 2 49602 49880
0 49882 7 1 2 49235 49881
0 49883 5 1 1 49882
0 49884 7 1 2 70431 49883
0 49885 5 1 1 49884
0 49886 7 1 2 73819 95239
0 49887 5 1 1 49886
0 49888 7 1 2 11630 49887
0 49889 5 1 1 49888
0 49890 7 1 2 58356 49889
0 49891 5 1 1 49890
0 49892 7 1 2 85766 49891
0 49893 5 1 1 49892
0 49894 7 1 2 73553 49893
0 49895 5 1 1 49894
0 49896 7 1 2 78976 77543
0 49897 5 1 1 49896
0 49898 7 1 2 76709 94663
0 49899 7 1 2 49897 49898
0 49900 5 1 1 49899
0 49901 7 1 2 49895 49900
0 49902 5 1 1 49901
0 49903 7 1 2 71086 49902
0 49904 5 1 1 49903
0 49905 7 1 2 70432 67488
0 49906 7 1 2 86242 95578
0 49907 7 1 2 49905 49906
0 49908 5 1 1 49907
0 49909 7 1 2 49904 49908
0 49910 5 1 1 49909
0 49911 7 1 2 66370 49910
0 49912 5 1 1 49911
0 49913 7 1 2 63411 86221
0 49914 5 1 1 49913
0 49915 7 2 2 76477 49914
0 49916 7 1 2 95551 95581
0 49917 5 1 1 49916
0 49918 7 1 2 49912 49917
0 49919 5 1 1 49918
0 49920 7 1 2 63649 49919
0 49921 5 1 1 49920
0 49922 7 1 2 66998 95582
0 49923 5 1 1 49922
0 49924 7 1 2 76585 81722
0 49925 7 1 2 80242 49924
0 49926 5 1 1 49925
0 49927 7 1 2 49923 49926
0 49928 5 1 1 49927
0 49929 7 1 2 82584 49928
0 49930 5 1 1 49929
0 49931 7 1 2 76861 94548
0 49932 7 1 2 95126 49931
0 49933 7 1 2 83630 49932
0 49934 5 1 1 49933
0 49935 7 1 2 49930 49934
0 49936 5 1 1 49935
0 49937 7 1 2 68667 49936
0 49938 5 1 1 49937
0 49939 7 1 2 49921 49938
0 49940 5 1 1 49939
0 49941 7 1 2 57797 49940
0 49942 5 1 1 49941
0 49943 7 1 2 72570 89382
0 49944 5 1 1 49943
0 49945 7 1 2 71352 93927
0 49946 5 1 1 49945
0 49947 7 1 2 95349 49946
0 49948 5 1 1 49947
0 49949 7 1 2 58896 49948
0 49950 5 1 1 49949
0 49951 7 1 2 63650 71376
0 49952 7 1 2 93928 49951
0 49953 5 1 1 49952
0 49954 7 1 2 49950 49953
0 49955 5 2 1 49954
0 49956 7 1 2 59174 72421
0 49957 7 1 2 95583 49956
0 49958 5 1 1 49957
0 49959 7 1 2 49944 49958
0 49960 5 1 1 49959
0 49961 7 1 2 65337 49960
0 49962 5 1 1 49961
0 49963 7 1 2 72422 83651
0 49964 7 1 2 92245 49963
0 49965 5 1 1 49964
0 49966 7 1 2 49962 49965
0 49967 5 1 1 49966
0 49968 7 1 2 67383 49967
0 49969 5 1 1 49968
0 49970 7 1 2 85298 95584
0 49971 5 1 1 49970
0 49972 7 1 2 61985 70433
0 49973 7 1 2 73985 91428
0 49974 7 1 2 49972 49973
0 49975 5 1 1 49974
0 49976 7 1 2 49971 49975
0 49977 5 1 1 49976
0 49978 7 1 2 62130 49977
0 49979 5 1 1 49978
0 49980 7 1 2 49969 49979
0 49981 7 1 2 49942 49980
0 49982 5 1 1 49981
0 49983 7 1 2 66947 49982
0 49984 5 1 1 49983
0 49985 7 1 2 65338 86675
0 49986 7 1 2 69249 49985
0 49987 7 1 2 89349 49986
0 49988 5 1 1 49987
0 49989 7 1 2 95315 95401
0 49990 5 1 1 49989
0 49991 7 1 2 57516 92354
0 49992 5 1 1 49991
0 49993 7 1 2 49990 49992
0 49994 5 1 1 49993
0 49995 7 1 2 76429 70549
0 49996 7 1 2 49994 49995
0 49997 5 1 1 49996
0 49998 7 1 2 49988 49997
0 49999 5 1 1 49998
0 50000 7 1 2 94493 49999
0 50001 5 1 1 50000
0 50002 7 1 2 83667 88106
0 50003 5 1 1 50002
0 50004 7 1 2 85282 82353
0 50005 5 1 1 50004
0 50006 7 1 2 18856 50005
0 50007 5 1 1 50006
0 50008 7 1 2 63651 50007
0 50009 5 1 1 50008
0 50010 7 1 2 50003 50009
0 50011 5 1 1 50010
0 50012 7 1 2 66726 50011
0 50013 5 1 1 50012
0 50014 7 1 2 76417 95537
0 50015 7 1 2 83106 50014
0 50016 5 1 1 50015
0 50017 7 1 2 50013 50016
0 50018 5 1 1 50017
0 50019 7 1 2 64745 50018
0 50020 5 1 1 50019
0 50021 7 2 2 62131 70434
0 50022 7 1 2 76587 95585
0 50023 5 1 1 50022
0 50024 7 1 2 85299 69581
0 50025 5 1 1 50024
0 50026 7 1 2 50023 50025
0 50027 5 1 1 50026
0 50028 7 1 2 59935 50027
0 50029 5 1 1 50028
0 50030 7 1 2 88171 94521
0 50031 5 1 1 50030
0 50032 7 1 2 63549 50031
0 50033 7 1 2 50029 50032
0 50034 5 1 1 50033
0 50035 7 1 2 58802 6383
0 50036 5 1 1 50035
0 50037 7 1 2 60062 50036
0 50038 7 1 2 50034 50037
0 50039 5 1 1 50038
0 50040 7 1 2 50020 50039
0 50041 5 1 1 50040
0 50042 7 1 2 74298 50041
0 50043 5 1 1 50042
0 50044 7 1 2 50001 50043
0 50045 5 1 1 50044
0 50046 7 1 2 61726 50045
0 50047 5 1 1 50046
0 50048 7 1 2 83608 82723
0 50049 7 1 2 95380 50048
0 50050 5 1 1 50049
0 50051 7 1 2 50047 50050
0 50052 5 1 1 50051
0 50053 7 1 2 68412 50052
0 50054 5 1 1 50053
0 50055 7 2 2 81121 83556
0 50056 7 1 2 84160 95587
0 50057 5 1 1 50056
0 50058 7 2 2 79030 81530
0 50059 7 1 2 82535 95589
0 50060 5 1 1 50059
0 50061 7 1 2 58803 76478
0 50062 7 1 2 81362 50061
0 50063 5 1 1 50062
0 50064 7 1 2 78973 95451
0 50065 7 1 2 80245 50064
0 50066 5 1 1 50065
0 50067 7 1 2 50063 50066
0 50068 5 1 1 50067
0 50069 7 1 2 57798 50068
0 50070 5 1 1 50069
0 50071 7 1 2 50060 50070
0 50072 5 1 1 50071
0 50073 7 1 2 70581 50072
0 50074 5 1 1 50073
0 50075 7 1 2 50057 50074
0 50076 5 1 1 50075
0 50077 7 1 2 64746 50076
0 50078 5 1 1 50077
0 50079 7 1 2 73971 69141
0 50080 7 1 2 83520 50079
0 50081 7 1 2 93929 50080
0 50082 5 1 1 50081
0 50083 7 1 2 50078 50082
0 50084 5 1 1 50083
0 50085 7 1 2 95580 50084
0 50086 5 1 1 50085
0 50087 7 1 2 69219 92611
0 50088 7 1 2 95588 50087
0 50089 5 1 1 50088
0 50090 7 1 2 50086 50089
0 50091 5 1 1 50090
0 50092 7 1 2 62132 50091
0 50093 5 1 1 50092
0 50094 7 2 2 83367 82421
0 50095 5 1 1 95591
0 50096 7 1 2 69195 82118
0 50097 5 1 1 50096
0 50098 7 1 2 50095 50097
0 50099 5 1 1 50098
0 50100 7 1 2 79835 50099
0 50101 5 1 1 50100
0 50102 7 2 2 79309 94441
0 50103 7 1 2 76101 82720
0 50104 7 1 2 95593 50103
0 50105 5 1 1 50104
0 50106 7 1 2 50101 50105
0 50107 5 1 1 50106
0 50108 7 1 2 76479 50107
0 50109 5 1 1 50108
0 50110 7 1 2 92230 94534
0 50111 5 1 1 50110
0 50112 7 1 2 81884 94537
0 50113 5 1 1 50112
0 50114 7 1 2 50111 50113
0 50115 5 3 1 50114
0 50116 7 1 2 62805 83824
0 50117 5 1 1 50116
0 50118 7 1 2 95595 50117
0 50119 5 1 1 50118
0 50120 7 1 2 83652 89335
0 50121 5 1 1 50120
0 50122 7 1 2 50119 50121
0 50123 5 1 1 50122
0 50124 7 1 2 58804 50123
0 50125 5 1 1 50124
0 50126 7 2 2 66636 91529
0 50127 7 1 2 76333 79042
0 50128 7 1 2 95598 50127
0 50129 5 1 1 50128
0 50130 7 1 2 50125 50129
0 50131 5 1 1 50130
0 50132 7 1 2 62133 50131
0 50133 5 1 1 50132
0 50134 7 1 2 50109 50133
0 50135 5 1 1 50134
0 50136 7 1 2 81046 50135
0 50137 5 1 1 50136
0 50138 7 2 2 76792 82119
0 50139 7 1 2 71124 95427
0 50140 7 1 2 95600 50139
0 50141 5 1 1 50140
0 50142 7 1 2 50137 50141
0 50143 5 1 1 50142
0 50144 7 1 2 72248 50143
0 50145 5 1 1 50144
0 50146 7 1 2 72710 95596
0 50147 5 1 1 50146
0 50148 7 1 2 70538 95592
0 50149 5 1 1 50148
0 50150 7 1 2 50147 50149
0 50151 5 1 1 50150
0 50152 7 1 2 57517 50151
0 50153 5 1 1 50152
0 50154 7 2 2 64747 89571
0 50155 5 1 1 95602
0 50156 7 1 2 81569 79814
0 50157 5 1 1 50156
0 50158 7 1 2 50155 50157
0 50159 5 1 1 50158
0 50160 7 1 2 58897 50159
0 50161 5 1 1 50160
0 50162 7 1 2 65095 90308
0 50163 7 1 2 92231 50162
0 50164 5 1 1 50163
0 50165 7 1 2 50161 50164
0 50166 5 1 1 50165
0 50167 7 1 2 74299 50166
0 50168 5 1 1 50167
0 50169 7 1 2 50153 50168
0 50170 5 1 1 50169
0 50171 7 1 2 74891 86320
0 50172 7 1 2 50170 50171
0 50173 5 1 1 50172
0 50174 7 1 2 84270 91658
0 50175 7 1 2 95457 50174
0 50176 5 1 1 50175
0 50177 7 1 2 50173 50176
0 50178 5 1 1 50177
0 50179 7 1 2 72211 50178
0 50180 5 1 1 50179
0 50181 7 1 2 76480 72670
0 50182 7 1 2 88290 50181
0 50183 7 1 2 61096 70725
0 50184 5 1 1 50183
0 50185 7 1 2 50184 95186
0 50186 7 1 2 50182 50185
0 50187 7 1 2 82324 50186
0 50188 5 1 1 50187
0 50189 7 1 2 50180 50188
0 50190 7 1 2 50145 50189
0 50191 7 1 2 50093 50190
0 50192 7 1 2 50054 50191
0 50193 7 1 2 49984 50192
0 50194 5 1 1 50193
0 50195 7 1 2 88307 50194
0 50196 5 1 1 50195
0 50197 7 1 2 72571 89389
0 50198 5 1 1 50197
0 50199 7 1 2 66637 94432
0 50200 7 1 2 95462 50199
0 50201 5 1 1 50200
0 50202 7 1 2 50198 50201
0 50203 5 1 1 50202
0 50204 7 1 2 67384 50203
0 50205 5 1 1 50204
0 50206 7 1 2 73358 90353
0 50207 7 1 2 95177 50206
0 50208 7 1 2 85300 50207
0 50209 5 1 1 50208
0 50210 7 1 2 50205 50209
0 50211 5 1 1 50210
0 50212 7 1 2 79915 50211
0 50213 5 1 1 50212
0 50214 7 1 2 73879 95452
0 50215 7 1 2 70560 50214
0 50216 5 1 1 50215
0 50217 7 1 2 67445 76053
0 50218 7 1 2 76862 50217
0 50219 7 1 2 81126 50218
0 50220 5 1 1 50219
0 50221 7 1 2 50216 50220
0 50222 5 1 1 50221
0 50223 7 1 2 70061 82646
0 50224 7 1 2 50222 50223
0 50225 5 1 1 50224
0 50226 7 1 2 50213 50225
0 50227 5 1 1 50226
0 50228 7 1 2 88308 50227
0 50229 5 1 1 50228
0 50230 7 1 2 66371 77375
0 50231 7 2 2 94737 50230
0 50232 7 1 2 81542 89152
0 50233 7 1 2 94867 50232
0 50234 7 1 2 95604 50233
0 50235 5 1 1 50234
0 50236 7 1 2 50229 50235
0 50237 5 1 1 50236
0 50238 7 1 2 94853 50237
0 50239 5 1 1 50238
0 50240 7 1 2 64637 72430
0 50241 7 1 2 90286 50240
0 50242 5 1 1 50241
0 50243 7 1 2 49400 50242
0 50244 5 1 1 50243
0 50245 7 1 2 63652 50244
0 50246 5 1 1 50245
0 50247 7 1 2 90313 95553
0 50248 5 1 1 50247
0 50249 7 1 2 50246 50248
0 50250 5 1 1 50249
0 50251 7 1 2 76481 50250
0 50252 5 1 1 50251
0 50253 7 1 2 82721 90211
0 50254 7 1 2 95374 50253
0 50255 5 1 1 50254
0 50256 7 1 2 50252 50255
0 50257 5 1 1 50256
0 50258 7 1 2 85301 50257
0 50259 5 1 1 50258
0 50260 7 1 2 80089 94854
0 50261 5 1 1 50260
0 50262 7 3 2 80462 69250
0 50263 5 3 1 95606
0 50264 7 1 2 50261 95609
0 50265 5 1 1 50264
0 50266 7 1 2 67385 50265
0 50267 5 1 1 50266
0 50268 7 1 2 72260 72444
0 50269 7 1 2 95586 50268
0 50270 5 1 1 50269
0 50271 7 1 2 50267 50270
0 50272 5 1 1 50271
0 50273 7 1 2 61727 50272
0 50274 5 1 1 50273
0 50275 7 1 2 66372 78974
0 50276 7 1 2 83428 50275
0 50277 5 1 1 50276
0 50278 7 1 2 50274 50277
0 50279 5 1 1 50278
0 50280 7 1 2 91411 50279
0 50281 5 1 1 50280
0 50282 7 1 2 50259 50281
0 50283 5 1 1 50282
0 50284 7 1 2 66948 50283
0 50285 5 1 1 50284
0 50286 7 1 2 74002 95428
0 50287 7 1 2 95601 50286
0 50288 5 1 1 50287
0 50289 7 1 2 74892 81047
0 50290 7 1 2 94855 50289
0 50291 7 1 2 95597 50290
0 50292 5 1 1 50291
0 50293 7 1 2 50288 50292
0 50294 5 1 1 50293
0 50295 7 1 2 67386 50294
0 50296 5 1 1 50295
0 50297 7 1 2 86926 87668
0 50298 5 1 1 50297
0 50299 7 1 2 82367 91118
0 50300 7 1 2 82828 50299
0 50301 5 1 1 50300
0 50302 7 1 2 50298 50301
0 50303 5 1 1 50302
0 50304 7 1 2 79836 50303
0 50305 5 1 1 50304
0 50306 7 1 2 67446 95590
0 50307 7 1 2 95594 50306
0 50308 5 1 1 50307
0 50309 7 1 2 50305 50308
0 50310 5 1 1 50309
0 50311 7 1 2 76482 50310
0 50312 5 1 1 50311
0 50313 7 1 2 76581 76854
0 50314 5 1 1 50313
0 50315 7 1 2 72126 50314
0 50316 5 1 1 50315
0 50317 7 1 2 68047 50316
0 50318 5 1 1 50317
0 50319 7 1 2 76573 50318
0 50320 5 1 1 50319
0 50321 7 1 2 64748 94435
0 50322 7 1 2 50320 50321
0 50323 5 1 1 50322
0 50324 7 1 2 50312 50323
0 50325 5 1 1 50324
0 50326 7 1 2 58671 50325
0 50327 5 1 1 50326
0 50328 7 1 2 50296 50327
0 50329 7 1 2 50285 50328
0 50330 5 1 1 50329
0 50331 7 1 2 88309 50330
0 50332 5 1 1 50331
0 50333 7 1 2 76437 89153
0 50334 7 1 2 94029 94553
0 50335 7 1 2 50333 50334
0 50336 7 1 2 95605 50335
0 50337 5 1 1 50336
0 50338 7 1 2 50332 50337
0 50339 5 1 1 50338
0 50340 7 1 2 71916 50339
0 50341 5 1 1 50340
0 50342 7 1 2 50239 50341
0 50343 7 1 2 50196 50342
0 50344 5 1 1 50343
0 50345 7 1 2 93830 50344
0 50346 5 1 1 50345
0 50347 7 1 2 88616 49519
0 50348 5 1 1 50347
0 50349 7 1 2 86927 50348
0 50350 5 1 1 50349
0 50351 7 1 2 87433 95273
0 50352 5 1 1 50351
0 50353 7 1 2 94455 50352
0 50354 7 1 2 50350 50353
0 50355 5 1 1 50354
0 50356 7 1 2 73057 50355
0 50357 5 1 1 50356
0 50358 7 1 2 59031 79461
0 50359 7 1 2 91450 50358
0 50360 5 1 1 50359
0 50361 7 1 2 50357 50360
0 50362 5 1 1 50361
0 50363 7 1 2 61097 50362
0 50364 5 1 1 50363
0 50365 7 1 2 74157 92735
0 50366 7 1 2 94755 50365
0 50367 5 1 1 50366
0 50368 7 1 2 50364 50367
0 50369 5 1 1 50368
0 50370 7 1 2 66638 50369
0 50371 5 1 1 50370
0 50372 7 1 2 74137 84579
0 50373 7 1 2 81742 50372
0 50374 7 1 2 94883 50373
0 50375 5 1 1 50374
0 50376 7 1 2 50371 50375
0 50377 5 1 1 50376
0 50378 7 1 2 60063 50377
0 50379 5 1 1 50378
0 50380 7 1 2 74546 74490
0 50381 7 1 2 86525 50380
0 50382 7 1 2 94665 50381
0 50383 5 1 1 50382
0 50384 7 1 2 50379 50383
0 50385 5 1 1 50384
0 50386 7 1 2 62134 50385
0 50387 5 1 1 50386
0 50388 7 2 2 94532 94879
0 50389 7 1 2 92309 94672
0 50390 7 1 2 95612 50389
0 50391 5 1 1 50390
0 50392 7 1 2 50387 50391
0 50393 5 1 1 50392
0 50394 7 1 2 70539 50393
0 50395 5 1 1 50394
0 50396 7 1 2 69582 89207
0 50397 5 1 1 50396
0 50398 7 1 2 5974 50397
0 50399 5 1 1 50398
0 50400 7 1 2 92105 50399
0 50401 5 1 1 50400
0 50402 7 1 2 67939 74429
0 50403 7 1 2 85112 50402
0 50404 7 1 2 95204 50403
0 50405 5 1 1 50404
0 50406 7 1 2 50401 50405
0 50407 5 1 1 50406
0 50408 7 1 2 85302 50407
0 50409 5 1 1 50408
0 50410 7 1 2 64749 95555
0 50411 5 1 1 50410
0 50412 7 1 2 63653 60064
0 50413 7 1 2 80442 50412
0 50414 7 1 2 95175 50413
0 50415 7 1 2 95136 50414
0 50416 5 1 1 50415
0 50417 7 1 2 50411 50416
0 50418 5 1 1 50417
0 50419 7 1 2 94658 50418
0 50420 5 1 1 50419
0 50421 7 1 2 79867 95556
0 50422 5 1 1 50421
0 50423 7 1 2 61728 74491
0 50424 7 1 2 80022 50423
0 50425 7 1 2 94303 50424
0 50426 5 1 1 50425
0 50427 7 1 2 50422 50426
0 50428 7 1 2 50420 50427
0 50429 7 1 2 50409 50428
0 50430 5 1 1 50429
0 50431 7 1 2 74161 50430
0 50432 5 1 1 50431
0 50433 7 1 2 86095 94844
0 50434 7 1 2 85283 50433
0 50435 5 1 1 50434
0 50436 7 1 2 50432 50435
0 50437 5 1 1 50436
0 50438 7 1 2 61986 50437
0 50439 5 1 1 50438
0 50440 7 1 2 74138 89188
0 50441 7 1 2 80122 50440
0 50442 5 1 1 50441
0 50443 7 1 2 73703 83536
0 50444 7 1 2 93831 50443
0 50445 5 1 1 50444
0 50446 7 1 2 50442 50445
0 50447 5 1 1 50446
0 50448 7 1 2 61729 95430
0 50449 7 1 2 50447 50448
0 50450 5 1 1 50449
0 50451 7 1 2 50439 50450
0 50452 7 1 2 50395 50451
0 50453 5 1 1 50452
0 50454 7 1 2 76483 50453
0 50455 5 1 1 50454
0 50456 7 1 2 59032 94393
0 50457 5 1 1 50456
0 50458 7 1 2 50457 47745
0 50459 5 1 1 50458
0 50460 7 1 2 58898 50459
0 50461 5 1 1 50460
0 50462 7 1 2 40204 50461
0 50463 5 1 1 50462
0 50464 7 1 2 59678 94856
0 50465 7 1 2 50463 50464
0 50466 5 2 1 50465
0 50467 7 1 2 70582 95546
0 50468 5 1 1 50467
0 50469 7 1 2 86112 74300
0 50470 7 1 2 76850 50469
0 50471 5 1 1 50470
0 50472 7 1 2 50468 50471
0 50473 5 1 1 50472
0 50474 7 1 2 66373 50473
0 50475 5 1 1 50474
0 50476 7 1 2 95614 50475
0 50477 5 1 1 50476
0 50478 7 1 2 62135 50477
0 50479 5 1 1 50478
0 50480 7 3 2 66079 70878
0 50481 5 1 1 95616
0 50482 7 1 2 59679 72203
0 50483 5 1 1 50482
0 50484 7 2 2 50481 50483
0 50485 5 2 1 95619
0 50486 7 1 2 90287 95548
0 50487 7 1 2 95621 50486
0 50488 5 1 1 50487
0 50489 7 1 2 50479 50488
0 50490 5 1 1 50489
0 50491 7 1 2 85303 50490
0 50492 5 1 1 50491
0 50493 7 1 2 74080 95620
0 50494 5 1 1 50493
0 50495 7 1 2 70561 94916
0 50496 5 1 1 50495
0 50497 7 1 2 82885 72573
0 50498 5 1 1 50497
0 50499 7 1 2 50496 50498
0 50500 5 1 1 50499
0 50501 7 1 2 50494 50500
0 50502 5 1 1 50501
0 50503 7 1 2 90251 95599
0 50504 5 1 1 50503
0 50505 7 2 2 61987 85304
0 50506 7 1 2 81512 67940
0 50507 7 1 2 95623 50506
0 50508 5 1 1 50507
0 50509 7 1 2 50504 50508
0 50510 5 1 1 50509
0 50511 7 1 2 75790 50510
0 50512 5 1 1 50511
0 50513 7 1 2 81570 84606
0 50514 5 1 1 50513
0 50515 7 1 2 66080 94917
0 50516 5 1 1 50515
0 50517 7 1 2 50514 50516
0 50518 5 1 1 50517
0 50519 7 1 2 72608 50518
0 50520 5 1 1 50519
0 50521 7 1 2 50512 50520
0 50522 7 1 2 95615 50521
0 50523 5 1 1 50522
0 50524 7 1 2 62136 50523
0 50525 5 1 1 50524
0 50526 7 1 2 50502 50525
0 50527 5 1 1 50526
0 50528 7 1 2 59936 50527
0 50529 5 1 1 50528
0 50530 7 1 2 83169 82107
0 50531 7 1 2 95558 50530
0 50532 5 1 1 50531
0 50533 7 1 2 85325 82663
0 50534 7 1 2 95522 50533
0 50535 5 1 1 50534
0 50536 7 1 2 50532 50535
0 50537 5 1 1 50536
0 50538 7 1 2 90549 50537
0 50539 5 1 1 50538
0 50540 7 1 2 50529 50539
0 50541 7 1 2 50492 50540
0 50542 5 1 1 50541
0 50543 7 1 2 66949 50542
0 50544 5 1 1 50543
0 50545 7 1 2 72204 79989
0 50546 7 1 2 90637 50545
0 50547 5 1 1 50546
0 50548 7 1 2 74076 82422
0 50549 7 1 2 94444 50548
0 50550 7 1 2 95624 50549
0 50551 5 1 1 50550
0 50552 7 1 2 50547 50551
0 50553 5 1 1 50552
0 50554 7 1 2 79978 50553
0 50555 5 1 1 50554
0 50556 7 1 2 82281 95014
0 50557 5 1 1 50556
0 50558 7 1 2 66639 72205
0 50559 7 1 2 95408 50558
0 50560 5 1 1 50559
0 50561 7 1 2 50557 50560
0 50562 5 1 1 50561
0 50563 7 1 2 70540 50562
0 50564 5 1 1 50563
0 50565 7 1 2 79189 74488
0 50566 5 1 1 50565
0 50567 7 1 2 87107 86676
0 50568 7 1 2 76588 50567
0 50569 5 1 1 50568
0 50570 7 1 2 50566 50569
0 50571 5 1 1 50570
0 50572 7 1 2 83051 50571
0 50573 5 1 1 50572
0 50574 7 1 2 50564 50573
0 50575 5 1 1 50574
0 50576 7 1 2 83170 50575
0 50577 5 1 1 50576
0 50578 7 1 2 50555 50577
0 50579 5 1 1 50578
0 50580 7 1 2 59680 50579
0 50581 5 1 1 50580
0 50582 7 1 2 87511 82423
0 50583 7 1 2 92042 50582
0 50584 5 1 1 50583
0 50585 7 1 2 61470 93994
0 50586 5 1 1 50585
0 50587 7 1 2 86334 67941
0 50588 7 1 2 50586 50587
0 50589 5 1 1 50588
0 50590 7 1 2 50584 50589
0 50591 5 1 1 50590
0 50592 7 1 2 58805 50591
0 50593 5 1 1 50592
0 50594 7 1 2 84607 94955
0 50595 5 1 1 50594
0 50596 7 1 2 91385 94511
0 50597 5 1 1 50596
0 50598 7 1 2 50595 50597
0 50599 5 1 1 50598
0 50600 7 1 2 67942 50599
0 50601 5 1 1 50600
0 50602 7 1 2 50593 50601
0 50603 5 1 1 50602
0 50604 7 1 2 83171 50603
0 50605 5 1 1 50604
0 50606 7 1 2 58899 76611
0 50607 7 1 2 68804 79561
0 50608 7 1 2 50606 50607
0 50609 7 1 2 91201 50608
0 50610 5 1 1 50609
0 50611 7 1 2 50605 50610
0 50612 5 1 1 50611
0 50613 7 1 2 61988 50612
0 50614 5 1 1 50613
0 50615 7 1 2 87108 82263
0 50616 5 1 1 50615
0 50617 7 1 2 75741 84590
0 50618 5 1 1 50617
0 50619 7 1 2 50616 50618
0 50620 5 1 1 50619
0 50621 7 1 2 94528 50620
0 50622 5 1 1 50621
0 50623 7 1 2 73269 82108
0 50624 7 1 2 91330 50623
0 50625 5 1 1 50624
0 50626 7 1 2 50622 50625
0 50627 5 1 1 50626
0 50628 7 1 2 70541 50627
0 50629 5 1 1 50628
0 50630 7 2 2 83947 86297
0 50631 7 2 2 91412 95625
0 50632 7 1 2 59033 95627
0 50633 5 1 1 50632
0 50634 7 1 2 61098 94649
0 50635 5 1 1 50634
0 50636 7 1 2 50633 50635
0 50637 5 1 1 50636
0 50638 7 1 2 87580 84537
0 50639 7 1 2 50637 50638
0 50640 5 1 1 50639
0 50641 7 1 2 50629 50640
0 50642 5 1 1 50641
0 50643 7 1 2 94857 50642
0 50644 5 1 1 50643
0 50645 7 1 2 50614 50644
0 50646 7 1 2 50581 50645
0 50647 5 1 1 50646
0 50648 7 1 2 62137 50647
0 50649 5 1 1 50648
0 50650 7 1 2 70940 74197
0 50651 5 1 1 50650
0 50652 7 1 2 77998 84919
0 50653 5 1 1 50652
0 50654 7 1 2 50651 50653
0 50655 5 1 1 50654
0 50656 7 2 2 87269 67541
0 50657 7 1 2 50655 95629
0 50658 5 1 1 50657
0 50659 7 1 2 83172 82435
0 50660 7 1 2 91157 50659
0 50661 5 1 1 50660
0 50662 7 1 2 50658 50661
0 50663 5 1 1 50662
0 50664 7 1 2 66081 50663
0 50665 5 1 1 50664
0 50666 7 1 2 67601 92601
0 50667 7 1 2 86657 50666
0 50668 5 1 1 50667
0 50669 7 1 2 50665 50668
0 50670 5 1 1 50669
0 50671 7 1 2 86073 50670
0 50672 5 1 1 50671
0 50673 7 1 2 73983 87429
0 50674 7 1 2 82120 94673
0 50675 7 1 2 50673 50674
0 50676 5 1 1 50675
0 50677 7 1 2 74815 87554
0 50678 7 1 2 95617 50677
0 50679 5 1 1 50678
0 50680 7 1 2 82334 82424
0 50681 7 1 2 95622 50680
0 50682 5 1 1 50681
0 50683 7 1 2 50679 50682
0 50684 5 1 1 50683
0 50685 7 1 2 63550 50684
0 50686 5 1 1 50685
0 50687 7 1 2 94965 95533
0 50688 5 1 1 50687
0 50689 7 1 2 50686 50688
0 50690 5 1 1 50689
0 50691 7 1 2 61989 83173
0 50692 7 1 2 50690 50691
0 50693 5 1 1 50692
0 50694 7 1 2 50676 50693
0 50695 5 1 1 50694
0 50696 7 1 2 69282 50695
0 50697 5 1 1 50696
0 50698 7 1 2 50672 50697
0 50699 7 1 2 50649 50698
0 50700 7 1 2 50544 50699
0 50701 7 1 2 50455 50700
0 50702 5 1 1 50701
0 50703 7 1 2 88310 50702
0 50704 5 1 1 50703
0 50705 7 1 2 76484 72585
0 50706 7 1 2 86324 50705
0 50707 7 1 2 82285 88154
0 50708 7 1 2 50706 50707
0 50709 7 1 2 94298 50708
0 50710 5 1 1 50709
0 50711 7 1 2 50704 50710
0 50712 5 1 1 50711
0 50713 7 1 2 71917 50712
0 50714 5 1 1 50713
0 50715 7 1 2 83099 88751
0 50716 7 1 2 95566 50715
0 50717 7 1 2 94839 50716
0 50718 5 1 1 50717
0 50719 7 1 2 57799 92497
0 50720 7 1 2 89347 50719
0 50721 5 1 1 50720
0 50722 7 1 2 50718 50721
0 50723 5 1 1 50722
0 50724 7 1 2 83394 50723
0 50725 5 1 1 50724
0 50726 7 1 2 17741 92722
0 50727 5 1 1 50726
0 50728 7 1 2 94699 50727
0 50729 5 1 1 50728
0 50730 7 1 2 68643 95447
0 50731 5 1 1 50730
0 50732 7 1 2 57518 95384
0 50733 5 1 1 50732
0 50734 7 1 2 50731 50733
0 50735 5 1 1 50734
0 50736 7 1 2 83174 50735
0 50737 5 1 1 50736
0 50738 7 1 2 50729 50737
0 50739 5 1 1 50738
0 50740 7 1 2 72711 70542
0 50741 7 1 2 94768 50740
0 50742 7 1 2 50739 50741
0 50743 5 1 1 50742
0 50744 7 1 2 50725 50743
0 50745 5 1 1 50744
0 50746 7 1 2 66640 50745
0 50747 5 1 1 50746
0 50748 7 1 2 83025 88311
0 50749 7 1 2 87392 50748
0 50750 7 1 2 72748 94356
0 50751 7 1 2 50749 50750
0 50752 5 1 1 50751
0 50753 7 1 2 50747 50752
0 50754 5 1 1 50753
0 50755 7 1 2 73447 50754
0 50756 5 1 1 50755
0 50757 7 1 2 59034 89478
0 50758 7 1 2 91659 50757
0 50759 7 1 2 95458 50758
0 50760 5 1 1 50759
0 50761 7 2 2 83007 95207
0 50762 7 1 2 64844 72405
0 50763 5 1 1 50762
0 50764 7 1 2 71967 94885
0 50765 7 1 2 50763 50764
0 50766 7 1 2 95631 50765
0 50767 5 1 1 50766
0 50768 7 1 2 50760 50767
0 50769 5 1 1 50768
0 50770 7 1 2 63654 50769
0 50771 5 1 1 50770
0 50772 7 1 2 87837 94668
0 50773 5 1 1 50772
0 50774 7 1 2 76034 95632
0 50775 5 1 1 50774
0 50776 7 1 2 50773 50775
0 50777 5 1 1 50776
0 50778 7 1 2 66374 82038
0 50779 7 1 2 50777 50778
0 50780 5 1 1 50779
0 50781 7 1 2 50771 50780
0 50782 5 1 1 50781
0 50783 7 1 2 88312 50782
0 50784 5 1 1 50783
0 50785 7 1 2 81757 83008
0 50786 7 1 2 95438 50785
0 50787 5 1 1 50786
0 50788 7 1 2 50784 50787
0 50789 5 1 1 50788
0 50790 7 1 2 76485 50789
0 50791 5 1 1 50790
0 50792 7 1 2 84023 95064
0 50793 5 1 1 50792
0 50794 7 1 2 85197 18574
0 50795 5 1 1 50794
0 50796 7 1 2 83175 50795
0 50797 5 1 1 50796
0 50798 7 1 2 79916 87838
0 50799 5 1 1 50798
0 50800 7 1 2 50797 50799
0 50801 5 1 1 50800
0 50802 7 1 2 58900 50801
0 50803 5 1 1 50802
0 50804 7 1 2 76612 74168
0 50805 7 1 2 94868 50804
0 50806 5 1 1 50805
0 50807 7 1 2 50803 50806
0 50808 5 1 1 50807
0 50809 7 1 2 76569 82425
0 50810 7 1 2 50808 50809
0 50811 5 1 1 50810
0 50812 7 1 2 50793 50811
0 50813 5 1 1 50812
0 50814 7 1 2 62138 50813
0 50815 5 1 1 50814
0 50816 7 1 2 76570 80035
0 50817 5 1 1 50816
0 50818 7 1 2 79933 92362
0 50819 5 1 1 50818
0 50820 7 1 2 50817 50819
0 50821 5 1 1 50820
0 50822 7 1 2 66375 50821
0 50823 5 1 1 50822
0 50824 7 1 2 79190 91596
0 50825 5 1 1 50824
0 50826 7 1 2 50823 50825
0 50827 5 1 1 50826
0 50828 7 1 2 94700 50827
0 50829 5 1 1 50828
0 50830 7 1 2 78914 80463
0 50831 7 1 2 95449 50830
0 50832 5 1 1 50831
0 50833 7 1 2 50829 50832
0 50834 7 1 2 50815 50833
0 50835 5 1 1 50834
0 50836 7 1 2 61990 50835
0 50837 5 1 1 50836
0 50838 7 1 2 94784 95466
0 50839 5 1 1 50838
0 50840 7 1 2 95464 50839
0 50841 5 1 1 50840
0 50842 7 1 2 61730 50841
0 50843 5 1 1 50842
0 50844 7 1 2 83026 73407
0 50845 7 1 2 79815 50844
0 50846 7 1 2 94324 50845
0 50847 5 1 1 50846
0 50848 7 1 2 50843 50847
0 50849 5 1 1 50848
0 50850 7 1 2 66641 70879
0 50851 7 1 2 50849 50850
0 50852 5 1 1 50851
0 50853 7 1 2 50837 50852
0 50854 5 1 1 50853
0 50855 7 1 2 88313 50854
0 50856 5 1 1 50855
0 50857 7 1 2 50791 50856
0 50858 5 1 1 50857
0 50859 7 1 2 64414 76285
0 50860 5 1 1 50859
0 50861 7 1 2 50858 50860
0 50862 5 1 1 50861
0 50863 7 1 2 50756 50862
0 50864 7 1 2 50714 50863
0 50865 7 1 2 50346 50864
0 50866 7 1 2 49885 50865
0 50867 7 1 2 48798 50866
0 50868 7 1 2 46668 50867
0 50869 7 1 2 44098 50868
0 50870 5 1 1 50869
0 50871 7 1 2 66534 50870
0 50872 5 1 1 50871
0 50873 7 2 2 84787 79462
0 50874 7 1 2 94326 95633
0 50875 5 1 1 50874
0 50876 7 1 2 88275 93776
0 50877 5 1 1 50876
0 50878 7 1 2 90556 95030
0 50879 5 1 1 50878
0 50880 7 1 2 50877 50879
0 50881 5 1 1 50880
0 50882 7 1 2 80870 50881
0 50883 5 1 1 50882
0 50884 7 1 2 50875 50883
0 50885 5 1 1 50884
0 50886 7 1 2 63412 50885
0 50887 5 1 1 50886
0 50888 7 1 2 88249 91607
0 50889 7 1 2 93016 50888
0 50890 5 1 1 50889
0 50891 7 1 2 50887 50890
0 50892 5 1 1 50891
0 50893 7 1 2 64638 50892
0 50894 5 1 1 50893
0 50895 7 1 2 86653 94721
0 50896 5 1 1 50895
0 50897 7 1 2 50894 50896
0 50898 5 1 1 50897
0 50899 7 1 2 80523 50898
0 50900 5 1 1 50899
0 50901 7 1 2 80308 94632
0 50902 5 1 1 50901
0 50903 7 1 2 65096 85715
0 50904 5 1 1 50903
0 50905 7 1 2 89034 50904
0 50906 5 1 1 50905
0 50907 7 1 2 73327 50906
0 50908 5 1 1 50907
0 50909 7 1 2 38275 50908
0 50910 5 1 1 50909
0 50911 7 1 2 76887 50910
0 50912 5 1 1 50911
0 50913 7 1 2 50902 50912
0 50914 5 1 1 50913
0 50915 7 1 2 72800 87270
0 50916 7 1 2 50914 50915
0 50917 5 1 1 50916
0 50918 7 1 2 50900 50917
0 50919 5 1 1 50918
0 50920 7 1 2 75965 50919
0 50921 5 1 1 50920
0 50922 7 1 2 63108 93241
0 50923 5 1 1 50922
0 50924 7 1 2 57519 50923
0 50925 5 1 1 50924
0 50926 7 2 2 75879 73179
0 50927 5 1 1 95635
0 50928 7 1 2 71752 95636
0 50929 5 1 1 50928
0 50930 7 1 2 70259 92756
0 50931 5 1 1 50930
0 50932 7 1 2 73180 81282
0 50933 5 2 1 50932
0 50934 7 1 2 50931 95637
0 50935 7 1 2 50929 50934
0 50936 7 1 2 50925 50935
0 50937 5 1 1 50936
0 50938 7 1 2 58672 50937
0 50939 5 1 1 50938
0 50940 7 1 2 57520 81531
0 50941 7 1 2 72416 50940
0 50942 5 1 1 50941
0 50943 7 1 2 50939 50942
0 50944 5 1 1 50943
0 50945 7 1 2 61731 50944
0 50946 5 1 1 50945
0 50947 7 1 2 70247 50927
0 50948 5 1 1 50947
0 50949 7 1 2 77159 50948
0 50950 5 1 1 50949
0 50951 7 1 2 70972 70260
0 50952 5 1 1 50951
0 50953 7 1 2 95638 50952
0 50954 7 1 2 50950 50953
0 50955 5 1 1 50954
0 50956 7 1 2 82218 50955
0 50957 5 1 1 50956
0 50958 7 1 2 50946 50957
0 50959 5 1 1 50958
0 50960 7 1 2 58076 50959
0 50961 5 1 1 50960
0 50962 7 2 2 59385 80948
0 50963 5 1 1 95639
0 50964 7 1 2 65727 95640
0 50965 5 2 1 50964
0 50966 7 1 2 76271 95641
0 50967 5 1 1 50966
0 50968 7 1 2 58077 50967
0 50969 5 1 1 50968
0 50970 7 1 2 86914 50969
0 50971 5 1 1 50970
0 50972 7 1 2 78615 50971
0 50973 5 1 1 50972
0 50974 7 1 2 82485 81635
0 50975 5 1 1 50974
0 50976 7 1 2 61732 87074
0 50977 7 1 2 50975 50976
0 50978 7 1 2 50973 50977
0 50979 5 1 1 50978
0 50980 7 1 2 68271 80530
0 50981 5 1 1 50980
0 50982 7 1 2 3363 50981
0 50983 5 1 1 50982
0 50984 7 1 2 62273 50983
0 50985 5 1 1 50984
0 50986 7 1 2 66376 5800
0 50987 7 1 2 50985 50986
0 50988 5 1 1 50987
0 50989 7 1 2 59937 50988
0 50990 7 1 2 50979 50989
0 50991 5 1 1 50990
0 50992 7 1 2 86917 81264
0 50993 5 1 1 50992
0 50994 7 1 2 94319 43542
0 50995 5 1 1 50994
0 50996 7 1 2 50993 50995
0 50997 5 1 1 50996
0 50998 7 1 2 73181 50997
0 50999 5 1 1 50998
0 51000 7 1 2 71753 87440
0 51001 5 1 1 51000
0 51002 7 1 2 17716 51001
0 51003 5 1 1 51002
0 51004 7 1 2 75880 51003
0 51005 5 1 1 51004
0 51006 7 1 2 87292 80580
0 51007 5 1 1 51006
0 51008 7 1 2 81265 51007
0 51009 5 1 1 51008
0 51010 7 1 2 51005 51009
0 51011 5 1 1 51010
0 51012 7 1 2 70261 51011
0 51013 5 1 1 51012
0 51014 7 1 2 73182 94320
0 51015 5 1 1 51014
0 51016 7 1 2 86850 95496
0 51017 7 1 2 70262 51016
0 51018 5 1 1 51017
0 51019 7 1 2 51015 51018
0 51020 5 1 1 51019
0 51021 7 1 2 81604 51020
0 51022 5 1 1 51021
0 51023 7 1 2 70263 84341
0 51024 5 1 1 51023
0 51025 7 1 2 70242 81192
0 51026 7 1 2 51024 51025
0 51027 5 1 1 51026
0 51028 7 1 2 86808 82433
0 51029 7 1 2 51027 51028
0 51030 5 1 1 51029
0 51031 7 1 2 51022 51030
0 51032 7 1 2 51013 51031
0 51033 7 1 2 50999 51032
0 51034 7 1 2 50991 51033
0 51035 7 1 2 50961 51034
0 51036 5 1 1 51035
0 51037 7 1 2 59681 51036
0 51038 5 1 1 51037
0 51039 7 1 2 6113 81544
0 51040 5 2 1 51039
0 51041 7 1 2 75493 95643
0 51042 5 1 1 51041
0 51043 7 1 2 84920 84904
0 51044 5 1 1 51043
0 51045 7 1 2 51042 51044
0 51046 5 1 1 51045
0 51047 7 1 2 58357 51046
0 51048 5 1 1 51047
0 51049 7 1 2 84921 84911
0 51050 5 1 1 51049
0 51051 7 1 2 51048 51050
0 51052 5 1 1 51051
0 51053 7 1 2 75597 51052
0 51054 5 1 1 51053
0 51055 7 1 2 75494 73907
0 51056 5 1 1 51055
0 51057 7 1 2 65097 93992
0 51058 5 1 1 51057
0 51059 7 1 2 68175 72498
0 51060 7 1 2 51058 51059
0 51061 7 1 2 51056 51060
0 51062 5 1 1 51061
0 51063 7 1 2 76662 51062
0 51064 5 1 1 51063
0 51065 7 1 2 61733 51064
0 51066 7 1 2 51054 51065
0 51067 5 1 1 51066
0 51068 7 1 2 77238 95644
0 51069 5 1 1 51068
0 51070 7 1 2 73908 94513
0 51071 5 1 1 51070
0 51072 7 1 2 51069 51071
0 51073 5 1 1 51072
0 51074 7 1 2 75791 51073
0 51075 5 1 1 51074
0 51076 7 1 2 77836 27945
0 51077 5 1 1 51076
0 51078 7 1 2 68805 51077
0 51079 5 1 1 51078
0 51080 7 1 2 94419 51079
0 51081 5 1 1 51080
0 51082 7 1 2 65728 51081
0 51083 5 1 1 51082
0 51084 7 1 2 68048 94514
0 51085 5 1 1 51084
0 51086 7 1 2 66377 51085
0 51087 7 1 2 51083 51086
0 51088 7 1 2 51075 51087
0 51089 5 1 1 51088
0 51090 7 1 2 51067 51089
0 51091 5 1 1 51090
0 51092 7 1 2 73941 82347
0 51093 5 1 1 51092
0 51094 7 1 2 83962 51093
0 51095 5 1 1 51094
0 51096 7 1 2 80771 51095
0 51097 5 1 1 51096
0 51098 7 1 2 67225 82349
0 51099 5 1 1 51098
0 51100 7 1 2 76663 51099
0 51101 5 1 1 51100
0 51102 7 1 2 61734 51101
0 51103 7 1 2 51097 51102
0 51104 5 1 1 51103
0 51105 7 1 2 85566 75719
0 51106 5 1 1 51105
0 51107 7 1 2 81078 51106
0 51108 5 1 1 51107
0 51109 7 1 2 77239 51108
0 51110 5 1 1 51109
0 51111 7 1 2 64108 83088
0 51112 5 1 1 51111
0 51113 7 1 2 94515 51112
0 51114 5 1 1 51113
0 51115 7 1 2 66378 51114
0 51116 7 1 2 51110 51115
0 51117 5 1 1 51116
0 51118 7 1 2 71918 51117
0 51119 7 1 2 51104 51118
0 51120 5 1 1 51119
0 51121 7 1 2 85305 82608
0 51122 5 1 1 51121
0 51123 7 2 2 91887 51122
0 51124 5 1 1 95645
0 51125 7 1 2 43617 95646
0 51126 5 1 1 51125
0 51127 7 1 2 65729 51126
0 51128 5 1 1 51127
0 51129 7 1 2 82604 91790
0 51130 5 1 1 51129
0 51131 7 1 2 75881 94186
0 51132 7 1 2 51130 51131
0 51133 5 1 1 51132
0 51134 7 1 2 82614 91884
0 51135 7 1 2 51133 51134
0 51136 5 1 1 51135
0 51137 7 1 2 86144 51136
0 51138 5 1 1 51137
0 51139 7 1 2 51128 51138
0 51140 5 1 1 51139
0 51141 7 1 2 68644 51140
0 51142 5 1 1 51141
0 51143 7 1 2 65730 90755
0 51144 5 1 1 51143
0 51145 7 1 2 63109 51144
0 51146 5 1 1 51145
0 51147 7 1 2 95515 51146
0 51148 5 1 1 51147
0 51149 7 1 2 51142 51148
0 51150 7 1 2 51120 51149
0 51151 7 1 2 51091 51150
0 51152 7 1 2 51038 51151
0 51153 5 1 1 51152
0 51154 7 1 2 66082 51153
0 51155 5 1 1 51154
0 51156 7 1 2 87516 91875
0 51157 5 1 1 51156
0 51158 7 1 2 68806 51157
0 51159 5 1 1 51158
0 51160 7 1 2 94429 51159
0 51161 5 1 1 51160
0 51162 7 1 2 82972 51161
0 51163 5 1 1 51162
0 51164 7 1 2 85764 84068
0 51165 5 1 1 51164
0 51166 7 1 2 79650 91965
0 51167 5 1 1 51166
0 51168 7 1 2 51165 51167
0 51169 5 1 1 51168
0 51170 7 1 2 65339 51169
0 51171 5 1 1 51170
0 51172 7 1 2 51163 51171
0 51173 5 1 1 51172
0 51174 7 1 2 68413 51173
0 51175 5 1 1 51174
0 51176 7 1 2 81218 94981
0 51177 5 1 1 51176
0 51178 7 1 2 94430 51177
0 51179 5 1 1 51178
0 51180 7 1 2 82973 51179
0 51181 5 1 1 51180
0 51182 7 1 2 84483 90356
0 51183 5 1 1 51182
0 51184 7 2 2 85808 81475
0 51185 5 1 1 95647
0 51186 7 1 2 93955 95648
0 51187 5 1 1 51186
0 51188 7 1 2 51183 51187
0 51189 7 1 2 51181 51188
0 51190 5 1 1 51189
0 51191 7 1 2 68807 51190
0 51192 5 1 1 51191
0 51193 7 1 2 69430 82585
0 51194 5 1 1 51193
0 51195 7 1 2 87517 51194
0 51196 5 2 1 51195
0 51197 7 1 2 85921 95649
0 51198 5 1 1 51197
0 51199 7 1 2 83043 95234
0 51200 5 1 1 51199
0 51201 7 1 2 70103 51200
0 51202 5 1 1 51201
0 51203 7 1 2 51198 51202
0 51204 7 1 2 51192 51203
0 51205 7 1 2 51175 51204
0 51206 5 1 1 51205
0 51207 7 1 2 67387 51206
0 51208 5 1 1 51207
0 51209 7 1 2 82974 87346
0 51210 5 1 1 51209
0 51211 7 1 2 95235 51210
0 51212 5 1 1 51211
0 51213 7 1 2 68414 51212
0 51214 5 1 1 51213
0 51215 7 2 2 85809 87434
0 51216 7 1 2 72530 95651
0 51217 5 1 1 51216
0 51218 7 1 2 91876 51217
0 51219 5 1 1 51218
0 51220 7 1 2 59682 51219
0 51221 5 1 1 51220
0 51222 7 1 2 81450 91786
0 51223 5 1 1 51222
0 51224 7 1 2 59683 95485
0 51225 5 1 1 51224
0 51226 7 1 2 51223 51225
0 51227 5 1 1 51226
0 51228 7 1 2 65340 51227
0 51229 5 1 1 51228
0 51230 7 1 2 51221 51229
0 51231 5 1 1 51230
0 51232 7 1 2 58358 51231
0 51233 5 1 1 51232
0 51234 7 1 2 51214 51233
0 51235 5 1 1 51234
0 51236 7 1 2 68049 51235
0 51237 5 1 1 51236
0 51238 7 1 2 73234 90357
0 51239 5 1 1 51238
0 51240 7 1 2 51185 51239
0 51241 5 1 1 51240
0 51242 7 1 2 85267 51241
0 51243 5 1 1 51242
0 51244 7 1 2 84685 95434
0 51245 5 1 1 51244
0 51246 7 1 2 58673 95650
0 51247 5 1 1 51246
0 51248 7 1 2 51245 51247
0 51249 7 1 2 51243 51248
0 51250 5 1 1 51249
0 51251 7 1 2 70435 51250
0 51252 5 1 1 51251
0 51253 7 1 2 85268 86280
0 51254 5 1 1 51253
0 51255 7 1 2 94420 51254
0 51256 5 1 1 51255
0 51257 7 1 2 66379 51256
0 51258 5 1 1 51257
0 51259 7 1 2 69431 89362
0 51260 5 1 1 51259
0 51261 7 1 2 51258 51260
0 51262 5 1 1 51261
0 51263 7 1 2 59684 51262
0 51264 5 1 1 51263
0 51265 7 1 2 85137 87347
0 51266 5 1 1 51265
0 51267 7 1 2 82426 92887
0 51268 5 1 1 51267
0 51269 7 1 2 51266 51268
0 51270 5 1 1 51269
0 51271 7 1 2 90756 51270
0 51272 5 1 1 51271
0 51273 7 1 2 83822 91901
0 51274 7 1 2 95128 51273
0 51275 5 1 1 51274
0 51276 7 1 2 51272 51275
0 51277 7 1 2 51264 51276
0 51278 7 1 2 51252 51277
0 51279 7 1 2 51237 51278
0 51280 7 1 2 51208 51279
0 51281 5 1 1 51280
0 51282 7 1 2 65731 51281
0 51283 5 1 1 51282
0 51284 7 1 2 72824 95237
0 51285 5 1 1 51284
0 51286 7 1 2 85184 51285
0 51287 5 1 1 51286
0 51288 7 1 2 61735 51287
0 51289 5 1 1 51288
0 51290 7 3 2 71543 87207
0 51291 5 1 1 95653
0 51292 7 1 2 51289 51291
0 51293 5 1 1 51292
0 51294 7 1 2 57800 51293
0 51295 5 1 1 51294
0 51296 7 1 2 68808 87208
0 51297 5 1 1 51296
0 51298 7 1 2 86825 51297
0 51299 5 1 1 51298
0 51300 7 1 2 71544 51299
0 51301 5 1 1 51300
0 51302 7 1 2 51295 51301
0 51303 5 1 1 51302
0 51304 7 1 2 59938 51303
0 51305 5 1 1 51304
0 51306 7 2 2 75792 84591
0 51307 7 1 2 85138 95656
0 51308 5 1 1 51307
0 51309 7 1 2 51305 51308
0 51310 5 1 1 51309
0 51311 7 1 2 72249 51310
0 51312 5 1 1 51311
0 51313 7 3 2 65098 84686
0 51314 5 2 1 95658
0 51315 7 1 2 78090 95659
0 51316 5 2 1 51315
0 51317 7 1 2 91885 95663
0 51318 5 1 1 51317
0 51319 7 1 2 70436 51318
0 51320 5 1 1 51319
0 51321 7 1 2 59685 51124
0 51322 5 1 1 51321
0 51323 7 1 2 51320 51322
0 51324 5 1 1 51323
0 51325 7 1 2 65732 51324
0 51326 5 1 1 51325
0 51327 7 1 2 82599 94399
0 51328 5 2 1 51327
0 51329 7 1 2 71545 95665
0 51330 5 1 1 51329
0 51331 7 1 2 70062 74139
0 51332 7 1 2 81349 51331
0 51333 5 1 1 51332
0 51334 7 1 2 51330 51333
0 51335 5 1 1 51334
0 51336 7 1 2 58674 51335
0 51337 5 1 1 51336
0 51338 7 2 2 72848 87209
0 51339 7 1 2 71546 95667
0 51340 5 1 1 51339
0 51341 7 1 2 51337 51340
0 51342 5 1 1 51341
0 51343 7 1 2 67388 51342
0 51344 5 1 1 51343
0 51345 7 1 2 82975 82609
0 51346 5 1 1 51345
0 51347 7 1 2 51346 95664
0 51348 5 1 1 51347
0 51349 7 1 2 73880 51348
0 51350 5 1 1 51349
0 51351 7 1 2 78274 95668
0 51352 5 1 1 51351
0 51353 7 1 2 68050 82976
0 51354 5 1 1 51353
0 51355 7 2 2 85185 51354
0 51356 5 3 1 95669
0 51357 7 1 2 95671 95666
0 51358 5 1 1 51357
0 51359 7 1 2 51352 51358
0 51360 7 1 2 51350 51359
0 51361 5 1 1 51360
0 51362 7 1 2 75882 51361
0 51363 5 1 1 51362
0 51364 7 1 2 51344 51363
0 51365 7 1 2 51326 51364
0 51366 5 1 1 51365
0 51367 7 1 2 68645 51366
0 51368 5 1 1 51367
0 51369 7 1 2 57801 84592
0 51370 5 1 1 51369
0 51371 7 1 2 91877 51370
0 51372 5 1 1 51371
0 51373 7 1 2 68809 51372
0 51374 5 1 1 51373
0 51375 7 1 2 72849 95497
0 51376 5 2 1 51375
0 51377 7 1 2 51374 95674
0 51378 5 1 1 51377
0 51379 7 1 2 51378 95672
0 51380 5 1 1 51379
0 51381 7 1 2 81272 87218
0 51382 5 2 1 51381
0 51383 7 1 2 84292 95676
0 51384 5 1 1 51383
0 51385 7 1 2 75720 84593
0 51386 7 1 2 78275 51385
0 51387 5 1 1 51386
0 51388 7 1 2 51384 51387
0 51389 5 1 1 51388
0 51390 7 1 2 59939 51389
0 51391 5 1 1 51390
0 51392 7 1 2 67389 85139
0 51393 7 1 2 84594 51392
0 51394 5 1 1 51393
0 51395 7 1 2 51391 51394
0 51396 7 1 2 51380 51395
0 51397 5 1 1 51396
0 51398 7 1 2 71919 51397
0 51399 5 1 1 51398
0 51400 7 1 2 57802 94942
0 51401 5 1 1 51400
0 51402 7 1 2 91878 51401
0 51403 5 1 1 51402
0 51404 7 1 2 58078 51403
0 51405 5 1 1 51404
0 51406 7 1 2 58079 87210
0 51407 5 1 1 51406
0 51408 7 1 2 95675 51407
0 51409 5 1 1 51408
0 51410 7 1 2 68810 51409
0 51411 5 1 1 51410
0 51412 7 1 2 51405 51411
0 51413 5 1 1 51412
0 51414 7 1 2 82977 72007
0 51415 5 1 1 51414
0 51416 7 1 2 85186 51415
0 51417 5 1 1 51416
0 51418 7 1 2 51413 51417
0 51419 5 1 1 51418
0 51420 7 1 2 71226 95516
0 51421 5 1 1 51420
0 51422 7 1 2 80638 95654
0 51423 5 1 1 51422
0 51424 7 1 2 78186 95657
0 51425 5 1 1 51424
0 51426 7 1 2 83432 95677
0 51427 5 1 1 51426
0 51428 7 1 2 51425 51427
0 51429 5 1 1 51428
0 51430 7 1 2 59940 51429
0 51431 5 1 1 51430
0 51432 7 1 2 51423 51431
0 51433 5 1 1 51432
0 51434 7 1 2 58080 51433
0 51435 5 1 1 51434
0 51436 7 1 2 51421 51435
0 51437 7 1 2 51419 51436
0 51438 7 1 2 51399 51437
0 51439 7 1 2 51368 51438
0 51440 7 1 2 51312 51439
0 51441 7 1 2 51283 51440
0 51442 7 1 2 51155 51441
0 51443 5 1 1 51442
0 51444 7 1 2 63551 51443
0 51445 5 1 1 51444
0 51446 7 1 2 58081 86768
0 51447 5 1 1 51446
0 51448 7 1 2 3410 51447
0 51449 5 1 1 51448
0 51450 7 1 2 82496 51449
0 51451 5 1 1 51450
0 51452 7 1 2 85578 77531
0 51453 5 1 1 51452
0 51454 7 1 2 78690 68904
0 51455 5 1 1 51454
0 51456 7 1 2 80153 51455
0 51457 5 1 1 51456
0 51458 7 1 2 68051 51457
0 51459 5 1 1 51458
0 51460 7 1 2 51453 51459
0 51461 7 1 2 51451 51460
0 51462 5 1 1 51461
0 51463 7 1 2 84788 94133
0 51464 7 1 2 51462 51463
0 51465 5 1 1 51464
0 51466 7 1 2 51445 51465
0 51467 5 1 1 51466
0 51468 7 1 2 61991 51467
0 51469 5 1 1 51468
0 51470 7 1 2 80547 91119
0 51471 5 2 1 51470
0 51472 7 1 2 84316 91772
0 51473 7 1 2 90603 51472
0 51474 5 1 1 51473
0 51475 7 1 2 95678 51474
0 51476 5 1 1 51475
0 51477 7 1 2 76230 51476
0 51478 5 1 1 51477
0 51479 7 2 2 74301 89298
0 51480 7 1 2 84400 95680
0 51481 5 1 1 51480
0 51482 7 1 2 51478 51481
0 51483 5 1 1 51482
0 51484 7 1 2 63552 51483
0 51485 5 1 1 51484
0 51486 7 1 2 74921 94636
0 51487 5 3 1 51486
0 51488 7 1 2 73393 94637
0 51489 5 1 1 51488
0 51490 7 1 2 84214 90396
0 51491 7 1 2 51489 51490
0 51492 7 1 2 95682 51491
0 51493 5 2 1 51492
0 51494 7 1 2 51485 95685
0 51495 5 1 1 51494
0 51496 7 1 2 78418 51495
0 51497 5 1 1 51496
0 51498 7 1 2 87692 89818
0 51499 5 1 1 51498
0 51500 7 1 2 76891 51499
0 51501 5 1 1 51500
0 51502 7 1 2 75559 51501
0 51503 5 1 1 51502
0 51504 7 1 2 80844 85956
0 51505 5 1 1 51504
0 51506 7 1 2 75560 93451
0 51507 5 1 1 51506
0 51508 7 1 2 51505 51507
0 51509 5 1 1 51508
0 51510 7 1 2 61099 51509
0 51511 5 1 1 51510
0 51512 7 1 2 51503 51511
0 51513 5 1 1 51512
0 51514 7 1 2 64415 51513
0 51515 5 1 1 51514
0 51516 7 1 2 71699 80310
0 51517 5 1 1 51516
0 51518 7 1 2 80293 51517
0 51519 5 1 1 51518
0 51520 7 1 2 89412 51519
0 51521 5 1 1 51520
0 51522 7 1 2 51515 51521
0 51523 5 1 1 51522
0 51524 7 1 2 61471 51523
0 51525 5 1 1 51524
0 51526 7 1 2 85641 91437
0 51527 5 1 1 51526
0 51528 7 1 2 51525 51527
0 51529 5 1 1 51528
0 51530 7 1 2 91811 51529
0 51531 5 1 1 51530
0 51532 7 1 2 51497 51531
0 51533 7 1 2 51469 51532
0 51534 5 1 1 51533
0 51535 7 1 2 64750 51534
0 51536 5 1 1 51535
0 51537 7 1 2 50921 51536
0 51538 5 1 1 51537
0 51539 7 1 2 66727 51538
0 51540 5 1 1 51539
0 51541 7 2 2 61736 73806
0 51542 7 1 2 69013 95687
0 51543 5 1 1 51542
0 51544 7 1 2 64109 87095
0 51545 5 1 1 51544
0 51546 7 2 2 84687 51545
0 51547 5 1 1 95689
0 51548 7 1 2 51543 51547
0 51549 5 2 1 51548
0 51550 7 1 2 57803 95691
0 51551 5 1 1 51550
0 51552 7 1 2 67602 95688
0 51553 5 1 1 51552
0 51554 7 2 2 67390 84688
0 51555 5 3 1 95693
0 51556 7 1 2 51553 95695
0 51557 5 1 1 51556
0 51558 7 1 2 71754 51557
0 51559 5 1 1 51558
0 51560 7 1 2 67391 94931
0 51561 5 2 1 51560
0 51562 7 1 2 51559 95698
0 51563 7 1 2 51551 51562
0 51564 5 1 1 51563
0 51565 7 1 2 59941 51564
0 51566 5 2 1 51565
0 51567 7 1 2 82635 78375
0 51568 7 1 2 94347 51567
0 51569 5 1 1 51568
0 51570 7 1 2 95700 51569
0 51571 5 1 1 51570
0 51572 7 1 2 59686 51571
0 51573 5 1 1 51572
0 51574 7 1 2 76596 94837
0 51575 7 1 2 95660 51574
0 51576 5 2 1 51575
0 51577 7 1 2 51573 95702
0 51578 5 1 1 51577
0 51579 7 1 2 58359 51578
0 51580 5 1 1 51579
0 51581 7 2 2 69825 84689
0 51582 5 1 1 95704
0 51583 7 1 2 59942 95705
0 51584 7 1 2 85932 51583
0 51585 5 2 1 51584
0 51586 7 1 2 51580 95706
0 51587 5 1 1 51586
0 51588 7 1 2 71920 51587
0 51589 5 1 1 51588
0 51590 7 1 2 70794 82586
0 51591 7 2 2 74158 51590
0 51592 5 2 1 95708
0 51593 7 1 2 76091 87581
0 51594 5 1 1 51593
0 51595 7 1 2 73505 51594
0 51596 5 1 1 51595
0 51597 7 2 2 66380 51596
0 51598 7 1 2 57521 95712
0 51599 5 1 1 51598
0 51600 7 1 2 95710 51599
0 51601 5 1 1 51600
0 51602 7 1 2 58082 51601
0 51603 5 1 1 51602
0 51604 7 1 2 59943 72250
0 51605 7 1 2 94932 51604
0 51606 5 2 1 51605
0 51607 7 1 2 51603 95714
0 51608 5 1 1 51607
0 51609 7 1 2 71227 51608
0 51610 5 1 1 51609
0 51611 7 1 2 71547 80401
0 51612 7 2 2 82427 51611
0 51613 7 2 2 68052 73857
0 51614 7 1 2 95716 95718
0 51615 5 2 1 51614
0 51616 7 1 2 51610 95720
0 51617 5 1 1 51616
0 51618 7 1 2 78328 51617
0 51619 5 1 1 51618
0 51620 7 1 2 57522 95709
0 51621 5 2 1 51620
0 51622 7 1 2 57804 95713
0 51623 5 1 1 51622
0 51624 7 1 2 95722 51623
0 51625 5 1 1 51624
0 51626 7 1 2 58083 51625
0 51627 5 1 1 51626
0 51628 7 1 2 75918 91966
0 51629 5 2 1 51628
0 51630 7 1 2 51627 95724
0 51631 5 1 1 51630
0 51632 7 1 2 71228 51631
0 51633 5 1 1 51632
0 51634 7 1 2 82445 95717
0 51635 5 2 1 51634
0 51636 7 1 2 51633 95726
0 51637 5 1 1 51636
0 51638 7 1 2 71755 51637
0 51639 5 1 1 51638
0 51640 7 1 2 51619 51639
0 51641 7 1 2 51589 51640
0 51642 5 1 1 51641
0 51643 7 1 2 58806 51642
0 51644 5 1 1 51643
0 51645 7 1 2 78376 79401
0 51646 7 1 2 94348 51645
0 51647 5 1 1 51646
0 51648 7 1 2 95701 51647
0 51649 5 1 1 51648
0 51650 7 1 2 59687 51649
0 51651 5 1 1 51650
0 51652 7 1 2 95703 51651
0 51653 5 1 1 51652
0 51654 7 1 2 58360 51653
0 51655 5 1 1 51654
0 51656 7 1 2 95707 51655
0 51657 5 1 1 51656
0 51658 7 1 2 71921 51657
0 51659 5 1 1 51658
0 51660 7 1 2 76092 73519
0 51661 5 1 1 51660
0 51662 7 1 2 73506 51661
0 51663 5 1 1 51662
0 51664 7 2 2 66381 51663
0 51665 7 1 2 57523 95728
0 51666 5 1 1 51665
0 51667 7 1 2 95711 51666
0 51668 5 1 1 51667
0 51669 7 1 2 58084 51668
0 51670 5 1 1 51669
0 51671 7 1 2 95715 51670
0 51672 5 1 1 51671
0 51673 7 1 2 71229 51672
0 51674 5 1 1 51673
0 51675 7 1 2 95721 51674
0 51676 5 1 1 51675
0 51677 7 1 2 78329 51676
0 51678 5 1 1 51677
0 51679 7 1 2 57805 95729
0 51680 5 1 1 51679
0 51681 7 1 2 95723 51680
0 51682 5 1 1 51681
0 51683 7 1 2 58085 51682
0 51684 5 1 1 51683
0 51685 7 1 2 95725 51684
0 51686 5 1 1 51685
0 51687 7 1 2 71230 51686
0 51688 5 1 1 51687
0 51689 7 1 2 95727 51688
0 51690 5 1 1 51689
0 51691 7 1 2 71756 51690
0 51692 5 1 1 51691
0 51693 7 1 2 51678 51692
0 51694 7 1 2 51659 51693
0 51695 5 1 1 51694
0 51696 7 1 2 60065 51695
0 51697 5 1 1 51696
0 51698 7 1 2 51644 51697
0 51699 5 1 1 51698
0 51700 7 1 2 65733 51699
0 51701 5 1 1 51700
0 51702 7 1 2 67392 86172
0 51703 5 1 1 51702
0 51704 7 1 2 68053 94364
0 51705 5 1 1 51704
0 51706 7 1 2 65734 80329
0 51707 5 1 1 51706
0 51708 7 1 2 51705 51707
0 51709 7 1 2 51703 51708
0 51710 5 1 1 51709
0 51711 7 1 2 66803 84690
0 51712 7 1 2 83830 51711
0 51713 7 1 2 51710 51712
0 51714 5 1 1 51713
0 51715 7 1 2 51701 51714
0 51716 5 1 1 51715
0 51717 7 1 2 58675 51716
0 51718 5 1 1 51717
0 51719 7 3 2 71453 70227
0 51720 5 1 1 95730
0 51721 7 1 2 58086 51720
0 51722 5 1 1 51721
0 51723 7 1 2 90983 51722
0 51724 5 1 1 51723
0 51725 7 1 2 80918 51724
0 51726 5 1 1 51725
0 51727 7 1 2 83963 36955
0 51728 5 1 1 51727
0 51729 7 1 2 58361 51728
0 51730 5 1 1 51729
0 51731 7 3 2 36963 51730
0 51732 5 1 1 95733
0 51733 7 1 2 82931 90987
0 51734 5 1 1 51733
0 51735 7 2 2 58676 86448
0 51736 5 1 1 95736
0 51737 7 1 2 81297 51736
0 51738 5 1 1 51737
0 51739 7 1 2 51734 51738
0 51740 5 1 1 51739
0 51741 7 1 2 95734 51740
0 51742 7 1 2 51726 51741
0 51743 5 2 1 51742
0 51744 7 1 2 64639 95738
0 51745 5 1 1 51744
0 51746 7 1 2 84967 86019
0 51747 5 1 1 51746
0 51748 7 1 2 86298 88065
0 51749 5 1 1 51748
0 51750 7 1 2 51747 51749
0 51751 5 1 1 51750
0 51752 7 1 2 68272 78010
0 51753 7 1 2 76394 51752
0 51754 5 1 1 51753
0 51755 7 1 2 75040 51754
0 51756 7 1 2 51751 51755
0 51757 5 1 1 51756
0 51758 7 1 2 59944 51757
0 51759 5 1 1 51758
0 51760 7 1 2 66382 51759
0 51761 7 1 2 51745 51760
0 51762 5 1 1 51761
0 51763 7 1 2 84908 85218
0 51764 5 1 1 51763
0 51765 7 1 2 82239 51764
0 51766 5 1 1 51765
0 51767 7 1 2 95735 51766
0 51768 5 1 1 51767
0 51769 7 1 2 75598 51768
0 51770 5 1 1 51769
0 51771 7 1 2 70177 80985
0 51772 7 1 2 88027 51771
0 51773 5 1 1 51772
0 51774 7 1 2 80783 51773
0 51775 5 1 1 51774
0 51776 7 1 2 73183 26031
0 51777 5 1 1 51776
0 51778 7 1 2 70228 88031
0 51779 7 1 2 51777 51778
0 51780 5 1 1 51779
0 51781 7 1 2 51775 51780
0 51782 5 1 1 51781
0 51783 7 1 2 13276 51782
0 51784 5 1 1 51783
0 51785 7 1 2 71922 51784
0 51786 5 1 1 51785
0 51787 7 1 2 84912 80986
0 51788 7 1 2 82240 51787
0 51789 5 1 1 51788
0 51790 7 1 2 59945 95737
0 51791 5 1 1 51790
0 51792 7 1 2 61737 51791
0 51793 7 1 2 51789 51792
0 51794 7 1 2 51786 51793
0 51795 7 1 2 51770 51794
0 51796 5 1 1 51795
0 51797 7 1 2 66083 51796
0 51798 7 1 2 51762 51797
0 51799 5 1 1 51798
0 51800 7 1 2 80185 92666
0 51801 5 2 1 51800
0 51802 7 1 2 75561 95740
0 51803 5 1 1 51802
0 51804 7 1 2 84691 51803
0 51805 5 1 1 51804
0 51806 7 1 2 76710 93210
0 51807 5 1 1 51806
0 51808 7 1 2 91787 93267
0 51809 7 1 2 51807 51808
0 51810 5 1 1 51809
0 51811 7 1 2 51805 51810
0 51812 5 1 1 51811
0 51813 7 1 2 71548 51812
0 51814 5 1 1 51813
0 51815 7 4 2 67393 76371
0 51816 5 1 1 95742
0 51817 7 1 2 78616 75254
0 51818 5 1 1 51817
0 51819 7 1 2 68176 42125
0 51820 7 1 2 51818 51819
0 51821 5 1 1 51820
0 51822 7 2 2 84554 51821
0 51823 5 1 1 95746
0 51824 7 1 2 51816 51823
0 51825 5 1 1 51824
0 51826 7 1 2 61738 85222
0 51827 7 1 2 51825 51826
0 51828 5 1 1 51827
0 51829 7 1 2 51814 51828
0 51830 5 1 1 51829
0 51831 7 1 2 68415 51830
0 51832 5 1 1 51831
0 51833 7 1 2 73942 81964
0 51834 5 1 1 51833
0 51835 7 1 2 83964 51834
0 51836 5 1 1 51835
0 51837 7 1 2 85223 51836
0 51838 5 1 1 51837
0 51839 7 1 2 93310 51838
0 51840 5 1 1 51839
0 51841 7 1 2 61739 51840
0 51842 5 1 1 51841
0 51843 7 1 2 69469 82397
0 51844 5 1 1 51843
0 51845 7 1 2 75255 84069
0 51846 5 1 1 51845
0 51847 7 1 2 51844 51846
0 51848 5 1 1 51847
0 51849 7 1 2 67697 51848
0 51850 5 1 1 51849
0 51851 7 1 2 71549 84692
0 51852 5 2 1 51851
0 51853 7 1 2 51850 95748
0 51854 5 1 1 51853
0 51855 7 1 2 75599 51854
0 51856 5 1 1 51855
0 51857 7 1 2 71550 89390
0 51858 5 1 1 51857
0 51859 7 2 2 80987 84693
0 51860 7 1 2 85900 95750
0 51861 5 1 1 51860
0 51862 7 1 2 81965 89391
0 51863 5 1 1 51862
0 51864 7 1 2 51861 51863
0 51865 5 1 1 51864
0 51866 7 1 2 67698 51865
0 51867 5 1 1 51866
0 51868 7 1 2 51858 51867
0 51869 7 1 2 51856 51868
0 51870 5 1 1 51869
0 51871 7 1 2 78617 51870
0 51872 5 1 1 51871
0 51873 7 1 2 51842 51872
0 51874 7 1 2 51832 51873
0 51875 7 1 2 84706 19422
0 51876 5 1 1 51875
0 51877 7 1 2 75600 51876
0 51878 5 1 1 51877
0 51879 7 1 2 89546 94084
0 51880 5 1 1 51879
0 51881 7 1 2 89365 51880
0 51882 7 1 2 51878 51881
0 51883 5 1 1 51882
0 51884 7 1 2 68811 51883
0 51885 5 1 1 51884
0 51886 7 1 2 70355 83350
0 51887 5 2 1 51886
0 51888 7 1 2 75562 95752
0 51889 5 1 1 51888
0 51890 7 1 2 65341 95445
0 51891 7 1 2 51889 51890
0 51892 5 1 1 51891
0 51893 7 1 2 76711 95753
0 51894 5 1 1 51893
0 51895 7 1 2 78654 91788
0 51896 7 1 2 51894 51895
0 51897 5 1 1 51896
0 51898 7 1 2 51892 51897
0 51899 7 1 2 51885 51898
0 51900 5 1 1 51899
0 51901 7 1 2 71551 51900
0 51902 5 1 1 51901
0 51903 7 1 2 78768 94621
0 51904 5 1 1 51903
0 51905 7 1 2 73924 51904
0 51906 5 1 1 51905
0 51907 7 1 2 57524 95743
0 51908 5 1 1 51907
0 51909 7 1 2 51906 51908
0 51910 5 1 1 51909
0 51911 7 1 2 68416 51910
0 51912 5 1 1 51911
0 51913 7 1 2 70007 94137
0 51914 5 1 1 51913
0 51915 7 1 2 67897 91153
0 51916 5 1 1 51915
0 51917 7 1 2 59688 80772
0 51918 5 1 1 51917
0 51919 7 2 2 73925 76515
0 51920 5 1 1 95754
0 51921 7 1 2 80714 95755
0 51922 5 1 1 51921
0 51923 7 1 2 51918 51922
0 51924 7 1 2 51916 51923
0 51925 7 1 2 51914 51924
0 51926 7 1 2 51912 51925
0 51927 5 1 1 51926
0 51928 7 1 2 95751 51927
0 51929 5 1 1 51928
0 51930 7 1 2 51902 51929
0 51931 7 1 2 51874 51930
0 51932 7 1 2 51799 51931
0 51933 5 1 1 51932
0 51934 7 1 2 66872 51933
0 51935 5 1 1 51934
0 51936 7 1 2 51718 51935
0 51937 5 1 1 51936
0 51938 7 1 2 67489 51937
0 51939 5 1 1 51938
0 51940 7 1 2 68534 86254
0 51941 5 1 1 51940
0 51942 7 1 2 7096 51941
0 51943 5 1 1 51942
0 51944 7 1 2 77276 51943
0 51945 5 1 1 51944
0 51946 7 1 2 61100 72555
0 51947 5 1 1 51946
0 51948 7 1 2 58362 51947
0 51949 5 1 1 51948
0 51950 7 1 2 75666 51949
0 51951 5 1 1 51950
0 51952 7 1 2 51945 51951
0 51953 5 1 1 51952
0 51954 7 1 2 86605 51953
0 51955 5 1 1 51954
0 51956 7 1 2 61472 81813
0 51957 5 1 1 51956
0 51958 7 1 2 86127 74302
0 51959 7 1 2 81758 51958
0 51960 5 1 1 51959
0 51961 7 1 2 9230 51960
0 51962 5 1 1 51961
0 51963 7 1 2 63110 51962
0 51964 5 1 1 51963
0 51965 7 1 2 51957 51964
0 51966 5 1 1 51965
0 51967 7 1 2 87271 51966
0 51968 5 1 1 51967
0 51969 7 1 2 83855 82623
0 51970 7 1 2 92150 51969
0 51971 5 1 1 51970
0 51972 7 1 2 51968 51971
0 51973 5 1 1 51972
0 51974 7 1 2 68535 51973
0 51975 5 1 1 51974
0 51976 7 1 2 66084 80002
0 51977 5 1 1 51976
0 51978 7 1 2 75667 51977
0 51979 5 1 1 51978
0 51980 7 1 2 66795 93968
0 51981 5 1 1 51980
0 51982 7 1 2 51979 51981
0 51983 5 1 1 51982
0 51984 7 1 2 60678 51983
0 51985 5 1 1 51984
0 51986 7 1 2 87880 77277
0 51987 5 1 1 51986
0 51988 7 1 2 51985 51987
0 51989 5 1 1 51988
0 51990 7 1 2 87272 51989
0 51991 5 1 1 51990
0 51992 7 1 2 51975 51991
0 51993 5 1 1 51992
0 51994 7 1 2 68273 51993
0 51995 5 1 1 51994
0 51996 7 1 2 51955 51995
0 51997 5 1 1 51996
0 51998 7 1 2 64416 51997
0 51999 5 1 1 51998
0 52000 7 1 2 74998 75769
0 52001 5 1 1 52000
0 52002 7 1 2 81824 52001
0 52003 5 1 1 52002
0 52004 7 1 2 87273 52003
0 52005 5 1 1 52004
0 52006 7 1 2 82664 74910
0 52007 7 1 2 92571 52006
0 52008 5 1 1 52007
0 52009 7 1 2 52005 52008
0 52010 5 1 1 52009
0 52011 7 1 2 68274 52010
0 52012 5 1 1 52011
0 52013 7 1 2 68536 91759
0 52014 7 1 2 95221 52013
0 52015 5 1 1 52014
0 52016 7 1 2 52012 52015
0 52017 5 1 1 52016
0 52018 7 1 2 75470 52017
0 52019 5 1 1 52018
0 52020 7 1 2 51999 52019
0 52021 5 1 1 52020
0 52022 7 1 2 63413 52021
0 52023 5 1 1 52022
0 52024 7 2 2 68275 87705
0 52025 7 1 2 61101 95756
0 52026 5 1 1 52025
0 52027 7 1 2 87701 52026
0 52028 5 1 1 52027
0 52029 7 1 2 63111 52028
0 52030 5 1 1 52029
0 52031 7 2 2 72878 87794
0 52032 5 1 1 95758
0 52033 7 1 2 52030 52032
0 52034 5 2 1 52033
0 52035 7 4 2 82109 86677
0 52036 5 1 1 95762
0 52037 7 2 2 83668 95763
0 52038 7 1 2 95760 95766
0 52039 5 1 1 52038
0 52040 7 1 2 84197 90820
0 52041 5 1 1 52040
0 52042 7 1 2 58807 85810
0 52043 5 1 1 52042
0 52044 7 1 2 52041 52043
0 52045 5 1 1 52044
0 52046 7 1 2 63112 52045
0 52047 5 1 1 52046
0 52048 7 1 2 58808 87698
0 52049 5 1 1 52048
0 52050 7 1 2 52047 52049
0 52051 5 1 1 52050
0 52052 7 1 2 68276 93975
0 52053 7 1 2 52051 52052
0 52054 5 1 1 52053
0 52055 7 2 2 82690 87138
0 52056 7 1 2 77999 90322
0 52057 7 1 2 95768 52056
0 52058 5 1 1 52057
0 52059 7 2 2 74668 82428
0 52060 7 1 2 87582 95770
0 52061 7 1 2 93196 52060
0 52062 5 1 1 52061
0 52063 7 1 2 52058 52062
0 52064 7 1 2 52054 52063
0 52065 5 1 1 52064
0 52066 7 1 2 61992 52065
0 52067 5 1 1 52066
0 52068 7 1 2 52039 52067
0 52069 5 1 1 52068
0 52070 7 1 2 68886 52069
0 52071 5 1 1 52070
0 52072 7 2 2 58363 90562
0 52073 5 1 1 95772
0 52074 7 1 2 59689 52073
0 52075 5 1 1 52074
0 52076 7 1 2 78147 87746
0 52077 7 1 2 80375 52076
0 52078 5 1 1 52077
0 52079 7 1 2 52075 52078
0 52080 5 2 1 52079
0 52081 7 1 2 87688 91120
0 52082 7 1 2 95774 52081
0 52083 5 1 1 52082
0 52084 7 1 2 52071 52083
0 52085 7 1 2 52023 52084
0 52086 5 1 1 52085
0 52087 7 1 2 66728 52086
0 52088 5 1 1 52087
0 52089 7 1 2 65735 84959
0 52090 5 1 1 52089
0 52091 7 2 2 82436 92573
0 52092 7 1 2 78011 95776
0 52093 7 1 2 52090 52092
0 52094 5 1 1 52093
0 52095 7 1 2 68887 82437
0 52096 7 1 2 93860 93988
0 52097 7 1 2 52095 52096
0 52098 5 1 1 52097
0 52099 7 1 2 52094 52098
0 52100 7 1 2 52088 52099
0 52101 5 1 1 52100
0 52102 7 1 2 68177 52101
0 52103 5 1 1 52102
0 52104 7 1 2 67394 95773
0 52105 5 1 1 52104
0 52106 7 1 2 91670 52105
0 52107 5 1 1 52106
0 52108 7 1 2 85990 87800
0 52109 5 1 1 52108
0 52110 7 1 2 67226 85887
0 52111 7 1 2 52109 52110
0 52112 5 2 1 52111
0 52113 7 1 2 52107 95778
0 52114 5 1 1 52113
0 52115 7 1 2 95630 52114
0 52116 5 1 1 52115
0 52117 7 1 2 78012 78148
0 52118 7 1 2 91975 94971
0 52119 7 1 2 52117 52118
0 52120 5 1 1 52119
0 52121 7 1 2 52116 52120
0 52122 5 1 1 52121
0 52123 7 1 2 58809 52122
0 52124 5 1 1 52123
0 52125 7 2 2 62530 69927
0 52126 7 2 2 87760 95780
0 52127 7 1 2 89618 90097
0 52128 7 1 2 95782 52127
0 52129 5 1 1 52128
0 52130 7 1 2 52124 52129
0 52131 5 1 1 52130
0 52132 7 1 2 60066 52131
0 52133 5 1 1 52132
0 52134 7 1 2 61473 93397
0 52135 5 1 1 52134
0 52136 7 1 2 80294 52135
0 52137 5 1 1 52136
0 52138 7 1 2 63553 82110
0 52139 7 1 2 94880 52138
0 52140 7 1 2 80839 52139
0 52141 7 1 2 52137 52140
0 52142 5 1 1 52141
0 52143 7 1 2 52133 52142
0 52144 5 1 1 52143
0 52145 7 1 2 62274 52144
0 52146 5 1 1 52145
0 52147 7 2 2 84789 91660
0 52148 7 1 2 89481 95784
0 52149 5 1 1 52148
0 52150 7 1 2 87176 73368
0 52151 5 1 1 52150
0 52152 7 1 2 73683 79043
0 52153 5 1 1 52152
0 52154 7 1 2 52151 52153
0 52155 5 1 1 52154
0 52156 7 1 2 80944 82665
0 52157 7 1 2 52155 52156
0 52158 5 1 1 52157
0 52159 7 1 2 52149 52158
0 52160 5 1 1 52159
0 52161 7 1 2 61102 52160
0 52162 5 1 1 52161
0 52163 7 1 2 83002 91121
0 52164 7 1 2 95181 52163
0 52165 5 1 1 52164
0 52166 7 1 2 52162 52165
0 52167 5 1 1 52166
0 52168 7 1 2 66729 52167
0 52169 5 1 1 52168
0 52170 7 1 2 52146 52169
0 52171 5 1 1 52170
0 52172 7 1 2 69071 52171
0 52173 5 1 1 52172
0 52174 7 1 2 67970 81898
0 52175 7 1 2 82429 92567
0 52176 7 1 2 52174 52175
0 52177 5 1 1 52176
0 52178 7 1 2 73554 90212
0 52179 7 1 2 90402 52178
0 52180 5 1 1 52179
0 52181 7 1 2 52177 52180
0 52182 5 1 1 52181
0 52183 7 1 2 65099 52182
0 52184 5 1 1 52183
0 52185 7 1 2 69072 93836
0 52186 5 1 1 52185
0 52187 7 1 2 95194 52186
0 52188 5 1 1 52187
0 52189 7 1 2 58810 82438
0 52190 7 1 2 52188 52189
0 52191 5 1 1 52190
0 52192 7 1 2 52184 52191
0 52193 5 1 1 52192
0 52194 7 1 2 66085 52193
0 52195 5 1 1 52194
0 52196 7 2 2 64417 81079
0 52197 7 1 2 92807 95786
0 52198 5 1 1 52197
0 52199 7 2 2 87917 94192
0 52200 5 1 1 95788
0 52201 7 1 2 62806 94144
0 52202 7 1 2 95789 52201
0 52203 5 1 1 52202
0 52204 7 1 2 52198 52203
0 52205 5 1 1 52204
0 52206 7 1 2 63414 52205
0 52207 5 1 1 52206
0 52208 7 1 2 80443 79147
0 52209 7 1 2 79176 52208
0 52210 5 1 1 52209
0 52211 7 1 2 52207 52210
0 52212 5 1 1 52211
0 52213 7 1 2 69073 52212
0 52214 5 1 1 52213
0 52215 7 3 2 63415 92568
0 52216 7 1 2 70376 73369
0 52217 7 1 2 95790 52216
0 52218 5 1 1 52217
0 52219 7 1 2 52214 52218
0 52220 5 1 1 52219
0 52221 7 1 2 61740 52220
0 52222 5 1 1 52221
0 52223 7 1 2 80871 84267
0 52224 7 1 2 87211 91362
0 52225 7 1 2 52223 52224
0 52226 5 1 1 52225
0 52227 7 1 2 52222 52226
0 52228 5 1 1 52227
0 52229 7 1 2 92737 52228
0 52230 5 1 1 52229
0 52231 7 1 2 52195 52230
0 52232 5 1 1 52231
0 52233 7 1 2 60067 52232
0 52234 5 1 1 52233
0 52235 7 1 2 78256 6013
0 52236 5 1 1 52235
0 52237 7 1 2 93141 52236
0 52238 5 1 1 52237
0 52239 7 1 2 69443 95731
0 52240 5 1 1 52239
0 52241 7 1 2 52238 52240
0 52242 5 1 1 52241
0 52243 7 2 2 66642 92272
0 52244 7 1 2 52242 95793
0 52245 5 1 1 52244
0 52246 7 1 2 59690 76395
0 52247 5 1 1 52246
0 52248 7 1 2 65342 75025
0 52249 5 1 1 52248
0 52250 7 1 2 52247 52249
0 52251 5 1 1 52250
0 52252 7 1 2 84580 82430
0 52253 7 1 2 52251 52252
0 52254 5 1 1 52253
0 52255 7 1 2 52245 52254
0 52256 5 1 1 52255
0 52257 7 1 2 62807 52256
0 52258 5 1 1 52257
0 52259 7 1 2 59691 79341
0 52260 7 2 2 92151 52259
0 52261 5 1 1 95795
0 52262 7 1 2 71454 80076
0 52263 7 1 2 95794 52262
0 52264 5 1 1 52263
0 52265 7 2 2 63787 73845
0 52266 7 1 2 86128 82666
0 52267 7 1 2 95797 52266
0 52268 5 1 1 52267
0 52269 7 1 2 52264 52268
0 52270 5 1 1 52269
0 52271 7 1 2 60679 52270
0 52272 5 1 1 52271
0 52273 7 1 2 52261 52272
0 52274 5 1 1 52273
0 52275 7 1 2 64110 52274
0 52276 5 1 1 52275
0 52277 7 1 2 78393 90638
0 52278 7 1 2 89213 52277
0 52279 5 1 1 52278
0 52280 7 1 2 95679 52279
0 52281 5 1 1 52280
0 52282 7 1 2 71335 52281
0 52283 5 1 1 52282
0 52284 7 1 2 76383 95796
0 52285 5 1 1 52284
0 52286 7 3 2 60680 82111
0 52287 7 1 2 80683 95799
0 52288 5 1 1 52287
0 52289 7 1 2 92022 94442
0 52290 5 1 1 52289
0 52291 7 1 2 52288 52290
0 52292 5 1 1 52291
0 52293 7 1 2 61474 52292
0 52294 5 1 1 52293
0 52295 7 1 2 52285 52294
0 52296 7 1 2 52283 52295
0 52297 7 1 2 52276 52296
0 52298 7 1 2 52258 52297
0 52299 5 1 1 52298
0 52300 7 1 2 63554 52299
0 52301 5 1 1 52300
0 52302 7 1 2 95686 52301
0 52303 5 1 1 52302
0 52304 7 1 2 94881 52303
0 52305 5 1 1 52304
0 52306 7 1 2 52234 52305
0 52307 5 1 1 52306
0 52308 7 1 2 62275 52307
0 52309 5 1 1 52308
0 52310 7 1 2 64418 81278
0 52311 5 1 1 52310
0 52312 7 1 2 69444 91591
0 52313 5 1 1 52312
0 52314 7 1 2 52311 52313
0 52315 5 1 1 52314
0 52316 7 1 2 61475 52315
0 52317 5 1 1 52316
0 52318 7 1 2 81014 94093
0 52319 5 1 1 52318
0 52320 7 2 2 71336 70229
0 52321 5 2 1 95802
0 52322 7 1 2 78056 95803
0 52323 7 1 2 91443 52322
0 52324 5 1 1 52323
0 52325 7 1 2 52319 52324
0 52326 7 1 2 52317 52325
0 52327 5 1 1 52326
0 52328 7 1 2 95767 52327
0 52329 5 1 1 52328
0 52330 7 3 2 80301 89199
0 52331 5 1 1 95806
0 52332 7 1 2 70230 90323
0 52333 5 1 1 52332
0 52334 7 1 2 22651 52200
0 52335 5 1 1 52334
0 52336 7 1 2 76712 76384
0 52337 7 1 2 52335 52336
0 52338 5 1 1 52337
0 52339 7 1 2 52333 52338
0 52340 5 1 1 52339
0 52341 7 1 2 62808 52340
0 52342 5 1 1 52341
0 52343 7 1 2 76260 92813
0 52344 5 1 1 52343
0 52345 7 1 2 90324 52344
0 52346 5 1 1 52345
0 52347 7 1 2 52342 52346
0 52348 5 1 1 52347
0 52349 7 1 2 64419 52348
0 52350 5 1 1 52349
0 52351 7 1 2 52331 52350
0 52352 5 1 1 52351
0 52353 7 1 2 87555 52352
0 52354 5 1 1 52353
0 52355 7 1 2 79031 73749
0 52356 5 1 1 52355
0 52357 7 1 2 80872 82809
0 52358 5 1 1 52357
0 52359 7 1 2 52356 52358
0 52360 5 1 1 52359
0 52361 7 2 2 64751 95054
0 52362 7 1 2 52360 95809
0 52363 5 1 1 52362
0 52364 7 1 2 61476 52363
0 52365 7 1 2 52354 52364
0 52366 5 1 1 52365
0 52367 7 1 2 74470 95771
0 52368 5 1 1 52367
0 52369 7 1 2 79843 82368
0 52370 7 1 2 90236 52369
0 52371 7 1 2 80840 52370
0 52372 5 1 1 52371
0 52373 7 1 2 52368 52372
0 52374 5 1 1 52373
0 52375 7 1 2 62809 52374
0 52376 5 1 1 52375
0 52377 7 1 2 77350 81408
0 52378 7 1 2 92441 52377
0 52379 5 1 1 52378
0 52380 7 1 2 52376 52379
0 52381 5 1 1 52380
0 52382 7 1 2 72406 52381
0 52383 5 1 1 52382
0 52384 7 1 2 62810 92210
0 52385 5 1 1 52384
0 52386 7 1 2 86434 78455
0 52387 7 1 2 52385 52386
0 52388 5 1 1 52387
0 52389 7 1 2 74669 52388
0 52390 5 1 1 52389
0 52391 7 1 2 63555 85703
0 52392 5 1 1 52391
0 52393 7 1 2 67227 85078
0 52394 5 1 1 52393
0 52395 7 1 2 52392 52394
0 52396 5 1 1 52395
0 52397 7 1 2 69074 72486
0 52398 7 1 2 52396 52397
0 52399 5 1 1 52398
0 52400 7 1 2 52390 52399
0 52401 5 1 1 52400
0 52402 7 1 2 95229 52401
0 52403 5 1 1 52402
0 52404 7 1 2 87556 88063
0 52405 7 1 2 95807 52404
0 52406 5 1 1 52405
0 52407 7 1 2 87771 92299
0 52408 7 1 2 90403 52407
0 52409 5 1 1 52408
0 52410 7 1 2 66086 52409
0 52411 7 1 2 52406 52410
0 52412 7 1 2 52403 52411
0 52413 7 1 2 52383 52412
0 52414 5 1 1 52413
0 52415 7 1 2 61993 52414
0 52416 7 1 2 52366 52415
0 52417 5 1 1 52416
0 52418 7 1 2 52329 52417
0 52419 5 1 1 52418
0 52420 7 1 2 66730 52419
0 52421 5 1 1 52420
0 52422 7 1 2 74551 37458
0 52423 5 2 1 52422
0 52424 7 1 2 80524 95777
0 52425 7 1 2 95811 52424
0 52426 5 1 1 52425
0 52427 7 1 2 52421 52426
0 52428 7 1 2 52309 52427
0 52429 5 1 1 52428
0 52430 7 1 2 67796 52429
0 52431 5 1 1 52430
0 52432 7 1 2 52173 52431
0 52433 7 1 2 52103 52432
0 52434 7 1 2 51939 52433
0 52435 7 1 2 51540 52434
0 52436 5 1 1 52435
0 52437 7 1 2 70543 52436
0 52438 5 1 1 52437
0 52439 7 2 2 66873 81421
0 52440 5 1 1 95813
0 52441 7 1 2 79444 4803
0 52442 5 1 1 52441
0 52443 7 1 2 84433 81547
0 52444 7 1 2 52442 52443
0 52445 5 1 1 52444
0 52446 7 1 2 52440 52445
0 52447 5 1 1 52446
0 52448 7 1 2 57525 52447
0 52449 5 1 1 52448
0 52450 7 1 2 87566 39803
0 52451 5 1 1 52450
0 52452 7 1 2 59035 52451
0 52453 5 1 1 52452
0 52454 7 1 2 47306 52453
0 52455 5 1 1 52454
0 52456 7 1 2 74753 52455
0 52457 5 1 1 52456
0 52458 7 1 2 52449 52457
0 52459 5 1 1 52458
0 52460 7 1 2 58364 52459
0 52461 5 1 1 52460
0 52462 7 1 2 76516 72917
0 52463 7 1 2 95814 52462
0 52464 5 1 1 52463
0 52465 7 1 2 52461 52464
0 52466 5 1 1 52465
0 52467 7 1 2 73408 52466
0 52468 5 1 1 52467
0 52469 7 2 2 61741 86268
0 52470 7 1 2 73943 75177
0 52471 5 1 1 52470
0 52472 7 1 2 81080 52471
0 52473 5 1 1 52472
0 52474 7 1 2 95815 52473
0 52475 5 1 1 52474
0 52476 7 3 2 87373 93143
0 52477 5 1 1 95817
0 52478 7 2 2 84707 52477
0 52479 5 3 1 95820
0 52480 7 1 2 67228 75196
0 52481 5 1 1 52480
0 52482 7 1 2 95822 52481
0 52483 5 1 1 52482
0 52484 7 1 2 52475 52483
0 52485 5 1 1 52484
0 52486 7 1 2 60068 52485
0 52487 5 1 1 52486
0 52488 7 1 2 83645 95524
0 52489 5 1 1 52488
0 52490 7 1 2 85865 93122
0 52491 5 1 1 52490
0 52492 7 1 2 87143 52491
0 52493 5 1 1 52492
0 52494 7 1 2 95132 52493
0 52495 5 1 1 52494
0 52496 7 1 2 61477 72943
0 52497 5 1 1 52496
0 52498 7 1 2 58365 52497
0 52499 5 1 1 52498
0 52500 7 1 2 1233 52499
0 52501 5 1 1 52500
0 52502 7 1 2 95285 52501
0 52503 5 1 1 52502
0 52504 7 1 2 52495 52503
0 52505 5 1 1 52504
0 52506 7 1 2 65343 52505
0 52507 5 1 1 52506
0 52508 7 1 2 52489 52507
0 52509 7 1 2 52487 52508
0 52510 5 1 1 52509
0 52511 7 1 2 58811 52510
0 52512 5 1 1 52511
0 52513 7 1 2 52468 52512
0 52514 5 1 1 52513
0 52515 7 1 2 67699 52514
0 52516 5 1 1 52515
0 52517 7 1 2 72359 94383
0 52518 5 1 1 52517
0 52519 7 1 2 57526 93699
0 52520 5 1 1 52519
0 52521 7 1 2 80576 52520
0 52522 5 1 1 52521
0 52523 7 1 2 86269 52522
0 52524 5 1 1 52523
0 52525 7 1 2 52518 52524
0 52526 5 1 1 52525
0 52527 7 1 2 87557 52526
0 52528 5 1 1 52527
0 52529 7 1 2 83646 87583
0 52530 5 1 1 52529
0 52531 7 1 2 87144 52530
0 52532 5 1 1 52531
0 52533 7 3 2 66383 52532
0 52534 7 1 2 69470 95825
0 52535 5 1 1 52534
0 52536 7 1 2 52528 52535
0 52537 5 1 1 52536
0 52538 7 1 2 65736 52537
0 52539 5 1 1 52538
0 52540 7 1 2 94379 95037
0 52541 5 2 1 52540
0 52542 7 2 2 87558 95828
0 52543 5 1 1 95830
0 52544 7 1 2 57527 95826
0 52545 5 1 1 52544
0 52546 7 1 2 52543 52545
0 52547 5 1 1 52546
0 52548 7 1 2 65737 52547
0 52549 5 1 1 52548
0 52550 7 1 2 82779 95823
0 52551 5 1 1 52550
0 52552 7 1 2 52549 52551
0 52553 5 1 1 52552
0 52554 7 1 2 71757 52553
0 52555 5 1 1 52554
0 52556 7 1 2 52539 52555
0 52557 5 1 1 52556
0 52558 7 1 2 57806 52557
0 52559 5 1 1 52558
0 52560 7 1 2 69974 75206
0 52561 7 1 2 95816 52560
0 52562 5 1 1 52561
0 52563 7 1 2 48602 52562
0 52564 5 1 1 52563
0 52565 7 1 2 59175 52564
0 52566 5 1 1 52565
0 52567 7 1 2 69471 75256
0 52568 5 1 1 52567
0 52569 7 2 2 76358 52568
0 52570 5 1 1 95832
0 52571 7 1 2 84694 52570
0 52572 5 1 1 52571
0 52573 7 1 2 52566 52572
0 52574 5 1 1 52573
0 52575 7 1 2 58087 52574
0 52576 5 1 1 52575
0 52577 7 1 2 88890 95833
0 52578 5 1 1 52577
0 52579 7 1 2 59386 52578
0 52580 5 1 1 52579
0 52581 7 1 2 71455 52580
0 52582 5 1 1 52581
0 52583 7 1 2 84695 52582
0 52584 5 1 1 52583
0 52585 7 1 2 2908 95824
0 52586 5 1 1 52585
0 52587 7 1 2 76305 84304
0 52588 7 1 2 95829 52587
0 52589 5 1 1 52588
0 52590 7 1 2 52586 52589
0 52591 5 1 1 52590
0 52592 7 1 2 57807 52591
0 52593 5 1 1 52592
0 52594 7 1 2 79618 86270
0 52595 5 1 1 52594
0 52596 7 1 2 61742 94380
0 52597 7 1 2 52595 52596
0 52598 5 1 1 52597
0 52599 7 1 2 80330 15901
0 52600 7 1 2 52598 52599
0 52601 5 1 1 52600
0 52602 7 1 2 79619 94384
0 52603 5 1 1 52602
0 52604 7 1 2 90017 52603
0 52605 5 1 1 52604
0 52606 7 1 2 61743 52605
0 52607 5 1 1 52606
0 52608 7 1 2 75207 95818
0 52609 5 1 1 52608
0 52610 7 1 2 17362 52609
0 52611 5 1 1 52610
0 52612 7 1 2 73909 52611
0 52613 5 1 1 52612
0 52614 7 1 2 52607 52613
0 52615 7 1 2 52601 52614
0 52616 7 1 2 52593 52615
0 52617 7 1 2 52584 52616
0 52618 7 1 2 52576 52617
0 52619 5 1 1 52618
0 52620 7 1 2 60069 52619
0 52621 5 1 1 52620
0 52622 7 1 2 88480 95827
0 52623 5 1 1 52622
0 52624 7 1 2 82780 95819
0 52625 5 1 1 52624
0 52626 7 1 2 65738 95831
0 52627 5 1 1 52626
0 52628 7 1 2 52625 52627
0 52629 5 1 1 52628
0 52630 7 1 2 76517 52629
0 52631 5 1 1 52630
0 52632 7 1 2 52623 52631
0 52633 5 1 1 52632
0 52634 7 1 2 71923 52633
0 52635 5 1 1 52634
0 52636 7 1 2 87537 80548
0 52637 7 1 2 93405 52636
0 52638 5 1 1 52637
0 52639 7 1 2 52635 52638
0 52640 7 1 2 52621 52639
0 52641 7 1 2 52559 52640
0 52642 5 1 1 52641
0 52643 7 1 2 58812 52642
0 52644 5 1 1 52643
0 52645 7 1 2 52516 52644
0 52646 5 1 1 52645
0 52647 7 1 2 58677 52646
0 52648 5 1 1 52647
0 52649 7 1 2 84467 91953
0 52650 5 1 1 52649
0 52651 7 1 2 86394 81438
0 52652 5 1 1 52651
0 52653 7 1 2 86396 52652
0 52654 5 1 1 52653
0 52655 7 1 2 65344 52654
0 52656 5 1 1 52655
0 52657 7 1 2 65100 74643
0 52658 5 1 1 52657
0 52659 7 1 2 14999 52658
0 52660 5 1 1 52659
0 52661 7 1 2 68417 52660
0 52662 5 1 1 52661
0 52663 7 2 2 59387 86113
0 52664 7 1 2 83445 95834
0 52665 5 1 1 52664
0 52666 7 1 2 52662 52665
0 52667 7 1 2 52656 52666
0 52668 5 1 1 52667
0 52669 7 1 2 71552 52668
0 52670 5 1 1 52669
0 52671 7 1 2 69075 94586
0 52672 5 1 1 52671
0 52673 7 1 2 74756 52672
0 52674 5 1 1 52673
0 52675 7 2 2 69852 73270
0 52676 7 1 2 59388 83446
0 52677 7 1 2 95836 52676
0 52678 5 1 1 52677
0 52679 7 1 2 52674 52678
0 52680 7 1 2 52670 52679
0 52681 5 1 1 52680
0 52682 7 1 2 57528 52681
0 52683 5 1 1 52682
0 52684 7 1 2 69131 79315
0 52685 5 1 1 52684
0 52686 7 1 2 79317 52685
0 52687 5 1 1 52686
0 52688 7 1 2 71553 52687
0 52689 5 1 1 52688
0 52690 7 1 2 73295 73136
0 52691 7 1 2 83867 52690
0 52692 5 1 1 52691
0 52693 7 1 2 71231 52692
0 52694 5 1 1 52693
0 52695 7 1 2 52689 52694
0 52696 5 1 1 52695
0 52697 7 1 2 61478 52696
0 52698 5 1 1 52697
0 52699 7 1 2 57808 74644
0 52700 5 1 1 52699
0 52701 7 1 2 6104 52700
0 52702 5 1 1 52701
0 52703 7 1 2 74040 52702
0 52704 5 1 1 52703
0 52705 7 1 2 92916 52704
0 52706 5 1 1 52705
0 52707 7 1 2 71554 52706
0 52708 5 1 1 52707
0 52709 7 1 2 61479 74041
0 52710 7 1 2 90198 52709
0 52711 5 2 1 52710
0 52712 7 1 2 52708 95838
0 52713 7 1 2 52698 52712
0 52714 7 1 2 52683 52713
0 52715 5 1 1 52714
0 52716 7 1 2 58088 52715
0 52717 5 1 1 52716
0 52718 7 1 2 57529 86183
0 52719 5 1 1 52718
0 52720 7 1 2 70848 83868
0 52721 5 1 1 52720
0 52722 7 1 2 59389 52721
0 52723 5 1 1 52722
0 52724 7 1 2 52719 52723
0 52725 5 1 1 52724
0 52726 7 1 2 71232 52725
0 52727 5 1 1 52726
0 52728 7 2 2 59692 76430
0 52729 5 1 1 95840
0 52730 7 2 2 70795 71555
0 52731 7 1 2 95804 95842
0 52732 5 1 1 52731
0 52733 7 1 2 52729 52732
0 52734 5 1 1 52733
0 52735 7 1 2 57809 52734
0 52736 5 1 1 52735
0 52737 7 1 2 65345 93123
0 52738 5 1 1 52737
0 52739 7 1 2 52736 52738
0 52740 5 1 1 52739
0 52741 7 1 2 77160 52740
0 52742 5 1 1 52741
0 52743 7 1 2 52727 52742
0 52744 5 1 1 52743
0 52745 7 1 2 61480 52744
0 52746 5 1 1 52745
0 52747 7 1 2 65739 82241
0 52748 5 1 1 52747
0 52749 7 1 2 67104 52748
0 52750 5 1 1 52749
0 52751 7 1 2 74676 52750
0 52752 5 1 1 52751
0 52753 7 1 2 86159 73745
0 52754 7 1 2 78382 52753
0 52755 5 1 1 52754
0 52756 7 1 2 52752 52755
0 52757 5 1 1 52756
0 52758 7 1 2 71924 52757
0 52759 5 1 1 52758
0 52760 7 3 2 61103 88497
0 52761 5 1 1 95844
0 52762 7 1 2 95358 95845
0 52763 5 1 1 52762
0 52764 7 1 2 61481 95841
0 52765 5 1 1 52764
0 52766 7 1 2 52763 52765
0 52767 5 1 1 52766
0 52768 7 1 2 72251 52767
0 52769 5 1 1 52768
0 52770 7 1 2 73534 83433
0 52771 7 1 2 79756 52770
0 52772 5 1 1 52771
0 52773 7 1 2 52769 52772
0 52774 7 1 2 52759 52773
0 52775 7 1 2 52746 52774
0 52776 7 1 2 52717 52775
0 52777 5 1 1 52776
0 52778 7 1 2 66384 52777
0 52779 5 1 1 52778
0 52780 7 1 2 52650 52779
0 52781 5 1 1 52780
0 52782 7 1 2 66874 52781
0 52783 5 1 1 52782
0 52784 7 1 2 52648 52783
0 52785 5 1 1 52784
0 52786 7 1 2 61994 52785
0 52787 5 1 1 52786
0 52788 7 1 2 87227 83991
0 52789 5 1 1 52788
0 52790 7 1 2 95696 52789
0 52791 5 1 1 52790
0 52792 7 1 2 71758 52791
0 52793 5 1 1 52792
0 52794 7 1 2 65346 95692
0 52795 5 1 1 52794
0 52796 7 1 2 52793 52795
0 52797 5 1 1 52796
0 52798 7 1 2 65740 52797
0 52799 5 1 1 52798
0 52800 7 1 2 68054 84696
0 52801 5 1 1 52800
0 52802 7 1 2 52799 52801
0 52803 5 1 1 52802
0 52804 7 1 2 82978 52803
0 52805 5 1 1 52804
0 52806 7 1 2 63416 95741
0 52807 5 1 1 52806
0 52808 7 1 2 84697 52807
0 52809 5 1 1 52808
0 52810 7 1 2 86949 95747
0 52811 5 1 1 52810
0 52812 7 1 2 52809 52811
0 52813 5 1 1 52812
0 52814 7 1 2 71556 52813
0 52815 5 1 1 52814
0 52816 7 1 2 85140 95744
0 52817 5 1 1 52816
0 52818 7 1 2 84489 52817
0 52819 5 1 1 52818
0 52820 7 1 2 86503 52819
0 52821 5 1 1 52820
0 52822 7 1 2 82979 94933
0 52823 7 1 2 95745 52822
0 52824 5 1 1 52823
0 52825 7 1 2 52821 52824
0 52826 7 1 2 52815 52825
0 52827 7 1 2 52805 52826
0 52828 5 1 1 52827
0 52829 7 1 2 68418 52828
0 52830 5 1 1 52829
0 52831 7 1 2 84698 84334
0 52832 5 1 1 52831
0 52833 7 2 2 86504 78655
0 52834 5 1 1 95847
0 52835 7 1 2 68055 95848
0 52836 5 1 1 52835
0 52837 7 1 2 52832 52836
0 52838 5 1 1 52837
0 52839 7 1 2 58678 52838
0 52840 5 1 1 52839
0 52841 7 1 2 79632 94934
0 52842 5 1 1 52841
0 52843 7 1 2 93415 52842
0 52844 5 1 1 52843
0 52845 7 1 2 58089 52844
0 52846 5 1 1 52845
0 52847 7 1 2 59390 86950
0 52848 5 1 1 52847
0 52849 7 1 2 52846 52848
0 52850 5 1 1 52849
0 52851 7 1 2 69472 52850
0 52852 5 1 1 52851
0 52853 7 2 2 66087 86851
0 52854 7 1 2 81378 95849
0 52855 5 1 1 52854
0 52856 7 4 2 65347 84699
0 52857 5 1 1 95851
0 52858 7 1 2 82446 95852
0 52859 5 1 1 52858
0 52860 7 1 2 52855 52859
0 52861 5 1 1 52860
0 52862 7 1 2 71759 52861
0 52863 5 1 1 52862
0 52864 7 1 2 68178 79609
0 52865 5 1 1 52864
0 52866 7 1 2 86951 52865
0 52867 5 1 1 52866
0 52868 7 1 2 52863 52867
0 52869 7 1 2 52852 52868
0 52870 5 1 1 52869
0 52871 7 1 2 65741 52870
0 52872 5 1 1 52871
0 52873 7 1 2 52840 52872
0 52874 5 1 1 52873
0 52875 7 1 2 71557 52874
0 52876 5 1 1 52875
0 52877 7 1 2 21216 52857
0 52878 5 1 1 52877
0 52879 7 1 2 68646 52878
0 52880 5 1 1 52879
0 52881 7 1 2 86704 95661
0 52882 5 1 1 52881
0 52883 7 1 2 65348 52882
0 52884 5 1 1 52883
0 52885 7 1 2 52880 52884
0 52886 5 1 1 52885
0 52887 7 1 2 58679 52886
0 52888 5 1 1 52887
0 52889 7 1 2 73765 84700
0 52890 5 1 1 52889
0 52891 7 1 2 66088 86822
0 52892 5 1 1 52891
0 52893 7 1 2 52890 52892
0 52894 5 1 1 52893
0 52895 7 1 2 68647 52894
0 52896 5 1 1 52895
0 52897 7 1 2 93416 51582
0 52898 5 1 1 52897
0 52899 7 1 2 65349 52898
0 52900 5 1 1 52899
0 52901 7 1 2 52896 52900
0 52902 5 1 1 52901
0 52903 7 1 2 58366 52902
0 52904 5 1 1 52903
0 52905 7 1 2 52888 52904
0 52906 5 1 1 52905
0 52907 7 1 2 67700 52906
0 52908 5 1 1 52907
0 52909 7 1 2 28123 95749
0 52910 5 1 1 52909
0 52911 7 1 2 58680 52910
0 52912 5 1 1 52911
0 52913 7 1 2 52908 52912
0 52914 5 1 1 52913
0 52915 7 1 2 78618 52914
0 52916 5 1 1 52915
0 52917 7 1 2 84708 52834
0 52918 5 1 1 52917
0 52919 7 1 2 86299 52918
0 52920 5 1 1 52919
0 52921 7 1 2 82447 86505
0 52922 5 1 1 52921
0 52923 7 1 2 95699 52922
0 52924 5 1 1 52923
0 52925 7 1 2 69473 52924
0 52926 5 1 1 52925
0 52927 7 1 2 67878 95690
0 52928 5 1 1 52927
0 52929 7 1 2 52926 52928
0 52930 5 1 1 52929
0 52931 7 1 2 65742 52930
0 52932 5 1 1 52931
0 52933 7 1 2 11650 80577
0 52934 5 1 1 52933
0 52935 7 1 2 94935 52934
0 52936 5 1 1 52935
0 52937 7 1 2 73944 95853
0 52938 5 1 1 52937
0 52939 7 2 2 68056 89697
0 52940 5 2 1 95855
0 52941 7 1 2 74009 95856
0 52942 5 1 1 52941
0 52943 7 1 2 52938 52942
0 52944 5 1 1 52943
0 52945 7 1 2 71760 52944
0 52946 5 1 1 52945
0 52947 7 1 2 52936 52946
0 52948 7 1 2 52932 52947
0 52949 5 1 1 52948
0 52950 7 1 2 82980 52949
0 52951 5 1 1 52950
0 52952 7 1 2 52920 52951
0 52953 7 1 2 52916 52952
0 52954 7 1 2 52876 52953
0 52955 7 1 2 52830 52954
0 52956 5 1 1 52955
0 52957 7 1 2 75770 52956
0 52958 5 1 1 52957
0 52959 7 2 2 77430 82810
0 52960 7 1 2 80673 94479
0 52961 7 1 2 95859 52960
0 52962 5 1 1 52961
0 52963 7 1 2 52958 52962
0 52964 7 1 2 52787 52963
0 52965 5 1 1 52964
0 52966 7 1 2 62139 52965
0 52967 5 1 1 52966
0 52968 7 1 2 87689 95739
0 52969 5 1 1 52968
0 52970 7 2 2 61482 76396
0 52971 7 1 2 94717 95861
0 52972 5 1 1 52971
0 52973 7 1 2 66385 52972
0 52974 7 1 2 52969 52973
0 52975 5 1 1 52974
0 52976 7 1 2 71700 73568
0 52977 5 1 1 52976
0 52978 7 1 2 81819 52977
0 52979 5 1 1 52978
0 52980 7 1 2 62276 52979
0 52981 5 1 1 52980
0 52982 7 1 2 66089 84034
0 52983 5 1 1 52982
0 52984 7 1 2 52981 52983
0 52985 5 1 1 52984
0 52986 7 1 2 84887 52985
0 52987 5 1 1 52986
0 52988 7 1 2 86779 95256
0 52989 5 1 1 52988
0 52990 7 1 2 52987 52989
0 52991 5 1 1 52990
0 52992 7 1 2 60070 52991
0 52993 5 1 1 52992
0 52994 7 1 2 69402 74492
0 52995 7 1 2 95850 52994
0 52996 7 1 2 94115 52995
0 52997 5 1 1 52996
0 52998 7 1 2 52993 52997
0 52999 5 1 1 52998
0 53000 7 1 2 61104 52999
0 53001 5 1 1 53000
0 53002 7 1 2 80729 51732
0 53003 5 1 1 53002
0 53004 7 1 2 73945 93628
0 53005 5 1 1 53004
0 53006 7 1 2 83965 53005
0 53007 5 1 1 53006
0 53008 7 1 2 71233 53007
0 53009 5 1 1 53008
0 53010 7 1 2 53003 53009
0 53011 5 1 1 53010
0 53012 7 1 2 58681 74659
0 53013 7 1 2 53011 53012
0 53014 5 1 1 53013
0 53015 7 1 2 73342 94638
0 53016 5 3 1 53015
0 53017 7 4 2 80873 85096
0 53018 5 1 1 95866
0 53019 7 1 2 95863 95867
0 53020 5 1 1 53019
0 53021 7 1 2 61744 53020
0 53022 7 1 2 53014 53021
0 53023 7 1 2 53001 53022
0 53024 5 1 1 53023
0 53025 7 1 2 66643 53024
0 53026 7 1 2 52975 53025
0 53027 5 1 1 53026
0 53028 7 2 2 88481 95266
0 53029 7 1 2 59391 95870
0 53030 5 1 1 53029
0 53031 7 1 2 79395 75425
0 53032 5 1 1 53031
0 53033 7 1 2 53030 53032
0 53034 5 1 1 53033
0 53035 7 1 2 67863 53034
0 53036 5 1 1 53035
0 53037 7 1 2 83293 70125
0 53038 7 1 2 94599 53037
0 53039 5 1 1 53038
0 53040 7 1 2 71558 53039
0 53041 5 1 1 53040
0 53042 7 1 2 93343 53041
0 53043 5 1 1 53042
0 53044 7 1 2 58813 53043
0 53045 5 1 1 53044
0 53046 7 1 2 68419 95626
0 53047 5 1 1 53046
0 53048 7 1 2 82448 95267
0 53049 5 2 1 53048
0 53050 7 1 2 58814 90979
0 53051 5 1 1 53050
0 53052 7 1 2 95872 53051
0 53053 5 1 1 53052
0 53054 7 1 2 78639 53053
0 53055 5 1 1 53054
0 53056 7 1 2 53047 53055
0 53057 7 1 2 53045 53056
0 53058 7 1 2 53036 53057
0 53059 5 1 1 53058
0 53060 7 1 2 65350 53059
0 53061 5 1 1 53060
0 53062 7 1 2 75944 83993
0 53063 5 1 1 53062
0 53064 7 1 2 69196 95871
0 53065 5 1 1 53064
0 53066 7 1 2 53063 53065
0 53067 5 1 1 53066
0 53068 7 1 2 72252 53067
0 53069 5 1 1 53068
0 53070 7 1 2 77760 14514
0 53071 5 1 1 53070
0 53072 7 1 2 77161 53071
0 53073 5 1 1 53072
0 53074 7 1 2 87402 53073
0 53075 5 1 1 53074
0 53076 7 1 2 58815 53075
0 53077 5 1 1 53076
0 53078 7 1 2 59176 80285
0 53079 7 1 2 94525 53078
0 53080 5 1 1 53079
0 53081 7 1 2 95873 53080
0 53082 7 1 2 53077 53081
0 53083 5 1 1 53082
0 53084 7 1 2 65743 53083
0 53085 5 1 1 53084
0 53086 7 1 2 39512 53085
0 53087 7 1 2 53069 53086
0 53088 7 1 2 53061 53087
0 53089 5 1 1 53088
0 53090 7 1 2 87613 53089
0 53091 5 1 1 53090
0 53092 7 1 2 53027 53091
0 53093 5 1 1 53092
0 53094 7 1 2 62140 53093
0 53095 5 1 1 53094
0 53096 7 2 2 67490 93931
0 53097 7 1 2 86689 95874
0 53098 5 1 1 53097
0 53099 7 1 2 74474 81127
0 53100 5 1 1 53099
0 53101 7 1 2 53098 53100
0 53102 5 1 1 53101
0 53103 7 1 2 63417 53102
0 53104 5 1 1 53103
0 53105 7 2 2 74471 89619
0 53106 7 1 2 90304 95876
0 53107 5 1 1 53106
0 53108 7 1 2 53104 53107
0 53109 5 1 1 53108
0 53110 7 1 2 68277 53109
0 53111 5 1 1 53110
0 53112 7 2 2 87847 90213
0 53113 5 1 1 95878
0 53114 7 1 2 61483 95879
0 53115 5 1 1 53114
0 53116 7 1 2 53111 53115
0 53117 5 1 1 53116
0 53118 7 1 2 62277 53117
0 53119 5 1 1 53118
0 53120 7 1 2 82811 88250
0 53121 7 1 2 95875 53120
0 53122 5 1 1 53121
0 53123 7 1 2 53119 53122
0 53124 5 1 1 53123
0 53125 7 1 2 80874 53124
0 53126 5 1 1 53125
0 53127 7 1 2 64420 75370
0 53128 7 1 2 92528 53127
0 53129 7 1 2 95613 53128
0 53130 5 1 1 53129
0 53131 7 1 2 53126 53130
0 53132 5 1 1 53131
0 53133 7 1 2 69076 53132
0 53134 5 1 1 53133
0 53135 7 1 2 87848 74499
0 53136 5 1 1 53135
0 53137 7 1 2 66875 84028
0 53138 5 1 1 53137
0 53139 7 1 2 53136 53138
0 53140 5 1 1 53139
0 53141 7 1 2 68278 53140
0 53142 5 1 1 53141
0 53143 7 1 2 82889 88281
0 53144 5 2 1 53143
0 53145 7 1 2 61105 74800
0 53146 7 1 2 95880 53145
0 53147 5 1 1 53146
0 53148 7 1 2 53142 53147
0 53149 5 1 1 53148
0 53150 7 1 2 61484 53149
0 53151 5 1 1 53150
0 53152 7 1 2 53151 53113
0 53153 5 1 1 53152
0 53154 7 1 2 80875 53153
0 53155 5 1 1 53154
0 53156 7 1 2 84029 90109
0 53157 7 1 2 93098 53156
0 53158 5 1 1 53157
0 53159 7 1 2 53155 53158
0 53160 5 1 1 53159
0 53161 7 1 2 64421 53160
0 53162 5 1 1 53161
0 53163 7 1 2 74750 89698
0 53164 7 1 2 95783 53163
0 53165 5 1 1 53164
0 53166 7 1 2 53162 53165
0 53167 5 1 1 53166
0 53168 7 1 2 79088 53167
0 53169 5 1 1 53168
0 53170 7 1 2 63418 95759
0 53171 5 1 1 53170
0 53172 7 1 2 95779 53171
0 53173 5 1 1 53172
0 53174 7 1 2 80525 53173
0 53175 5 1 1 53174
0 53176 7 1 2 63922 91286
0 53177 5 1 1 53176
0 53178 7 1 2 53175 53177
0 53179 5 1 1 53178
0 53180 7 1 2 81122 74308
0 53181 7 1 2 53179 53180
0 53182 5 1 1 53181
0 53183 7 1 2 53169 53182
0 53184 7 1 2 53134 53183
0 53185 7 1 2 53095 53184
0 53186 5 1 1 53185
0 53187 7 1 2 64640 53186
0 53188 5 1 1 53187
0 53189 7 1 2 93085 95877
0 53190 5 1 1 53189
0 53191 7 1 2 81476 74751
0 53192 7 1 2 78884 53191
0 53193 5 1 1 53192
0 53194 7 1 2 53190 53193
0 53195 5 1 1 53194
0 53196 7 1 2 63556 94715
0 53197 7 1 2 53195 53196
0 53198 5 1 1 53197
0 53199 7 1 2 53188 53198
0 53200 7 1 2 52967 53199
0 53201 5 1 1 53200
0 53202 7 1 2 67943 53201
0 53203 5 1 1 53202
0 53204 7 3 2 79184 90265
0 53205 5 1 1 95882
0 53206 7 2 2 86335 71377
0 53207 5 1 1 95885
0 53208 7 1 2 53205 53207
0 53209 5 1 1 53208
0 53210 7 1 2 58682 53209
0 53211 5 1 1 53210
0 53212 7 1 2 86805 87153
0 53213 5 1 1 53212
0 53214 7 1 2 87538 80261
0 53215 5 1 1 53214
0 53216 7 1 2 53213 53215
0 53217 5 1 1 53216
0 53218 7 1 2 64641 53217
0 53219 5 1 1 53218
0 53220 7 4 2 59946 88251
0 53221 5 2 1 95887
0 53222 7 1 2 64752 95888
0 53223 5 1 1 53222
0 53224 7 1 2 53219 53223
0 53225 5 1 1 53224
0 53226 7 1 2 69077 53225
0 53227 5 1 1 53226
0 53228 7 4 2 93935 95487
0 53229 7 1 2 78739 95893
0 53230 5 1 1 53229
0 53231 7 1 2 92656 94218
0 53232 5 1 1 53231
0 53233 7 1 2 53230 53232
0 53234 5 1 1 53233
0 53235 7 1 2 61106 53234
0 53236 5 1 1 53235
0 53237 7 1 2 64753 86002
0 53238 7 1 2 86598 53237
0 53239 5 1 1 53238
0 53240 7 1 2 53236 53239
0 53241 7 1 2 53227 53240
0 53242 5 1 1 53241
0 53243 7 1 2 60681 53242
0 53244 5 1 1 53243
0 53245 7 2 2 87795 90595
0 53246 5 1 1 95897
0 53247 7 1 2 64754 95898
0 53248 5 1 1 53247
0 53249 7 1 2 53244 53248
0 53250 5 1 1 53249
0 53251 7 1 2 76231 53250
0 53252 5 1 1 53251
0 53253 7 1 2 68279 78406
0 53254 5 1 1 53253
0 53255 7 1 2 58367 53254
0 53256 5 1 1 53255
0 53257 7 1 2 95894 53256
0 53258 5 1 1 53257
0 53259 7 1 2 85204 87539
0 53260 5 1 1 53259
0 53261 7 1 2 53258 53260
0 53262 5 1 1 53261
0 53263 7 1 2 61107 53262
0 53264 5 1 1 53263
0 53265 7 1 2 75883 93555
0 53266 5 1 1 53265
0 53267 7 1 2 92313 53266
0 53268 5 1 1 53267
0 53269 7 1 2 53264 53268
0 53270 5 1 1 53269
0 53271 7 1 2 68179 53270
0 53272 5 1 1 53271
0 53273 7 1 2 80876 82219
0 53274 5 1 1 53273
0 53275 7 1 2 88621 53274
0 53276 5 1 1 53275
0 53277 7 1 2 64755 53276
0 53278 5 1 1 53277
0 53279 7 1 2 53272 53278
0 53280 7 1 2 53252 53279
0 53281 5 1 1 53280
0 53282 7 1 2 60168 53281
0 53283 5 1 1 53282
0 53284 7 1 2 53211 53283
0 53285 5 1 1 53284
0 53286 7 1 2 58816 53285
0 53287 5 1 1 53286
0 53288 7 1 2 72061 80748
0 53289 5 1 1 53288
0 53290 7 1 2 90596 53289
0 53291 5 1 1 53290
0 53292 7 1 2 95891 53291
0 53293 5 1 1 53292
0 53294 7 1 2 63113 53293
0 53295 5 1 1 53294
0 53296 7 1 2 87296 95119
0 53297 5 1 1 53296
0 53298 7 1 2 66386 85205
0 53299 5 1 1 53298
0 53300 7 1 2 53297 53299
0 53301 5 1 1 53300
0 53302 7 1 2 62531 95116
0 53303 7 1 2 53301 53302
0 53304 5 1 1 53303
0 53305 7 1 2 53295 53304
0 53306 5 1 1 53305
0 53307 7 1 2 68180 53306
0 53308 5 1 1 53307
0 53309 7 2 2 70928 95108
0 53310 5 1 1 95899
0 53311 7 1 2 95892 53310
0 53312 5 1 1 53311
0 53313 7 1 2 69078 53312
0 53314 5 1 1 53313
0 53315 7 1 2 90597 92940
0 53316 7 1 2 42593 53315
0 53317 5 1 1 53316
0 53318 7 1 2 78740 95889
0 53319 5 1 1 53318
0 53320 7 1 2 53317 53319
0 53321 7 1 2 53314 53320
0 53322 5 1 1 53321
0 53323 7 1 2 60682 53322
0 53324 5 1 1 53323
0 53325 7 1 2 53246 53324
0 53326 5 1 1 53325
0 53327 7 1 2 76232 53326
0 53328 5 1 1 53327
0 53329 7 1 2 66387 80845
0 53330 5 1 1 53329
0 53331 7 1 2 25340 53330
0 53332 7 1 2 53328 53331
0 53333 7 1 2 53308 53332
0 53334 5 1 1 53333
0 53335 7 1 2 60071 53334
0 53336 5 1 1 53335
0 53337 7 1 2 87653 53336
0 53338 5 1 1 53337
0 53339 7 1 2 88054 53338
0 53340 5 1 1 53339
0 53341 7 1 2 53287 53340
0 53342 5 1 1 53341
0 53343 7 1 2 58901 53342
0 53344 5 1 1 53343
0 53345 7 1 2 94300 95564
0 53346 5 1 1 53345
0 53347 7 1 2 53344 53346
0 53348 5 1 1 53347
0 53349 7 1 2 67491 53348
0 53350 5 1 1 53349
0 53351 7 1 2 67608 90598
0 53352 5 1 1 53351
0 53353 7 1 2 82600 53352
0 53354 5 2 1 53353
0 53355 7 1 2 67080 95901
0 53356 5 1 1 53355
0 53357 7 2 2 62811 82112
0 53358 7 1 2 79185 95903
0 53359 5 1 1 53358
0 53360 7 1 2 53356 53359
0 53361 5 1 1 53360
0 53362 7 1 2 60072 53361
0 53363 5 1 1 53362
0 53364 7 2 2 75563 76063
0 53365 5 1 1 95905
0 53366 7 1 2 95906 95904
0 53367 5 1 1 53366
0 53368 7 1 2 53363 53367
0 53369 5 1 1 53368
0 53370 7 1 2 64111 53369
0 53371 5 1 1 53370
0 53372 7 1 2 87192 94538
0 53373 5 1 1 53372
0 53374 7 1 2 53371 53373
0 53375 5 1 1 53374
0 53376 7 1 2 70849 53375
0 53377 5 1 1 53376
0 53378 7 1 2 92127 94539
0 53379 5 1 1 53378
0 53380 7 3 2 76713 88456
0 53381 7 1 2 60073 95907
0 53382 5 1 1 53381
0 53383 7 1 2 5212 53365
0 53384 5 1 1 53383
0 53385 7 5 2 61745 53384
0 53386 7 1 2 62532 66644
0 53387 7 1 2 95910 53386
0 53388 5 1 1 53387
0 53389 7 1 2 53382 53388
0 53390 5 1 1 53389
0 53391 7 1 2 64112 53390
0 53392 5 1 1 53391
0 53393 7 1 2 53379 53392
0 53394 5 1 1 53393
0 53395 7 1 2 74877 53394
0 53396 5 1 1 53395
0 53397 7 2 2 64113 90599
0 53398 5 1 1 95915
0 53399 7 2 2 87947 95916
0 53400 5 1 1 95917
0 53401 7 1 2 62533 69809
0 53402 5 1 1 53401
0 53403 7 1 2 63788 85365
0 53404 5 1 1 53403
0 53405 7 2 2 53402 53404
0 53406 7 1 2 67395 95919
0 53407 5 1 1 53406
0 53408 7 1 2 82587 53407
0 53409 5 1 1 53408
0 53410 7 1 2 53400 53409
0 53411 5 1 1 53410
0 53412 7 1 2 77018 53411
0 53413 5 1 1 53412
0 53414 7 1 2 53396 53413
0 53415 7 1 2 53377 53414
0 53416 5 1 1 53415
0 53417 7 1 2 61108 53416
0 53418 5 1 1 53417
0 53419 7 1 2 80526 95900
0 53420 5 1 1 53419
0 53421 7 1 2 76385 95113
0 53422 5 1 1 53421
0 53423 7 1 2 53420 53422
0 53424 5 1 1 53423
0 53425 7 1 2 77019 53424
0 53426 5 1 1 53425
0 53427 7 1 2 57810 94148
0 53428 5 1 1 53427
0 53429 7 1 2 80581 53428
0 53430 5 1 1 53429
0 53431 7 1 2 71925 53430
0 53432 5 1 1 53431
0 53433 7 1 2 95908 53432
0 53434 5 1 1 53433
0 53435 7 1 2 64845 91907
0 53436 7 1 2 95800 53435
0 53437 5 1 1 53436
0 53438 7 1 2 53434 53437
0 53439 5 1 1 53438
0 53440 7 1 2 60074 53439
0 53441 5 1 1 53440
0 53442 7 1 2 63923 84459
0 53443 7 1 2 76936 53442
0 53444 7 1 2 95764 53443
0 53445 5 1 1 53444
0 53446 7 1 2 53441 53445
0 53447 5 1 1 53446
0 53448 7 1 2 62812 53447
0 53449 5 1 1 53448
0 53450 7 1 2 53426 53449
0 53451 7 1 2 53418 53450
0 53452 5 1 1 53451
0 53453 7 1 2 70231 53452
0 53454 5 1 1 53453
0 53455 7 1 2 62534 81100
0 53456 5 1 1 53455
0 53457 7 1 2 73483 53456
0 53458 5 1 1 53457
0 53459 7 1 2 53458 95909
0 53460 5 1 1 53459
0 53461 7 1 2 68280 95142
0 53462 5 1 1 53461
0 53463 7 1 2 68944 53462
0 53464 5 1 1 53463
0 53465 7 1 2 59947 91474
0 53466 7 1 2 53464 53465
0 53467 5 1 1 53466
0 53468 7 1 2 53460 53467
0 53469 5 1 1 53468
0 53470 7 1 2 60075 53469
0 53471 5 1 1 53470
0 53472 7 2 2 70929 86678
0 53473 7 1 2 87194 84135
0 53474 7 1 2 95921 53473
0 53475 5 1 1 53474
0 53476 7 1 2 53471 53475
0 53477 5 1 1 53476
0 53478 7 1 2 62813 53477
0 53479 5 1 1 53478
0 53480 7 2 2 66388 92414
0 53481 5 1 1 95923
0 53482 7 1 2 95104 53481
0 53483 5 1 1 53482
0 53484 7 1 2 70126 53483
0 53485 5 1 1 53484
0 53486 7 1 2 60683 95101
0 53487 5 1 1 53486
0 53488 7 1 2 53398 53487
0 53489 5 1 1 53488
0 53490 7 1 2 67797 53489
0 53491 5 1 1 53490
0 53492 7 1 2 53485 53491
0 53493 5 1 1 53492
0 53494 7 1 2 61109 53493
0 53495 5 1 1 53494
0 53496 7 1 2 84603 95924
0 53497 5 1 1 53496
0 53498 7 1 2 53495 53497
0 53499 5 1 1 53498
0 53500 7 1 2 77020 53499
0 53501 5 1 1 53500
0 53502 7 1 2 53479 53501
0 53503 5 1 1 53502
0 53504 7 1 2 69079 53503
0 53505 5 1 1 53504
0 53506 7 1 2 58683 84424
0 53507 5 1 1 53506
0 53508 7 1 2 66999 53507
0 53509 5 1 1 53508
0 53510 7 1 2 70897 92793
0 53511 5 2 1 53510
0 53512 7 1 2 61995 67798
0 53513 7 1 2 80335 53512
0 53514 7 1 2 95925 53513
0 53515 5 1 1 53514
0 53516 7 1 2 53509 53515
0 53517 5 1 1 53516
0 53518 7 1 2 82588 53517
0 53519 5 1 1 53518
0 53520 7 1 2 76714 74945
0 53521 7 1 2 32870 53520
0 53522 5 1 1 53521
0 53523 7 1 2 75601 53522
0 53524 5 1 1 53523
0 53525 7 1 2 88457 53524
0 53526 5 1 1 53525
0 53527 7 1 2 53519 53526
0 53528 5 1 1 53527
0 53529 7 1 2 60076 53528
0 53530 5 1 1 53529
0 53531 7 1 2 76064 91122
0 53532 5 1 1 53531
0 53533 7 1 2 87629 67000
0 53534 5 1 1 53533
0 53535 7 1 2 53532 53534
0 53536 5 1 1 53535
0 53537 7 1 2 58684 53536
0 53538 5 1 1 53537
0 53539 7 2 2 84877 78709
0 53540 7 1 2 69220 95765
0 53541 7 1 2 95927 53540
0 53542 5 1 1 53541
0 53543 7 1 2 63655 53542
0 53544 7 1 2 53538 53543
0 53545 7 1 2 53530 53544
0 53546 7 1 2 53505 53545
0 53547 7 1 2 53454 53546
0 53548 5 1 1 53547
0 53549 7 1 2 74947 32915
0 53550 5 1 1 53549
0 53551 7 1 2 67799 53550
0 53552 5 1 1 53551
0 53553 7 1 2 77682 94788
0 53554 5 1 1 53553
0 53555 7 1 2 84418 53554
0 53556 7 1 2 53552 53555
0 53557 5 1 1 53556
0 53558 7 1 2 90600 53557
0 53559 5 1 1 53558
0 53560 7 1 2 67800 76559
0 53561 7 1 2 89824 53560
0 53562 5 1 1 53561
0 53563 7 1 2 53559 53562
0 53564 5 1 1 53563
0 53565 7 1 2 76035 53564
0 53566 5 1 1 53565
0 53567 7 1 2 84393 86833
0 53568 7 1 2 95886 53567
0 53569 5 1 1 53568
0 53570 7 1 2 53566 53569
0 53571 5 1 1 53570
0 53572 7 1 2 70232 53571
0 53573 5 1 1 53572
0 53574 7 1 2 95926 95911
0 53575 5 1 1 53574
0 53576 7 5 2 82715 93167
0 53577 7 1 2 83905 95929
0 53578 5 1 1 53577
0 53579 7 1 2 53575 53578
0 53580 5 1 1 53579
0 53581 7 1 2 75841 53580
0 53582 5 1 1 53581
0 53583 7 2 2 62535 95930
0 53584 5 1 1 95934
0 53585 7 2 2 68537 75133
0 53586 7 1 2 95935 95936
0 53587 5 1 1 53586
0 53588 7 1 2 53582 53587
0 53589 5 1 1 53588
0 53590 7 1 2 60420 53589
0 53591 5 1 1 53590
0 53592 7 1 2 76715 78057
0 53593 7 1 2 91994 53592
0 53594 5 1 1 53593
0 53595 7 1 2 60077 75602
0 53596 7 1 2 53594 53595
0 53597 5 1 1 53596
0 53598 7 1 2 82716 94222
0 53599 7 1 2 53597 53598
0 53600 5 1 1 53599
0 53601 7 1 2 53591 53600
0 53602 7 1 2 53573 53601
0 53603 5 1 1 53602
0 53604 7 1 2 61996 53603
0 53605 5 1 1 53604
0 53606 7 1 2 68181 95931
0 53607 5 1 1 53606
0 53608 7 1 2 70930 95912
0 53609 5 1 1 53608
0 53610 7 1 2 53607 53609
0 53611 5 1 1 53610
0 53612 7 1 2 70850 53611
0 53613 5 1 1 53612
0 53614 7 1 2 62278 95913
0 53615 5 1 1 53614
0 53616 7 1 2 53584 53615
0 53617 5 1 1 53616
0 53618 7 1 2 87119 53617
0 53619 5 1 1 53618
0 53620 7 1 2 53613 53619
0 53621 5 1 1 53620
0 53622 7 1 2 61110 53621
0 53623 5 1 1 53622
0 53624 7 1 2 62536 92770
0 53625 5 1 1 53624
0 53626 7 1 2 73910 53625
0 53627 5 1 1 53626
0 53628 7 1 2 95932 53627
0 53629 5 1 1 53628
0 53630 7 1 2 53623 53629
0 53631 5 1 1 53630
0 53632 7 1 2 61997 53631
0 53633 5 1 1 53632
0 53634 7 1 2 67229 86547
0 53635 7 1 2 95542 53634
0 53636 7 1 2 95922 53635
0 53637 5 1 1 53636
0 53638 7 1 2 53633 53637
0 53639 5 1 1 53638
0 53640 7 1 2 69080 53639
0 53641 5 1 1 53640
0 53642 7 1 2 80321 95920
0 53643 5 1 1 53642
0 53644 7 1 2 95914 53643
0 53645 5 1 1 53644
0 53646 7 1 2 76036 95902
0 53647 5 1 1 53646
0 53648 7 2 2 76065 92273
0 53649 5 1 1 95938
0 53650 7 1 2 53647 53649
0 53651 5 1 1 53650
0 53652 7 1 2 72225 53651
0 53653 5 1 1 53652
0 53654 7 1 2 76037 95918
0 53655 5 1 1 53654
0 53656 7 1 2 53653 53655
0 53657 7 1 2 53645 53656
0 53658 5 1 1 53657
0 53659 7 1 2 61998 53658
0 53660 5 1 1 53659
0 53661 7 1 2 87677 95144
0 53662 5 1 1 53661
0 53663 7 1 2 76038 91413
0 53664 5 1 1 53663
0 53665 7 1 2 53662 53664
0 53666 5 1 1 53665
0 53667 7 1 2 89803 53666
0 53668 5 1 1 53667
0 53669 7 1 2 84215 95933
0 53670 5 1 1 53669
0 53671 7 1 2 53668 53670
0 53672 5 1 1 53671
0 53673 7 1 2 74878 53672
0 53674 5 1 1 53673
0 53675 7 1 2 70851 82113
0 53676 7 1 2 79304 53675
0 53677 7 1 2 91531 53676
0 53678 5 1 1 53677
0 53679 7 1 2 53674 53678
0 53680 7 1 2 53660 53679
0 53681 5 1 1 53680
0 53682 7 1 2 61111 53681
0 53683 5 1 1 53682
0 53684 7 1 2 70233 77476
0 53685 7 1 2 79305 53684
0 53686 7 1 2 89434 95801
0 53687 7 1 2 53685 53686
0 53688 5 1 1 53687
0 53689 7 1 2 82114 86685
0 53690 7 1 2 95928 53689
0 53691 5 1 1 53690
0 53692 7 1 2 58902 53691
0 53693 7 1 2 53688 53692
0 53694 7 1 2 53683 53693
0 53695 7 1 2 53641 53694
0 53696 7 1 2 53605 53695
0 53697 5 1 1 53696
0 53698 7 1 2 53548 53697
0 53699 5 1 1 53698
0 53700 7 1 2 63557 53699
0 53701 5 1 1 53700
0 53702 7 1 2 29062 52036
0 53703 5 1 1 53702
0 53704 7 1 2 58685 53703
0 53705 5 1 1 53704
0 53706 7 1 2 63924 84086
0 53707 5 1 1 53706
0 53708 7 1 2 65744 53707
0 53709 5 1 1 53708
0 53710 7 1 2 64114 76252
0 53711 7 1 2 53709 53710
0 53712 5 1 1 53711
0 53713 7 1 2 93261 53712
0 53714 5 1 1 53713
0 53715 7 1 2 62814 53714
0 53716 5 1 1 53715
0 53717 7 1 2 77814 93672
0 53718 7 1 2 53716 53717
0 53719 5 1 1 53718
0 53720 7 1 2 66645 95895
0 53721 7 1 2 53719 53720
0 53722 5 1 1 53721
0 53723 7 1 2 53705 53722
0 53724 5 1 1 53723
0 53725 7 1 2 69561 53724
0 53726 5 1 1 53725
0 53727 7 1 2 1544 95106
0 53728 5 1 1 53727
0 53729 7 2 2 85191 92839
0 53730 7 1 2 63419 95940
0 53731 5 1 1 53730
0 53732 7 1 2 53728 53731
0 53733 5 1 1 53732
0 53734 7 1 2 60684 53733
0 53735 5 1 1 53734
0 53736 7 1 2 76716 78604
0 53737 5 1 1 53736
0 53738 7 1 2 75603 53737
0 53739 7 1 2 53735 53738
0 53740 5 1 1 53739
0 53741 7 1 2 66389 53740
0 53742 5 1 1 53741
0 53743 7 1 2 67230 95890
0 53744 5 1 1 53743
0 53745 7 1 2 53742 53744
0 53746 5 1 1 53745
0 53747 7 1 2 64756 53746
0 53748 5 1 1 53747
0 53749 7 1 2 31367 47058
0 53750 5 1 1 53749
0 53751 7 1 2 63420 53750
0 53752 5 1 1 53751
0 53753 7 1 2 64757 89837
0 53754 5 1 1 53753
0 53755 7 1 2 53752 53754
0 53756 5 2 1 53755
0 53757 7 1 2 93187 95942
0 53758 5 1 1 53757
0 53759 7 2 2 76717 87540
0 53760 7 1 2 90729 95944
0 53761 5 1 1 53760
0 53762 7 1 2 53758 53761
0 53763 5 1 1 53762
0 53764 7 1 2 61112 53763
0 53765 5 1 1 53764
0 53766 7 1 2 66390 86679
0 53767 7 1 2 95941 53766
0 53768 5 1 1 53767
0 53769 7 1 2 53765 53768
0 53770 5 1 1 53769
0 53771 7 1 2 70852 53770
0 53772 5 1 1 53771
0 53773 7 1 2 61113 93265
0 53774 5 1 1 53773
0 53775 7 1 2 85104 53774
0 53776 5 1 1 53775
0 53777 7 1 2 87541 53776
0 53778 5 1 1 53777
0 53779 7 1 2 69403 83966
0 53780 7 1 2 95896 53779
0 53781 5 1 1 53780
0 53782 7 1 2 53778 53781
0 53783 5 1 1 53782
0 53784 7 1 2 67801 53783
0 53785 5 1 1 53784
0 53786 7 1 2 95293 47313
0 53787 5 1 1 53786
0 53788 7 1 2 63421 53787
0 53789 5 1 1 53788
0 53790 7 1 2 89829 91913
0 53791 5 1 1 53790
0 53792 7 1 2 64758 53791
0 53793 5 1 1 53792
0 53794 7 1 2 53789 53793
0 53795 5 1 1 53794
0 53796 7 1 2 93317 53795
0 53797 5 1 1 53796
0 53798 7 1 2 95121 95945
0 53799 5 1 1 53798
0 53800 7 1 2 53797 53799
0 53801 7 1 2 53785 53800
0 53802 5 1 1 53801
0 53803 7 1 2 68888 53802
0 53804 5 1 1 53803
0 53805 7 1 2 93281 95943
0 53806 5 1 1 53805
0 53807 7 1 2 71837 93266
0 53808 5 1 1 53807
0 53809 7 1 2 85105 53808
0 53810 5 1 1 53809
0 53811 7 1 2 92556 53810
0 53812 5 1 1 53811
0 53813 7 1 2 53806 53812
0 53814 5 1 1 53813
0 53815 7 1 2 70651 53814
0 53816 5 1 1 53815
0 53817 7 1 2 63422 78605
0 53818 7 1 2 87630 53817
0 53819 5 1 1 53818
0 53820 7 1 2 53816 53819
0 53821 7 1 2 53804 53820
0 53822 7 1 2 53772 53821
0 53823 7 1 2 53748 53822
0 53824 5 1 1 53823
0 53825 7 1 2 61999 69565
0 53826 7 1 2 53824 53825
0 53827 5 1 1 53826
0 53828 7 1 2 53726 53827
0 53829 5 1 1 53828
0 53830 7 1 2 67947 53829
0 53831 5 1 1 53830
0 53832 7 1 2 58817 53831
0 53833 5 1 1 53832
0 53834 7 1 2 63114 53833
0 53835 7 1 2 53701 53834
0 53836 5 1 1 53835
0 53837 7 4 2 79831 94287
0 53838 7 1 2 93027 95946
0 53839 5 1 1 53838
0 53840 7 2 2 77179 88252
0 53841 7 1 2 64115 77243
0 53842 7 1 2 87160 53841
0 53843 7 1 2 95950 53842
0 53844 5 1 1 53843
0 53845 7 1 2 53839 53844
0 53846 5 1 1 53845
0 53847 7 1 2 60685 53846
0 53848 5 1 1 53847
0 53849 7 2 2 61114 91236
0 53850 7 1 2 85385 95781
0 53851 7 1 2 95952 53850
0 53852 5 1 1 53851
0 53853 7 1 2 95482 53852
0 53854 5 1 1 53853
0 53855 7 1 2 62815 53854
0 53856 5 1 1 53855
0 53857 7 1 2 63558 85627
0 53858 7 1 2 87642 53857
0 53859 5 1 1 53858
0 53860 7 1 2 53856 53859
0 53861 7 1 2 53848 53860
0 53862 5 1 1 53861
0 53863 7 1 2 70544 53862
0 53864 5 1 1 53863
0 53865 7 1 2 66391 79610
0 53866 7 1 2 93925 53865
0 53867 5 1 1 53866
0 53868 7 1 2 67231 88061
0 53869 7 1 2 95951 53868
0 53870 5 1 1 53869
0 53871 7 1 2 53867 53870
0 53872 5 1 1 53871
0 53873 7 1 2 60686 53872
0 53874 5 1 1 53873
0 53875 7 1 2 94301 95883
0 53876 5 1 1 53875
0 53877 7 1 2 89342 90751
0 53878 7 1 2 95953 53877
0 53879 5 1 1 53878
0 53880 7 1 2 53876 53879
0 53881 5 1 1 53880
0 53882 7 1 2 68182 53881
0 53883 5 1 1 53882
0 53884 7 1 2 53874 53883
0 53885 7 1 2 53864 53884
0 53886 5 1 1 53885
0 53887 7 1 2 62000 53886
0 53888 5 1 1 53887
0 53889 7 1 2 86431 70895
0 53890 7 1 2 95111 53889
0 53891 5 1 1 53890
0 53892 7 1 2 87449 53891
0 53893 5 1 1 53892
0 53894 7 1 2 62537 53893
0 53895 5 1 1 53894
0 53896 7 1 2 77484 90841
0 53897 5 1 1 53896
0 53898 7 1 2 87450 53897
0 53899 5 1 1 53898
0 53900 7 1 2 69081 53899
0 53901 5 1 1 53900
0 53902 7 1 2 31865 53901
0 53903 7 1 2 53895 53902
0 53904 5 1 1 53903
0 53905 7 1 2 70853 53904
0 53906 5 1 1 53905
0 53907 7 1 2 70738 93206
0 53908 5 1 1 53907
0 53909 7 1 2 75604 53908
0 53910 5 1 1 53909
0 53911 7 1 2 66392 78353
0 53912 7 1 2 53910 53911
0 53913 5 1 1 53912
0 53914 7 1 2 70739 92535
0 53915 7 1 2 77739 53914
0 53916 5 1 1 53915
0 53917 7 1 2 87120 88562
0 53918 5 1 1 53917
0 53919 7 1 2 53916 53918
0 53920 7 1 2 19684 53919
0 53921 7 1 2 53913 53920
0 53922 7 1 2 53906 53921
0 53923 5 1 1 53922
0 53924 7 1 2 72749 53923
0 53925 5 1 1 53924
0 53926 7 1 2 23426 92922
0 53927 7 1 2 94675 53926
0 53928 5 1 1 53927
0 53929 7 1 2 72756 88018
0 53930 7 1 2 53928 53929
0 53931 5 1 1 53930
0 53932 7 1 2 53925 53931
0 53933 5 1 1 53932
0 53934 7 1 2 66950 53933
0 53935 5 1 1 53934
0 53936 7 1 2 53888 53935
0 53937 7 1 2 53836 53936
0 53938 5 1 1 53937
0 53939 7 1 2 66731 53938
0 53940 5 1 1 53939
0 53941 7 1 2 53350 53940
0 53942 5 1 1 53941
0 53943 7 1 2 73704 53942
0 53944 5 1 1 53943
0 53945 7 1 2 84878 86424
0 53946 5 1 1 53945
0 53947 7 1 2 60687 91439
0 53948 7 1 2 86780 53947
0 53949 5 1 1 53948
0 53950 7 1 2 53946 53949
0 53951 5 1 1 53950
0 53952 7 1 2 64422 53951
0 53953 5 1 1 53952
0 53954 7 2 2 87761 80674
0 53955 5 1 1 95954
0 53956 7 1 2 53953 53955
0 53957 5 1 1 53956
0 53958 7 1 2 62279 53957
0 53959 5 1 1 53958
0 53960 7 1 2 70884 84268
0 53961 5 1 1 53960
0 53962 7 1 2 88073 53961
0 53963 5 1 1 53962
0 53964 7 1 2 84888 53963
0 53965 5 1 1 53964
0 53966 7 1 2 53959 53965
0 53967 5 1 1 53966
0 53968 7 1 2 61115 53967
0 53969 5 1 1 53968
0 53970 7 1 2 85052 95955
0 53971 5 1 1 53970
0 53972 7 1 2 53969 53971
0 53973 5 1 1 53972
0 53974 7 1 2 66876 53973
0 53975 5 1 1 53974
0 53976 7 1 2 70796 69716
0 53977 7 1 2 85811 93708
0 53978 7 1 2 53976 53977
0 53979 7 1 2 95124 53978
0 53980 5 1 1 53979
0 53981 7 1 2 53975 53980
0 53982 5 1 1 53981
0 53983 7 1 2 61746 53982
0 53984 5 1 1 53983
0 53985 7 1 2 71559 94002
0 53986 5 1 1 53985
0 53987 7 1 2 65745 82981
0 53988 7 1 2 94170 53987
0 53989 5 1 1 53988
0 53990 7 1 2 53986 53989
0 53991 5 1 1 53990
0 53992 7 1 2 67396 53991
0 53993 5 1 1 53992
0 53994 7 1 2 85306 81451
0 53995 5 1 1 53994
0 53996 7 1 2 87407 53995
0 53997 5 1 1 53996
0 53998 7 1 2 65351 53997
0 53999 5 1 1 53998
0 54000 7 1 2 58686 87010
0 54001 5 1 1 54000
0 54002 7 1 2 53999 54001
0 54003 5 1 1 54002
0 54004 7 1 2 72918 54003
0 54005 5 1 1 54004
0 54006 7 1 2 86884 95673
0 54007 5 1 1 54006
0 54008 7 1 2 72659 4851
0 54009 5 1 1 54008
0 54010 7 1 2 54007 54009
0 54011 5 1 1 54010
0 54012 7 1 2 66090 54011
0 54013 5 1 1 54012
0 54014 7 1 2 54005 54013
0 54015 7 1 2 82982 93887
0 54016 5 1 1 54015
0 54017 7 1 2 63423 73809
0 54018 5 1 1 54017
0 54019 7 1 2 82293 54018
0 54020 5 1 1 54019
0 54021 7 2 2 54016 54020
0 54022 5 1 1 95956
0 54023 7 1 2 81636 54022
0 54024 5 1 1 54023
0 54025 7 1 2 79603 80246
0 54026 5 1 1 54025
0 54027 7 1 2 86929 54026
0 54028 5 2 1 54027
0 54029 7 1 2 65352 95958
0 54030 5 1 1 54029
0 54031 7 1 2 7037 54030
0 54032 5 1 1 54031
0 54033 7 1 2 85538 54032
0 54034 5 1 1 54033
0 54035 7 1 2 54024 54034
0 54036 7 1 2 54014 54035
0 54037 7 1 2 53993 54036
0 54038 5 1 1 54037
0 54039 7 1 2 82189 54038
0 54040 5 1 1 54039
0 54041 7 1 2 53984 54040
0 54042 5 1 1 54041
0 54043 7 1 2 66646 54042
0 54044 5 1 1 54043
0 54045 7 1 2 73807 83597
0 54046 5 1 1 54045
0 54047 7 1 2 80595 54046
0 54048 5 1 1 54047
0 54049 7 1 2 71560 54048
0 54050 5 1 1 54049
0 54051 7 3 2 85534 85973
0 54052 5 6 1 95960
0 54053 7 1 2 85232 95963
0 54054 5 1 1 54053
0 54055 7 1 2 90803 54054
0 54056 5 1 1 54055
0 54057 7 1 2 67397 54056
0 54058 5 1 1 54057
0 54059 7 1 2 35473 35748
0 54060 5 1 1 54059
0 54061 7 1 2 82983 54060
0 54062 5 1 1 54061
0 54063 7 1 2 54058 54062
0 54064 7 1 2 54050 54063
0 54065 5 1 1 54064
0 54066 7 1 2 68420 54065
0 54067 5 1 1 54066
0 54068 7 1 2 71616 81307
0 54069 5 1 1 54068
0 54070 7 1 2 82984 82150
0 54071 7 1 2 54069 54070
0 54072 5 1 1 54071
0 54073 7 1 2 71561 71628
0 54074 7 1 2 92923 54073
0 54075 5 1 1 54074
0 54076 7 1 2 85187 54075
0 54077 7 1 2 54072 54076
0 54078 5 1 1 54077
0 54079 7 1 2 66091 54078
0 54080 5 1 1 54079
0 54081 7 1 2 66092 84846
0 54082 5 1 1 54081
0 54083 7 1 2 73881 95964
0 54084 5 1 1 54083
0 54085 7 1 2 54082 54084
0 54086 5 1 1 54085
0 54087 7 1 2 75884 54086
0 54088 5 1 1 54087
0 54089 7 1 2 95957 54088
0 54090 5 1 1 54089
0 54091 7 1 2 78640 54090
0 54092 5 1 1 54091
0 54093 7 1 2 85915 67898
0 54094 5 1 1 54093
0 54095 7 1 2 85141 94127
0 54096 5 1 1 54095
0 54097 7 1 2 54094 54096
0 54098 5 1 1 54097
0 54099 7 1 2 65746 54098
0 54100 5 1 1 54099
0 54101 7 1 2 15301 54100
0 54102 7 1 2 54092 54101
0 54103 7 1 2 54080 54102
0 54104 7 1 2 54067 54103
0 54105 5 1 1 54104
0 54106 7 1 2 95389 54105
0 54107 5 1 1 54106
0 54108 7 1 2 54044 54107
0 54109 5 1 1 54108
0 54110 7 1 2 64642 54109
0 54111 5 1 1 54110
0 54112 7 1 2 84425 89772
0 54113 5 1 1 54112
0 54114 7 1 2 80746 94049
0 54115 5 1 1 54114
0 54116 7 1 2 67398 54115
0 54117 5 1 1 54116
0 54118 7 1 2 85844 78137
0 54119 5 1 1 54118
0 54120 7 1 2 54117 54119
0 54121 5 1 1 54120
0 54122 7 1 2 71761 54121
0 54123 5 1 1 54122
0 54124 7 1 2 57811 73955
0 54125 5 1 1 54124
0 54126 7 1 2 83967 54125
0 54127 5 1 1 54126
0 54128 7 1 2 71762 54127
0 54129 5 1 1 54128
0 54130 7 1 2 67701 84138
0 54131 5 1 1 54130
0 54132 7 1 2 92868 54131
0 54133 7 1 2 54129 54132
0 54134 5 1 1 54133
0 54135 7 1 2 65353 54134
0 54136 5 1 1 54135
0 54137 7 1 2 54123 54136
0 54138 5 1 1 54137
0 54139 7 1 2 57530 54138
0 54140 5 1 1 54139
0 54141 7 2 2 65354 94596
0 54142 5 1 1 95969
0 54143 7 1 2 87035 54142
0 54144 5 1 1 54143
0 54145 7 1 2 69901 54144
0 54146 5 1 1 54145
0 54147 7 1 2 17822 54146
0 54148 7 1 2 54140 54147
0 54149 5 1 1 54148
0 54150 7 1 2 61747 54149
0 54151 5 1 1 54150
0 54152 7 1 2 54113 54151
0 54153 5 1 1 54152
0 54154 7 1 2 71234 54153
0 54155 5 1 1 54154
0 54156 7 1 2 72531 87212
0 54157 5 2 1 54156
0 54158 7 1 2 86705 95971
0 54159 5 1 1 54158
0 54160 7 1 2 57812 54159
0 54161 5 1 1 54160
0 54162 7 2 2 73766 86506
0 54163 5 1 1 95973
0 54164 7 1 2 54161 54163
0 54165 5 1 1 54164
0 54166 7 1 2 67399 54165
0 54167 5 1 1 54166
0 54168 7 1 2 57813 94811
0 54169 5 1 1 54168
0 54170 7 1 2 12186 54169
0 54171 5 1 1 54170
0 54172 7 1 2 81513 54171
0 54173 5 1 1 54172
0 54174 7 1 2 54167 54173
0 54175 5 1 1 54174
0 54176 7 1 2 58368 54175
0 54177 5 1 1 54176
0 54178 7 1 2 75346 94982
0 54179 5 1 1 54178
0 54180 7 1 2 95857 54179
0 54181 5 1 1 54180
0 54182 7 1 2 74162 54181
0 54183 5 1 1 54182
0 54184 7 1 2 54177 54183
0 54185 5 1 1 54184
0 54186 7 1 2 74042 54185
0 54187 5 1 1 54186
0 54188 7 1 2 72532 95655
0 54189 5 1 1 54188
0 54190 7 1 2 84070 95509
0 54191 5 1 1 54190
0 54192 7 1 2 54189 54191
0 54193 5 1 1 54192
0 54194 7 1 2 58090 54193
0 54195 5 1 1 54194
0 54196 7 2 2 86507 70447
0 54197 7 1 2 71235 95975
0 54198 5 1 1 54197
0 54199 7 1 2 54195 54198
0 54200 5 1 1 54199
0 54201 7 1 2 69095 54200
0 54202 5 1 1 54201
0 54203 7 1 2 90495 95376
0 54204 5 1 1 54203
0 54205 7 1 2 89773 54204
0 54206 5 1 1 54205
0 54207 7 1 2 68421 54206
0 54208 5 1 1 54207
0 54209 7 1 2 66093 75257
0 54210 7 1 2 94245 54209
0 54211 5 1 1 54210
0 54212 7 1 2 54208 54211
0 54213 5 1 1 54212
0 54214 7 1 2 68057 54213
0 54215 5 1 1 54214
0 54216 7 1 2 74226 89699
0 54217 5 1 1 54216
0 54218 7 1 2 89774 54217
0 54219 5 1 1 54218
0 54220 7 1 2 59036 54219
0 54221 5 1 1 54220
0 54222 7 1 2 74520 84595
0 54223 5 1 1 54222
0 54224 7 1 2 54221 54223
0 54225 5 1 1 54224
0 54226 7 1 2 67899 54225
0 54227 5 1 1 54226
0 54228 7 1 2 71337 69903
0 54229 5 1 1 54228
0 54230 7 1 2 58091 95976
0 54231 5 1 1 54230
0 54232 7 1 2 95972 54231
0 54233 5 1 1 54232
0 54234 7 1 2 54229 54233
0 54235 5 1 1 54234
0 54236 7 1 2 54227 54235
0 54237 7 1 2 54215 54236
0 54238 5 1 1 54237
0 54239 7 1 2 71562 54238
0 54240 5 1 1 54239
0 54241 7 1 2 54202 54240
0 54242 7 1 2 54187 54241
0 54243 7 1 2 54155 54242
0 54244 5 1 1 54243
0 54245 7 1 2 76931 54244
0 54246 5 1 1 54245
0 54247 7 1 2 72937 88259
0 54248 5 1 1 54247
0 54249 7 1 2 90935 54248
0 54250 5 1 1 54249
0 54251 7 1 2 70797 54250
0 54252 5 1 1 54251
0 54253 7 1 2 59392 95501
0 54254 5 1 1 54253
0 54255 7 1 2 54252 54254
0 54256 5 1 1 54255
0 54257 7 1 2 57531 54256
0 54258 5 1 1 54257
0 54259 7 1 2 73491 74077
0 54260 5 1 1 54259
0 54261 7 1 2 54258 54260
0 54262 5 1 1 54261
0 54263 7 1 2 58092 54262
0 54264 5 1 1 54263
0 54265 7 1 2 70359 91220
0 54266 5 1 1 54265
0 54267 7 2 2 70798 74159
0 54268 7 1 2 54266 95977
0 54269 5 1 1 54268
0 54270 7 1 2 54264 54269
0 54271 5 1 1 54270
0 54272 7 1 2 61748 54271
0 54273 5 1 1 54272
0 54274 7 1 2 73946 86508
0 54275 5 1 1 54274
0 54276 7 1 2 94926 54275
0 54277 5 1 1 54276
0 54278 7 1 2 75885 54277
0 54279 5 1 1 54278
0 54280 7 1 2 74181 95694
0 54281 5 1 1 54280
0 54282 7 1 2 95858 54281
0 54283 7 1 2 54279 54282
0 54284 5 1 1 54283
0 54285 7 1 2 71763 54284
0 54286 5 1 1 54285
0 54287 7 1 2 73947 78337
0 54288 5 1 1 54287
0 54289 7 1 2 81081 54288
0 54290 5 1 1 54289
0 54291 7 1 2 86509 54290
0 54292 5 1 1 54291
0 54293 7 1 2 84596 94277
0 54294 5 1 1 54293
0 54295 7 1 2 54292 54294
0 54296 5 1 1 54295
0 54297 7 1 2 71926 54296
0 54298 5 1 1 54297
0 54299 7 1 2 68812 77196
0 54300 5 1 1 54299
0 54301 7 1 2 36336 54300
0 54302 5 1 1 54301
0 54303 7 1 2 84701 54302
0 54304 5 1 1 54303
0 54305 7 1 2 57814 95241
0 54306 5 1 1 54305
0 54307 7 1 2 78330 84597
0 54308 5 1 1 54307
0 54309 7 1 2 54306 54308
0 54310 5 1 1 54309
0 54311 7 1 2 73911 54310
0 54312 5 1 1 54311
0 54313 7 1 2 54304 54312
0 54314 7 1 2 54298 54313
0 54315 7 1 2 54286 54314
0 54316 7 1 2 54273 54315
0 54317 5 1 1 54316
0 54318 7 1 2 71563 54317
0 54319 5 1 1 54318
0 54320 7 1 2 81637 43017
0 54321 5 1 1 54320
0 54322 7 1 2 90936 95642
0 54323 5 1 1 54322
0 54324 7 1 2 58093 54323
0 54325 5 1 1 54324
0 54326 7 1 2 78619 94171
0 54327 5 1 1 54326
0 54328 7 1 2 87054 54327
0 54329 7 1 2 54325 54328
0 54330 7 1 2 54321 54329
0 54331 5 1 1 54330
0 54332 7 1 2 84071 54331
0 54333 5 1 1 54332
0 54334 7 1 2 54319 54333
0 54335 5 1 1 54334
0 54336 7 1 2 58687 54335
0 54337 5 1 1 54336
0 54338 7 1 2 73926 73820
0 54339 7 1 2 77075 54338
0 54340 5 1 1 54339
0 54341 7 1 2 85563 54340
0 54342 5 1 1 54341
0 54343 7 1 2 59037 54342
0 54344 5 1 1 54343
0 54345 7 1 2 84893 93667
0 54346 5 1 1 54345
0 54347 7 1 2 54344 54346
0 54348 5 1 1 54347
0 54349 7 1 2 57815 54348
0 54350 5 1 1 54349
0 54351 7 1 2 77076 92904
0 54352 5 1 1 54351
0 54353 7 1 2 59177 88223
0 54354 5 1 1 54353
0 54355 7 1 2 54352 54354
0 54356 5 1 1 54355
0 54357 7 1 2 68058 54356
0 54358 5 1 1 54357
0 54359 7 1 2 54350 54358
0 54360 5 1 1 54359
0 54361 7 1 2 57532 54360
0 54362 5 1 1 54361
0 54363 7 1 2 83977 80060
0 54364 5 1 1 54363
0 54365 7 1 2 54362 54364
0 54366 5 1 1 54365
0 54367 7 1 2 84702 54366
0 54368 5 1 1 54367
0 54369 7 1 2 83125 89700
0 54370 7 1 2 82522 54369
0 54371 5 1 1 54370
0 54372 7 1 2 54368 54371
0 54373 7 1 2 54337 54372
0 54374 5 1 1 54373
0 54375 7 1 2 75966 94292
0 54376 7 1 2 54374 54375
0 54377 5 1 1 54376
0 54378 7 1 2 54246 54377
0 54379 7 1 2 54111 54378
0 54380 5 1 1 54379
0 54381 7 1 2 69283 54380
0 54382 5 1 1 54381
0 54383 7 2 2 94741 94886
0 54384 7 1 2 68059 76520
0 54385 5 1 1 54384
0 54386 7 1 2 95979 54385
0 54387 5 1 1 54386
0 54388 7 1 2 79196 94976
0 54389 5 1 1 54388
0 54390 7 1 2 61116 86754
0 54391 5 1 1 54390
0 54392 7 1 2 33903 54391
0 54393 5 1 1 54392
0 54394 7 1 2 62816 54393
0 54395 5 1 1 54394
0 54396 7 1 2 64116 93094
0 54397 5 1 1 54396
0 54398 7 1 2 54395 54397
0 54399 5 1 1 54398
0 54400 7 1 2 90237 54399
0 54401 5 1 1 54400
0 54402 7 1 2 66393 33905
0 54403 5 1 1 54402
0 54404 7 1 2 80877 54403
0 54405 5 1 1 54404
0 54406 7 1 2 44117 54405
0 54407 5 1 1 54406
0 54408 7 1 2 95787 54407
0 54409 5 1 1 54408
0 54410 7 1 2 54401 54409
0 54411 5 1 1 54410
0 54412 7 1 2 60688 54411
0 54413 5 1 1 54412
0 54414 7 1 2 78013 76892
0 54415 5 1 1 54414
0 54416 7 1 2 61749 85837
0 54417 7 1 2 54415 54416
0 54418 5 1 1 54417
0 54419 7 1 2 54413 54418
0 54420 5 1 1 54419
0 54421 7 1 2 75564 54420
0 54422 5 1 1 54421
0 54423 7 1 2 54389 54422
0 54424 5 1 1 54423
0 54425 7 1 2 79945 94219
0 54426 7 1 2 54424 54425
0 54427 5 1 1 54426
0 54428 7 1 2 54387 54427
0 54429 5 1 1 54428
0 54430 7 1 2 67944 54429
0 54431 5 1 1 54430
0 54432 7 2 2 76113 79270
0 54433 7 2 2 73423 95981
0 54434 7 1 2 90605 95983
0 54435 5 1 1 54434
0 54436 7 1 2 64117 95603
0 54437 7 1 2 87842 54436
0 54438 5 1 1 54437
0 54439 7 1 2 54435 54438
0 54440 5 1 1 54439
0 54441 7 1 2 62817 54440
0 54442 5 1 1 54441
0 54443 7 1 2 14703 91195
0 54444 5 1 1 54443
0 54445 7 1 2 59693 54444
0 54446 5 1 1 54445
0 54447 7 1 2 74116 54446
0 54448 5 1 1 54447
0 54449 7 1 2 76114 95884
0 54450 7 1 2 54448 54449
0 54451 5 1 1 54450
0 54452 7 1 2 54442 54451
0 54453 5 1 1 54452
0 54454 7 1 2 66732 54453
0 54455 5 1 1 54454
0 54456 7 1 2 82431 93381
0 54457 7 2 2 83430 54456
0 54458 5 2 1 95985
0 54459 7 1 2 60689 95986
0 54460 5 1 1 54459
0 54461 7 1 2 54455 54460
0 54462 5 1 1 54461
0 54463 7 1 2 75193 54462
0 54464 5 1 1 54463
0 54465 7 2 2 86953 95984
0 54466 5 2 1 95989
0 54467 7 1 2 66733 81082
0 54468 7 1 2 51920 54467
0 54469 7 1 2 95990 54468
0 54470 5 1 1 54469
0 54471 7 1 2 62001 54470
0 54472 7 1 2 54464 54471
0 54473 7 1 2 54431 54472
0 54474 5 1 1 54473
0 54475 7 1 2 90354 93785
0 54476 5 1 1 54475
0 54477 7 1 2 80881 43107
0 54478 5 1 1 54477
0 54479 7 1 2 72879 95881
0 54480 7 1 2 54478 54479
0 54481 5 1 1 54480
0 54482 7 1 2 54476 54481
0 54483 5 1 1 54482
0 54484 7 1 2 69082 54483
0 54485 5 1 1 54484
0 54486 7 1 2 72787 91441
0 54487 5 1 1 54486
0 54488 7 1 2 63424 54487
0 54489 5 1 1 54488
0 54490 7 1 2 85648 5740
0 54491 5 1 1 54490
0 54492 7 1 2 54489 54491
0 54493 5 1 1 54492
0 54494 7 1 2 62818 54493
0 54495 5 1 1 54494
0 54496 7 1 2 72808 12144
0 54497 5 1 1 54496
0 54498 7 1 2 61485 85188
0 54499 7 1 2 54497 54498
0 54500 5 1 1 54499
0 54501 7 1 2 54495 54500
0 54502 5 1 1 54501
0 54503 7 1 2 88276 54502
0 54504 5 1 1 54503
0 54505 7 1 2 87762 95060
0 54506 5 1 1 54505
0 54507 7 1 2 54504 54506
0 54508 5 1 1 54507
0 54509 7 1 2 60690 54508
0 54510 5 1 1 54509
0 54511 7 1 2 54485 54510
0 54512 5 1 1 54511
0 54513 7 1 2 84019 54512
0 54514 5 1 1 54513
0 54515 7 1 2 38084 53018
0 54516 5 1 1 54515
0 54517 7 1 2 63559 54516
0 54518 5 1 1 54517
0 54519 7 1 2 67232 93944
0 54520 5 1 1 54519
0 54521 7 1 2 85592 94557
0 54522 5 1 1 54521
0 54523 7 1 2 54520 54522
0 54524 5 1 1 54523
0 54525 7 1 2 63115 93274
0 54526 7 1 2 54524 54525
0 54527 5 1 1 54526
0 54528 7 1 2 54518 54527
0 54529 5 1 1 54528
0 54530 7 1 2 66394 54529
0 54531 5 1 1 54530
0 54532 7 1 2 85386 88639
0 54533 7 1 2 82853 54532
0 54534 5 1 1 54533
0 54535 7 1 2 54531 54534
0 54536 5 1 1 54535
0 54537 7 1 2 63789 54536
0 54538 5 1 1 54537
0 54539 7 1 2 60691 85366
0 54540 5 1 1 54539
0 54541 7 1 2 59694 54540
0 54542 5 1 1 54541
0 54543 7 1 2 90325 54542
0 54544 5 1 1 54543
0 54545 7 1 2 84720 31908
0 54546 7 1 2 87380 54545
0 54547 5 1 1 54546
0 54548 7 1 2 54544 54547
0 54549 5 1 1 54548
0 54550 7 1 2 61750 54549
0 54551 5 1 1 54550
0 54552 7 1 2 84889 90886
0 54553 5 1 1 54552
0 54554 7 1 2 54551 54553
0 54555 5 1 1 54554
0 54556 7 1 2 87139 54555
0 54557 5 1 1 54556
0 54558 7 1 2 74916 94241
0 54559 5 1 1 54558
0 54560 7 1 2 74018 80878
0 54561 7 1 2 95247 54560
0 54562 5 1 1 54561
0 54563 7 1 2 54559 54562
0 54564 5 1 1 54563
0 54565 7 1 2 66094 54564
0 54566 5 1 1 54565
0 54567 7 1 2 54557 54566
0 54568 7 1 2 54538 54567
0 54569 5 1 1 54568
0 54570 7 1 2 62280 54569
0 54571 5 1 1 54570
0 54572 7 1 2 86048 95052
0 54573 5 1 1 54572
0 54574 7 1 2 83338 94642
0 54575 5 1 1 54574
0 54576 7 1 2 32904 54575
0 54577 5 1 1 54576
0 54578 7 3 2 60078 84790
0 54579 7 1 2 80764 95993
0 54580 7 1 2 54577 54579
0 54581 5 1 1 54580
0 54582 7 1 2 54573 54581
0 54583 5 1 1 54582
0 54584 7 1 2 59948 54583
0 54585 5 1 1 54584
0 54586 7 1 2 54571 54585
0 54587 7 1 2 54514 54586
0 54588 5 1 1 54587
0 54589 7 1 2 61117 54588
0 54590 5 1 1 54589
0 54591 7 1 2 69748 87507
0 54592 5 1 1 54591
0 54593 7 1 2 94639 54592
0 54594 5 3 1 54593
0 54595 7 1 2 80822 95996
0 54596 5 1 1 54595
0 54597 7 1 2 73390 86046
0 54598 5 1 1 54597
0 54599 7 1 2 54596 54598
0 54600 5 1 1 54599
0 54601 7 1 2 87542 84087
0 54602 7 1 2 54600 54601
0 54603 5 1 1 54602
0 54604 7 1 2 63116 95864
0 54605 5 1 1 54604
0 54606 7 1 2 40724 54605
0 54607 5 1 1 54606
0 54608 7 1 2 78769 93976
0 54609 7 1 2 54607 54608
0 54610 5 1 1 54609
0 54611 7 1 2 54603 54610
0 54612 5 1 1 54611
0 54613 7 1 2 68183 54612
0 54614 5 1 1 54613
0 54615 7 1 2 73555 93786
0 54616 5 1 1 54615
0 54617 7 1 2 72880 87918
0 54618 7 1 2 80846 54617
0 54619 5 1 1 54618
0 54620 7 1 2 54616 54619
0 54621 5 1 1 54620
0 54622 7 1 2 60079 84317
0 54623 7 1 2 80936 54622
0 54624 7 1 2 54621 54623
0 54625 5 1 1 54624
0 54626 7 1 2 54614 54625
0 54627 7 1 2 54590 54626
0 54628 5 1 1 54627
0 54629 7 1 2 69684 54628
0 54630 5 1 1 54629
0 54631 7 1 2 74385 90994
0 54632 5 1 1 54631
0 54633 7 1 2 93663 54632
0 54634 5 1 1 54633
0 54635 7 1 2 66095 54634
0 54636 5 1 1 54635
0 54637 7 1 2 16696 54636
0 54638 5 1 1 54637
0 54639 7 1 2 95947 54638
0 54640 5 1 1 54639
0 54641 7 1 2 64423 78885
0 54642 5 1 1 54641
0 54643 7 1 2 29162 54642
0 54644 5 1 1 54643
0 54645 7 1 2 60692 54644
0 54646 5 1 1 54645
0 54647 7 1 2 61486 80937
0 54648 5 1 1 54647
0 54649 7 1 2 54646 54648
0 54650 5 1 1 54649
0 54651 7 1 2 63117 54650
0 54652 5 1 1 54651
0 54653 7 1 2 79089 72881
0 54654 5 1 1 54653
0 54655 7 1 2 54652 54654
0 54656 5 1 1 54655
0 54657 7 1 2 61118 54656
0 54658 5 1 1 54657
0 54659 7 1 2 85655 54658
0 54660 5 1 1 54659
0 54661 7 1 2 89324 54660
0 54662 5 1 1 54661
0 54663 7 1 2 54640 54662
0 54664 5 1 1 54663
0 54665 7 1 2 68184 54664
0 54666 5 1 1 54665
0 54667 7 2 2 91542 92028
0 54668 5 1 1 95999
0 54669 7 1 2 61487 96000
0 54670 5 1 1 54669
0 54671 7 1 2 77595 87631
0 54672 7 1 2 95860 54671
0 54673 5 1 1 54672
0 54674 7 1 2 54670 54673
0 54675 5 1 1 54674
0 54676 7 1 2 69083 54675
0 54677 5 1 1 54676
0 54678 7 1 2 85552 79499
0 54679 7 1 2 75081 54678
0 54680 7 1 2 95230 54679
0 54681 5 1 1 54680
0 54682 7 1 2 54677 54681
0 54683 5 1 1 54682
0 54684 7 1 2 62281 54683
0 54685 5 1 1 54684
0 54686 7 1 2 85860 95791
0 54687 7 1 2 91815 54686
0 54688 5 1 1 54687
0 54689 7 1 2 90255 34017
0 54690 5 1 1 54689
0 54691 7 1 2 95480 54690
0 54692 5 1 1 54691
0 54693 7 1 2 75194 95994
0 54694 7 1 2 95808 54693
0 54695 5 1 1 54694
0 54696 7 1 2 54692 54695
0 54697 7 1 2 54688 54696
0 54698 7 1 2 54685 54697
0 54699 5 1 1 54698
0 54700 7 1 2 60693 54699
0 54701 5 1 1 54700
0 54702 7 1 2 78000 93870
0 54703 7 1 2 95810 54702
0 54704 5 1 1 54703
0 54705 7 1 2 5963 44171
0 54706 5 1 1 54705
0 54707 7 1 2 81409 87886
0 54708 7 1 2 54706 54707
0 54709 5 1 1 54708
0 54710 7 1 2 54704 54709
0 54711 7 1 2 54701 54710
0 54712 7 1 2 54666 54711
0 54713 5 1 1 54712
0 54714 7 1 2 69284 54713
0 54715 5 1 1 54714
0 54716 7 1 2 66647 54715
0 54717 7 1 2 54630 54716
0 54718 5 1 1 54717
0 54719 7 1 2 67802 54718
0 54720 7 1 2 54474 54719
0 54721 5 1 1 54720
0 54722 7 1 2 13631 33956
0 54723 5 1 1 54722
0 54724 7 1 2 58688 54723
0 54725 5 1 1 54724
0 54726 7 1 2 65101 87796
0 54727 5 1 1 54726
0 54728 7 1 2 75155 54727
0 54729 5 1 1 54728
0 54730 7 1 2 85873 54729
0 54731 5 1 1 54730
0 54732 7 1 2 54725 54731
0 54733 5 1 1 54732
0 54734 7 1 2 95948 54733
0 54735 5 1 1 54734
0 54736 7 1 2 89325 95761
0 54737 5 1 1 54736
0 54738 7 1 2 54735 54737
0 54739 5 1 1 54738
0 54740 7 1 2 69285 54739
0 54741 5 1 1 54740
0 54742 7 1 2 68281 95089
0 54743 5 1 1 54742
0 54744 7 1 2 65747 91451
0 54745 5 1 1 54744
0 54746 7 1 2 54743 54745
0 54747 5 1 1 54746
0 54748 7 1 2 60080 54747
0 54749 5 1 1 54748
0 54750 7 1 2 87488 82624
0 54751 5 1 1 54750
0 54752 7 1 2 54749 54751
0 54753 5 1 1 54752
0 54754 7 1 2 64424 54753
0 54755 5 1 1 54754
0 54756 7 1 2 93777 95248
0 54757 5 1 1 54756
0 54758 7 1 2 44928 54757
0 54759 5 1 1 54758
0 54760 7 1 2 58818 54759
0 54761 5 1 1 54760
0 54762 7 1 2 54755 54761
0 54763 5 1 1 54762
0 54764 7 1 2 63425 54763
0 54765 5 1 1 54764
0 54766 7 1 2 58819 90375
0 54767 7 1 2 94962 54766
0 54768 5 1 1 54767
0 54769 7 1 2 54765 54768
0 54770 5 1 1 54769
0 54771 7 1 2 63118 54770
0 54772 5 1 1 54771
0 54773 7 1 2 87161 95634
0 54774 5 3 1 54773
0 54775 7 1 2 86129 82536
0 54776 7 1 2 92442 54775
0 54777 5 1 1 54776
0 54778 7 1 2 96001 54777
0 54779 7 1 2 54772 54778
0 54780 5 1 1 54779
0 54781 7 1 2 76938 54780
0 54782 5 1 1 54781
0 54783 7 1 2 54741 54782
0 54784 5 1 1 54783
0 54785 7 1 2 68889 54784
0 54786 5 1 1 54785
0 54787 7 1 2 80068 83493
0 54788 5 1 1 54787
0 54789 7 3 2 61488 95607
0 54790 5 1 1 96004
0 54791 7 1 2 54788 96005
0 54792 5 1 1 54791
0 54793 7 1 2 84045 93679
0 54794 5 1 1 54793
0 54795 7 1 2 75458 54794
0 54796 5 1 1 54795
0 54797 7 1 2 69286 54796
0 54798 5 1 1 54797
0 54799 7 1 2 7875 54798
0 54800 5 1 1 54799
0 54801 7 1 2 61119 54800
0 54802 5 1 1 54801
0 54803 7 2 2 75450 69287
0 54804 7 1 2 60421 96007
0 54805 5 1 1 54804
0 54806 7 1 2 70675 68686
0 54807 5 1 1 54806
0 54808 7 1 2 54805 54807
0 54809 5 1 1 54808
0 54810 7 1 2 68538 54809
0 54811 5 1 1 54810
0 54812 7 1 2 84385 96008
0 54813 5 1 1 54812
0 54814 7 1 2 68282 72120
0 54815 5 1 1 54814
0 54816 7 1 2 54813 54815
0 54817 7 1 2 54811 54816
0 54818 7 1 2 54802 54817
0 54819 5 1 1 54818
0 54820 7 1 2 66096 54819
0 54821 5 1 1 54820
0 54822 7 1 2 54792 54821
0 54823 5 1 1 54822
0 54824 7 1 2 95949 54823
0 54825 5 1 1 54824
0 54826 7 1 2 85594 90378
0 54827 5 1 1 54826
0 54828 7 1 2 68539 54827
0 54829 5 1 1 54828
0 54830 7 1 2 59695 83936
0 54831 5 1 1 54830
0 54832 7 1 2 61489 54831
0 54833 5 1 1 54832
0 54834 7 1 2 54829 54833
0 54835 5 1 1 54834
0 54836 7 1 2 89326 54835
0 54837 5 1 1 54836
0 54838 7 4 2 83003 94972
0 54839 7 1 2 69432 96009
0 54840 5 1 1 54839
0 54841 7 1 2 54837 54840
0 54842 5 1 1 54841
0 54843 7 1 2 69288 54842
0 54844 5 1 1 54843
0 54845 7 1 2 81820 35076
0 54846 5 1 1 54845
0 54847 7 1 2 92274 54846
0 54848 5 1 1 54847
0 54849 7 1 2 88622 94456
0 54850 5 1 1 54849
0 54851 7 1 2 72556 72882
0 54852 7 1 2 54850 54851
0 54853 5 1 1 54852
0 54854 7 1 2 54848 54853
0 54855 5 1 1 54854
0 54856 7 1 2 60081 68687
0 54857 7 1 2 84046 54856
0 54858 7 1 2 54855 54857
0 54859 5 1 1 54858
0 54860 7 1 2 54844 54859
0 54861 5 1 1 54860
0 54862 7 1 2 61120 54861
0 54863 5 1 1 54862
0 54864 7 1 2 64425 69583
0 54865 5 1 1 54864
0 54866 7 1 2 69227 54865
0 54867 5 1 1 54866
0 54868 7 1 2 94633 54867
0 54869 5 1 1 54868
0 54870 7 1 2 69488 90924
0 54871 5 1 1 54870
0 54872 7 1 2 54869 54871
0 54873 5 1 1 54872
0 54874 7 1 2 93977 54873
0 54875 5 1 1 54874
0 54876 7 1 2 80648 90717
0 54877 7 1 2 82625 88081
0 54878 7 1 2 54876 54877
0 54879 5 1 1 54878
0 54880 7 1 2 54875 54879
0 54881 5 1 1 54880
0 54882 7 1 2 72557 54881
0 54883 5 1 1 54882
0 54884 7 1 2 87635 87545
0 54885 5 1 1 54884
0 54886 7 1 2 94634 54885
0 54887 5 1 1 54886
0 54888 7 1 2 87649 73338
0 54889 5 1 1 54888
0 54890 7 1 2 54887 54889
0 54891 5 1 1 54890
0 54892 7 1 2 80962 54891
0 54893 5 1 1 54892
0 54894 7 1 2 63426 81818
0 54895 7 1 2 91378 54894
0 54896 7 1 2 95769 54895
0 54897 5 1 1 54896
0 54898 7 1 2 49238 54897
0 54899 5 1 1 54898
0 54900 7 1 2 69289 54899
0 54901 5 1 1 54900
0 54902 7 1 2 54893 54901
0 54903 5 1 1 54902
0 54904 7 1 2 68283 54903
0 54905 5 1 1 54904
0 54906 7 2 2 62141 90309
0 54907 7 1 2 64759 80959
0 54908 7 1 2 76900 54907
0 54909 7 1 2 96013 54908
0 54910 7 1 2 95997 54909
0 54911 5 1 1 54910
0 54912 7 1 2 54905 54911
0 54913 7 1 2 54883 54912
0 54914 7 1 2 54863 54913
0 54915 5 1 1 54914
0 54916 7 1 2 63119 54915
0 54917 5 1 1 54916
0 54918 7 1 2 3295 76940
0 54919 5 1 1 54918
0 54920 7 1 2 60422 54919
0 54921 5 1 1 54920
0 54922 7 1 2 72564 90284
0 54923 5 1 1 54922
0 54924 7 1 2 68696 54923
0 54925 5 1 1 54924
0 54926 7 1 2 78419 54925
0 54927 5 1 1 54926
0 54928 7 1 2 54921 54927
0 54929 5 1 1 54928
0 54930 7 1 2 64426 54929
0 54931 5 1 1 54930
0 54932 7 1 2 59696 12969
0 54933 5 1 1 54932
0 54934 7 1 2 83537 54933
0 54935 5 1 1 54934
0 54936 7 1 2 84198 69290
0 54937 7 1 2 85000 54936
0 54938 5 1 1 54937
0 54939 7 1 2 54935 54938
0 54940 7 1 2 54931 54939
0 54941 5 1 1 54940
0 54942 7 1 2 94635 54941
0 54943 5 1 1 54942
0 54944 7 1 2 58903 93645
0 54945 7 1 2 87802 54944
0 54946 7 2 2 60169 90550
0 54947 7 1 2 92522 96015
0 54948 7 1 2 54945 54947
0 54949 5 1 1 54948
0 54950 7 1 2 54943 54949
0 54951 5 1 1 54950
0 54952 7 1 2 93978 54951
0 54953 5 1 1 54952
0 54954 7 1 2 66648 54953
0 54955 7 1 2 54917 54954
0 54956 7 1 2 54825 54955
0 54957 7 1 2 54786 54956
0 54958 5 1 1 54957
0 54959 7 1 2 79962 95939
0 54960 7 1 2 92937 54959
0 54961 5 1 1 54960
0 54962 7 1 2 95991 54961
0 54963 5 1 1 54962
0 54964 7 1 2 68284 54963
0 54965 5 1 1 54964
0 54966 7 1 2 64643 85985
0 54967 7 1 2 79925 89572
0 54968 7 1 2 54966 54967
0 54969 7 1 2 74917 54968
0 54970 5 1 1 54969
0 54971 7 1 2 95992 54970
0 54972 5 1 1 54971
0 54973 7 1 2 61121 54972
0 54974 5 1 1 54973
0 54975 7 1 2 54965 54974
0 54976 5 1 1 54975
0 54977 7 1 2 66734 54976
0 54978 5 1 1 54977
0 54979 7 1 2 54978 95987
0 54980 5 1 1 54979
0 54981 7 1 2 68890 54980
0 54982 5 1 1 54981
0 54983 7 1 2 82009 95980
0 54984 5 1 1 54983
0 54985 7 1 2 85974 95757
0 54986 5 1 1 54985
0 54987 7 1 2 14744 54986
0 54988 5 1 1 54987
0 54989 7 1 2 72558 54988
0 54990 5 1 1 54989
0 54991 7 1 2 86271 54990
0 54992 5 1 1 54991
0 54993 7 1 2 74309 92275
0 54994 7 1 2 54992 54993
0 54995 5 1 1 54994
0 54996 7 1 2 54984 54995
0 54997 5 1 1 54996
0 54998 7 1 2 67945 54997
0 54999 5 1 1 54998
0 55000 7 1 2 90143 95982
0 55001 7 1 2 95775 55000
0 55002 5 1 1 55001
0 55003 7 1 2 62002 55002
0 55004 7 1 2 54999 55003
0 55005 7 1 2 54982 55004
0 55006 5 1 1 55005
0 55007 7 1 2 68185 55006
0 55008 7 1 2 54958 55007
0 55009 5 1 1 55008
0 55010 7 1 2 73020 93838
0 55011 5 1 1 55010
0 55012 7 1 2 58820 95862
0 55013 5 1 1 55012
0 55014 7 1 2 55011 55013
0 55015 5 1 1 55014
0 55016 7 1 2 62282 55015
0 55017 5 1 1 55016
0 55018 7 1 2 80077 95683
0 55019 5 1 1 55018
0 55020 7 1 2 55017 55019
0 55021 5 1 1 55020
0 55022 7 1 2 87274 55021
0 55023 5 1 1 55022
0 55024 7 1 2 82509 92401
0 55025 5 1 1 55024
0 55026 7 1 2 55023 55025
0 55027 5 1 1 55026
0 55028 7 1 2 60082 55027
0 55029 5 1 1 55028
0 55030 7 1 2 68540 79832
0 55031 7 1 2 77566 55030
0 55032 7 1 2 90606 55031
0 55033 5 1 1 55032
0 55034 7 1 2 55029 55033
0 55035 5 1 1 55034
0 55036 7 1 2 67803 55035
0 55037 5 1 1 55036
0 55038 7 1 2 85903 92708
0 55039 7 1 2 95865 55038
0 55040 5 1 1 55039
0 55041 7 1 2 61122 78420
0 55042 7 1 2 95684 55041
0 55043 5 1 1 55042
0 55044 7 1 2 47155 55043
0 55045 7 1 2 55040 55044
0 55046 5 1 1 55045
0 55047 7 1 2 95249 55046
0 55048 5 1 1 55047
0 55049 7 1 2 87070 95291
0 55050 7 1 2 95998 55049
0 55051 5 1 1 55050
0 55052 7 1 2 55048 55051
0 55053 7 1 2 55037 55052
0 55054 5 1 1 55053
0 55055 7 1 2 80963 55054
0 55056 5 1 1 55055
0 55057 7 1 2 63790 95527
0 55058 5 1 1 55057
0 55059 7 1 2 96002 55058
0 55060 5 1 1 55059
0 55061 7 1 2 62283 55060
0 55062 5 1 1 55061
0 55063 7 2 2 84020 84791
0 55064 7 1 2 72801 92569
0 55065 7 1 2 96017 55064
0 55066 5 1 1 55065
0 55067 7 1 2 70676 96010
0 55068 5 1 1 55067
0 55069 7 1 2 55066 55068
0 55070 7 1 2 55062 55069
0 55071 5 1 1 55070
0 55072 7 1 2 68285 55071
0 55073 5 1 1 55072
0 55074 7 1 2 72156 96011
0 55075 5 1 1 55074
0 55076 7 1 2 87140 84318
0 55077 7 1 2 92212 55076
0 55078 5 1 1 55077
0 55079 7 1 2 55075 55078
0 55080 5 1 1 55079
0 55081 7 1 2 76967 55080
0 55082 5 1 1 55081
0 55083 7 1 2 91665 92213
0 55084 5 1 1 55083
0 55085 7 1 2 67804 66796
0 55086 7 1 2 72342 55085
0 55087 7 1 2 87489 95798
0 55088 7 1 2 55086 55087
0 55089 5 1 1 55088
0 55090 7 1 2 55084 55089
0 55091 7 1 2 55082 55090
0 55092 7 1 2 55073 55091
0 55093 5 1 1 55092
0 55094 7 1 2 60423 55093
0 55095 5 1 1 55094
0 55096 7 1 2 93691 96012
0 55097 5 1 1 55096
0 55098 7 2 2 87187 90326
0 55099 7 1 2 87141 37353
0 55100 7 1 2 96019 55099
0 55101 5 1 1 55100
0 55102 7 1 2 55097 55101
0 55103 5 1 1 55102
0 55104 7 1 2 68891 55103
0 55105 5 1 1 55104
0 55106 7 1 2 82137 89755
0 55107 5 1 1 55106
0 55108 7 1 2 96003 55107
0 55109 5 1 1 55108
0 55110 7 1 2 70854 55109
0 55111 5 1 1 55110
0 55112 7 1 2 84460 79463
0 55113 7 1 2 96018 55112
0 55114 5 1 1 55113
0 55115 7 1 2 86954 81051
0 55116 7 1 2 74852 55115
0 55117 5 1 1 55116
0 55118 7 1 2 55114 55117
0 55119 7 1 2 55111 55118
0 55120 5 1 1 55119
0 55121 7 1 2 61123 55120
0 55122 5 1 1 55121
0 55123 7 1 2 82647 94969
0 55124 5 1 1 55123
0 55125 7 1 2 64644 71112
0 55126 7 1 2 95792 95995
0 55127 7 1 2 55125 55126
0 55128 5 1 1 55127
0 55129 7 1 2 55124 55128
0 55130 5 1 1 55129
0 55131 7 1 2 83840 55130
0 55132 5 1 1 55131
0 55133 7 1 2 67570 77297
0 55134 7 1 2 96020 55133
0 55135 5 1 1 55134
0 55136 7 1 2 54668 55135
0 55137 5 1 1 55136
0 55138 7 1 2 61490 55137
0 55139 5 1 1 55138
0 55140 7 1 2 55132 55139
0 55141 7 1 2 55122 55140
0 55142 7 1 2 55105 55141
0 55143 7 1 2 55095 55142
0 55144 5 1 1 55143
0 55145 7 1 2 69291 55144
0 55146 5 1 1 55145
0 55147 7 1 2 66649 55146
0 55148 7 1 2 55056 55147
0 55149 5 1 1 55148
0 55150 7 1 2 78532 81456
0 55151 5 1 1 55150
0 55152 7 1 2 65748 94130
0 55153 5 1 1 55152
0 55154 7 1 2 55151 55153
0 55155 5 1 1 55154
0 55156 7 2 2 76115 89479
0 55157 7 1 2 82693 96021
0 55158 7 1 2 55155 55157
0 55159 5 1 1 55158
0 55160 7 1 2 92743 95785
0 55161 5 1 1 55160
0 55162 7 1 2 83669 91680
0 55163 5 1 1 55162
0 55164 7 1 2 55161 55163
0 55165 5 1 1 55164
0 55166 7 1 2 69489 55165
0 55167 5 1 1 55166
0 55168 7 1 2 87154 82356
0 55169 7 1 2 89756 55168
0 55170 5 1 1 55169
0 55171 7 1 2 55167 55170
0 55172 7 1 2 55159 55171
0 55173 5 1 1 55172
0 55174 7 1 2 66735 55173
0 55175 5 1 1 55174
0 55176 7 1 2 62003 95988
0 55177 7 1 2 55175 55176
0 55178 5 1 1 55177
0 55179 7 1 2 76233 55178
0 55180 7 1 2 55149 55179
0 55181 5 1 1 55180
0 55182 7 1 2 55009 55181
0 55183 7 1 2 54721 55182
0 55184 7 1 2 54382 55183
0 55185 7 1 2 53944 55184
0 55186 7 1 2 73858 69853
0 55187 5 1 1 55186
0 55188 7 1 2 67400 95403
0 55189 5 1 1 55188
0 55190 7 1 2 55187 55189
0 55191 5 1 1 55190
0 55192 7 1 2 73271 55191
0 55193 5 1 1 55192
0 55194 7 1 2 61491 69882
0 55195 7 1 2 93018 55194
0 55196 5 1 1 55195
0 55197 7 1 2 55193 55196
0 55198 5 1 1 55197
0 55199 7 1 2 71564 55198
0 55200 5 1 1 55199
0 55201 7 1 2 72360 92119
0 55202 5 1 1 55201
0 55203 7 1 2 57533 73409
0 55204 7 1 2 86217 55203
0 55205 5 1 1 55204
0 55206 7 1 2 55202 55205
0 55207 5 1 1 55206
0 55208 7 1 2 59178 55207
0 55209 5 1 1 55208
0 55210 7 1 2 55200 55209
0 55211 5 1 1 55210
0 55212 7 1 2 59038 55211
0 55213 5 1 1 55212
0 55214 7 1 2 70310 95618
0 55215 7 1 2 84293 55214
0 55216 5 1 1 55215
0 55217 7 1 2 55213 55216
0 55218 5 1 1 55217
0 55219 7 1 2 57816 55218
0 55220 5 1 1 55219
0 55221 7 1 2 86409 95359
0 55222 5 1 1 55221
0 55223 7 1 2 74679 55222
0 55224 5 1 1 55223
0 55225 7 1 2 73859 55224
0 55226 5 1 1 55225
0 55227 7 1 2 95839 55226
0 55228 5 1 1 55227
0 55229 7 1 2 67401 55228
0 55230 5 1 1 55229
0 55231 7 1 2 93514 55230
0 55232 7 1 2 55220 55231
0 55233 5 1 1 55232
0 55234 7 1 2 83030 55233
0 55235 5 1 1 55234
0 55236 7 1 2 74227 85713
0 55237 5 1 1 55236
0 55238 7 1 2 85863 55237
0 55239 5 1 1 55238
0 55240 7 1 2 84703 55239
0 55241 5 1 1 55240
0 55242 7 1 2 81418 90656
0 55243 5 1 1 55242
0 55244 7 1 2 55241 55243
0 55245 5 1 1 55244
0 55246 7 1 2 69685 55245
0 55247 5 1 1 55246
0 55248 7 1 2 73767 83100
0 55249 7 1 2 84598 55248
0 55250 7 1 2 80026 55249
0 55251 5 1 1 55250
0 55252 7 1 2 55247 55251
0 55253 5 1 1 55252
0 55254 7 1 2 71764 55253
0 55255 5 1 1 55254
0 55256 7 1 2 86163 74060
0 55257 5 1 1 55256
0 55258 7 1 2 76836 55257
0 55259 5 1 1 55258
0 55260 7 1 2 79248 84760
0 55261 7 1 2 88028 55260
0 55262 5 1 1 55261
0 55263 7 1 2 55259 55262
0 55264 5 1 1 55263
0 55265 7 1 2 58369 55264
0 55266 5 1 1 55265
0 55267 7 1 2 80607 82706
0 55268 7 1 2 76776 55267
0 55269 7 1 2 83538 55268
0 55270 5 1 1 55269
0 55271 7 1 2 55266 55270
0 55272 5 1 1 55271
0 55273 7 1 2 66395 55272
0 55274 5 1 1 55273
0 55275 7 1 2 72179 89518
0 55276 7 1 2 83102 55275
0 55277 5 1 1 55276
0 55278 7 1 2 55274 55277
0 55279 5 1 1 55278
0 55280 7 1 2 71927 55279
0 55281 5 1 1 55280
0 55282 7 1 2 95719 95974
0 55283 5 1 1 55282
0 55284 7 1 2 73602 73788
0 55285 5 1 1 55284
0 55286 7 1 2 66396 67402
0 55287 7 1 2 55285 55286
0 55288 5 1 1 55287
0 55289 7 1 2 55283 55288
0 55290 5 1 1 55289
0 55291 7 1 2 69686 55290
0 55292 5 1 1 55291
0 55293 7 1 2 79745 90718
0 55294 7 1 2 85758 95570
0 55295 7 1 2 55293 55294
0 55296 5 1 1 55295
0 55297 7 1 2 55292 55296
0 55298 5 1 1 55297
0 55299 7 1 2 58370 55298
0 55300 5 1 1 55299
0 55301 7 1 2 66097 81877
0 55302 7 1 2 77743 55301
0 55303 7 1 2 76837 55302
0 55304 5 1 1 55303
0 55305 7 1 2 55300 55304
0 55306 5 1 1 55305
0 55307 7 1 2 78331 55306
0 55308 5 1 1 55307
0 55309 7 1 2 55281 55308
0 55310 7 1 2 55255 55309
0 55311 7 1 2 55235 55310
0 55312 5 1 1 55311
0 55313 7 1 2 58689 55312
0 55314 5 1 1 55313
0 55315 7 1 2 83027 71135
0 55316 7 1 2 95837 55315
0 55317 7 1 2 72840 55316
0 55318 5 1 1 55317
0 55319 7 1 2 55314 55318
0 55320 5 1 1 55319
0 55321 7 1 2 66804 55320
0 55322 5 1 1 55321
0 55323 7 1 2 85307 81638
0 55324 5 1 1 55323
0 55325 7 1 2 70880 95317
0 55326 5 1 1 55325
0 55327 7 1 2 38342 55326
0 55328 5 1 1 55327
0 55329 7 1 2 67403 55328
0 55330 5 1 1 55329
0 55331 7 1 2 87408 55330
0 55332 7 1 2 55324 55331
0 55333 5 1 1 55332
0 55334 7 1 2 61751 55333
0 55335 5 1 1 55334
0 55336 7 1 2 58371 82886
0 55337 5 1 1 55336
0 55338 7 1 2 55335 55337
0 55339 5 1 1 55338
0 55340 7 1 2 72919 55339
0 55341 5 1 1 55340
0 55342 7 1 2 74744 94278
0 55343 5 1 1 55342
0 55344 7 1 2 92775 95835
0 55345 5 1 1 55344
0 55346 7 1 2 55343 55345
0 55347 5 1 1 55346
0 55348 7 1 2 71928 55347
0 55349 5 1 1 55348
0 55350 7 1 2 74745 73912
0 55351 5 1 1 55350
0 55352 7 1 2 80402 83351
0 55353 5 1 1 55352
0 55354 7 1 2 55351 55353
0 55355 5 1 1 55354
0 55356 7 1 2 78332 55355
0 55357 5 1 1 55356
0 55358 7 1 2 68060 74701
0 55359 5 1 1 55358
0 55360 7 1 2 68286 84627
0 55361 5 1 1 55360
0 55362 7 1 2 14867 55361
0 55363 5 1 1 55362
0 55364 7 1 2 59697 55363
0 55365 5 1 1 55364
0 55366 7 1 2 55359 55365
0 55367 7 1 2 55357 55366
0 55368 7 1 2 55349 55367
0 55369 5 1 1 55368
0 55370 7 1 2 81410 55369
0 55371 5 1 1 55370
0 55372 7 2 2 61752 85539
0 55373 5 1 1 96023
0 55374 7 1 2 94927 55373
0 55375 5 1 1 55374
0 55376 7 1 2 70437 55375
0 55377 5 1 1 55376
0 55378 7 1 2 74182 84401
0 55379 5 1 1 55378
0 55380 7 1 2 55377 55379
0 55381 5 1 1 55380
0 55382 7 1 2 75886 55381
0 55383 5 1 1 55382
0 55384 7 1 2 92080 94928
0 55385 5 1 1 55384
0 55386 7 1 2 59698 55385
0 55387 5 1 1 55386
0 55388 7 1 2 57534 81411
0 55389 7 1 2 74702 55388
0 55390 5 1 1 55389
0 55391 7 1 2 93561 55390
0 55392 7 1 2 55387 55391
0 55393 5 1 1 55392
0 55394 7 1 2 67404 55393
0 55395 5 1 1 55394
0 55396 7 1 2 55383 55395
0 55397 5 1 1 55396
0 55398 7 1 2 71765 55397
0 55399 5 1 1 55398
0 55400 7 1 2 57535 86385
0 55401 5 1 1 55400
0 55402 7 1 2 1211 55401
0 55403 5 1 1 55402
0 55404 7 1 2 72253 55403
0 55405 5 1 1 55404
0 55406 7 1 2 59699 85553
0 55407 5 1 1 55406
0 55408 7 1 2 86930 55407
0 55409 7 1 2 55405 55408
0 55410 7 1 2 69200 78225
0 55411 5 1 1 55410
0 55412 7 1 2 72212 55411
0 55413 5 1 1 55412
0 55414 7 1 2 70438 78338
0 55415 5 1 1 55414
0 55416 7 1 2 76234 55415
0 55417 5 1 1 55416
0 55418 7 1 2 71929 55417
0 55419 5 1 1 55418
0 55420 7 1 2 55413 55419
0 55421 7 1 2 55409 55420
0 55422 5 1 1 55421
0 55423 7 1 2 96024 55422
0 55424 5 1 1 55423
0 55425 7 1 2 55399 55424
0 55426 7 1 2 55371 55425
0 55427 7 1 2 55341 55426
0 55428 5 1 1 55427
0 55429 7 1 2 69292 55428
0 55430 5 1 1 55429
0 55431 7 2 2 67405 81300
0 55432 5 1 1 96025
0 55433 7 1 2 71565 96026
0 55434 5 1 1 55433
0 55435 7 1 2 80906 55434
0 55436 5 1 1 55435
0 55437 7 1 2 78276 55436
0 55438 5 1 1 55437
0 55439 7 1 2 61753 84844
0 55440 7 1 2 55438 55439
0 55441 5 1 1 55440
0 55442 7 1 2 60424 84963
0 55443 5 1 1 55442
0 55444 7 1 2 68287 76550
0 55445 5 1 1 55444
0 55446 7 1 2 66397 72660
0 55447 7 1 2 91154 55446
0 55448 7 1 2 55445 55447
0 55449 7 1 2 55443 55448
0 55450 5 1 1 55449
0 55451 7 1 2 66098 55450
0 55452 7 1 2 55441 55451
0 55453 5 1 1 55452
0 55454 7 1 2 95470 95662
0 55455 5 1 1 55454
0 55456 7 1 2 75340 55455
0 55457 5 1 1 55456
0 55458 7 1 2 67702 94798
0 55459 5 1 1 55458
0 55460 7 1 2 55457 55459
0 55461 5 1 1 55460
0 55462 7 1 2 65355 55461
0 55463 5 1 1 55462
0 55464 7 1 2 67406 95469
0 55465 5 1 1 55464
0 55466 7 1 2 95697 55465
0 55467 5 2 1 55466
0 55468 7 1 2 68422 96027
0 55469 5 1 1 55468
0 55470 7 1 2 55463 55469
0 55471 5 1 1 55470
0 55472 7 1 2 68648 55471
0 55473 5 1 1 55472
0 55474 7 1 2 85911 95471
0 55475 5 1 1 55474
0 55476 7 1 2 85913 96028
0 55477 7 1 2 55475 55476
0 55478 5 1 1 55477
0 55479 7 1 2 65102 84847
0 55480 7 1 2 81199 55479
0 55481 5 1 1 55480
0 55482 7 1 2 95670 55481
0 55483 5 1 1 55482
0 55484 7 1 2 61754 55483
0 55485 5 1 1 55484
0 55486 7 2 2 68813 75341
0 55487 5 1 1 96029
0 55488 7 1 2 69433 96030
0 55489 5 1 1 55488
0 55490 7 1 2 71456 93275
0 55491 7 1 2 55489 55490
0 55492 5 1 1 55491
0 55493 7 1 2 84704 55492
0 55494 5 1 1 55493
0 55495 7 1 2 55485 55494
0 55496 7 1 2 55478 55495
0 55497 7 1 2 55473 55496
0 55498 7 1 2 55453 55497
0 55499 5 1 1 55498
0 55500 7 1 2 69687 55499
0 55501 5 1 1 55500
0 55502 7 1 2 55430 55501
0 55503 5 1 1 55502
0 55504 7 1 2 66877 55503
0 55505 5 1 1 55504
0 55506 7 1 2 62004 55505
0 55507 7 1 2 55322 55506
0 55508 5 1 1 55507
0 55509 7 1 2 58690 92050
0 55510 5 1 1 55509
0 55511 7 1 2 58691 41587
0 55512 5 1 1 55511
0 55513 7 1 2 85704 55512
0 55514 7 1 2 16353 55513
0 55515 5 1 1 55514
0 55516 7 1 2 60694 55515
0 55517 5 1 1 55516
0 55518 7 1 2 55510 55517
0 55519 5 1 1 55518
0 55520 7 1 2 80444 55519
0 55521 5 1 1 55520
0 55522 7 1 2 65356 16204
0 55523 5 1 1 55522
0 55524 7 1 2 93803 95410
0 55525 5 1 1 55524
0 55526 7 1 2 55523 55525
0 55527 5 1 1 55526
0 55528 7 1 2 59700 55527
0 55529 5 1 1 55528
0 55530 7 1 2 69434 83311
0 55531 5 1 1 55530
0 55532 7 1 2 78403 78428
0 55533 7 1 2 55531 55532
0 55534 5 1 1 55533
0 55535 7 1 2 66099 55534
0 55536 5 1 1 55535
0 55537 7 1 2 55529 55536
0 55538 5 1 1 55537
0 55539 7 1 2 63427 55538
0 55540 5 1 1 55539
0 55541 7 1 2 55521 55540
0 55542 5 1 1 55541
0 55543 7 1 2 69293 55542
0 55544 5 1 1 55543
0 55545 7 1 2 73272 93705
0 55546 5 1 1 55545
0 55547 7 1 2 75473 94362
0 55548 5 1 1 55547
0 55549 7 1 2 85558 55548
0 55550 5 1 1 55549
0 55551 7 1 2 55546 55550
0 55552 5 1 1 55551
0 55553 7 1 2 59701 55552
0 55554 5 1 1 55553
0 55555 7 1 2 77931 84330
0 55556 5 1 1 55555
0 55557 7 1 2 83312 55556
0 55558 5 1 1 55557
0 55559 7 1 2 76306 80352
0 55560 5 1 1 55559
0 55561 7 1 2 76235 55560
0 55562 7 1 2 55558 55561
0 55563 5 1 1 55562
0 55564 7 1 2 61492 55563
0 55565 5 1 1 55564
0 55566 7 1 2 55554 55565
0 55567 5 1 1 55566
0 55568 7 1 2 69688 55567
0 55569 5 1 1 55568
0 55570 7 1 2 66100 82250
0 55571 5 1 1 55570
0 55572 7 1 2 65357 96006
0 55573 5 1 1 55572
0 55574 7 1 2 55571 55573
0 55575 5 1 1 55574
0 55576 7 1 2 63120 55575
0 55577 5 1 1 55576
0 55578 7 1 2 66398 55577
0 55579 7 1 2 55569 55578
0 55580 7 1 2 55544 55579
0 55581 5 1 1 55580
0 55582 7 1 2 86150 69294
0 55583 5 1 1 55582
0 55584 7 1 2 68697 55583
0 55585 5 1 1 55584
0 55586 7 1 2 85892 55585
0 55587 5 1 1 55586
0 55588 7 1 2 80024 88838
0 55589 5 1 1 55588
0 55590 7 1 2 84856 69689
0 55591 5 1 1 55590
0 55592 7 1 2 55589 55591
0 55593 5 1 1 55592
0 55594 7 1 2 95965 55593
0 55595 5 1 1 55594
0 55596 7 1 2 55587 55595
0 55597 5 1 1 55596
0 55598 7 1 2 77162 55597
0 55599 5 1 1 55598
0 55600 7 1 2 57817 80090
0 55601 5 1 1 55600
0 55602 7 1 2 95610 55601
0 55603 5 1 1 55602
0 55604 7 1 2 72920 55603
0 55605 5 1 1 55604
0 55606 7 1 2 910 72264
0 55607 5 1 1 55606
0 55608 7 1 2 85540 55607
0 55609 5 1 1 55608
0 55610 7 1 2 55605 55609
0 55611 5 1 1 55610
0 55612 7 1 2 80331 55611
0 55613 5 1 1 55612
0 55614 7 1 2 67421 69295
0 55615 5 1 1 55614
0 55616 7 1 2 68698 55615
0 55617 5 1 1 55616
0 55618 7 1 2 85893 55617
0 55619 5 1 1 55618
0 55620 7 1 2 83053 95966
0 55621 5 1 1 55620
0 55622 7 1 2 55619 55621
0 55623 5 1 1 55622
0 55624 7 1 2 71930 55623
0 55625 5 1 1 55624
0 55626 7 1 2 69705 344
0 55627 5 2 1 55626
0 55628 7 1 2 94385 96031
0 55629 5 1 1 55628
0 55630 7 1 2 84569 85656
0 55631 7 1 2 69690 55630
0 55632 5 1 1 55631
0 55633 7 1 2 55629 55632
0 55634 5 1 1 55633
0 55635 7 1 2 58692 55634
0 55636 5 1 1 55635
0 55637 7 1 2 84570 69353
0 55638 7 1 2 90011 55637
0 55639 5 1 1 55638
0 55640 7 1 2 61755 55639
0 55641 7 1 2 55636 55640
0 55642 7 1 2 55625 55641
0 55643 7 1 2 55613 55642
0 55644 7 1 2 55599 55643
0 55645 5 1 1 55644
0 55646 7 1 2 66797 55645
0 55647 7 1 2 55581 55646
0 55648 5 1 1 55647
0 55649 7 1 2 77937 79014
0 55650 5 1 1 55649
0 55651 7 1 2 80403 95959
0 55652 5 1 1 55651
0 55653 7 1 2 55650 55652
0 55654 5 1 1 55653
0 55655 7 1 2 69296 55654
0 55656 5 1 1 55655
0 55657 7 1 2 79245 80715
0 55658 7 1 2 82343 55657
0 55659 5 1 1 55658
0 55660 7 1 2 48369 55659
0 55661 5 1 1 55660
0 55662 7 1 2 80302 83864
0 55663 5 1 1 55662
0 55664 7 1 2 95419 55663
0 55665 5 1 1 55664
0 55666 7 1 2 83875 55665
0 55667 5 1 1 55666
0 55668 7 1 2 55661 55667
0 55669 5 1 1 55668
0 55670 7 1 2 55656 55669
0 55671 5 1 1 55670
0 55672 7 1 2 82190 55671
0 55673 5 1 1 55672
0 55674 7 1 2 89308 90144
0 55675 5 1 1 55674
0 55676 7 1 2 84792 69691
0 55677 7 1 2 95868 55676
0 55678 5 1 1 55677
0 55679 7 1 2 55675 55678
0 55680 5 2 1 55679
0 55681 7 1 2 77077 96033
0 55682 5 1 1 55681
0 55683 7 1 2 85986 69562
0 55684 7 1 2 72314 91475
0 55685 7 1 2 55683 55684
0 55686 7 1 2 85861 92846
0 55687 7 1 2 55685 55686
0 55688 5 1 1 55687
0 55689 7 1 2 55682 55688
0 55690 5 1 1 55689
0 55691 7 1 2 68288 55690
0 55692 5 1 1 55691
0 55693 7 1 2 86654 80337
0 55694 7 1 2 95869 55693
0 55695 5 1 1 55694
0 55696 7 1 2 55692 55695
0 55697 7 1 2 55673 55696
0 55698 5 1 1 55697
0 55699 7 1 2 64427 55698
0 55700 5 1 1 55699
0 55701 7 1 2 66650 55700
0 55702 7 1 2 55648 55701
0 55703 5 1 1 55702
0 55704 7 1 2 55508 55703
0 55705 5 1 1 55704
0 55706 7 1 2 80907 78260
0 55707 7 1 2 55432 55706
0 55708 5 1 1 55707
0 55709 7 1 2 80036 55708
0 55710 5 1 1 55709
0 55711 7 1 2 72883 86918
0 55712 5 1 1 55711
0 55713 7 1 2 78167 80949
0 55714 5 1 1 55713
0 55715 7 1 2 55712 55714
0 55716 5 1 1 55715
0 55717 7 1 2 67407 55716
0 55718 5 1 1 55717
0 55719 7 1 2 81639 94179
0 55720 5 1 1 55719
0 55721 7 1 2 92888 93436
0 55722 5 1 1 55721
0 55723 7 1 2 55720 55722
0 55724 7 1 2 55718 55723
0 55725 5 1 1 55724
0 55726 7 1 2 69297 55725
0 55727 5 1 1 55726
0 55728 7 1 2 55710 55727
0 55729 5 1 1 55728
0 55730 7 1 2 63560 55729
0 55731 5 1 1 55730
0 55732 7 1 2 83395 88082
0 55733 5 1 1 55732
0 55734 7 1 2 72802 69692
0 55735 5 1 1 55734
0 55736 7 1 2 55733 55735
0 55737 5 1 1 55736
0 55738 7 1 2 63121 55737
0 55739 5 1 1 55738
0 55740 7 1 2 7459 55739
0 55741 5 1 1 55740
0 55742 7 1 2 67233 55741
0 55743 5 1 1 55742
0 55744 7 1 2 63122 95046
0 55745 7 1 2 50963 55744
0 55746 7 1 2 81631 55745
0 55747 5 1 1 55746
0 55748 7 1 2 69584 83670
0 55749 7 1 2 55747 55748
0 55750 5 1 1 55749
0 55751 7 1 2 55743 55750
0 55752 5 1 1 55751
0 55753 7 1 2 66101 55752
0 55754 5 1 1 55753
0 55755 7 1 2 73784 68688
0 55756 5 1 1 55755
0 55757 7 1 2 54790 55756
0 55758 5 1 1 55757
0 55759 7 1 2 63561 55758
0 55760 5 1 1 55759
0 55761 7 1 2 80960 90552
0 55762 7 1 2 89537 55761
0 55763 5 1 1 55762
0 55764 7 1 2 55760 55763
0 55765 5 1 1 55764
0 55766 7 1 2 78886 55765
0 55767 5 1 1 55766
0 55768 7 1 2 79246 80222
0 55769 7 1 2 89301 55768
0 55770 5 1 1 55769
0 55771 7 1 2 55767 55770
0 55772 5 1 1 55771
0 55773 7 1 2 68289 55772
0 55774 5 1 1 55773
0 55775 7 1 2 55754 55774
0 55776 7 1 2 55731 55775
0 55777 5 1 1 55776
0 55778 7 1 2 66399 55777
0 55779 5 1 1 55778
0 55780 7 1 2 72396 72565
0 55781 7 1 2 94197 55780
0 55782 5 1 1 55781
0 55783 7 1 2 76420 55782
0 55784 5 1 1 55783
0 55785 7 1 2 57536 55784
0 55786 5 1 1 55785
0 55787 7 1 2 69474 69693
0 55788 5 1 1 55787
0 55789 7 1 2 55786 55788
0 55790 5 1 1 55789
0 55791 7 1 2 66102 55790
0 55792 5 1 1 55791
0 55793 7 1 2 95611 55792
0 55794 5 1 1 55793
0 55795 7 1 2 67408 55794
0 55796 5 1 1 55795
0 55797 7 1 2 67805 84355
0 55798 5 1 1 55797
0 55799 7 1 2 69298 55798
0 55800 5 1 1 55799
0 55801 7 1 2 68699 55800
0 55802 5 1 1 55801
0 55803 7 1 2 58693 55802
0 55804 5 1 1 55803
0 55805 7 1 2 69500 48598
0 55806 5 2 1 55805
0 55807 7 1 2 68061 96035
0 55808 5 1 1 55807
0 55809 7 1 2 73569 68689
0 55810 5 1 1 55809
0 55811 7 1 2 55808 55810
0 55812 5 1 1 55811
0 55813 7 1 2 67703 55812
0 55814 5 1 1 55813
0 55815 7 1 2 58094 72176
0 55816 7 1 2 96016 55815
0 55817 5 1 1 55816
0 55818 7 1 2 55814 55817
0 55819 7 1 2 55804 55818
0 55820 7 1 2 55796 55819
0 55821 5 1 1 55820
0 55822 7 1 2 71566 55821
0 55823 5 1 1 55822
0 55824 7 1 2 95038 95961
0 55825 5 3 1 55824
0 55826 7 1 2 69496 96037
0 55827 5 1 1 55826
0 55828 7 1 2 85308 72921
0 55829 5 1 1 55828
0 55830 7 1 2 70439 85541
0 55831 5 1 1 55830
0 55832 7 1 2 55829 55831
0 55833 5 1 1 55832
0 55834 7 1 2 69299 55833
0 55835 5 1 1 55834
0 55836 7 1 2 55827 55835
0 55837 5 1 1 55836
0 55838 7 1 2 68423 55837
0 55839 5 1 1 55838
0 55840 7 1 2 82932 47766
0 55841 7 1 2 95039 55840
0 55842 5 1 1 55841
0 55843 7 1 2 69354 55842
0 55844 5 1 1 55843
0 55845 7 1 2 82985 80716
0 55846 7 1 2 69300 55845
0 55847 5 1 1 55846
0 55848 7 1 2 55844 55847
0 55849 5 1 1 55848
0 55850 7 1 2 67704 55849
0 55851 5 1 1 55850
0 55852 7 1 2 55839 55851
0 55853 5 1 1 55852
0 55854 7 1 2 77163 55853
0 55855 5 1 1 55854
0 55856 7 1 2 68700 3037
0 55857 5 1 1 55856
0 55858 7 1 2 58095 55857
0 55859 5 1 1 55858
0 55860 7 1 2 72185 55859
0 55861 5 2 1 55860
0 55862 7 1 2 95967 96040
0 55863 5 1 1 55862
0 55864 7 1 2 85894 76840
0 55865 5 1 1 55864
0 55866 7 1 2 55863 55865
0 55867 5 1 1 55866
0 55868 7 1 2 72277 55867
0 55869 5 1 1 55868
0 55870 7 1 2 78641 96041
0 55871 5 1 1 55870
0 55872 7 1 2 67705 69301
0 55873 5 1 1 55872
0 55874 7 1 2 69706 55873
0 55875 5 1 1 55874
0 55876 7 1 2 85845 55875
0 55877 5 1 1 55876
0 55878 7 1 2 70799 80028
0 55879 5 1 1 55878
0 55880 7 1 2 67409 96036
0 55881 5 1 1 55880
0 55882 7 1 2 55879 55881
0 55883 7 1 2 55877 55882
0 55884 7 1 2 55871 55883
0 55885 5 1 1 55884
0 55886 7 1 2 82986 55885
0 55887 5 1 1 55886
0 55888 7 1 2 69197 68690
0 55889 7 1 2 95978 55888
0 55890 5 1 1 55889
0 55891 7 1 2 55887 55890
0 55892 7 1 2 55869 55891
0 55893 7 1 2 55855 55892
0 55894 7 1 2 55823 55893
0 55895 5 1 1 55894
0 55896 7 1 2 90299 55895
0 55897 5 1 1 55896
0 55898 7 1 2 55779 55897
0 55899 5 1 1 55898
0 55900 7 1 2 75742 55899
0 55901 5 1 1 55900
0 55902 7 1 2 85660 94613
0 55903 5 1 1 55902
0 55904 7 1 2 95962 55903
0 55905 5 1 1 55904
0 55906 7 1 2 95498 55905
0 55907 5 1 1 55906
0 55908 7 1 2 69014 84705
0 55909 5 2 1 55908
0 55910 7 1 2 55907 96042
0 55911 5 1 1 55910
0 55912 7 1 2 71931 55911
0 55913 5 1 1 55912
0 55914 7 1 2 66400 95334
0 55915 5 1 1 55914
0 55916 7 2 2 61756 96038
0 55917 5 1 1 96044
0 55918 7 1 2 57537 96045
0 55919 5 1 1 55918
0 55920 7 1 2 55915 55919
0 55921 5 1 1 55920
0 55922 7 1 2 81605 55921
0 55923 5 1 1 55922
0 55924 7 1 2 81273 95821
0 55925 5 1 1 55924
0 55926 7 1 2 73913 55925
0 55927 5 1 1 55926
0 55928 7 1 2 55923 55927
0 55929 7 1 2 55913 55928
0 55930 7 1 2 57818 96039
0 55931 5 1 1 55930
0 55932 7 1 2 70800 85657
0 55933 7 1 2 92763 55932
0 55934 5 1 1 55933
0 55935 7 1 2 55931 55934
0 55936 5 1 1 55935
0 55937 7 1 2 57538 55936
0 55938 5 1 1 55937
0 55939 7 2 2 65358 86272
0 55940 7 1 2 83352 96046
0 55941 5 1 1 55940
0 55942 7 1 2 55938 55941
0 55943 5 1 1 55942
0 55944 7 1 2 61757 55943
0 55945 5 1 1 55944
0 55946 7 1 2 85661 94246
0 55947 5 1 1 55946
0 55948 7 1 2 94936 55917
0 55949 5 1 1 55948
0 55950 7 1 2 70973 55949
0 55951 5 1 1 55950
0 55952 7 1 2 55947 55951
0 55953 5 1 1 55952
0 55954 7 1 2 71766 55953
0 55955 5 1 1 55954
0 55956 7 1 2 55945 55955
0 55957 7 1 2 55929 55956
0 55958 5 1 1 55957
0 55959 7 1 2 69694 55958
0 55960 5 1 1 55959
0 55961 7 1 2 78736 77083
0 55962 5 1 1 55961
0 55963 7 1 2 57539 91859
0 55964 5 1 1 55963
0 55965 7 1 2 80053 55964
0 55966 5 1 1 55965
0 55967 7 1 2 57819 55966
0 55968 5 1 1 55967
0 55969 7 1 2 63123 95117
0 55970 7 1 2 55968 55969
0 55971 5 1 1 55970
0 55972 7 1 2 64428 55971
0 55973 5 1 1 55972
0 55974 7 1 2 55962 55973
0 55975 5 1 1 55974
0 55976 7 1 2 61493 55975
0 55977 5 1 1 55976
0 55978 7 1 2 86991 55977
0 55979 5 1 1 55978
0 55980 7 1 2 67410 55979
0 55981 5 1 1 55980
0 55982 7 1 2 69509 3377
0 55983 5 1 1 55982
0 55984 7 1 2 57540 55983
0 55985 5 1 1 55984
0 55986 7 1 2 80066 55985
0 55987 5 1 1 55986
0 55988 7 1 2 85855 55987
0 55989 5 1 1 55988
0 55990 7 1 2 71629 80376
0 55991 5 1 1 55990
0 55992 7 1 2 84037 55991
0 55993 5 1 1 55992
0 55994 7 1 2 73098 55993
0 55995 5 1 1 55994
0 55996 7 1 2 86987 92872
0 55997 5 1 1 55996
0 55998 7 1 2 66401 55997
0 55999 7 1 2 55995 55998
0 56000 7 1 2 55989 55999
0 56001 7 1 2 55981 56000
0 56002 5 1 1 56001
0 56003 7 1 2 68062 85962
0 56004 5 1 1 56003
0 56005 7 1 2 86911 56004
0 56006 7 1 2 81642 56005
0 56007 5 1 1 56006
0 56008 7 1 2 95968 56007
0 56009 5 1 1 56008
0 56010 7 1 2 85022 96047
0 56011 5 1 1 56010
0 56012 7 1 2 85895 94902
0 56013 5 1 1 56012
0 56014 7 1 2 61758 56013
0 56015 7 1 2 56011 56014
0 56016 7 1 2 56009 56015
0 56017 5 1 1 56016
0 56018 7 1 2 69585 56017
0 56019 7 1 2 56002 56018
0 56020 5 1 1 56019
0 56021 7 1 2 55960 56020
0 56022 5 1 1 56021
0 56023 7 1 2 66878 56022
0 56024 5 1 1 56023
0 56025 7 1 2 86696 87290
0 56026 5 1 1 56025
0 56027 7 1 2 17720 94937
0 56028 5 1 1 56027
0 56029 7 1 2 71767 56028
0 56030 5 1 1 56029
0 56031 7 1 2 57541 87480
0 56032 5 1 1 56031
0 56033 7 1 2 96043 56032
0 56034 7 1 2 56030 56033
0 56035 5 1 1 56034
0 56036 7 1 2 70801 56035
0 56037 5 1 1 56036
0 56038 7 1 2 56026 56037
0 56039 5 1 1 56038
0 56040 7 1 2 58372 56039
0 56041 5 1 1 56040
0 56042 7 1 2 73230 95854
0 56043 7 1 2 75286 56042
0 56044 5 1 1 56043
0 56045 7 1 2 56041 56044
0 56046 5 1 1 56045
0 56047 7 1 2 57820 56046
0 56048 5 1 1 56047
0 56049 7 1 2 65103 87228
0 56050 7 1 2 74557 56049
0 56051 5 1 1 56050
0 56052 7 1 2 84709 56051
0 56053 5 1 1 56052
0 56054 7 1 2 71236 56053
0 56055 5 1 1 56054
0 56056 7 1 2 56048 56055
0 56057 5 1 1 56056
0 56058 7 1 2 69695 56057
0 56059 5 1 1 56058
0 56060 7 1 2 74581 73424
0 56061 7 1 2 72566 56060
0 56062 7 1 2 95243 95652
0 56063 7 1 2 56061 56062
0 56064 5 1 1 56063
0 56065 7 1 2 56059 56064
0 56066 5 1 1 56065
0 56067 7 1 2 67411 56066
0 56068 5 1 1 56067
0 56069 7 2 2 61494 78892
0 56070 7 1 2 83031 96048
0 56071 5 1 1 56070
0 56072 7 1 2 81606 69696
0 56073 5 1 1 56072
0 56074 7 1 2 57821 80342
0 56075 7 1 2 72433 56074
0 56076 5 1 1 56075
0 56077 7 1 2 56073 56076
0 56078 5 1 1 56077
0 56079 7 1 2 57542 56078
0 56080 5 1 1 56079
0 56081 7 1 2 78837 67609
0 56082 7 1 2 81291 56081
0 56083 5 1 1 56082
0 56084 7 1 2 69697 56083
0 56085 5 1 1 56084
0 56086 7 1 2 56080 56085
0 56087 5 1 1 56086
0 56088 7 1 2 86510 56087
0 56089 5 1 1 56088
0 56090 7 1 2 57543 94983
0 56091 7 1 2 72220 56090
0 56092 5 1 1 56091
0 56093 7 1 2 56089 56092
0 56094 5 1 1 56093
0 56095 7 1 2 59702 56094
0 56096 5 1 1 56095
0 56097 7 1 2 56071 56096
0 56098 5 1 1 56097
0 56099 7 1 2 78915 56098
0 56100 5 1 1 56099
0 56101 7 1 2 70440 82244
0 56102 7 1 2 96014 56101
0 56103 7 1 2 96049 56102
0 56104 5 1 1 56103
0 56105 7 1 2 56100 56104
0 56106 7 1 2 56068 56105
0 56107 5 1 1 56106
0 56108 7 1 2 58694 66805
0 56109 7 1 2 56107 56108
0 56110 5 1 1 56109
0 56111 7 1 2 56024 56110
0 56112 5 1 1 56111
0 56113 7 1 2 62005 56112
0 56114 5 1 1 56113
0 56115 7 1 2 55901 56114
0 56116 5 1 1 56115
0 56117 7 1 2 65749 56116
0 56118 5 1 1 56117
0 56119 7 1 2 77298 83331
0 56120 7 1 2 90288 96022
0 56121 7 1 2 56119 56120
0 56122 5 1 1 56121
0 56123 7 1 2 64429 66651
0 56124 7 1 2 78149 56123
0 56125 7 1 2 96034 56124
0 56126 5 1 1 56125
0 56127 7 1 2 56122 56126
0 56128 5 1 1 56127
0 56129 7 1 2 84331 56128
0 56130 5 1 1 56129
0 56131 7 1 2 56118 56130
0 56132 7 1 2 55705 56131
0 56133 5 1 1 56132
0 56134 7 1 2 59949 56133
0 56135 5 1 1 56134
0 56136 7 1 2 70335 71338
0 56137 5 1 1 56136
0 56138 7 1 2 93218 56137
0 56139 5 1 1 56138
0 56140 7 1 2 63428 56139
0 56141 5 1 1 56140
0 56142 7 1 2 93193 56141
0 56143 5 1 1 56142
0 56144 7 1 2 64645 56143
0 56145 5 1 1 56144
0 56146 7 1 2 93223 56145
0 56147 5 1 1 56146
0 56148 7 1 2 91773 56147
0 56149 5 1 1 56148
0 56150 7 1 2 65359 77183
0 56151 5 1 1 56150
0 56152 7 1 2 86154 56151
0 56153 5 1 1 56152
0 56154 7 1 2 67412 74303
0 56155 7 1 2 91746 56154
0 56156 7 1 2 56153 56155
0 56157 5 1 1 56156
0 56158 7 1 2 68063 72661
0 56159 7 1 2 95681 56158
0 56160 5 1 1 56159
0 56161 7 2 2 92074 93969
0 56162 5 1 1 96050
0 56163 7 1 2 56160 56162
0 56164 7 1 2 56157 56163
0 56165 5 1 1 56164
0 56166 7 1 2 58373 56165
0 56167 5 1 1 56166
0 56168 7 1 2 92873 95628
0 56169 5 1 1 56168
0 56170 7 1 2 68541 90752
0 56171 5 1 1 56170
0 56172 7 1 2 96051 56171
0 56173 5 1 1 56172
0 56174 7 1 2 56169 56173
0 56175 7 1 2 56167 56174
0 56176 7 1 2 56149 56175
0 56177 5 1 1 56176
0 56178 7 1 2 63656 56177
0 56179 5 1 1 56178
0 56180 7 1 2 70465 56179
0 56181 5 1 1 56180
0 56182 7 1 2 58695 17342
0 56183 5 2 1 56182
0 56184 7 4 2 94145 96052
0 56185 7 1 2 62819 91223
0 56186 5 1 1 56185
0 56187 7 1 2 70234 71772
0 56188 5 1 1 56187
0 56189 7 1 2 67413 76261
0 56190 5 1 1 56189
0 56191 7 1 2 84932 56190
0 56192 5 1 1 56191
0 56193 7 1 2 56188 56192
0 56194 7 1 2 56186 56193
0 56195 5 1 1 56194
0 56196 7 1 2 96054 56195
0 56197 5 1 1 56196
0 56198 7 1 2 76664 72922
0 56199 5 2 1 56198
0 56200 7 2 2 61124 96058
0 56201 7 1 2 64118 95075
0 56202 7 1 2 96060 56201
0 56203 5 1 1 56202
0 56204 7 1 2 56197 56203
0 56205 5 1 1 56204
0 56206 7 1 2 70855 56205
0 56207 5 1 1 56206
0 56208 7 1 2 81101 96055
0 56209 5 1 1 56208
0 56210 7 1 2 94831 96061
0 56211 5 1 1 56210
0 56212 7 1 2 56209 56211
0 56213 5 1 1 56212
0 56214 7 1 2 62820 56213
0 56215 5 1 1 56214
0 56216 7 1 2 81314 87757
0 56217 5 1 1 56216
0 56218 7 1 2 96056 56217
0 56219 5 1 1 56218
0 56220 7 1 2 56215 56219
0 56221 5 1 1 56220
0 56222 7 1 2 78354 56221
0 56223 5 1 1 56222
0 56224 7 1 2 64646 91671
0 56225 5 1 1 56224
0 56226 7 1 2 70264 74862
0 56227 5 1 1 56226
0 56228 7 1 2 76272 56227
0 56229 5 1 1 56228
0 56230 7 1 2 21478 56229
0 56231 5 1 1 56230
0 56232 7 1 2 96057 56231
0 56233 5 1 1 56232
0 56234 7 1 2 56225 56233
0 56235 7 1 2 56223 56234
0 56236 7 1 2 56207 56235
0 56237 5 1 1 56236
0 56238 7 1 2 62006 56237
0 56239 5 1 1 56238
0 56240 7 1 2 69566 56239
0 56241 5 1 1 56240
0 56242 7 1 2 66736 56241
0 56243 7 1 2 56181 56242
0 56244 5 1 1 56243
0 56245 7 1 2 12943 87972
0 56246 5 1 1 56245
0 56247 7 1 2 69563 93296
0 56248 5 1 1 56247
0 56249 7 1 2 56246 56248
0 56250 5 1 1 56249
0 56251 7 1 2 66652 56250
0 56252 5 1 1 56251
0 56253 7 1 2 71567 94597
0 56254 7 1 2 77164 56253
0 56255 5 1 1 56254
0 56256 7 1 2 82297 56255
0 56257 5 1 1 56256
0 56258 7 1 2 71932 56257
0 56259 5 1 1 56258
0 56260 7 1 2 82242 95843
0 56261 5 1 1 56260
0 56262 7 1 2 71339 56261
0 56263 5 1 1 56262
0 56264 7 1 2 75945 56263
0 56265 5 1 1 56264
0 56266 7 1 2 56259 56265
0 56267 5 1 1 56266
0 56268 7 1 2 95608 56267
0 56269 5 1 1 56268
0 56270 7 1 2 71933 78642
0 56271 5 1 1 56270
0 56272 7 1 2 87360 56271
0 56273 5 1 1 56272
0 56274 7 1 2 58096 56273
0 56275 5 1 1 56274
0 56276 7 1 2 86892 56275
0 56277 5 1 1 56276
0 56278 7 1 2 65750 56277
0 56279 5 1 1 56278
0 56280 7 1 2 86310 95970
0 56281 5 1 1 56280
0 56282 7 1 2 56279 56281
0 56283 5 1 1 56282
0 56284 7 1 2 82987 56283
0 56285 5 1 1 56284
0 56286 7 1 2 85142 92876
0 56287 5 1 1 56286
0 56288 7 1 2 56285 56287
0 56289 5 1 1 56288
0 56290 7 1 2 69698 56289
0 56291 5 1 1 56290
0 56292 7 1 2 56269 56291
0 56293 5 1 1 56292
0 56294 7 1 2 59393 56293
0 56295 5 1 1 56294
0 56296 7 1 2 71934 80129
0 56297 5 1 1 56296
0 56298 7 1 2 80015 72265
0 56299 7 1 2 56297 56298
0 56300 5 1 1 56299
0 56301 7 1 2 75287 56300
0 56302 5 1 1 56301
0 56303 7 1 2 86140 69699
0 56304 5 1 1 56303
0 56305 7 1 2 56302 56304
0 56306 5 1 1 56305
0 56307 7 1 2 65751 56306
0 56308 5 1 1 56307
0 56309 7 1 2 69201 81680
0 56310 5 1 1 56309
0 56311 7 1 2 69497 56310
0 56312 5 1 1 56311
0 56313 7 1 2 56308 56312
0 56314 5 1 1 56313
0 56315 7 1 2 71568 56314
0 56316 5 1 1 56315
0 56317 7 1 2 69302 82299
0 56318 5 1 1 56317
0 56319 7 1 2 69198 72121
0 56320 5 1 1 56319
0 56321 7 1 2 56318 56320
0 56322 5 1 1 56321
0 56323 7 1 2 77165 56322
0 56324 5 1 1 56323
0 56325 7 1 2 72171 74163
0 56326 5 1 1 56325
0 56327 7 1 2 6553 68701
0 56328 5 1 1 56327
0 56329 7 1 2 58097 56328
0 56330 5 1 1 56329
0 56331 7 1 2 72127 56330
0 56332 5 1 1 56331
0 56333 7 1 2 71569 56332
0 56334 5 1 1 56333
0 56335 7 1 2 56326 56334
0 56336 7 1 2 56324 56335
0 56337 5 1 1 56336
0 56338 7 1 2 72254 56337
0 56339 5 1 1 56338
0 56340 7 1 2 73296 75935
0 56341 5 1 1 56340
0 56342 7 1 2 75288 56341
0 56343 5 1 1 56342
0 56344 7 1 2 70974 75946
0 56345 5 1 1 56344
0 56346 7 1 2 76344 69357
0 56347 7 1 2 56345 56346
0 56348 7 1 2 56343 56347
0 56349 5 1 1 56348
0 56350 7 1 2 71237 96032
0 56351 7 1 2 56349 56350
0 56352 5 1 1 56351
0 56353 7 1 2 56339 56352
0 56354 7 1 2 56316 56353
0 56355 5 1 1 56354
0 56356 7 1 2 58696 56355
0 56357 5 1 1 56356
0 56358 7 1 2 58904 76334
0 56359 7 1 2 94567 56358
0 56360 7 1 2 75919 56359
0 56361 7 1 2 84099 56360
0 56362 5 1 1 56361
0 56363 7 1 2 56357 56362
0 56364 7 1 2 56295 56363
0 56365 5 1 1 56364
0 56366 7 1 2 91414 56365
0 56367 5 1 1 56366
0 56368 7 1 2 56252 56367
0 56369 5 1 1 56368
0 56370 7 1 2 66103 56369
0 56371 5 1 1 56370
0 56372 7 1 2 84207 10979
0 56373 5 1 1 56372
0 56374 7 1 2 68186 56373
0 56375 5 1 1 56374
0 56376 7 1 2 85319 21674
0 56377 5 1 1 56376
0 56378 7 1 2 61125 56377
0 56379 5 1 1 56378
0 56380 7 1 2 56375 56379
0 56381 5 1 1 56380
0 56382 7 1 2 61495 56381
0 56383 5 1 1 56382
0 56384 7 1 2 38783 56383
0 56385 5 1 1 56384
0 56386 7 1 2 76718 56385
0 56387 5 1 1 56386
0 56388 7 1 2 85649 79382
0 56389 5 1 1 56388
0 56390 7 1 2 75605 56389
0 56391 5 1 1 56390
0 56392 7 1 2 68542 56391
0 56393 5 1 1 56392
0 56394 7 1 2 28633 56393
0 56395 5 1 1 56394
0 56396 7 1 2 68187 56395
0 56397 5 1 1 56396
0 56398 7 1 2 84815 85650
0 56399 5 1 1 56398
0 56400 7 1 2 68649 89933
0 56401 5 1 1 56400
0 56402 7 1 2 64647 56401
0 56403 7 1 2 85488 56402
0 56404 5 1 1 56403
0 56405 7 1 2 56399 56404
0 56406 5 1 1 56405
0 56407 7 1 2 61126 56406
0 56408 5 1 1 56407
0 56409 7 1 2 56397 56408
0 56410 7 1 2 56387 56409
0 56411 5 1 1 56410
0 56412 7 1 2 67806 56411
0 56413 5 1 1 56412
0 56414 7 1 2 85838 79500
0 56415 5 1 1 56414
0 56416 7 1 2 71340 84725
0 56417 5 1 1 56416
0 56418 7 1 2 85981 93144
0 56419 7 1 2 94166 56418
0 56420 7 1 2 56417 56419
0 56421 5 1 1 56420
0 56422 7 1 2 61127 56421
0 56423 5 1 1 56422
0 56424 7 1 2 56415 56423
0 56425 5 1 1 56424
0 56426 7 1 2 76719 56425
0 56427 5 1 1 56426
0 56428 7 1 2 15258 25630
0 56429 5 1 1 56428
0 56430 7 1 2 81083 56429
0 56431 5 1 1 56430
0 56432 7 1 2 56427 56431
0 56433 5 1 1 56432
0 56434 7 1 2 84353 56433
0 56435 5 1 1 56434
0 56436 7 1 2 76720 26368
0 56437 5 1 1 56436
0 56438 7 1 2 85658 56437
0 56439 5 1 1 56438
0 56440 7 1 2 73919 56439
0 56441 5 1 1 56440
0 56442 7 1 2 72884 89677
0 56443 5 1 1 56442
0 56444 7 1 2 34535 56443
0 56445 5 1 1 56444
0 56446 7 1 2 60425 56445
0 56447 5 1 1 56446
0 56448 7 1 2 56441 56447
0 56449 5 1 1 56448
0 56450 7 1 2 70953 56449
0 56451 5 1 1 56450
0 56452 7 1 2 56435 56451
0 56453 5 1 1 56452
0 56454 7 1 2 68892 56453
0 56455 5 1 1 56454
0 56456 7 1 2 68424 80379
0 56457 5 1 1 56456
0 56458 7 1 2 89678 56457
0 56459 5 1 1 56458
0 56460 7 2 2 81659 90730
0 56461 5 1 1 96062
0 56462 7 1 2 80377 96063
0 56463 5 1 1 56462
0 56464 7 1 2 93268 56463
0 56465 7 1 2 56459 56464
0 56466 5 1 1 56465
0 56467 7 1 2 72885 56466
0 56468 5 1 1 56467
0 56469 7 1 2 68543 95122
0 56470 5 1 1 56469
0 56471 7 1 2 90757 56470
0 56472 5 1 1 56471
0 56473 7 1 2 85206 56472
0 56474 5 1 1 56473
0 56475 7 1 2 76910 68427
0 56476 5 1 1 56475
0 56477 7 1 2 75565 56476
0 56478 5 1 1 56477
0 56479 7 1 2 56474 56478
0 56480 7 1 2 56468 56479
0 56481 5 1 1 56480
0 56482 7 1 2 61128 56481
0 56483 5 1 1 56482
0 56484 7 1 2 68544 92935
0 56485 5 1 1 56484
0 56486 7 1 2 72923 85595
0 56487 7 1 2 56485 56486
0 56488 5 1 1 56487
0 56489 7 1 2 76721 85826
0 56490 7 1 2 56488 56489
0 56491 5 1 1 56490
0 56492 7 1 2 75606 56491
0 56493 5 1 1 56492
0 56494 7 1 2 93044 56493
0 56495 5 1 1 56494
0 56496 7 1 2 68443 96053
0 56497 5 1 1 56496
0 56498 7 1 2 77431 84604
0 56499 5 1 1 56498
0 56500 7 1 2 56497 56499
0 56501 5 1 1 56500
0 56502 7 1 2 76901 94146
0 56503 7 1 2 56501 56502
0 56504 5 1 1 56503
0 56505 7 1 2 56495 56504
0 56506 7 1 2 56483 56505
0 56507 7 1 2 56455 56506
0 56508 7 1 2 56413 56507
0 56509 5 1 1 56508
0 56510 7 1 2 72689 56509
0 56511 5 1 1 56510
0 56512 7 1 2 66402 56511
0 56513 7 1 2 56371 56512
0 56514 7 1 2 56244 56513
0 56515 5 1 1 56514
0 56516 7 1 2 61129 84088
0 56517 5 1 1 56516
0 56518 7 1 2 67807 92479
0 56519 5 1 1 56518
0 56520 7 1 2 30455 56519
0 56521 7 1 2 56517 56520
0 56522 5 1 1 56521
0 56523 7 1 2 63429 56522
0 56524 5 1 1 56523
0 56525 7 1 2 78574 84047
0 56526 5 1 1 56525
0 56527 7 1 2 56524 56526
0 56528 5 1 1 56527
0 56529 7 1 2 68188 56528
0 56530 5 1 1 56529
0 56531 7 1 2 76888 83586
0 56532 5 1 1 56531
0 56533 7 1 2 80826 92739
0 56534 5 1 1 56533
0 56535 7 1 2 93790 56534
0 56536 5 1 1 56535
0 56537 7 1 2 56532 56536
0 56538 7 1 2 56530 56537
0 56539 5 1 1 56538
0 56540 7 1 2 59950 56539
0 56541 5 1 1 56540
0 56542 7 1 2 67808 93624
0 56543 5 1 1 56542
0 56544 7 1 2 11938 56543
0 56545 5 1 1 56544
0 56546 7 1 2 60695 56545
0 56547 5 1 1 56546
0 56548 7 1 2 78001 70116
0 56549 5 1 1 56548
0 56550 7 1 2 85143 56549
0 56551 7 1 2 56547 56550
0 56552 5 1 1 56551
0 56553 7 1 2 68189 56552
0 56554 5 1 1 56553
0 56555 7 1 2 76156 79735
0 56556 5 1 1 56555
0 56557 7 1 2 64430 56556
0 56558 5 1 1 56557
0 56559 7 1 2 72515 81238
0 56560 5 1 1 56559
0 56561 7 1 2 84975 56461
0 56562 7 1 2 56560 56561
0 56563 7 1 2 56558 56562
0 56564 5 1 1 56563
0 56565 7 1 2 78887 56564
0 56566 5 1 1 56565
0 56567 7 1 2 67414 85561
0 56568 5 1 1 56567
0 56569 7 1 2 78002 56568
0 56570 5 1 1 56569
0 56571 7 1 2 85489 70117
0 56572 5 1 1 56571
0 56573 7 1 2 59951 56572
0 56574 7 1 2 56570 56573
0 56575 7 1 2 56566 56574
0 56576 7 1 2 56554 56575
0 56577 5 1 1 56576
0 56578 7 1 2 61496 56577
0 56579 5 1 1 56578
0 56580 7 1 2 56541 56579
0 56581 5 1 1 56580
0 56582 7 1 2 81022 93795
0 56583 5 1 1 56582
0 56584 7 1 2 58374 56583
0 56585 5 1 1 56584
0 56586 7 1 2 68064 86885
0 56587 5 1 1 56586
0 56588 7 1 2 56585 56587
0 56589 7 1 2 86038 56588
0 56590 5 1 1 56589
0 56591 7 1 2 60696 56590
0 56592 5 1 1 56591
0 56593 7 1 2 74100 86815
0 56594 5 1 1 56593
0 56595 7 1 2 87250 94921
0 56596 5 1 1 56595
0 56597 7 1 2 59703 56596
0 56598 5 1 1 56597
0 56599 7 1 2 65752 56598
0 56600 7 1 2 56594 56599
0 56601 7 1 2 56592 56600
0 56602 5 1 1 56601
0 56603 7 1 2 78277 81640
0 56604 5 1 1 56603
0 56605 7 1 2 71570 85963
0 56606 5 1 1 56605
0 56607 7 1 2 86912 56606
0 56608 5 1 1 56607
0 56609 7 1 2 67415 56608
0 56610 5 1 1 56609
0 56611 7 1 2 84841 78050
0 56612 7 1 2 56610 56611
0 56613 7 1 2 56604 56612
0 56614 5 1 1 56613
0 56615 7 1 2 56602 56614
0 56616 5 1 1 56615
0 56617 7 1 2 64648 8892
0 56618 7 1 2 56616 56617
0 56619 5 1 1 56618
0 56620 7 1 2 56581 56619
0 56621 5 1 1 56620
0 56622 7 1 2 78770 93619
0 56623 5 1 1 56622
0 56624 7 1 2 74605 56623
0 56625 5 1 1 56624
0 56626 7 1 2 67234 56625
0 56627 5 1 1 56626
0 56628 7 1 2 85354 94679
0 56629 5 1 1 56628
0 56630 7 1 2 56627 56629
0 56631 5 1 1 56630
0 56632 7 1 2 85189 56631
0 56633 5 1 1 56632
0 56634 7 1 2 84842 69435
0 56635 5 1 1 56634
0 56636 7 1 2 94989 56635
0 56637 5 1 1 56636
0 56638 7 1 2 82933 56637
0 56639 5 1 1 56638
0 56640 7 1 2 56633 56639
0 56641 5 1 1 56640
0 56642 7 1 2 65753 56641
0 56643 5 1 1 56642
0 56644 7 2 2 65104 84867
0 56645 5 3 1 96064
0 56646 7 1 2 91566 96066
0 56647 5 1 1 56646
0 56648 7 1 2 62538 56647
0 56649 5 1 1 56648
0 56650 7 1 2 59704 90814
0 56651 5 1 1 56650
0 56652 7 1 2 96067 56651
0 56653 5 1 1 56652
0 56654 7 1 2 68893 56653
0 56655 5 1 1 56654
0 56656 7 1 2 56649 56655
0 56657 5 1 1 56656
0 56658 7 1 2 70856 56657
0 56659 5 1 1 56658
0 56660 7 1 2 65360 80214
0 56661 5 1 1 56660
0 56662 7 1 2 74552 56661
0 56663 5 1 1 56662
0 56664 7 1 2 62821 56663
0 56665 5 1 1 56664
0 56666 7 1 2 65361 81487
0 56667 5 1 1 56666
0 56668 7 1 2 79411 56667
0 56669 7 1 2 56665 56668
0 56670 5 1 1 56669
0 56671 7 1 2 76968 56670
0 56672 5 1 1 56671
0 56673 7 1 2 59705 91431
0 56674 5 1 1 56673
0 56675 7 1 2 96068 56674
0 56676 5 1 1 56675
0 56677 7 1 2 71838 56676
0 56678 5 1 1 56677
0 56679 7 1 2 78178 56678
0 56680 7 1 2 56672 56679
0 56681 7 1 2 85144 82848
0 56682 5 1 1 56681
0 56683 7 1 2 65754 56682
0 56684 5 1 1 56683
0 56685 7 1 2 94328 56684
0 56686 5 1 1 56685
0 56687 7 1 2 69436 56686
0 56688 5 1 1 56687
0 56689 7 1 2 62539 96065
0 56690 5 1 1 56689
0 56691 7 1 2 85007 56690
0 56692 5 1 1 56691
0 56693 7 1 2 68894 56692
0 56694 5 1 1 56693
0 56695 7 1 2 56688 56694
0 56696 7 1 2 56680 56695
0 56697 7 1 2 56659 56696
0 56698 7 1 2 65755 74603
0 56699 5 1 1 56698
0 56700 7 1 2 86943 56699
0 56701 5 1 1 56700
0 56702 7 1 2 75842 56701
0 56703 5 1 1 56702
0 56704 7 1 2 95195 56703
0 56705 5 1 1 56704
0 56706 7 1 2 68895 56705
0 56707 5 1 1 56706
0 56708 7 1 2 84048 84736
0 56709 5 1 1 56708
0 56710 7 1 2 77751 56709
0 56711 7 1 2 56707 56710
0 56712 5 1 1 56711
0 56713 7 1 2 68190 56712
0 56714 5 1 1 56713
0 56715 7 1 2 70862 94987
0 56716 5 1 1 56715
0 56717 7 1 2 59394 76819
0 56718 5 1 1 56717
0 56719 7 1 2 62822 56718
0 56720 5 1 1 56719
0 56721 7 1 2 77620 91995
0 56722 5 1 1 56721
0 56723 7 1 2 56720 56722
0 56724 5 1 1 56723
0 56725 7 1 2 61130 78426
0 56726 7 1 2 87414 56725
0 56727 7 1 2 56724 56726
0 56728 5 1 1 56727
0 56729 7 1 2 64431 56728
0 56730 7 1 2 56716 56729
0 56731 5 1 1 56730
0 56732 7 1 2 56714 56731
0 56733 7 1 2 56697 56732
0 56734 5 1 1 56733
0 56735 7 1 2 64649 56734
0 56736 5 1 1 56735
0 56737 7 1 2 56643 56736
0 56738 5 1 1 56737
0 56739 7 1 2 66104 56738
0 56740 5 1 1 56739
0 56741 7 2 2 76722 91486
0 56742 7 1 2 67235 96069
0 56743 5 1 1 56742
0 56744 7 1 2 73520 87945
0 56745 5 1 1 56744
0 56746 7 1 2 56743 56745
0 56747 5 1 1 56746
0 56748 7 1 2 77078 56747
0 56749 5 1 1 56748
0 56750 7 1 2 72487 80900
0 56751 5 1 1 56750
0 56752 7 1 2 78945 87830
0 56753 5 1 1 56752
0 56754 7 1 2 56751 56753
0 56755 7 1 2 56749 56754
0 56756 7 1 2 56740 56755
0 56757 7 1 2 56621 56756
0 56758 5 1 1 56757
0 56759 7 1 2 72750 56758
0 56760 5 1 1 56759
0 56761 7 1 2 79716 70009
0 56762 5 1 1 56761
0 56763 7 1 2 57822 56762
0 56764 5 1 1 56763
0 56765 7 1 2 80718 56764
0 56766 5 1 1 56765
0 56767 7 1 2 92874 56766
0 56768 5 1 1 56767
0 56769 7 1 2 70377 56768
0 56770 5 1 1 56769
0 56771 7 1 2 63430 56770
0 56772 5 1 1 56771
0 56773 7 1 2 66105 93045
0 56774 5 1 1 56773
0 56775 7 1 2 79757 87594
0 56776 5 1 1 56775
0 56777 7 1 2 56774 56776
0 56778 5 1 1 56777
0 56779 7 1 2 60697 56778
0 56780 5 1 1 56779
0 56781 7 1 2 66106 85042
0 56782 5 1 1 56781
0 56783 7 1 2 56780 56782
0 56784 5 1 1 56783
0 56785 7 1 2 61131 56784
0 56786 5 1 1 56785
0 56787 7 1 2 62823 87599
0 56788 5 1 1 56787
0 56789 7 1 2 87574 56788
0 56790 5 1 1 56789
0 56791 7 1 2 66107 56790
0 56792 5 1 1 56791
0 56793 7 2 2 87595 94314
0 56794 5 1 1 96071
0 56795 7 1 2 63431 82261
0 56796 5 1 1 56795
0 56797 7 1 2 56794 56796
0 56798 5 1 1 56797
0 56799 7 1 2 57544 56798
0 56800 5 1 1 56799
0 56801 7 1 2 63432 94439
0 56802 5 1 1 56801
0 56803 7 1 2 56800 56802
0 56804 5 1 1 56803
0 56805 7 1 2 71935 56804
0 56806 5 1 1 56805
0 56807 7 1 2 61497 95846
0 56808 5 1 1 56807
0 56809 7 1 2 74203 56808
0 56810 5 1 1 56809
0 56811 7 1 2 73914 56810
0 56812 5 1 1 56811
0 56813 7 1 2 56806 56812
0 56814 7 1 2 56792 56813
0 56815 7 1 2 56786 56814
0 56816 7 1 2 56772 56815
0 56817 5 1 1 56816
0 56818 7 1 2 59706 56817
0 56819 5 1 1 56818
0 56820 7 1 2 64432 94919
0 56821 5 1 1 56820
0 56822 7 1 2 69759 52761
0 56823 5 1 1 56822
0 56824 7 1 2 58098 56823
0 56825 5 1 1 56824
0 56826 7 1 2 61498 56825
0 56827 7 1 2 56821 56826
0 56828 5 1 1 56827
0 56829 7 1 2 72213 85559
0 56830 7 1 2 56828 56829
0 56831 5 1 1 56830
0 56832 7 1 2 78014 85596
0 56833 5 1 1 56832
0 56834 7 1 2 58697 56833
0 56835 5 1 1 56834
0 56836 7 1 2 75887 6766
0 56837 5 1 1 56836
0 56838 7 1 2 73684 94188
0 56839 7 1 2 56837 56838
0 56840 5 1 1 56839
0 56841 7 1 2 56835 56840
0 56842 5 1 1 56841
0 56843 7 1 2 68545 56842
0 56844 5 1 1 56843
0 56845 7 1 2 67422 77746
0 56846 5 1 1 56845
0 56847 7 1 2 428 56846
0 56848 5 1 1 56847
0 56849 7 1 2 74691 56848
0 56850 5 1 1 56849
0 56851 7 1 2 64650 56850
0 56852 7 1 2 56844 56851
0 56853 7 1 2 56831 56852
0 56854 7 1 2 75342 86735
0 56855 5 1 1 56854
0 56856 7 1 2 38622 56855
0 56857 5 1 1 56856
0 56858 7 1 2 72545 56857
0 56859 5 1 1 56858
0 56860 7 1 2 60698 75304
0 56861 7 1 2 74703 56860
0 56862 5 1 1 56861
0 56863 7 1 2 93737 56862
0 56864 5 1 1 56863
0 56865 7 1 2 71659 56864
0 56866 5 1 1 56865
0 56867 7 1 2 56859 56866
0 56868 5 1 1 56867
0 56869 7 1 2 65105 56868
0 56870 5 1 1 56869
0 56871 7 1 2 80482 86745
0 56872 5 1 1 56871
0 56873 7 1 2 75947 56872
0 56874 5 1 1 56873
0 56875 7 1 2 77521 88482
0 56876 5 1 1 56875
0 56877 7 1 2 69717 82160
0 56878 5 1 1 56877
0 56879 7 1 2 56876 56878
0 56880 5 1 1 56879
0 56881 7 1 2 95335 56880
0 56882 5 1 1 56881
0 56883 7 1 2 56874 56882
0 56884 5 1 1 56883
0 56885 7 1 2 72255 56884
0 56886 5 1 1 56885
0 56887 7 1 2 56870 56886
0 56888 7 1 2 56853 56887
0 56889 7 1 2 67425 55487
0 56890 5 1 1 56889
0 56891 7 1 2 65362 56890
0 56892 5 1 1 56891
0 56893 7 1 2 65756 83090
0 56894 5 1 1 56893
0 56895 7 1 2 56892 56894
0 56896 5 1 1 56895
0 56897 7 1 2 63433 56896
0 56898 5 1 1 56897
0 56899 7 1 2 84199 75305
0 56900 7 1 2 83138 56899
0 56901 5 1 1 56900
0 56902 7 1 2 56898 56901
0 56903 5 1 1 56902
0 56904 7 1 2 66108 56903
0 56905 5 1 1 56904
0 56906 7 1 2 86746 93434
0 56907 5 1 1 56906
0 56908 7 1 2 75793 56907
0 56909 5 1 1 56908
0 56910 7 1 2 77933 94998
0 56911 5 1 1 56910
0 56912 7 1 2 56909 56911
0 56913 5 1 1 56912
0 56914 7 1 2 65757 56913
0 56915 5 1 1 56914
0 56916 7 1 2 76579 96072
0 56917 5 1 1 56916
0 56918 7 1 2 56915 56917
0 56919 5 1 1 56918
0 56920 7 1 2 71936 56919
0 56921 5 1 1 56920
0 56922 7 1 2 56905 56921
0 56923 7 1 2 56888 56922
0 56924 7 1 2 56819 56923
0 56925 5 1 1 56924
0 56926 7 1 2 68290 86795
0 56927 5 1 1 56926
0 56928 7 1 2 71571 56927
0 56929 5 1 1 56928
0 56930 7 1 2 61499 56929
0 56931 5 1 1 56930
0 56932 7 1 2 80827 56931
0 56933 5 1 1 56932
0 56934 7 1 2 83968 56933
0 56935 5 1 1 56934
0 56936 7 1 2 63124 80938
0 56937 5 1 1 56936
0 56938 7 1 2 90379 56937
0 56939 5 1 1 56938
0 56940 7 1 2 61500 56939
0 56941 5 1 1 56940
0 56942 7 1 2 63434 71666
0 56943 5 1 1 56942
0 56944 7 1 2 56941 56943
0 56945 5 1 1 56944
0 56946 7 1 2 85575 56945
0 56947 5 1 1 56946
0 56948 7 1 2 70740 87881
0 56949 5 1 1 56948
0 56950 7 1 2 80828 56949
0 56951 5 1 1 56950
0 56952 7 1 2 62540 56951
0 56953 5 1 1 56952
0 56954 7 1 2 85816 81661
0 56955 5 1 1 56954
0 56956 7 1 2 63435 56955
0 56957 5 1 1 56956
0 56958 7 1 2 56953 56957
0 56959 5 1 1 56958
0 56960 7 1 2 68546 56959
0 56961 5 1 1 56960
0 56962 7 1 2 78620 93215
0 56963 5 1 1 56962
0 56964 7 1 2 85885 56963
0 56965 5 1 1 56964
0 56966 7 1 2 56961 56965
0 56967 7 1 2 56947 56966
0 56968 7 1 2 56935 56967
0 56969 5 1 1 56968
0 56970 7 1 2 60699 56969
0 56971 5 1 1 56970
0 56972 7 1 2 79501 93046
0 56973 5 1 1 56972
0 56974 7 1 2 85477 92782
0 56975 5 1 1 56974
0 56976 7 1 2 81169 56975
0 56977 5 1 1 56976
0 56978 7 1 2 56973 56977
0 56979 5 1 1 56978
0 56980 7 1 2 61132 56979
0 56981 5 1 1 56980
0 56982 7 1 2 85473 76803
0 56983 5 1 1 56982
0 56984 7 1 2 56981 56983
0 56985 5 1 1 56984
0 56986 7 1 2 61501 56985
0 56987 5 1 1 56986
0 56988 7 1 2 83587 90061
0 56989 5 1 1 56988
0 56990 7 1 2 80829 56989
0 56991 5 1 1 56990
0 56992 7 1 2 70235 56991
0 56993 5 1 1 56992
0 56994 7 1 2 84880 34098
0 56995 5 1 1 56994
0 56996 7 1 2 76273 56995
0 56997 5 1 1 56996
0 56998 7 1 2 44777 56997
0 56999 7 1 2 56993 56998
0 57000 5 1 1 56999
0 57001 7 1 2 76969 57000
0 57002 5 1 1 57001
0 57003 7 1 2 74841 86548
0 57004 5 1 1 57003
0 57005 7 1 2 85889 57004
0 57006 5 1 1 57005
0 57007 7 1 2 85576 57006
0 57008 5 1 1 57007
0 57009 7 1 2 72924 28362
0 57010 5 1 1 57009
0 57011 7 1 2 63436 57010
0 57012 5 1 1 57011
0 57013 7 1 2 59952 57012
0 57014 7 1 2 57008 57013
0 57015 7 1 2 57002 57014
0 57016 7 1 2 56987 57015
0 57017 7 1 2 56971 57016
0 57018 5 1 1 57017
0 57019 7 1 2 56925 57018
0 57020 5 1 1 57019
0 57021 7 1 2 85817 14769
0 57022 5 1 1 57021
0 57023 7 1 2 75843 94173
0 57024 5 2 1 57023
0 57025 7 1 2 58698 45190
0 57026 5 1 1 57025
0 57027 7 1 2 79342 57026
0 57028 5 1 1 57027
0 57029 7 1 2 96073 57028
0 57030 5 1 1 57029
0 57031 7 1 2 57022 57030
0 57032 5 1 1 57031
0 57033 7 1 2 77843 95085
0 57034 5 1 1 57033
0 57035 7 1 2 61133 57034
0 57036 5 1 1 57035
0 57037 7 1 2 96074 57036
0 57038 5 1 1 57037
0 57039 7 1 2 87706 57038
0 57040 5 1 1 57039
0 57041 7 1 2 73730 86160
0 57042 5 1 1 57041
0 57043 7 1 2 72062 93532
0 57044 5 1 1 57043
0 57045 7 1 2 72925 15964
0 57046 5 1 1 57045
0 57047 7 1 2 59953 57046
0 57048 7 1 2 57044 57047
0 57049 5 1 1 57048
0 57050 7 1 2 57042 57049
0 57051 5 1 1 57050
0 57052 7 1 2 76236 57051
0 57053 5 1 1 57052
0 57054 7 1 2 85839 90098
0 57055 5 1 1 57054
0 57056 7 1 2 60426 94189
0 57057 7 1 2 96070 57056
0 57058 5 1 1 57057
0 57059 7 1 2 57055 57058
0 57060 5 1 1 57059
0 57061 7 1 2 81090 57060
0 57062 5 1 1 57061
0 57063 7 1 2 60427 70378
0 57064 7 1 2 91487 96059
0 57065 7 1 2 57063 57064
0 57066 5 1 1 57065
0 57067 7 1 2 57062 57066
0 57068 7 1 2 57053 57067
0 57069 7 1 2 57040 57068
0 57070 5 1 1 57069
0 57071 7 1 2 68896 57070
0 57072 5 1 1 57071
0 57073 7 1 2 57032 57072
0 57074 7 1 2 57020 57073
0 57075 5 1 1 57074
0 57076 7 1 2 84225 57075
0 57077 5 1 1 57076
0 57078 7 1 2 56760 57077
0 57079 5 1 1 57078
0 57080 7 1 2 66737 57079
0 57081 5 1 1 57080
0 57082 7 1 2 79611 95812
0 57083 5 1 1 57082
0 57084 7 1 2 59395 83323
0 57085 5 1 1 57084
0 57086 7 1 2 60428 57085
0 57087 5 1 1 57086
0 57088 7 1 2 89071 57087
0 57089 5 1 1 57088
0 57090 7 1 2 65758 57089
0 57091 5 1 1 57090
0 57092 7 1 2 57083 57091
0 57093 5 1 1 57092
0 57094 7 1 2 60700 57093
0 57095 5 1 1 57094
0 57096 7 1 2 74553 93606
0 57097 5 1 1 57096
0 57098 7 1 2 68191 57097
0 57099 5 1 1 57098
0 57100 7 1 2 61134 94131
0 57101 5 1 1 57100
0 57102 7 1 2 60701 94315
0 57103 5 1 1 57102
0 57104 7 1 2 69510 57103
0 57105 5 1 1 57104
0 57106 7 1 2 57545 57105
0 57107 5 1 1 57106
0 57108 7 1 2 59707 6545
0 57109 5 1 1 57108
0 57110 7 1 2 65759 70943
0 57111 7 1 2 86811 57110
0 57112 5 1 1 57111
0 57113 7 1 2 57109 57112
0 57114 7 1 2 93743 57113
0 57115 7 1 2 57107 57114
0 57116 7 1 2 57101 57115
0 57117 7 1 2 57099 57116
0 57118 7 1 2 57095 57117
0 57119 5 1 1 57118
0 57120 7 1 2 64651 57119
0 57121 5 1 1 57120
0 57122 7 2 2 70677 75404
0 57123 7 1 2 95937 96075
0 57124 5 1 1 57123
0 57125 7 1 2 83906 96076
0 57126 5 1 1 57125
0 57127 7 1 2 76495 81308
0 57128 5 1 1 57127
0 57129 7 1 2 94128 57128
0 57130 5 1 1 57129
0 57131 7 1 2 70336 77523
0 57132 7 1 2 57130 57131
0 57133 5 1 1 57132
0 57134 7 1 2 57126 57133
0 57135 5 1 1 57134
0 57136 7 1 2 62541 57135
0 57137 5 1 1 57136
0 57138 7 1 2 57124 57137
0 57139 5 1 1 57138
0 57140 7 1 2 71341 57139
0 57141 5 1 1 57140
0 57142 7 1 2 58099 86166
0 57143 5 1 1 57142
0 57144 7 1 2 60702 57143
0 57145 5 1 1 57144
0 57146 7 1 2 92818 57145
0 57147 5 1 1 57146
0 57148 7 1 2 62542 57147
0 57149 5 1 1 57148
0 57150 7 1 2 60703 95188
0 57151 5 1 1 57150
0 57152 7 1 2 67416 57151
0 57153 7 1 2 57149 57152
0 57154 5 1 1 57153
0 57155 7 1 2 90796 57154
0 57156 5 1 1 57155
0 57157 7 1 2 72160 93596
0 57158 5 1 1 57157
0 57159 7 1 2 85490 93603
0 57160 7 1 2 57158 57159
0 57161 5 1 1 57160
0 57162 7 1 2 57156 57161
0 57163 7 1 2 57141 57162
0 57164 7 1 2 57121 57163
0 57165 5 1 1 57164
0 57166 7 1 2 66109 57165
0 57167 5 1 1 57166
0 57168 7 1 2 30263 93216
0 57169 5 1 1 57168
0 57170 7 1 2 88777 57169
0 57171 5 1 1 57170
0 57172 7 1 2 93615 57171
0 57173 5 1 1 57172
0 57174 7 1 2 84551 57173
0 57175 5 1 1 57174
0 57176 7 1 2 81457 95007
0 57177 5 1 1 57176
0 57178 7 1 2 34580 57177
0 57179 7 1 2 57175 57178
0 57180 5 1 1 57179
0 57181 7 1 2 61135 57180
0 57182 5 1 1 57181
0 57183 7 1 2 80830 57182
0 57184 5 1 1 57183
0 57185 7 1 2 59954 57184
0 57186 5 1 1 57185
0 57187 7 1 2 85705 89077
0 57188 5 1 1 57187
0 57189 7 1 2 78003 81458
0 57190 5 1 1 57189
0 57191 7 1 2 57188 57190
0 57192 5 1 1 57191
0 57193 7 1 2 60704 57192
0 57194 5 1 1 57193
0 57195 7 1 2 73221 83896
0 57196 7 1 2 93541 57195
0 57197 5 1 1 57196
0 57198 7 1 2 84282 57197
0 57199 5 1 1 57198
0 57200 7 1 2 60429 57199
0 57201 5 1 1 57200
0 57202 7 1 2 84279 79612
0 57203 5 1 1 57202
0 57204 7 1 2 78015 57203
0 57205 7 1 2 57201 57204
0 57206 5 1 1 57205
0 57207 7 1 2 68192 57206
0 57208 5 1 1 57207
0 57209 7 1 2 4256 95805
0 57210 5 1 1 57209
0 57211 7 1 2 93604 57210
0 57212 5 1 1 57211
0 57213 7 1 2 85706 86878
0 57214 5 1 1 57213
0 57215 7 1 2 85430 57214
0 57216 7 1 2 57212 57215
0 57217 7 1 2 57208 57216
0 57218 7 1 2 57194 57217
0 57219 5 1 1 57218
0 57220 7 1 2 61502 57219
0 57221 5 1 1 57220
0 57222 7 1 2 57186 57221
0 57223 5 1 1 57222
0 57224 7 1 2 7730 95732
0 57225 5 1 1 57224
0 57226 7 1 2 58375 90398
0 57227 5 1 1 57226
0 57228 7 1 2 78249 88643
0 57229 5 1 1 57228
0 57230 7 1 2 59708 57229
0 57231 5 1 1 57230
0 57232 7 1 2 75278 57231
0 57233 7 1 2 57227 57232
0 57234 5 1 1 57233
0 57235 7 1 2 57225 57234
0 57236 5 1 1 57235
0 57237 7 1 2 58100 36371
0 57238 5 1 1 57237
0 57239 7 1 2 64652 81104
0 57240 7 1 2 57238 57239
0 57241 7 1 2 57236 57240
0 57242 5 1 1 57241
0 57243 7 1 2 57223 57242
0 57244 5 1 1 57243
0 57245 7 1 2 57167 57244
0 57246 5 1 1 57245
0 57247 7 1 2 72690 57246
0 57248 5 1 1 57247
0 57249 7 1 2 61759 57248
0 57250 7 1 2 57081 57249
0 57251 5 1 1 57250
0 57252 7 1 2 56515 57251
0 57253 5 1 1 57252
0 57254 7 1 2 66653 69586
0 57255 7 1 2 93152 57254
0 57256 5 1 1 57255
0 57257 7 1 2 57253 57256
0 57258 5 1 1 57257
0 57259 7 1 2 66951 57258
0 57260 5 1 1 57259
0 57261 7 1 2 56135 57260
0 57262 7 1 2 55185 57261
0 57263 7 1 2 53203 57262
0 57264 7 1 2 52438 57263
0 57265 5 1 1 57264
0 57266 7 1 2 61873 88314
0 57267 7 1 2 57265 57266
0 57268 5 1 1 57267
0 57269 7 1 2 50872 57268
0 57270 7 1 2 41474 57269
0 57271 5 1 1 57270
0 57272 7 1 2 62143 57271
0 57273 5 1 1 57272
0 57274 7 1 2 32684 57273
3 129999 5 0 1 57274
