1 0 0 2 0
2 49 1 0
2 734 1 0
1 1 0 2 0
2 735 1 1
2 736 1 1
1 2 0 2 0
2 737 1 2
2 738 1 2
1 3 0 2 0
2 739 1 3
2 740 1 3
1 4 0 2 0
2 741 1 4
2 742 1 4
1 5 0 2 0
2 743 1 5
2 744 1 5
1 6 0 2 0
2 745 1 6
2 746 1 6
1 7 0 2 0
2 747 1 7
2 748 1 7
1 8 0 2 0
2 749 1 8
2 750 1 8
1 9 0 2 0
2 751 1 9
2 752 1 9
1 10 0 2 0
2 753 1 10
2 754 1 10
1 11 0 2 0
2 755 1 11
2 756 1 11
1 12 0 2 0
2 757 1 12
2 758 1 12
1 13 0 2 0
2 759 1 13
2 760 1 13
1 14 0 2 0
2 761 1 14
2 762 1 14
1 15 0 2 0
2 763 1 15
2 764 1 15
1 16 0 2 0
2 765 1 16
2 766 1 16
1 17 0 2 0
2 767 1 17
2 768 1 17
1 18 0 2 0
2 769 1 18
2 770 1 18
1 19 0 2 0
2 771 1 19
2 772 1 19
1 20 0 2 0
2 773 1 20
2 774 1 20
1 21 0 2 0
2 775 1 21
2 776 1 21
1 22 0 2 0
2 777 1 22
2 778 1 22
1 23 0 2 0
2 779 1 23
2 780 1 23
1 24 0 2 0
2 781 1 24
2 782 1 24
1 25 0 2 0
2 783 1 25
2 784 1 25
1 26 0 2 0
2 785 1 26
2 786 1 26
1 27 0 2 0
2 787 1 27
2 788 1 27
1 28 0 2 0
2 789 1 28
2 790 1 28
1 29 0 2 0
2 791 1 29
2 792 1 29
1 30 0 2 0
2 793 1 30
2 794 1 30
1 31 0 2 0
2 795 1 31
2 796 1 31
1 32 0 2 0
2 797 1 32
2 798 1 32
1 33 0 2 0
2 799 1 33
2 800 1 33
1 34 0 3 0
2 801 1 34
2 802 1 34
2 803 1 34
1 35 0 2 0
2 804 1 35
2 805 1 35
1 36 0 2 0
2 806 1 36
2 807 1 36
1 37 0 2 0
2 808 1 37
2 809 1 37
1 38 0 2 0
2 810 1 38
2 811 1 38
1 39 0 2 0
2 812 1 39
2 813 1 39
1 40 0 2 0
2 814 1 40
2 815 1 40
1 41 0 2 0
2 816 1 41
2 817 1 41
1 42 0 2 0
2 818 1 42
2 819 1 42
1 43 0 2 0
2 820 1 43
2 821 1 43
1 44 0 2 0
2 822 1 44
2 823 1 44
1 45 0 2 0
2 824 1 45
2 825 1 45
1 46 0 2 0
2 826 1 46
2 827 1 46
1 47 0 2 0
2 828 1 47
2 829 1 47
1 48 0 2 0
2 830 1 48
2 831 1 48
2 832 1 69
2 833 1 69
2 834 1 70
2 835 1 70
2 836 1 71
2 837 1 71
2 838 1 72
2 839 1 72
2 840 1 73
2 841 1 73
2 842 1 74
2 843 1 74
2 844 1 75
2 845 1 75
2 846 1 76
2 847 1 76
2 848 1 77
2 849 1 77
2 850 1 78
2 851 1 78
2 852 1 79
2 853 1 79
2 854 1 80
2 855 1 80
2 856 1 81
2 857 1 81
2 858 1 100
2 859 1 100
2 860 1 102
2 861 1 102
2 862 1 104
2 863 1 104
2 864 1 106
2 865 1 106
2 866 1 107
2 867 1 107
2 868 1 108
2 869 1 108
2 870 1 108
2 871 1 111
2 872 1 111
2 873 1 112
2 874 1 112
2 875 1 115
2 876 1 115
2 877 1 118
2 878 1 118
2 879 1 120
2 880 1 120
2 881 1 123
2 882 1 123
2 883 1 126
2 884 1 126
2 885 1 128
2 886 1 128
2 887 1 131
2 888 1 131
2 889 1 134
2 890 1 134
2 891 1 136
2 892 1 136
2 893 1 139
2 894 1 139
2 895 1 142
2 896 1 142
2 897 1 144
2 898 1 144
2 899 1 147
2 900 1 147
2 901 1 150
2 902 1 150
2 903 1 152
2 904 1 152
2 905 1 155
2 906 1 155
2 907 1 158
2 908 1 158
2 909 1 160
2 910 1 160
2 911 1 163
2 912 1 163
2 913 1 166
2 914 1 166
2 915 1 168
2 916 1 168
2 917 1 171
2 918 1 171
2 919 1 174
2 920 1 174
2 921 1 176
2 922 1 176
2 923 1 179
2 924 1 179
2 925 1 182
2 926 1 182
2 927 1 184
2 928 1 184
2 929 1 187
2 930 1 187
2 931 1 190
2 932 1 190
2 933 1 192
2 934 1 192
2 935 1 195
2 936 1 195
2 937 1 198
2 938 1 198
2 939 1 200
2 940 1 200
2 941 1 203
2 942 1 203
2 943 1 206
2 944 1 206
2 945 1 208
2 946 1 208
2 947 1 211
2 948 1 211
2 949 1 214
2 950 1 214
2 951 1 216
2 952 1 216
2 953 1 219
2 954 1 219
2 955 1 221
2 956 1 221
2 957 1 222
2 958 1 222
2 959 1 223
2 960 1 223
2 961 1 224
2 962 1 224
2 963 1 225
2 964 1 225
2 965 1 231
2 966 1 231
2 967 1 233
2 968 1 233
2 969 1 234
2 970 1 234
2 971 1 234
2 972 1 235
2 973 1 235
2 974 1 241
2 975 1 241
2 976 1 244
2 977 1 244
2 978 1 244
2 979 1 244
2 980 1 246
2 981 1 246
2 982 1 246
2 983 1 247
2 984 1 247
2 985 1 253
2 986 1 253
2 987 1 256
2 988 1 256
2 989 1 256
2 990 1 256
2 991 1 257
2 992 1 257
2 993 1 263
2 994 1 263
2 995 1 266
2 996 1 266
2 997 1 266
2 998 1 267
2 999 1 267
2 1000 1 273
2 1001 1 273
2 1002 1 276
2 1003 1 276
2 1004 1 276
2 1005 1 278
2 1006 1 278
2 1007 1 278
2 1008 1 279
2 1009 1 279
2 1010 1 285
2 1011 1 285
2 1012 1 288
2 1013 1 288
2 1014 1 288
2 1015 1 288
2 1016 1 290
2 1017 1 290
2 1018 1 290
2 1019 1 291
2 1020 1 291
2 1021 1 297
2 1022 1 297
2 1023 1 300
2 1024 1 300
2 1025 1 300
2 1026 1 300
2 1027 1 301
2 1028 1 301
2 1029 1 307
2 1030 1 307
2 1031 1 310
2 1032 1 310
2 1033 1 310
2 1034 1 312
2 1035 1 312
2 1036 1 312
2 1037 1 313
2 1038 1 313
2 1039 1 319
2 1040 1 319
2 1041 1 322
2 1042 1 322
2 1043 1 322
2 1044 1 323
2 1045 1 323
2 1046 1 324
2 1047 1 324
2 1048 1 324
2 1049 1 325
2 1050 1 325
2 1051 1 331
2 1052 1 331
2 1053 1 334
2 1054 1 334
2 1055 1 334
2 1056 1 334
2 1057 1 336
2 1058 1 336
2 1059 1 336
2 1060 1 337
2 1061 1 337
2 1062 1 343
2 1063 1 343
2 1064 1 346
2 1065 1 346
2 1066 1 346
2 1067 1 346
2 1068 1 348
2 1069 1 348
2 1070 1 348
2 1071 1 349
2 1072 1 349
2 1073 1 355
2 1074 1 355
2 1075 1 358
2 1076 1 358
2 1077 1 358
2 1078 1 358
2 1079 1 359
2 1080 1 359
2 1081 1 365
2 1082 1 365
2 1083 1 368
2 1084 1 368
2 1085 1 368
2 1086 1 368
2 1087 1 370
2 1088 1 370
2 1089 1 370
2 1090 1 371
2 1091 1 371
2 1092 1 377
2 1093 1 377
2 1094 1 380
2 1095 1 380
2 1096 1 380
2 1097 1 380
2 1098 1 382
2 1099 1 382
2 1100 1 382
2 1101 1 383
2 1102 1 383
2 1103 1 389
2 1104 1 389
2 1105 1 392
2 1106 1 392
2 1107 1 394
2 1108 1 394
2 1109 1 397
2 1110 1 397
2 1111 1 403
2 1112 1 403
2 1113 1 405
2 1114 1 405
2 1115 1 408
2 1116 1 408
2 1117 1 412
2 1118 1 412
2 1119 1 416
2 1120 1 416
2 1121 1 416
2 1122 1 416
2 1123 1 418
2 1124 1 418
2 1125 1 420
2 1126 1 420
2 1127 1 421
2 1128 1 421
2 1129 1 425
2 1130 1 425
2 1131 1 428
2 1132 1 428
2 1133 1 429
2 1134 1 429
2 1135 1 432
2 1136 1 432
2 1137 1 436
2 1138 1 436
2 1139 1 436
2 1140 1 436
2 1141 1 438
2 1142 1 438
2 1143 1 440
2 1144 1 440
2 1145 1 441
2 1146 1 441
2 1147 1 444
2 1148 1 444
2 1149 1 446
2 1150 1 446
2 1151 1 450
2 1152 1 450
2 1153 1 451
2 1154 1 451
2 1155 1 451
2 1156 1 453
2 1157 1 453
2 1158 1 455
2 1159 1 455
2 1160 1 455
2 1161 1 455
2 1162 1 462
2 1163 1 462
2 1164 1 463
2 1165 1 463
2 1166 1 464
2 1167 1 464
2 1168 1 464
2 1169 1 467
2 1170 1 467
2 1171 1 471
2 1172 1 471
2 1173 1 475
2 1174 1 475
2 1175 1 481
2 1176 1 481
2 1177 1 481
2 1178 1 487
2 1179 1 487
2 1180 1 487
2 1181 1 493
2 1182 1 493
2 1183 1 494
2 1184 1 494
2 1185 1 497
2 1186 1 497
2 1187 1 497
2 1188 1 498
2 1189 1 498
2 1190 1 503
2 1191 1 503
2 1192 1 504
2 1193 1 504
2 1194 1 508
2 1195 1 508
2 1196 1 511
2 1197 1 511
2 1198 1 512
2 1199 1 512
2 1200 1 512
2 1201 1 519
2 1202 1 519
2 1203 1 520
2 1204 1 520
2 1205 1 523
2 1206 1 523
2 1207 1 524
2 1208 1 524
2 1209 1 527
2 1210 1 527
2 1211 1 528
2 1212 1 528
2 1213 1 534
2 1214 1 534
2 1215 1 537
2 1216 1 537
2 1217 1 538
2 1218 1 538
2 1219 1 547
2 1220 1 547
2 1221 1 547
2 1222 1 549
2 1223 1 549
2 1224 1 550
2 1225 1 550
2 1226 1 590
2 1227 1 590
2 1228 1 592
2 1229 1 592
2 1230 1 594
2 1231 1 594
2 1232 1 598
2 1233 1 598
2 1234 1 602
2 1235 1 602
2 1236 1 607
2 1237 1 607
2 1238 1 610
2 1239 1 610
2 1240 1 611
2 1241 1 611
2 1242 1 615
2 1243 1 615
2 1244 1 618
2 1245 1 618
2 1246 1 622
2 1247 1 622
2 1248 1 623
2 1249 1 623
2 1250 1 626
2 1251 1 626
2 1252 1 627
2 1253 1 627
2 1254 1 630
2 1255 1 630
2 1256 1 631
2 1257 1 631
2 1258 1 634
2 1259 1 634
2 1260 1 635
2 1261 1 635
2 1262 1 638
2 1263 1 638
2 1264 1 638
0 50 5 1 1 49
0 51 5 1 1 735
0 52 5 1 1 737
0 53 5 1 1 739
0 54 5 1 1 741
0 55 5 1 1 743
0 56 5 1 1 745
0 57 5 1 1 747
0 58 5 1 1 749
0 59 5 1 1 751
0 60 5 1 1 753
0 61 5 1 1 755
0 62 5 1 1 757
0 63 5 1 1 759
0 64 5 1 1 761
0 65 5 1 1 763
0 66 5 1 1 765
0 67 5 1 1 767
0 68 5 1 1 769
0 69 5 2 1 771
0 70 5 2 1 773
0 71 5 2 1 775
0 72 5 2 1 777
0 73 5 2 1 779
0 74 5 2 1 781
0 75 5 2 1 783
0 76 5 2 1 785
0 77 5 2 1 787
0 78 5 2 1 789
0 79 5 2 1 791
0 80 5 2 1 793
0 81 5 2 1 795
0 82 5 1 1 797
0 83 5 1 1 799
0 84 5 1 1 801
0 85 5 1 1 804
0 86 5 1 1 806
0 87 5 1 1 808
0 88 5 1 1 810
0 89 5 1 1 812
0 90 5 1 1 814
0 91 5 1 1 816
0 92 5 1 1 818
0 93 5 1 1 820
0 94 5 1 1 822
0 95 5 1 1 824
0 96 5 1 1 826
0 97 5 1 1 828
0 98 5 1 1 830
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 738 770
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 736 768
0 106 5 2 1 105
0 107 7 2 2 734 766
0 108 5 3 1 866
0 109 7 1 2 864 868
0 110 5 1 1 109
0 111 7 2 2 862 110
0 112 5 2 1 871
0 113 7 1 2 860 873
0 114 5 1 1 113
0 115 7 2 2 858 114
0 116 5 1 1 875
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 740 876
0 120 5 2 1 119
0 121 7 1 2 832 879
0 122 5 1 1 121
0 123 7 2 2 877 122
0 124 5 1 1 881
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 742 882
0 128 5 2 1 127
0 129 7 1 2 834 885
0 130 5 1 1 129
0 131 7 2 2 883 130
0 132 5 1 1 887
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 744 888
0 136 5 2 1 135
0 137 7 1 2 836 891
0 138 5 1 1 137
0 139 7 2 2 889 138
0 140 5 1 1 893
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 746 894
0 144 5 2 1 143
0 145 7 1 2 838 897
0 146 5 1 1 145
0 147 7 2 2 895 146
0 148 5 1 1 899
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 748 900
0 152 5 2 1 151
0 153 7 1 2 840 903
0 154 5 1 1 153
0 155 7 2 2 901 154
0 156 5 1 1 905
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 750 906
0 160 5 2 1 159
0 161 7 1 2 842 909
0 162 5 1 1 161
0 163 7 2 2 907 162
0 164 5 1 1 911
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 752 912
0 168 5 2 1 167
0 169 7 1 2 844 915
0 170 5 1 1 169
0 171 7 2 2 913 170
0 172 5 1 1 917
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 754 918
0 176 5 2 1 175
0 177 7 1 2 846 921
0 178 5 1 1 177
0 179 7 2 2 919 178
0 180 5 1 1 923
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 756 924
0 184 5 2 1 183
0 185 7 1 2 848 927
0 186 5 1 1 185
0 187 7 2 2 925 186
0 188 5 1 1 929
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 758 930
0 192 5 2 1 191
0 193 7 1 2 850 933
0 194 5 1 1 193
0 195 7 2 2 931 194
0 196 5 1 1 935
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 760 936
0 200 5 2 1 199
0 201 7 1 2 852 939
0 202 5 1 1 201
0 203 7 2 2 937 202
0 204 5 1 1 941
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 762 942
0 208 5 2 1 207
0 209 7 1 2 854 945
0 210 5 1 1 209
0 211 7 2 2 943 210
0 212 5 1 1 947
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 764 948
0 216 5 2 1 215
0 217 7 1 2 856 951
0 218 5 1 1 217
0 219 7 2 2 949 218
0 220 5 1 1 953
0 221 7 2 2 831 220
0 222 5 2 1 955
0 223 7 2 2 98 954
0 224 5 2 1 959
0 225 7 2 2 950 952
0 226 5 1 1 963
0 227 7 1 2 796 226
0 228 5 1 1 227
0 229 7 1 2 857 964
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 965
0 233 7 2 2 829 966
0 234 5 3 1 967
0 235 7 2 2 944 946
0 236 5 1 1 972
0 237 7 1 2 794 973
0 238 5 1 1 237
0 239 7 1 2 855 236
0 240 5 1 1 239
0 241 7 2 2 238 240
0 242 5 1 1 974
0 243 7 1 2 827 242
0 244 5 4 1 243
0 245 7 1 2 96 975
0 246 5 3 1 245
0 247 7 2 2 938 940
0 248 5 1 1 983
0 249 7 1 2 792 984
0 250 5 1 1 249
0 251 7 1 2 853 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 985
0 255 7 1 2 95 986
0 256 5 4 1 255
0 257 7 2 2 932 934
0 258 5 1 1 991
0 259 7 1 2 790 992
0 260 5 1 1 259
0 261 7 1 2 851 258
0 262 5 1 1 261
0 263 7 2 2 260 262
0 264 5 1 1 993
0 265 7 1 2 94 994
0 266 5 3 1 265
0 267 7 2 2 926 928
0 268 5 1 1 998
0 269 7 1 2 788 999
0 270 5 1 1 269
0 271 7 1 2 849 268
0 272 5 1 1 271
0 273 7 2 2 270 272
0 274 5 1 1 1000
0 275 7 1 2 821 274
0 276 5 3 1 275
0 277 7 1 2 93 1001
0 278 5 3 1 277
0 279 7 2 2 920 922
0 280 5 1 1 1008
0 281 7 1 2 786 1009
0 282 5 1 1 281
0 283 7 1 2 847 280
0 284 5 1 1 283
0 285 7 2 2 282 284
0 286 5 1 1 1010
0 287 7 1 2 819 286
0 288 5 4 1 287
0 289 7 1 2 92 1011
0 290 5 3 1 289
0 291 7 2 2 914 916
0 292 5 1 1 1019
0 293 7 1 2 784 1020
0 294 5 1 1 293
0 295 7 1 2 845 292
0 296 5 1 1 295
0 297 7 2 2 294 296
0 298 5 1 1 1021
0 299 7 1 2 817 298
0 300 5 4 1 299
0 301 7 2 2 908 910
0 302 5 1 1 1027
0 303 7 1 2 782 1028
0 304 5 1 1 303
0 305 7 1 2 843 302
0 306 5 1 1 305
0 307 7 2 2 304 306
0 308 5 1 1 1029
0 309 7 1 2 815 308
0 310 5 3 1 309
0 311 7 1 2 90 1030
0 312 5 3 1 311
0 313 7 2 2 902 904
0 314 5 1 1 1037
0 315 7 1 2 780 1038
0 316 5 1 1 315
0 317 7 1 2 841 314
0 318 5 1 1 317
0 319 7 2 2 316 318
0 320 5 1 1 1039
0 321 7 1 2 813 320
0 322 5 3 1 321
0 323 7 2 2 89 1040
0 324 5 3 1 1044
0 325 7 2 2 896 898
0 326 5 1 1 1049
0 327 7 1 2 778 1050
0 328 5 1 1 327
0 329 7 1 2 839 326
0 330 5 1 1 329
0 331 7 2 2 328 330
0 332 5 1 1 1051
0 333 7 1 2 811 332
0 334 5 4 1 333
0 335 7 1 2 88 1052
0 336 5 3 1 335
0 337 7 2 2 890 892
0 338 5 1 1 1060
0 339 7 1 2 776 1061
0 340 5 1 1 339
0 341 7 1 2 837 338
0 342 5 1 1 341
0 343 7 2 2 340 342
0 344 5 1 1 1062
0 345 7 1 2 809 344
0 346 5 4 1 345
0 347 7 1 2 87 1063
0 348 5 3 1 347
0 349 7 2 2 884 886
0 350 5 1 1 1071
0 351 7 1 2 774 1072
0 352 5 1 1 351
0 353 7 1 2 835 350
0 354 5 1 1 353
0 355 7 2 2 352 354
0 356 5 1 1 1073
0 357 7 1 2 807 356
0 358 5 4 1 357
0 359 7 2 2 878 880
0 360 5 1 1 1079
0 361 7 1 2 772 1080
0 362 5 1 1 361
0 363 7 1 2 833 360
0 364 5 1 1 363
0 365 7 2 2 362 364
0 366 5 1 1 1081
0 367 7 1 2 85 1082
0 368 5 4 1 367
0 369 7 1 2 805 366
0 370 5 3 1 369
0 371 7 2 2 859 861
0 372 5 1 1 1090
0 373 7 1 2 872 372
0 374 5 1 1 373
0 375 7 1 2 874 1091
0 376 5 1 1 375
0 377 7 2 2 374 376
0 378 5 1 1 1092
0 379 7 1 2 84 378
0 380 5 4 1 379
0 381 7 1 2 802 1093
0 382 5 3 1 381
0 383 7 2 2 863 865
0 384 5 1 1 1101
0 385 7 1 2 867 384
0 386 5 1 1 385
0 387 7 1 2 869 1102
0 388 5 1 1 387
0 389 7 2 2 386 388
0 390 5 1 1 1103
0 391 7 1 2 83 390
0 392 5 2 1 391
0 393 7 1 2 800 1104
0 394 5 2 1 393
0 395 7 1 2 50 66
0 396 5 1 1 395
0 397 7 2 2 870 396
0 398 5 1 1 1109
0 399 7 1 2 798 398
0 400 5 1 1 399
0 401 7 1 2 1107 400
0 402 5 1 1 401
0 403 7 2 2 1105 402
0 404 5 1 1 1111
0 405 7 2 2 1098 404
0 406 5 1 1 1113
0 407 7 1 2 1094 406
0 408 5 2 1 407
0 409 7 1 2 1087 1115
0 410 5 1 1 409
0 411 7 1 2 1083 410
0 412 5 2 1 411
0 413 7 1 2 1075 1117
0 414 5 1 1 413
0 415 7 1 2 86 1074
0 416 5 4 1 415
0 417 7 1 2 414 1119
0 418 7 2 2 1068 417
0 419 5 1 1 1123
0 420 7 2 2 1064 419
0 421 5 2 1 1125
0 422 7 1 2 1057 1127
0 423 5 1 1 422
0 424 7 1 2 1053 423
0 425 5 2 1 424
0 426 7 1 2 1046 1129
0 427 5 1 1 426
0 428 7 2 2 1041 427
0 429 5 2 1 1131
0 430 7 1 2 1034 1133
0 431 5 1 1 430
0 432 7 2 2 1031 431
0 433 7 1 2 1023 1135
0 434 5 1 1 433
0 435 7 1 2 91 1022
0 436 5 4 1 435
0 437 7 1 2 434 1137
0 438 7 2 2 1016 437
0 439 5 1 1 1141
0 440 7 2 2 1012 439
0 441 5 2 1 1143
0 442 7 1 2 1005 1145
0 443 5 1 1 442
0 444 7 2 2 1002 443
0 445 5 1 1 1147
0 446 7 2 2 995 445
0 447 5 1 1 1149
0 448 7 1 2 987 1150
0 449 5 1 1 448
0 450 7 2 2 823 264
0 451 5 3 1 1151
0 452 7 1 2 988 1152
0 453 5 2 1 452
0 454 7 1 2 825 254
0 455 5 4 1 454
0 456 7 1 2 1156 1158
0 457 7 1 2 449 456
0 458 5 1 1 457
0 459 7 1 2 980 458
0 460 5 1 1 459
0 461 7 1 2 976 460
0 462 5 2 1 461
0 463 7 2 2 97 232
0 464 5 3 1 1164
0 465 7 1 2 1162 1166
0 466 5 1 1 465
0 467 7 2 2 969 466
0 468 5 1 1 1169
0 469 7 1 2 961 468
0 470 5 1 1 469
0 471 7 2 2 957 470
0 472 5 1 1 1171
0 473 7 1 2 960 1170
0 474 5 1 1 473
0 475 7 2 2 1167 970
0 476 5 1 1 1173
0 477 7 1 2 977 476
0 478 5 1 1 477
0 479 7 1 2 1163 1174
0 480 5 1 1 479
0 481 7 3 2 978 981
0 482 5 1 1 1175
0 483 7 1 2 1157 1176
0 484 5 1 1 483
0 485 7 1 2 1159 484
0 486 5 1 1 485
0 487 7 3 2 989 1160
0 488 5 1 1 1178
0 489 7 1 2 447 1179
0 490 5 1 1 489
0 491 7 1 2 1153 490
0 492 5 1 1 491
0 493 7 2 2 1154 996
0 494 5 2 1 1181
0 495 7 1 2 1148 1183
0 496 5 1 1 495
0 497 7 3 2 1003 1006
0 498 5 2 1 1185
0 499 7 1 2 1144 1186
0 500 5 1 1 499
0 501 7 1 2 1013 1142
0 502 5 1 1 501
0 503 7 2 2 1014 1017
0 504 5 2 1 1190
0 505 7 1 2 1024 1192
0 506 5 1 1 505
0 507 7 1 2 1025 1138
0 508 5 2 1 507
0 509 7 1 2 1136 1194
0 510 5 1 1 509
0 511 7 2 2 1032 1035
0 512 5 3 1 1196
0 513 7 1 2 1045 1198
0 514 5 1 1 513
0 515 7 1 2 1132 514
0 516 5 1 1 515
0 517 7 1 2 1134 1199
0 518 5 1 1 517
0 519 7 2 2 1042 1047
0 520 5 2 1 1201
0 521 7 1 2 1130 1203
0 522 5 1 1 521
0 523 7 2 2 1054 1058
0 524 5 2 1 1205
0 525 7 1 2 1126 1206
0 526 5 1 1 525
0 527 7 2 2 1065 1069
0 528 5 2 1 1209
0 529 7 1 2 1076 1211
0 530 5 1 1 529
0 531 7 1 2 1066 1124
0 532 5 1 1 531
0 533 7 1 2 1077 1120
0 534 5 2 1 533
0 535 7 1 2 1118 1213
0 536 5 1 1 535
0 537 7 2 2 1084 1088
0 538 5 2 1 1215
0 539 7 1 2 1116 1217
0 540 5 1 1 539
0 541 7 1 2 803 1216
0 542 5 1 1 541
0 543 7 1 2 82 1110
0 544 5 1 1 543
0 545 7 1 2 1106 544
0 546 5 1 1 545
0 547 7 3 2 1108 546
0 548 5 1 1 1219
0 549 7 2 2 1095 1099
0 550 5 2 1 1222
0 551 7 1 2 548 1224
0 552 7 1 2 542 551
0 553 5 1 1 552
0 554 7 1 2 1096 1114
0 555 5 1 1 554
0 556 7 1 2 553 555
0 557 5 1 1 556
0 558 7 1 2 540 557
0 559 7 1 2 536 558
0 560 7 1 2 532 559
0 561 7 1 2 530 560
0 562 5 1 1 561
0 563 7 1 2 1128 1207
0 564 5 1 1 563
0 565 7 1 2 562 564
0 566 7 1 2 526 565
0 567 7 1 2 522 566
0 568 7 1 2 518 567
0 569 7 1 2 516 568
0 570 5 1 1 569
0 571 7 1 2 510 570
0 572 7 1 2 506 571
0 573 7 1 2 502 572
0 574 5 1 1 573
0 575 7 1 2 1146 1188
0 576 5 1 1 575
0 577 7 1 2 574 576
0 578 7 1 2 500 577
0 579 5 1 1 578
0 580 7 1 2 496 579
0 581 7 1 2 492 580
0 582 7 1 2 486 581
0 583 7 1 2 480 582
0 584 7 1 2 478 583
0 585 7 1 2 474 584
0 586 7 1 2 1172 585
0 587 5 1 1 586
0 588 7 1 2 1100 1220
0 589 5 1 1 588
0 590 7 2 2 1097 589
0 591 5 1 1 1226
0 592 7 2 2 1089 591
0 593 5 1 1 1228
0 594 7 2 2 1085 593
0 595 5 1 1 1230
0 596 7 1 2 1078 595
0 597 5 1 1 596
0 598 7 2 2 1121 597
0 599 5 1 1 1232
0 600 7 1 2 1070 1233
0 601 5 1 1 600
0 602 7 2 2 1067 601
0 603 5 1 1 1234
0 604 7 1 2 1059 603
0 605 5 1 1 604
0 606 7 1 2 1055 605
0 607 5 2 1 606
0 608 7 1 2 1048 1236
0 609 5 1 1 608
0 610 7 2 2 1043 609
0 611 5 2 1 1238
0 612 7 1 2 1036 1240
0 613 5 1 1 612
0 614 7 1 2 1033 613
0 615 5 2 1 614
0 616 7 1 2 1139 1242
0 617 5 1 1 616
0 618 7 2 2 1026 617
0 619 5 1 1 1244
0 620 7 1 2 1018 619
0 621 5 1 1 620
0 622 7 2 2 1015 621
0 623 5 2 1 1246
0 624 7 1 2 1007 1248
0 625 5 1 1 624
0 626 7 2 2 1004 625
0 627 5 2 1 1250
0 628 7 1 2 997 1252
0 629 5 1 1 628
0 630 7 2 2 1155 629
0 631 5 2 1 1254
0 632 7 1 2 990 1256
0 633 5 1 1 632
0 634 7 2 2 1161 633
0 635 5 2 1 1258
0 636 7 1 2 982 1260
0 637 5 1 1 636
0 638 7 3 2 979 637
0 639 5 1 1 1262
0 640 7 1 2 971 1263
0 641 5 1 1 640
0 642 7 1 2 958 641
0 643 5 1 1 642
0 644 7 1 2 1168 643
0 645 5 1 1 644
0 646 7 1 2 968 639
0 647 5 1 1 646
0 648 7 1 2 956 1264
0 649 5 1 1 648
0 650 7 1 2 1165 649
0 651 5 1 1 650
0 652 7 1 2 1180 1257
0 653 5 1 1 652
0 654 7 1 2 488 1255
0 655 5 1 1 654
0 656 7 1 2 653 655
0 657 5 1 1 656
0 658 7 1 2 1191 1245
0 659 5 1 1 658
0 660 7 1 2 1140 1193
0 661 5 1 1 660
0 662 7 1 2 1195 1243
0 663 5 1 1 662
0 664 7 1 2 1197 1241
0 665 5 1 1 664
0 666 7 1 2 1200 1239
0 667 5 1 1 666
0 668 7 1 2 1056 1204
0 669 5 1 1 668
0 670 7 1 2 1202 1237
0 671 5 1 1 670
0 672 7 1 2 1208 1235
0 673 5 1 1 672
0 674 7 1 2 1210 599
0 675 5 1 1 674
0 676 7 1 2 1122 1212
0 677 5 1 1 676
0 678 7 1 2 1214 1231
0 679 5 1 1 678
0 680 7 1 2 1218 1227
0 681 5 1 1 680
0 682 7 1 2 1086 1229
0 683 5 1 1 682
0 684 7 1 2 1221 1223
0 685 5 1 1 684
0 686 7 1 2 1112 1225
0 687 5 1 1 686
0 688 7 1 2 685 687
0 689 7 1 2 683 688
0 690 7 1 2 681 689
0 691 7 1 2 679 690
0 692 7 1 2 677 691
0 693 7 1 2 675 692
0 694 5 1 1 693
0 695 7 1 2 673 694
0 696 7 1 2 671 695
0 697 7 1 2 669 696
0 698 7 1 2 667 697
0 699 7 1 2 665 698
0 700 5 1 1 699
0 701 7 1 2 663 700
0 702 7 1 2 661 701
0 703 7 1 2 659 702
0 704 5 1 1 703
0 705 7 1 2 1189 1249
0 706 5 1 1 705
0 707 7 1 2 1187 1247
0 708 5 1 1 707
0 709 7 1 2 706 708
0 710 5 1 1 709
0 711 7 1 2 704 710
0 712 5 1 1 711
0 713 7 1 2 1182 1253
0 714 5 1 1 713
0 715 7 1 2 1184 1251
0 716 5 1 1 715
0 717 7 1 2 714 716
0 718 5 1 1 717
0 719 7 1 2 712 718
0 720 7 1 2 657 719
0 721 7 1 2 962 720
0 722 7 1 2 482 1261
0 723 5 1 1 722
0 724 7 1 2 1177 1259
0 725 5 1 1 724
0 726 7 1 2 723 725
0 727 7 1 2 721 726
0 728 7 1 2 651 727
0 729 7 1 2 647 728
0 730 7 1 2 645 729
0 731 7 1 2 472 730
0 732 5 1 1 731
0 733 7 1 2 587 732
3 2499 5 0 1 733
