1 0 0 2 0
2 49 1 0
2 720 1 0
1 1 0 2 0
2 721 1 1
2 722 1 1
1 2 0 2 0
2 723 1 2
2 724 1 2
1 3 0 2 0
2 725 1 3
2 726 1 3
1 4 0 2 0
2 727 1 4
2 728 1 4
1 5 0 2 0
2 729 1 5
2 730 1 5
1 6 0 2 0
2 731 1 6
2 732 1 6
1 7 0 2 0
2 733 1 7
2 734 1 7
1 8 0 2 0
2 735 1 8
2 736 1 8
1 9 0 2 0
2 737 1 9
2 738 1 9
1 10 0 2 0
2 739 1 10
2 740 1 10
1 11 0 2 0
2 741 1 11
2 742 1 11
1 12 0 2 0
2 743 1 12
2 744 1 12
1 13 0 2 0
2 745 1 13
2 746 1 13
1 14 0 2 0
2 747 1 14
2 748 1 14
1 15 0 2 0
2 749 1 15
2 750 1 15
1 16 0 2 0
2 751 1 16
2 752 1 16
1 17 0 2 0
2 753 1 17
2 754 1 17
1 18 0 2 0
2 755 1 18
2 756 1 18
1 19 0 2 0
2 757 1 19
2 758 1 19
1 20 0 2 0
2 759 1 20
2 760 1 20
1 21 0 2 0
2 761 1 21
2 762 1 21
1 22 0 2 0
2 763 1 22
2 764 1 22
1 23 0 2 0
2 765 1 23
2 766 1 23
1 24 0 2 0
2 767 1 24
2 768 1 24
1 25 0 2 0
2 769 1 25
2 770 1 25
1 26 0 2 0
2 771 1 26
2 772 1 26
1 27 0 2 0
2 773 1 27
2 774 1 27
1 28 0 2 0
2 775 1 28
2 776 1 28
1 29 0 2 0
2 777 1 29
2 778 1 29
1 30 0 2 0
2 779 1 30
2 780 1 30
1 31 0 2 0
2 781 1 31
2 782 1 31
1 32 0 2 0
2 783 1 32
2 784 1 32
1 33 0 2 0
2 785 1 33
2 786 1 33
1 34 0 2 0
2 787 1 34
2 788 1 34
1 35 0 2 0
2 789 1 35
2 790 1 35
1 36 0 2 0
2 791 1 36
2 792 1 36
1 37 0 2 0
2 793 1 37
2 794 1 37
1 38 0 2 0
2 795 1 38
2 796 1 38
1 39 0 2 0
2 797 1 39
2 798 1 39
1 40 0 2 0
2 799 1 40
2 800 1 40
1 41 0 2 0
2 801 1 41
2 802 1 41
1 42 0 2 0
2 803 1 42
2 804 1 42
1 43 0 2 0
2 805 1 43
2 806 1 43
1 44 0 2 0
2 807 1 44
2 808 1 44
1 45 0 2 0
2 809 1 45
2 810 1 45
1 46 0 2 0
2 811 1 46
2 812 1 46
1 47 0 2 0
2 813 1 47
2 814 1 47
1 48 0 2 0
2 815 1 48
2 816 1 48
2 817 1 69
2 818 1 69
2 819 1 70
2 820 1 70
2 821 1 71
2 822 1 71
2 823 1 72
2 824 1 72
2 825 1 73
2 826 1 73
2 827 1 74
2 828 1 74
2 829 1 75
2 830 1 75
2 831 1 76
2 832 1 76
2 833 1 77
2 834 1 77
2 835 1 78
2 836 1 78
2 837 1 79
2 838 1 79
2 839 1 80
2 840 1 80
2 841 1 81
2 842 1 81
2 843 1 100
2 844 1 100
2 845 1 102
2 846 1 102
2 847 1 104
2 848 1 104
2 849 1 106
2 850 1 106
2 851 1 107
2 852 1 107
2 853 1 108
2 854 1 108
2 855 1 108
2 856 1 111
2 857 1 111
2 858 1 112
2 859 1 112
2 860 1 115
2 861 1 115
2 862 1 118
2 863 1 118
2 864 1 120
2 865 1 120
2 866 1 123
2 867 1 123
2 868 1 126
2 869 1 126
2 870 1 128
2 871 1 128
2 872 1 131
2 873 1 131
2 874 1 134
2 875 1 134
2 876 1 136
2 877 1 136
2 878 1 139
2 879 1 139
2 880 1 142
2 881 1 142
2 882 1 144
2 883 1 144
2 884 1 147
2 885 1 147
2 886 1 150
2 887 1 150
2 888 1 152
2 889 1 152
2 890 1 155
2 891 1 155
2 892 1 158
2 893 1 158
2 894 1 160
2 895 1 160
2 896 1 163
2 897 1 163
2 898 1 166
2 899 1 166
2 900 1 168
2 901 1 168
2 902 1 171
2 903 1 171
2 904 1 174
2 905 1 174
2 906 1 176
2 907 1 176
2 908 1 179
2 909 1 179
2 910 1 182
2 911 1 182
2 912 1 184
2 913 1 184
2 914 1 187
2 915 1 187
2 916 1 190
2 917 1 190
2 918 1 192
2 919 1 192
2 920 1 195
2 921 1 195
2 922 1 198
2 923 1 198
2 924 1 200
2 925 1 200
2 926 1 203
2 927 1 203
2 928 1 206
2 929 1 206
2 930 1 208
2 931 1 208
2 932 1 211
2 933 1 211
2 934 1 214
2 935 1 214
2 936 1 216
2 937 1 216
2 938 1 219
2 939 1 219
2 940 1 221
2 941 1 221
2 942 1 222
2 943 1 222
2 944 1 223
2 945 1 223
2 946 1 224
2 947 1 224
2 948 1 225
2 949 1 225
2 950 1 231
2 951 1 231
2 952 1 233
2 953 1 233
2 954 1 234
2 955 1 234
2 956 1 234
2 957 1 235
2 958 1 235
2 959 1 241
2 960 1 241
2 961 1 244
2 962 1 244
2 963 1 244
2 964 1 244
2 965 1 246
2 966 1 246
2 967 1 246
2 968 1 247
2 969 1 247
2 970 1 253
2 971 1 253
2 972 1 256
2 973 1 256
2 974 1 256
2 975 1 256
2 976 1 258
2 977 1 258
2 978 1 258
2 979 1 259
2 980 1 259
2 981 1 265
2 982 1 265
2 983 1 268
2 984 1 268
2 985 1 268
2 986 1 268
2 987 1 269
2 988 1 269
2 989 1 275
2 990 1 275
2 991 1 278
2 992 1 278
2 993 1 278
2 994 1 278
2 995 1 280
2 996 1 280
2 997 1 280
2 998 1 281
2 999 1 281
2 1000 1 287
2 1001 1 287
2 1002 1 290
2 1003 1 290
2 1004 1 290
2 1005 1 290
2 1006 1 292
2 1007 1 292
2 1008 1 292
2 1009 1 293
2 1010 1 293
2 1011 1 299
2 1012 1 299
2 1013 1 302
2 1014 1 302
2 1015 1 302
2 1016 1 304
2 1017 1 304
2 1018 1 304
2 1019 1 305
2 1020 1 305
2 1021 1 311
2 1022 1 311
2 1023 1 314
2 1024 1 314
2 1025 1 314
2 1026 1 316
2 1027 1 316
2 1028 1 316
2 1029 1 317
2 1030 1 317
2 1031 1 323
2 1032 1 323
2 1033 1 326
2 1034 1 326
2 1035 1 326
2 1036 1 328
2 1037 1 328
2 1038 1 328
2 1039 1 328
2 1040 1 329
2 1041 1 329
2 1042 1 335
2 1043 1 335
2 1044 1 337
2 1045 1 337
2 1046 1 338
2 1047 1 338
2 1048 1 338
2 1049 1 339
2 1050 1 339
2 1051 1 340
2 1052 1 340
2 1053 1 340
2 1054 1 341
2 1055 1 341
2 1056 1 347
2 1057 1 347
2 1058 1 349
2 1059 1 349
2 1060 1 350
2 1061 1 350
2 1062 1 350
2 1063 1 350
2 1064 1 351
2 1065 1 351
2 1066 1 352
2 1067 1 352
2 1068 1 352
2 1069 1 353
2 1070 1 353
2 1071 1 359
2 1072 1 359
2 1073 1 362
2 1074 1 362
2 1075 1 362
2 1076 1 362
2 1077 1 364
2 1078 1 364
2 1079 1 364
2 1080 1 365
2 1081 1 365
2 1082 1 371
2 1083 1 371
2 1084 1 374
2 1085 1 374
2 1086 1 374
2 1087 1 376
2 1088 1 376
2 1089 1 376
2 1090 1 377
2 1091 1 377
2 1092 1 383
2 1093 1 383
2 1094 1 386
2 1095 1 386
2 1096 1 386
2 1097 1 388
2 1098 1 388
2 1099 1 388
2 1100 1 389
2 1101 1 389
2 1102 1 395
2 1103 1 395
2 1104 1 398
2 1105 1 398
2 1106 1 400
2 1107 1 400
2 1108 1 403
2 1109 1 403
2 1110 1 407
2 1111 1 407
2 1112 1 413
2 1113 1 413
2 1114 1 413
2 1115 1 417
2 1116 1 417
2 1117 1 419
2 1118 1 419
2 1119 1 421
2 1120 1 421
2 1121 1 422
2 1122 1 422
2 1123 1 429
2 1124 1 429
2 1125 1 432
2 1126 1 432
2 1127 1 433
2 1128 1 433
2 1129 1 436
2 1130 1 436
2 1131 1 437
2 1132 1 437
2 1133 1 440
2 1134 1 440
2 1135 1 443
2 1136 1 443
2 1137 1 447
2 1138 1 447
2 1139 1 452
2 1140 1 452
2 1141 1 452
2 1142 1 455
2 1143 1 455
2 1144 1 461
2 1145 1 461
2 1146 1 462
2 1147 1 462
2 1148 1 463
2 1149 1 463
2 1150 1 463
2 1151 1 466
2 1152 1 466
2 1153 1 470
2 1154 1 470
2 1155 1 474
2 1156 1 474
2 1157 1 480
2 1158 1 480
2 1159 1 480
2 1160 1 486
2 1161 1 486
2 1162 1 487
2 1163 1 487
2 1164 1 490
2 1165 1 490
2 1166 1 490
2 1167 1 496
2 1168 1 496
2 1169 1 496
2 1170 1 502
2 1171 1 502
2 1172 1 503
2 1173 1 503
2 1174 1 506
2 1175 1 506
2 1176 1 506
2 1177 1 507
2 1178 1 507
2 1179 1 512
2 1180 1 512
2 1181 1 512
2 1182 1 513
2 1183 1 513
2 1184 1 518
2 1185 1 518
2 1186 1 519
2 1187 1 519
2 1188 1 522
2 1189 1 522
2 1190 1 534
2 1191 1 534
2 1192 1 535
2 1193 1 535
2 1194 1 538
2 1195 1 538
2 1196 1 538
2 1197 1 539
2 1198 1 539
2 1199 1 545
2 1200 1 545
2 1201 1 549
2 1202 1 549
2 1203 1 581
2 1204 1 581
2 1205 1 582
2 1206 1 582
2 1207 1 585
2 1208 1 585
2 1209 1 586
2 1210 1 586
2 1211 1 589
2 1212 1 589
2 1213 1 593
2 1214 1 593
2 1215 1 600
2 1216 1 600
2 1217 1 603
2 1218 1 603
2 1219 1 604
2 1220 1 604
2 1221 1 607
2 1222 1 607
2 1223 1 608
2 1224 1 608
2 1225 1 611
2 1226 1 611
2 1227 1 612
2 1228 1 612
2 1229 1 615
2 1230 1 615
2 1231 1 616
2 1232 1 616
2 1233 1 619
2 1234 1 619
2 1235 1 620
2 1236 1 620
2 1237 1 623
2 1238 1 623
2 1239 1 624
2 1240 1 624
2 1241 1 627
2 1242 1 627
2 1243 1 628
2 1244 1 628
0 50 5 1 1 49
0 51 5 1 1 721
0 52 5 1 1 723
0 53 5 1 1 725
0 54 5 1 1 727
0 55 5 1 1 729
0 56 5 1 1 731
0 57 5 1 1 733
0 58 5 1 1 735
0 59 5 1 1 737
0 60 5 1 1 739
0 61 5 1 1 741
0 62 5 1 1 743
0 63 5 1 1 745
0 64 5 1 1 747
0 65 5 1 1 749
0 66 5 1 1 751
0 67 5 1 1 753
0 68 5 1 1 755
0 69 5 2 1 757
0 70 5 2 1 759
0 71 5 2 1 761
0 72 5 2 1 763
0 73 5 2 1 765
0 74 5 2 1 767
0 75 5 2 1 769
0 76 5 2 1 771
0 77 5 2 1 773
0 78 5 2 1 775
0 79 5 2 1 777
0 80 5 2 1 779
0 81 5 2 1 781
0 82 5 1 1 783
0 83 5 1 1 785
0 84 5 1 1 787
0 85 5 1 1 789
0 86 5 1 1 791
0 87 5 1 1 793
0 88 5 1 1 795
0 89 5 1 1 797
0 90 5 1 1 799
0 91 5 1 1 801
0 92 5 1 1 803
0 93 5 1 1 805
0 94 5 1 1 807
0 95 5 1 1 809
0 96 5 1 1 811
0 97 5 1 1 813
0 98 5 1 1 815
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 724 756
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 722 754
0 106 5 2 1 105
0 107 7 2 2 720 752
0 108 5 3 1 851
0 109 7 1 2 849 853
0 110 5 1 1 109
0 111 7 2 2 847 110
0 112 5 2 1 856
0 113 7 1 2 845 858
0 114 5 1 1 113
0 115 7 2 2 843 114
0 116 5 1 1 860
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 726 861
0 120 5 2 1 119
0 121 7 1 2 817 864
0 122 5 1 1 121
0 123 7 2 2 862 122
0 124 5 1 1 866
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 728 867
0 128 5 2 1 127
0 129 7 1 2 819 870
0 130 5 1 1 129
0 131 7 2 2 868 130
0 132 5 1 1 872
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 730 873
0 136 5 2 1 135
0 137 7 1 2 821 876
0 138 5 1 1 137
0 139 7 2 2 874 138
0 140 5 1 1 878
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 732 879
0 144 5 2 1 143
0 145 7 1 2 823 882
0 146 5 1 1 145
0 147 7 2 2 880 146
0 148 5 1 1 884
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 734 885
0 152 5 2 1 151
0 153 7 1 2 825 888
0 154 5 1 1 153
0 155 7 2 2 886 154
0 156 5 1 1 890
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 736 891
0 160 5 2 1 159
0 161 7 1 2 827 894
0 162 5 1 1 161
0 163 7 2 2 892 162
0 164 5 1 1 896
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 738 897
0 168 5 2 1 167
0 169 7 1 2 829 900
0 170 5 1 1 169
0 171 7 2 2 898 170
0 172 5 1 1 902
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 740 903
0 176 5 2 1 175
0 177 7 1 2 831 906
0 178 5 1 1 177
0 179 7 2 2 904 178
0 180 5 1 1 908
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 742 909
0 184 5 2 1 183
0 185 7 1 2 833 912
0 186 5 1 1 185
0 187 7 2 2 910 186
0 188 5 1 1 914
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 744 915
0 192 5 2 1 191
0 193 7 1 2 835 918
0 194 5 1 1 193
0 195 7 2 2 916 194
0 196 5 1 1 920
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 746 921
0 200 5 2 1 199
0 201 7 1 2 837 924
0 202 5 1 1 201
0 203 7 2 2 922 202
0 204 5 1 1 926
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 748 927
0 208 5 2 1 207
0 209 7 1 2 839 930
0 210 5 1 1 209
0 211 7 2 2 928 210
0 212 5 1 1 932
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 750 933
0 216 5 2 1 215
0 217 7 1 2 841 936
0 218 5 1 1 217
0 219 7 2 2 934 218
0 220 5 1 1 938
0 221 7 2 2 816 220
0 222 5 2 1 940
0 223 7 2 2 98 939
0 224 5 2 1 944
0 225 7 2 2 935 937
0 226 5 1 1 948
0 227 7 1 2 782 226
0 228 5 1 1 227
0 229 7 1 2 842 949
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 950
0 233 7 2 2 814 951
0 234 5 3 1 952
0 235 7 2 2 929 931
0 236 5 1 1 957
0 237 7 1 2 780 958
0 238 5 1 1 237
0 239 7 1 2 840 236
0 240 5 1 1 239
0 241 7 2 2 238 240
0 242 5 1 1 959
0 243 7 1 2 812 242
0 244 5 4 1 243
0 245 7 1 2 96 960
0 246 5 3 1 245
0 247 7 2 2 923 925
0 248 5 1 1 968
0 249 7 1 2 778 969
0 250 5 1 1 249
0 251 7 1 2 838 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 970
0 255 7 1 2 810 254
0 256 5 4 1 255
0 257 7 1 2 95 971
0 258 5 3 1 257
0 259 7 2 2 917 919
0 260 5 1 1 979
0 261 7 1 2 776 980
0 262 5 1 1 261
0 263 7 1 2 836 260
0 264 5 1 1 263
0 265 7 2 2 262 264
0 266 5 1 1 981
0 267 7 1 2 808 266
0 268 5 4 1 267
0 269 7 2 2 911 913
0 270 5 1 1 987
0 271 7 1 2 774 988
0 272 5 1 1 271
0 273 7 1 2 834 270
0 274 5 1 1 273
0 275 7 2 2 272 274
0 276 5 1 1 989
0 277 7 1 2 806 276
0 278 5 4 1 277
0 279 7 1 2 93 990
0 280 5 3 1 279
0 281 7 2 2 905 907
0 282 5 1 1 998
0 283 7 1 2 772 999
0 284 5 1 1 283
0 285 7 1 2 832 282
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 1000
0 289 7 1 2 804 288
0 290 5 4 1 289
0 291 7 1 2 92 1001
0 292 5 3 1 291
0 293 7 2 2 899 901
0 294 5 1 1 1009
0 295 7 1 2 770 1010
0 296 5 1 1 295
0 297 7 1 2 830 294
0 298 5 1 1 297
0 299 7 2 2 296 298
0 300 5 1 1 1011
0 301 7 1 2 91 1012
0 302 5 3 1 301
0 303 7 1 2 802 300
0 304 5 3 1 303
0 305 7 2 2 893 895
0 306 5 1 1 1019
0 307 7 1 2 768 1020
0 308 5 1 1 307
0 309 7 1 2 828 306
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 1021
0 313 7 1 2 90 1022
0 314 5 3 1 313
0 315 7 1 2 800 312
0 316 5 3 1 315
0 317 7 2 2 887 889
0 318 5 1 1 1029
0 319 7 1 2 766 1030
0 320 5 1 1 319
0 321 7 1 2 826 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1031
0 325 7 1 2 89 1032
0 326 5 3 1 325
0 327 7 1 2 798 324
0 328 5 4 1 327
0 329 7 2 2 881 883
0 330 5 1 1 1040
0 331 7 1 2 764 1041
0 332 5 1 1 331
0 333 7 1 2 824 330
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 1042
0 337 7 2 2 88 1043
0 338 5 3 1 1044
0 339 7 2 2 796 336
0 340 5 3 1 1049
0 341 7 2 2 875 877
0 342 5 1 1 1054
0 343 7 1 2 762 1055
0 344 5 1 1 343
0 345 7 1 2 822 342
0 346 5 1 1 345
0 347 7 2 2 344 346
0 348 5 1 1 1056
0 349 7 2 2 794 348
0 350 5 4 1 1058
0 351 7 2 2 87 1057
0 352 5 3 1 1064
0 353 7 2 2 869 871
0 354 5 1 1 1069
0 355 7 1 2 760 1070
0 356 5 1 1 355
0 357 7 1 2 820 354
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 1071
0 361 7 1 2 792 360
0 362 5 4 1 361
0 363 7 1 2 86 1072
0 364 5 3 1 363
0 365 7 2 2 863 865
0 366 5 1 1 1080
0 367 7 1 2 758 1081
0 368 5 1 1 367
0 369 7 1 2 818 366
0 370 5 1 1 369
0 371 7 2 2 368 370
0 372 5 1 1 1082
0 373 7 1 2 790 372
0 374 5 3 1 373
0 375 7 1 2 85 1083
0 376 5 3 1 375
0 377 7 2 2 844 846
0 378 5 1 1 1090
0 379 7 1 2 857 378
0 380 5 1 1 379
0 381 7 1 2 859 1091
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 1092
0 385 7 1 2 84 384
0 386 5 3 1 385
0 387 7 1 2 788 1093
0 388 5 3 1 387
0 389 7 2 2 848 850
0 390 5 1 1 1100
0 391 7 1 2 852 390
0 392 5 1 1 391
0 393 7 1 2 854 1101
0 394 5 1 1 393
0 395 7 2 2 392 394
0 396 5 1 1 1102
0 397 7 1 2 83 396
0 398 5 2 1 397
0 399 7 1 2 786 1103
0 400 5 2 1 399
0 401 7 1 2 50 66
0 402 5 1 1 401
0 403 7 2 2 855 402
0 404 5 1 1 1108
0 405 7 1 2 784 404
0 406 5 1 1 405
0 407 7 2 2 1106 406
0 408 5 1 1 1110
0 409 7 1 2 1104 408
0 410 5 1 1 409
0 411 7 1 2 1097 410
0 412 5 1 1 411
0 413 7 3 2 1094 412
0 414 5 1 1 1112
0 415 7 1 2 1087 1113
0 416 5 1 1 415
0 417 7 2 2 1084 416
0 418 5 1 1 1115
0 419 7 2 2 1077 418
0 420 5 1 1 1117
0 421 7 2 2 1073 420
0 422 5 2 1 1119
0 423 7 1 2 1066 1121
0 424 5 1 1 423
0 425 7 1 2 1060 424
0 426 7 1 2 1051 425
0 427 5 1 1 426
0 428 7 1 2 1046 427
0 429 5 2 1 428
0 430 7 1 2 1036 1123
0 431 5 1 1 430
0 432 7 2 2 1033 431
0 433 5 2 1 1125
0 434 7 1 2 1026 1127
0 435 5 1 1 434
0 436 7 2 2 1023 435
0 437 5 2 1 1129
0 438 7 1 2 1016 1131
0 439 5 1 1 438
0 440 7 2 2 1013 439
0 441 5 1 1 1133
0 442 7 1 2 1006 1134
0 443 5 2 1 442
0 444 7 1 2 1002 1135
0 445 5 1 1 444
0 446 7 1 2 995 445
0 447 5 2 1 446
0 448 7 1 2 991 1137
0 449 7 1 2 983 448
0 450 5 1 1 449
0 451 7 1 2 94 982
0 452 5 3 1 451
0 453 7 1 2 450 1139
0 454 7 1 2 976 453
0 455 5 2 1 454
0 456 7 1 2 972 1142
0 457 5 1 1 456
0 458 7 1 2 965 457
0 459 5 1 1 458
0 460 7 1 2 961 459
0 461 5 2 1 460
0 462 7 2 2 97 232
0 463 5 3 1 1146
0 464 7 1 2 1144 1148
0 465 5 1 1 464
0 466 7 2 2 954 465
0 467 5 1 1 1151
0 468 7 1 2 946 467
0 469 5 1 1 468
0 470 7 2 2 942 469
0 471 5 1 1 1153
0 472 7 1 2 945 1152
0 473 5 1 1 472
0 474 7 2 2 1149 955
0 475 5 1 1 1155
0 476 7 1 2 962 475
0 477 5 1 1 476
0 478 7 1 2 1145 1156
0 479 5 1 1 478
0 480 7 3 2 963 966
0 481 5 1 1 1157
0 482 7 1 2 1143 1158
0 483 5 1 1 482
0 484 7 1 2 973 483
0 485 5 1 1 484
0 486 7 2 2 974 977
0 487 5 2 1 1160
0 488 7 1 2 984 1162
0 489 5 1 1 488
0 490 7 3 2 985 1140
0 491 5 1 1 1164
0 492 7 1 2 1138 1165
0 493 5 1 1 492
0 494 7 1 2 992 493
0 495 5 1 1 494
0 496 7 3 2 993 996
0 497 5 1 1 1167
0 498 7 1 2 1136 1168
0 499 5 1 1 498
0 500 7 1 2 1003 499
0 501 5 1 1 500
0 502 7 2 2 1004 1007
0 503 5 2 1 1170
0 504 7 1 2 441 1172
0 505 5 1 1 504
0 506 7 3 2 1014 1017
0 507 5 2 1 1174
0 508 7 1 2 1132 1175
0 509 5 1 1 508
0 510 7 1 2 1130 1177
0 511 5 1 1 510
0 512 7 3 2 1024 1027
0 513 5 2 1 1179
0 514 7 1 2 1126 1182
0 515 5 1 1 514
0 516 7 1 2 1128 1180
0 517 5 1 1 516
0 518 7 2 2 1034 1037
0 519 5 2 1 1184
0 520 7 1 2 1124 1185
0 521 5 1 1 520
0 522 7 2 2 1065 1120
0 523 5 1 1 1188
0 524 7 1 2 1045 1189
0 525 5 1 1 524
0 526 7 1 2 1186 525
0 527 5 1 1 526
0 528 7 1 2 1050 523
0 529 5 1 1 528
0 530 7 1 2 1059 1122
0 531 5 1 1 530
0 532 7 1 2 1074 1118
0 533 5 1 1 532
0 534 7 2 2 1075 1078
0 535 5 2 1 1190
0 536 7 1 2 1116 1192
0 537 5 1 1 536
0 538 7 3 2 1085 1088
0 539 5 2 1 1194
0 540 7 1 2 414 1195
0 541 5 1 1 540
0 542 7 1 2 1095 1098
0 543 7 1 2 82 1109
0 544 5 1 1 543
0 545 7 2 2 1105 544
0 546 5 1 1 1199
0 547 7 1 2 1111 1200
0 548 7 1 2 542 547
0 549 5 2 1 548
0 550 7 1 2 1114 1197
0 551 5 1 1 550
0 552 7 1 2 1201 551
0 553 7 1 2 541 552
0 554 5 1 1 553
0 555 7 1 2 537 554
0 556 7 1 2 533 555
0 557 5 1 1 556
0 558 7 1 2 531 557
0 559 7 1 2 529 558
0 560 7 1 2 527 559
0 561 7 1 2 521 560
0 562 7 1 2 517 561
0 563 7 1 2 515 562
0 564 7 1 2 511 563
0 565 7 1 2 509 564
0 566 5 1 1 565
0 567 7 1 2 505 566
0 568 7 1 2 501 567
0 569 7 1 2 495 568
0 570 7 1 2 489 569
0 571 7 1 2 485 570
0 572 7 1 2 479 571
0 573 7 1 2 477 572
0 574 7 1 2 473 573
0 575 7 1 2 1154 574
0 576 5 1 1 575
0 577 7 1 2 1107 546
0 578 5 1 1 577
0 579 7 1 2 1096 578
0 580 5 1 1 579
0 581 7 2 2 1099 580
0 582 5 2 1 1203
0 583 7 1 2 1089 1205
0 584 5 1 1 583
0 585 7 2 2 1086 584
0 586 5 2 1 1207
0 587 7 1 2 1079 1209
0 588 5 1 1 587
0 589 7 2 2 1076 588
0 590 5 1 1 1211
0 591 7 1 2 1067 590
0 592 5 1 1 591
0 593 7 2 2 1052 592
0 594 7 1 2 1061 1213
0 595 5 1 1 594
0 596 7 1 2 1047 595
0 597 7 1 2 1035 596
0 598 5 1 1 597
0 599 7 1 2 1038 598
0 600 5 2 1 599
0 601 7 1 2 1025 1215
0 602 5 1 1 601
0 603 7 2 2 1028 602
0 604 5 2 1 1217
0 605 7 1 2 1015 1219
0 606 5 1 1 605
0 607 7 2 2 1018 606
0 608 5 2 1 1221
0 609 7 1 2 1008 1223
0 610 5 1 1 609
0 611 7 2 2 1005 610
0 612 5 2 1 1225
0 613 7 1 2 997 1227
0 614 5 1 1 613
0 615 7 2 2 994 614
0 616 5 2 1 1229
0 617 7 1 2 1141 1231
0 618 5 1 1 617
0 619 7 2 2 986 618
0 620 5 2 1 1233
0 621 7 1 2 978 1235
0 622 5 1 1 621
0 623 7 2 2 975 622
0 624 5 2 1 1237
0 625 7 1 2 967 1239
0 626 5 1 1 625
0 627 7 2 2 964 626
0 628 5 2 1 1241
0 629 7 1 2 1150 1243
0 630 5 1 1 629
0 631 7 1 2 956 943
0 632 7 1 2 630 631
0 633 5 1 1 632
0 634 7 1 2 1147 1242
0 635 5 1 1 634
0 636 7 1 2 941 635
0 637 5 1 1 636
0 638 7 1 2 953 1244
0 639 5 1 1 638
0 640 7 1 2 1159 1240
0 641 5 1 1 640
0 642 7 1 2 481 1238
0 643 5 1 1 642
0 644 7 1 2 641 643
0 645 5 1 1 644
0 646 7 1 2 1161 1236
0 647 5 1 1 646
0 648 7 1 2 1163 1234
0 649 5 1 1 648
0 650 7 1 2 647 649
0 651 5 1 1 650
0 652 7 1 2 1166 1230
0 653 5 1 1 652
0 654 7 1 2 491 1232
0 655 5 1 1 654
0 656 7 1 2 1169 1226
0 657 5 1 1 656
0 658 7 1 2 497 1228
0 659 5 1 1 658
0 660 7 1 2 1171 1224
0 661 5 1 1 660
0 662 7 1 2 1173 1222
0 663 5 1 1 662
0 664 7 1 2 661 663
0 665 5 1 1 664
0 666 7 1 2 1178 1218
0 667 5 1 1 666
0 668 7 1 2 1176 1220
0 669 5 1 1 668
0 670 7 1 2 1039 1183
0 671 5 1 1 670
0 672 7 1 2 1181 1216
0 673 5 1 1 672
0 674 7 1 2 1053 1187
0 675 5 1 1 674
0 676 7 1 2 1048 1214
0 677 5 1 1 676
0 678 7 1 2 1062 677
0 679 5 1 1 678
0 680 7 1 2 1063 1068
0 681 5 1 1 680
0 682 7 1 2 1212 681
0 683 5 1 1 682
0 684 7 1 2 1191 1208
0 685 5 1 1 684
0 686 7 1 2 1196 1206
0 687 5 1 1 686
0 688 7 1 2 1198 1204
0 689 5 1 1 688
0 690 7 1 2 1202 689
0 691 7 1 2 687 690
0 692 5 1 1 691
0 693 7 1 2 1193 1210
0 694 5 1 1 693
0 695 7 1 2 692 694
0 696 7 1 2 685 695
0 697 5 1 1 696
0 698 7 1 2 683 697
0 699 7 1 2 679 698
0 700 7 1 2 675 699
0 701 7 1 2 673 700
0 702 7 1 2 671 701
0 703 7 1 2 669 702
0 704 7 1 2 667 703
0 705 5 1 1 704
0 706 7 1 2 665 705
0 707 7 1 2 659 706
0 708 7 1 2 657 707
0 709 7 1 2 655 708
0 710 7 1 2 653 709
0 711 7 1 2 651 710
0 712 7 1 2 947 711
0 713 7 1 2 645 712
0 714 7 1 2 639 713
0 715 7 1 2 637 714
0 716 7 1 2 633 715
0 717 7 1 2 471 716
0 718 5 1 1 717
0 719 7 1 2 576 718
3 3499 5 0 1 719
