1 0 0 3 0
2 7 1 0
2 8 1 0
2 9 1 0
1 1 0 2 0
2 10 1 1
2 29 1 1
1 2 0 2 0
2 49 1 2
2 71 1 2
1 3 0 2 0
2 75 1 3
2 76 1 3
1 4 0 2 0
2 77 1 4
2 78 1 4
1 5 0 2 0
2 79 1 5
2 80 1 5
1 6 0 2 0
2 81 1 6
2 82 1 6
2 83 1 11
2 84 1 11
2 85 1 19
2 86 1 19
2 87 1 19
2 88 1 21
2 89 1 21
2 90 1 21
2 91 1 22
2 92 1 22
2 93 1 31
2 94 1 31
2 95 1 31
2 96 1 31
2 97 1 33
2 98 1 33
2 99 1 33
2 100 1 34
2 101 1 34
2 102 1 39
2 103 1 39
2 104 1 45
2 105 1 45
2 106 1 51
2 107 1 51
2 108 1 53
2 109 1 53
2 110 1 54
2 111 1 54
2 112 1 54
2 113 1 55
2 114 1 55
2 115 1 56
2 116 1 56
0 11 5 2 1 7
0 12 5 1 1 10
0 13 5 1 1 49
0 14 5 1 1 75
0 15 5 1 1 77
0 16 5 1 1 79
0 17 5 1 1 81
0 18 7 1 2 76 82
0 19 5 3 1 18
0 20 7 1 2 14 17
0 21 5 3 1 20
0 22 7 2 2 85 88
0 23 5 1 1 91
0 24 7 1 2 8 23
0 25 5 1 1 24
0 26 7 1 2 83 92
0 27 5 1 1 26
0 28 7 1 2 25 27
3 596 5 0 1 28
0 30 7 1 2 29 78
0 31 5 4 1 30
0 32 7 1 2 12 15
0 33 5 3 1 32
0 34 7 2 2 93 97
0 35 5 1 1 100
0 36 7 1 2 84 86
0 37 5 1 1 36
0 38 7 1 2 89 37
0 39 5 2 1 38
0 40 7 1 2 101 102
0 41 5 1 1 40
0 42 7 1 2 9 90
0 43 5 1 1 42
0 44 7 1 2 87 43
0 45 5 2 1 44
0 46 7 1 2 35 104
0 47 5 1 1 46
0 48 7 1 2 41 47
3 597 5 0 1 48
0 50 7 1 2 71 80
0 51 5 2 1 50
0 52 7 1 2 13 16
0 53 5 2 1 52
0 54 7 3 2 106 108
0 55 5 2 1 110
0 56 7 2 2 98 105
0 57 5 1 1 115
0 58 7 1 2 113 116
0 59 5 1 1 58
0 60 7 1 2 94 111
0 61 7 1 2 103 60
0 62 5 1 1 61
0 63 7 1 2 99 112
0 64 5 1 1 63
0 65 7 1 2 95 114
0 66 5 1 1 65
0 67 7 1 2 64 66
0 68 5 1 1 67
0 69 7 1 2 62 68
0 70 7 1 2 59 69
3 598 5 0 1 70
0 72 7 1 2 96 107
0 73 7 1 2 57 72
0 74 5 1 1 73
3 599 7 0 2 109 74
