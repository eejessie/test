1 0 0 4 0
2 49 1 0
2 3446 1 0
2 3447 1 0
2 3448 1 0
1 1 0 5 0
2 3449 1 1
2 3450 1 1
2 3451 1 1
2 3452 1 1
2 3453 1 1
1 2 0 6 0
2 3454 1 2
2 3455 1 2
2 3456 1 2
2 3457 1 2
2 3458 1 2
2 3459 1 2
1 3 0 6 0
2 3460 1 3
2 3461 1 3
2 3462 1 3
2 3463 1 3
2 3464 1 3
2 3465 1 3
1 4 0 6 0
2 3466 1 4
2 3467 1 4
2 3468 1 4
2 3469 1 4
2 3470 1 4
2 3471 1 4
1 5 0 7 0
2 3472 1 5
2 3473 1 5
2 3474 1 5
2 3475 1 5
2 3476 1 5
2 3477 1 5
2 3478 1 5
1 6 0 7 0
2 3479 1 6
2 3480 1 6
2 3481 1 6
2 3482 1 6
2 3483 1 6
2 3484 1 6
2 3485 1 6
1 7 0 6 0
2 3486 1 7
2 3487 1 7
2 3488 1 7
2 3489 1 7
2 3490 1 7
2 3491 1 7
1 8 0 7 0
2 3492 1 8
2 3493 1 8
2 3494 1 8
2 3495 1 8
2 3496 1 8
2 3497 1 8
2 3498 1 8
1 9 0 6 0
2 3499 1 9
2 3500 1 9
2 3501 1 9
2 3502 1 9
2 3503 1 9
2 3504 1 9
1 10 0 6 0
2 3505 1 10
2 3506 1 10
2 3507 1 10
2 3508 1 10
2 3509 1 10
2 3510 1 10
1 11 0 7 0
2 3511 1 11
2 3512 1 11
2 3513 1 11
2 3514 1 11
2 3515 1 11
2 3516 1 11
2 3517 1 11
1 12 0 7 0
2 3518 1 12
2 3519 1 12
2 3520 1 12
2 3521 1 12
2 3522 1 12
2 3523 1 12
2 3524 1 12
1 13 0 6 0
2 3525 1 13
2 3526 1 13
2 3527 1 13
2 3528 1 13
2 3529 1 13
2 3530 1 13
1 14 0 7 0
2 3531 1 14
2 3532 1 14
2 3533 1 14
2 3534 1 14
2 3535 1 14
2 3536 1 14
2 3537 1 14
1 15 0 6 0
2 3538 1 15
2 3539 1 15
2 3540 1 15
2 3541 1 15
2 3542 1 15
2 3543 1 15
1 16 0 6 0
2 3544 1 16
2 3545 1 16
2 3546 1 16
2 3547 1 16
2 3548 1 16
2 3549 1 16
1 17 0 7 0
2 3550 1 17
2 3551 1 17
2 3552 1 17
2 3553 1 17
2 3554 1 17
2 3555 1 17
2 3556 1 17
1 18 0 7 0
2 3557 1 18
2 3558 1 18
2 3559 1 18
2 3560 1 18
2 3561 1 18
2 3562 1 18
2 3563 1 18
1 19 0 6 0
2 3564 1 19
2 3565 1 19
2 3566 1 19
2 3567 1 19
2 3568 1 19
2 3569 1 19
1 20 0 7 0
2 3570 1 20
2 3571 1 20
2 3572 1 20
2 3573 1 20
2 3574 1 20
2 3575 1 20
2 3576 1 20
1 21 0 6 0
2 3577 1 21
2 3578 1 21
2 3579 1 21
2 3580 1 21
2 3581 1 21
2 3582 1 21
1 22 0 6 0
2 3583 1 22
2 3584 1 22
2 3585 1 22
2 3586 1 22
2 3587 1 22
2 3588 1 22
1 23 0 7 0
2 3589 1 23
2 3590 1 23
2 3591 1 23
2 3592 1 23
2 3593 1 23
2 3594 1 23
2 3595 1 23
1 24 0 7 0
2 3596 1 24
2 3597 1 24
2 3598 1 24
2 3599 1 24
2 3600 1 24
2 3601 1 24
2 3602 1 24
1 25 0 6 0
2 3603 1 25
2 3604 1 25
2 3605 1 25
2 3606 1 25
2 3607 1 25
2 3608 1 25
1 26 0 7 0
2 3609 1 26
2 3610 1 26
2 3611 1 26
2 3612 1 26
2 3613 1 26
2 3614 1 26
2 3615 1 26
1 27 0 6 0
2 3616 1 27
2 3617 1 27
2 3618 1 27
2 3619 1 27
2 3620 1 27
2 3621 1 27
1 28 0 6 0
2 3622 1 28
2 3623 1 28
2 3624 1 28
2 3625 1 28
2 3626 1 28
2 3627 1 28
1 29 0 7 0
2 3628 1 29
2 3629 1 29
2 3630 1 29
2 3631 1 29
2 3632 1 29
2 3633 1 29
2 3634 1 29
1 30 0 7 0
2 3635 1 30
2 3636 1 30
2 3637 1 30
2 3638 1 30
2 3639 1 30
2 3640 1 30
2 3641 1 30
1 31 0 6 0
2 3642 1 31
2 3643 1 31
2 3644 1 31
2 3645 1 31
2 3646 1 31
2 3647 1 31
1 32 0 7 0
2 3648 1 32
2 3649 1 32
2 3650 1 32
2 3651 1 32
2 3652 1 32
2 3653 1 32
2 3654 1 32
1 33 0 6 0
2 3655 1 33
2 3656 1 33
2 3657 1 33
2 3658 1 33
2 3659 1 33
2 3660 1 33
1 34 0 6 0
2 3661 1 34
2 3662 1 34
2 3663 1 34
2 3664 1 34
2 3665 1 34
2 3666 1 34
1 35 0 7 0
2 3667 1 35
2 3668 1 35
2 3669 1 35
2 3670 1 35
2 3671 1 35
2 3672 1 35
2 3673 1 35
1 36 0 7 0
2 3674 1 36
2 3675 1 36
2 3676 1 36
2 3677 1 36
2 3678 1 36
2 3679 1 36
2 3680 1 36
1 37 0 6 0
2 3681 1 37
2 3682 1 37
2 3683 1 37
2 3684 1 37
2 3685 1 37
2 3686 1 37
1 38 0 7 0
2 3687 1 38
2 3688 1 38
2 3689 1 38
2 3690 1 38
2 3691 1 38
2 3692 1 38
2 3693 1 38
1 39 0 6 0
2 3694 1 39
2 3695 1 39
2 3696 1 39
2 3697 1 39
2 3698 1 39
2 3699 1 39
1 40 0 6 0
2 3700 1 40
2 3701 1 40
2 3702 1 40
2 3703 1 40
2 3704 1 40
2 3705 1 40
1 41 0 7 0
2 3706 1 41
2 3707 1 41
2 3708 1 41
2 3709 1 41
2 3710 1 41
2 3711 1 41
2 3712 1 41
1 42 0 7 0
2 3713 1 42
2 3714 1 42
2 3715 1 42
2 3716 1 42
2 3717 1 42
2 3718 1 42
2 3719 1 42
1 43 0 7 0
2 3720 1 43
2 3721 1 43
2 3722 1 43
2 3723 1 43
2 3724 1 43
2 3725 1 43
2 3726 1 43
1 44 0 7 0
2 3727 1 44
2 3728 1 44
2 3729 1 44
2 3730 1 44
2 3731 1 44
2 3732 1 44
2 3733 1 44
1 45 0 8 0
2 3734 1 45
2 3735 1 45
2 3736 1 45
2 3737 1 45
2 3738 1 45
2 3739 1 45
2 3740 1 45
2 3741 1 45
1 46 0 8 0
2 3742 1 46
2 3743 1 46
2 3744 1 46
2 3745 1 46
2 3746 1 46
2 3747 1 46
2 3748 1 46
2 3749 1 46
1 47 0 7 0
2 3750 1 47
2 3751 1 47
2 3752 1 47
2 3753 1 47
2 3754 1 47
2 3755 1 47
2 3756 1 47
1 48 0 6 0
2 3757 1 48
2 3758 1 48
2 3759 1 48
2 3760 1 48
2 3761 1 48
2 3762 1 48
2 3763 1 50
2 3764 1 50
2 3765 1 50
2 3766 1 50
2 3767 1 50
2 3768 1 51
2 3769 1 51
2 3770 1 51
2 3771 1 51
2 3772 1 51
2 3773 1 51
2 3774 1 52
2 3775 1 52
2 3776 1 52
2 3777 1 52
2 3778 1 52
2 3779 1 52
2 3780 1 53
2 3781 1 53
2 3782 1 53
2 3783 1 53
2 3784 1 53
2 3785 1 53
2 3786 1 54
2 3787 1 54
2 3788 1 54
2 3789 1 54
2 3790 1 54
2 3791 1 54
2 3792 1 55
2 3793 1 55
2 3794 1 55
2 3795 1 55
2 3796 1 55
2 3797 1 56
2 3798 1 56
2 3799 1 56
2 3800 1 56
2 3801 1 56
2 3802 1 56
2 3803 1 57
2 3804 1 57
2 3805 1 57
2 3806 1 57
2 3807 1 57
2 3808 1 57
2 3809 1 58
2 3810 1 58
2 3811 1 58
2 3812 1 58
2 3813 1 58
2 3814 1 59
2 3815 1 59
2 3816 1 59
2 3817 1 59
2 3818 1 59
2 3819 1 59
2 3820 1 60
2 3821 1 60
2 3822 1 60
2 3823 1 60
2 3824 1 60
2 3825 1 60
2 3826 1 61
2 3827 1 61
2 3828 1 61
2 3829 1 61
2 3830 1 61
2 3831 1 62
2 3832 1 62
2 3833 1 62
2 3834 1 62
2 3835 1 62
2 3836 1 62
2 3837 1 63
2 3838 1 63
2 3839 1 63
2 3840 1 63
2 3841 1 63
2 3842 1 63
2 3843 1 64
2 3844 1 64
2 3845 1 64
2 3846 1 64
2 3847 1 64
2 3848 1 65
2 3849 1 65
2 3850 1 65
2 3851 1 65
2 3852 1 65
2 3853 1 65
2 3854 1 66
2 3855 1 66
2 3856 1 66
2 3857 1 66
2 3858 1 66
2 3859 1 66
2 3860 1 67
2 3861 1 67
2 3862 1 67
2 3863 1 67
2 3864 1 67
2 3865 1 68
2 3866 1 68
2 3867 1 68
2 3868 1 68
2 3869 1 68
2 3870 1 68
2 3871 1 69
2 3872 1 69
2 3873 1 69
2 3874 1 69
2 3875 1 69
2 3876 1 69
2 3877 1 69
2 3878 1 70
2 3879 1 70
2 3880 1 70
2 3881 1 70
2 3882 1 70
2 3883 1 70
2 3884 1 71
2 3885 1 71
2 3886 1 71
2 3887 1 71
2 3888 1 71
2 3889 1 71
2 3890 1 71
2 3891 1 72
2 3892 1 72
2 3893 1 72
2 3894 1 72
2 3895 1 72
2 3896 1 72
2 3897 1 72
2 3898 1 73
2 3899 1 73
2 3900 1 73
2 3901 1 73
2 3902 1 73
2 3903 1 73
2 3904 1 74
2 3905 1 74
2 3906 1 74
2 3907 1 74
2 3908 1 74
2 3909 1 74
2 3910 1 74
2 3911 1 75
2 3912 1 75
2 3913 1 75
2 3914 1 75
2 3915 1 75
2 3916 1 75
2 3917 1 75
2 3918 1 76
2 3919 1 76
2 3920 1 76
2 3921 1 76
2 3922 1 76
2 3923 1 76
2 3924 1 77
2 3925 1 77
2 3926 1 77
2 3927 1 77
2 3928 1 77
2 3929 1 77
2 3930 1 77
2 3931 1 78
2 3932 1 78
2 3933 1 78
2 3934 1 78
2 3935 1 78
2 3936 1 78
2 3937 1 78
2 3938 1 79
2 3939 1 79
2 3940 1 79
2 3941 1 79
2 3942 1 79
2 3943 1 79
2 3944 1 80
2 3945 1 80
2 3946 1 80
2 3947 1 80
2 3948 1 80
2 3949 1 80
2 3950 1 80
2 3951 1 81
2 3952 1 81
2 3953 1 81
2 3954 1 81
2 3955 1 81
2 3956 1 81
2 3957 1 81
2 3958 1 82
2 3959 1 82
2 3960 1 82
2 3961 1 82
2 3962 1 82
2 3963 1 83
2 3964 1 83
2 3965 1 83
2 3966 1 83
2 3967 1 83
2 3968 1 83
2 3969 1 84
2 3970 1 84
2 3971 1 84
2 3972 1 84
2 3973 1 84
2 3974 1 84
2 3975 1 85
2 3976 1 85
2 3977 1 85
2 3978 1 85
2 3979 1 85
2 3980 1 86
2 3981 1 86
2 3982 1 86
2 3983 1 86
2 3984 1 86
2 3985 1 86
2 3986 1 87
2 3987 1 87
2 3988 1 87
2 3989 1 87
2 3990 1 87
2 3991 1 87
2 3992 1 88
2 3993 1 88
2 3994 1 88
2 3995 1 88
2 3996 1 88
2 3997 1 89
2 3998 1 89
2 3999 1 89
2 4000 1 89
2 4001 1 89
2 4002 1 89
2 4003 1 90
2 4004 1 90
2 4005 1 90
2 4006 1 90
2 4007 1 90
2 4008 1 90
2 4009 1 91
2 4010 1 91
2 4011 1 91
2 4012 1 91
2 4013 1 91
2 4014 1 92
2 4015 1 92
2 4016 1 92
2 4017 1 92
2 4018 1 92
2 4019 1 92
2 4020 1 93
2 4021 1 93
2 4022 1 93
2 4023 1 93
2 4024 1 93
2 4025 1 94
2 4026 1 94
2 4027 1 94
2 4028 1 94
2 4029 1 94
2 4030 1 94
2 4031 1 95
2 4032 1 95
2 4033 1 95
2 4034 1 95
2 4035 1 95
2 4036 1 95
2 4037 1 96
2 4038 1 96
2 4039 1 96
2 4040 1 96
2 4041 1 96
2 4042 1 97
2 4043 1 97
2 4044 1 97
2 4045 1 98
2 4046 1 98
2 4047 1 98
2 4048 1 98
2 4049 1 103
2 4050 1 103
2 4051 1 104
2 4052 1 104
2 4053 1 105
2 4054 1 105
2 4055 1 109
2 4056 1 109
2 4057 1 111
2 4058 1 111
2 4059 1 112
2 4060 1 112
2 4061 1 115
2 4062 1 115
2 4063 1 116
2 4064 1 116
2 4065 1 120
2 4066 1 120
2 4067 1 123
2 4068 1 123
2 4069 1 126
2 4070 1 126
2 4071 1 128
2 4072 1 128
2 4073 1 129
2 4074 1 129
2 4075 1 132
2 4076 1 132
2 4077 1 133
2 4078 1 133
2 4079 1 134
2 4080 1 134
2 4081 1 138
2 4082 1 138
2 4083 1 141
2 4084 1 141
2 4085 1 142
2 4086 1 142
2 4087 1 145
2 4088 1 145
2 4089 1 148
2 4090 1 148
2 4091 1 150
2 4092 1 150
2 4093 1 151
2 4094 1 151
2 4095 1 156
2 4096 1 156
2 4097 1 159
2 4098 1 159
2 4099 1 164
2 4100 1 164
2 4101 1 164
2 4102 1 170
2 4103 1 170
2 4104 1 170
2 4105 1 172
2 4106 1 172
2 4107 1 175
2 4108 1 175
2 4109 1 178
2 4110 1 178
2 4111 1 180
2 4112 1 180
2 4113 1 181
2 4114 1 181
2 4115 1 186
2 4116 1 186
2 4117 1 189
2 4118 1 189
2 4119 1 190
2 4120 1 190
2 4121 1 193
2 4122 1 193
2 4123 1 196
2 4124 1 196
2 4125 1 198
2 4126 1 198
2 4127 1 199
2 4128 1 199
2 4129 1 204
2 4130 1 204
2 4131 1 207
2 4132 1 207
2 4133 1 212
2 4134 1 212
2 4135 1 212
2 4136 1 218
2 4137 1 218
2 4138 1 218
2 4139 1 220
2 4140 1 220
2 4141 1 223
2 4142 1 223
2 4143 1 226
2 4144 1 226
2 4145 1 228
2 4146 1 228
2 4147 1 229
2 4148 1 229
2 4149 1 234
2 4150 1 234
2 4151 1 237
2 4152 1 237
2 4153 1 238
2 4154 1 238
2 4155 1 241
2 4156 1 241
2 4157 1 244
2 4158 1 244
2 4159 1 246
2 4160 1 246
2 4161 1 247
2 4162 1 247
2 4163 1 252
2 4164 1 252
2 4165 1 255
2 4166 1 255
2 4167 1 260
2 4168 1 260
2 4169 1 260
2 4170 1 266
2 4171 1 266
2 4172 1 266
2 4173 1 268
2 4174 1 268
2 4175 1 271
2 4176 1 271
2 4177 1 274
2 4178 1 274
2 4179 1 276
2 4180 1 276
2 4181 1 277
2 4182 1 277
2 4183 1 282
2 4184 1 282
2 4185 1 285
2 4186 1 285
2 4187 1 286
2 4188 1 286
2 4189 1 289
2 4190 1 289
2 4191 1 292
2 4192 1 292
2 4193 1 294
2 4194 1 294
2 4195 1 295
2 4196 1 295
2 4197 1 300
2 4198 1 300
2 4199 1 303
2 4200 1 303
2 4201 1 308
2 4202 1 308
2 4203 1 308
2 4204 1 314
2 4205 1 314
2 4206 1 314
2 4207 1 316
2 4208 1 316
2 4209 1 319
2 4210 1 319
2 4211 1 322
2 4212 1 322
2 4213 1 324
2 4214 1 324
2 4215 1 325
2 4216 1 325
2 4217 1 330
2 4218 1 330
2 4219 1 333
2 4220 1 333
2 4221 1 334
2 4222 1 334
2 4223 1 337
2 4224 1 337
2 4225 1 340
2 4226 1 340
2 4227 1 342
2 4228 1 342
2 4229 1 343
2 4230 1 343
2 4231 1 348
2 4232 1 348
2 4233 1 351
2 4234 1 351
2 4235 1 356
2 4236 1 356
2 4237 1 356
2 4238 1 362
2 4239 1 362
2 4240 1 362
2 4241 1 364
2 4242 1 364
2 4243 1 367
2 4244 1 367
2 4245 1 370
2 4246 1 370
2 4247 1 372
2 4248 1 372
2 4249 1 373
2 4250 1 373
2 4251 1 378
2 4252 1 378
2 4253 1 381
2 4254 1 381
2 4255 1 382
2 4256 1 382
2 4257 1 385
2 4258 1 385
2 4259 1 388
2 4260 1 388
2 4261 1 390
2 4262 1 390
2 4263 1 391
2 4264 1 391
2 4265 1 396
2 4266 1 396
2 4267 1 399
2 4268 1 399
2 4269 1 404
2 4270 1 404
2 4271 1 404
2 4272 1 410
2 4273 1 410
2 4274 1 410
2 4275 1 412
2 4276 1 412
2 4277 1 415
2 4278 1 415
2 4279 1 418
2 4280 1 418
2 4281 1 420
2 4282 1 420
2 4283 1 421
2 4284 1 421
2 4285 1 426
2 4286 1 426
2 4287 1 429
2 4288 1 429
2 4289 1 430
2 4290 1 430
2 4291 1 433
2 4292 1 433
2 4293 1 436
2 4294 1 436
2 4295 1 438
2 4296 1 438
2 4297 1 439
2 4298 1 439
2 4299 1 444
2 4300 1 444
2 4301 1 447
2 4302 1 447
2 4303 1 452
2 4304 1 452
2 4305 1 452
2 4306 1 458
2 4307 1 458
2 4308 1 458
2 4309 1 460
2 4310 1 460
2 4311 1 463
2 4312 1 463
2 4313 1 466
2 4314 1 466
2 4315 1 468
2 4316 1 468
2 4317 1 469
2 4318 1 469
2 4319 1 474
2 4320 1 474
2 4321 1 477
2 4322 1 477
2 4323 1 478
2 4324 1 478
2 4325 1 481
2 4326 1 481
2 4327 1 484
2 4328 1 484
2 4329 1 486
2 4330 1 486
2 4331 1 487
2 4332 1 487
2 4333 1 492
2 4334 1 492
2 4335 1 495
2 4336 1 495
2 4337 1 500
2 4338 1 500
2 4339 1 500
2 4340 1 506
2 4341 1 506
2 4342 1 506
2 4343 1 508
2 4344 1 508
2 4345 1 511
2 4346 1 511
2 4347 1 514
2 4348 1 514
2 4349 1 516
2 4350 1 516
2 4351 1 517
2 4352 1 517
2 4353 1 522
2 4354 1 522
2 4355 1 525
2 4356 1 525
2 4357 1 526
2 4358 1 526
2 4359 1 529
2 4360 1 529
2 4361 1 532
2 4362 1 532
2 4363 1 534
2 4364 1 534
2 4365 1 535
2 4366 1 535
2 4367 1 540
2 4368 1 540
2 4369 1 543
2 4370 1 543
2 4371 1 548
2 4372 1 548
2 4373 1 548
2 4374 1 554
2 4375 1 554
2 4376 1 554
2 4377 1 556
2 4378 1 556
2 4379 1 559
2 4380 1 559
2 4381 1 562
2 4382 1 562
2 4383 1 564
2 4384 1 564
2 4385 1 565
2 4386 1 565
2 4387 1 570
2 4388 1 570
2 4389 1 573
2 4390 1 573
2 4391 1 574
2 4392 1 574
2 4393 1 577
2 4394 1 577
2 4395 1 580
2 4396 1 580
2 4397 1 582
2 4398 1 582
2 4399 1 583
2 4400 1 583
2 4401 1 588
2 4402 1 588
2 4403 1 591
2 4404 1 591
2 4405 1 596
2 4406 1 596
2 4407 1 596
2 4408 1 602
2 4409 1 602
2 4410 1 602
2 4411 1 604
2 4412 1 604
2 4413 1 607
2 4414 1 607
2 4415 1 610
2 4416 1 610
2 4417 1 612
2 4418 1 612
2 4419 1 613
2 4420 1 613
2 4421 1 618
2 4422 1 618
2 4423 1 621
2 4424 1 621
2 4425 1 622
2 4426 1 622
2 4427 1 625
2 4428 1 625
2 4429 1 628
2 4430 1 628
2 4431 1 630
2 4432 1 630
2 4433 1 631
2 4434 1 631
2 4435 1 636
2 4436 1 636
2 4437 1 639
2 4438 1 639
2 4439 1 644
2 4440 1 644
2 4441 1 644
2 4442 1 650
2 4443 1 650
2 4444 1 650
2 4445 1 652
2 4446 1 652
2 4447 1 655
2 4448 1 655
2 4449 1 658
2 4450 1 658
2 4451 1 660
2 4452 1 660
2 4453 1 661
2 4454 1 661
2 4455 1 666
2 4456 1 666
2 4457 1 669
2 4458 1 669
2 4459 1 670
2 4460 1 670
2 4461 1 673
2 4462 1 673
2 4463 1 676
2 4464 1 676
2 4465 1 678
2 4466 1 678
2 4467 1 679
2 4468 1 679
2 4469 1 684
2 4470 1 684
2 4471 1 687
2 4472 1 687
2 4473 1 692
2 4474 1 692
2 4475 1 692
2 4476 1 698
2 4477 1 698
2 4478 1 698
2 4479 1 700
2 4480 1 700
2 4481 1 703
2 4482 1 703
2 4483 1 706
2 4484 1 706
2 4485 1 708
2 4486 1 708
2 4487 1 709
2 4488 1 709
2 4489 1 714
2 4490 1 714
2 4491 1 717
2 4492 1 717
2 4493 1 718
2 4494 1 718
2 4495 1 721
2 4496 1 721
2 4497 1 724
2 4498 1 724
2 4499 1 726
2 4500 1 726
2 4501 1 727
2 4502 1 727
2 4503 1 732
2 4504 1 732
2 4505 1 735
2 4506 1 735
2 4507 1 740
2 4508 1 740
2 4509 1 740
2 4510 1 746
2 4511 1 746
2 4512 1 746
2 4513 1 748
2 4514 1 748
2 4515 1 751
2 4516 1 751
2 4517 1 754
2 4518 1 754
2 4519 1 756
2 4520 1 756
2 4521 1 757
2 4522 1 757
2 4523 1 762
2 4524 1 762
2 4525 1 765
2 4526 1 765
2 4527 1 766
2 4528 1 766
2 4529 1 769
2 4530 1 769
2 4531 1 772
2 4532 1 772
2 4533 1 774
2 4534 1 774
2 4535 1 775
2 4536 1 775
2 4537 1 780
2 4538 1 780
2 4539 1 783
2 4540 1 783
2 4541 1 788
2 4542 1 788
2 4543 1 788
2 4544 1 794
2 4545 1 794
2 4546 1 794
2 4547 1 796
2 4548 1 796
2 4549 1 799
2 4550 1 799
2 4551 1 802
2 4552 1 802
2 4553 1 804
2 4554 1 804
2 4555 1 805
2 4556 1 805
2 4557 1 810
2 4558 1 810
2 4559 1 813
2 4560 1 813
2 4561 1 814
2 4562 1 814
2 4563 1 817
2 4564 1 817
2 4565 1 820
2 4566 1 820
2 4567 1 822
2 4568 1 822
2 4569 1 823
2 4570 1 823
2 4571 1 828
2 4572 1 828
2 4573 1 831
2 4574 1 831
2 4575 1 836
2 4576 1 836
2 4577 1 836
2 4578 1 842
2 4579 1 842
2 4580 1 842
2 4581 1 844
2 4582 1 844
2 4583 1 847
2 4584 1 847
2 4585 1 850
2 4586 1 850
2 4587 1 852
2 4588 1 852
2 4589 1 853
2 4590 1 853
2 4591 1 858
2 4592 1 858
2 4593 1 861
2 4594 1 861
2 4595 1 862
2 4596 1 862
2 4597 1 865
2 4598 1 865
2 4599 1 868
2 4600 1 868
2 4601 1 870
2 4602 1 870
2 4603 1 871
2 4604 1 871
2 4605 1 876
2 4606 1 876
2 4607 1 879
2 4608 1 879
2 4609 1 884
2 4610 1 884
2 4611 1 884
2 4612 1 890
2 4613 1 890
2 4614 1 890
2 4615 1 892
2 4616 1 892
2 4617 1 895
2 4618 1 895
2 4619 1 898
2 4620 1 898
2 4621 1 900
2 4622 1 900
2 4623 1 901
2 4624 1 901
2 4625 1 906
2 4626 1 906
2 4627 1 909
2 4628 1 909
2 4629 1 910
2 4630 1 910
2 4631 1 913
2 4632 1 913
2 4633 1 916
2 4634 1 916
2 4635 1 918
2 4636 1 918
2 4637 1 919
2 4638 1 919
2 4639 1 924
2 4640 1 924
2 4641 1 927
2 4642 1 927
2 4643 1 932
2 4644 1 932
2 4645 1 932
2 4646 1 938
2 4647 1 938
2 4648 1 938
2 4649 1 940
2 4650 1 940
2 4651 1 943
2 4652 1 943
2 4653 1 946
2 4654 1 946
2 4655 1 948
2 4656 1 948
2 4657 1 949
2 4658 1 949
2 4659 1 954
2 4660 1 954
2 4661 1 957
2 4662 1 957
2 4663 1 958
2 4664 1 958
2 4665 1 961
2 4666 1 961
2 4667 1 964
2 4668 1 964
2 4669 1 966
2 4670 1 966
2 4671 1 967
2 4672 1 967
2 4673 1 972
2 4674 1 972
2 4675 1 975
2 4676 1 975
2 4677 1 980
2 4678 1 980
2 4679 1 980
2 4680 1 986
2 4681 1 986
2 4682 1 986
2 4683 1 988
2 4684 1 988
2 4685 1 991
2 4686 1 991
2 4687 1 994
2 4688 1 994
2 4689 1 996
2 4690 1 996
2 4691 1 997
2 4692 1 997
2 4693 1 1002
2 4694 1 1002
2 4695 1 1005
2 4696 1 1005
2 4697 1 1006
2 4698 1 1006
2 4699 1 1009
2 4700 1 1009
2 4701 1 1012
2 4702 1 1012
2 4703 1 1014
2 4704 1 1014
2 4705 1 1015
2 4706 1 1015
2 4707 1 1020
2 4708 1 1020
2 4709 1 1023
2 4710 1 1023
2 4711 1 1028
2 4712 1 1028
2 4713 1 1028
2 4714 1 1034
2 4715 1 1034
2 4716 1 1034
2 4717 1 1036
2 4718 1 1036
2 4719 1 1039
2 4720 1 1039
2 4721 1 1042
2 4722 1 1042
2 4723 1 1044
2 4724 1 1044
2 4725 1 1045
2 4726 1 1045
2 4727 1 1050
2 4728 1 1050
2 4729 1 1053
2 4730 1 1053
2 4731 1 1054
2 4732 1 1054
2 4733 1 1057
2 4734 1 1057
2 4735 1 1060
2 4736 1 1060
2 4737 1 1062
2 4738 1 1062
2 4739 1 1063
2 4740 1 1063
2 4741 1 1068
2 4742 1 1068
2 4743 1 1071
2 4744 1 1071
2 4745 1 1076
2 4746 1 1076
2 4747 1 1076
2 4748 1 1082
2 4749 1 1082
2 4750 1 1082
2 4751 1 1084
2 4752 1 1084
2 4753 1 1087
2 4754 1 1087
2 4755 1 1090
2 4756 1 1090
2 4757 1 1092
2 4758 1 1092
2 4759 1 1093
2 4760 1 1093
2 4761 1 1098
2 4762 1 1098
2 4763 1 1101
2 4764 1 1101
2 4765 1 1102
2 4766 1 1102
2 4767 1 1105
2 4768 1 1105
2 4769 1 1108
2 4770 1 1108
2 4771 1 1110
2 4772 1 1110
2 4773 1 1111
2 4774 1 1111
2 4775 1 1116
2 4776 1 1116
2 4777 1 1119
2 4778 1 1119
2 4779 1 1124
2 4780 1 1124
2 4781 1 1124
2 4782 1 1126
2 4783 1 1126
2 4784 1 1129
2 4785 1 1129
2 4786 1 1132
2 4787 1 1132
2 4788 1 1132
2 4789 1 1133
2 4790 1 1133
2 4791 1 1135
2 4792 1 1135
2 4793 1 1140
2 4794 1 1140
2 4795 1 1143
2 4796 1 1143
2 4797 1 1148
2 4798 1 1148
2 4799 1 1154
2 4800 1 1154
2 4801 1 1156
2 4802 1 1156
2 4803 1 1159
2 4804 1 1159
2 4805 1 1160
2 4806 1 1160
2 4807 1 1163
2 4808 1 1163
2 4809 1 1163
2 4810 1 1170
2 4811 1 1170
2 4812 1 1189
2 4813 1 1189
2 4814 1 1193
2 4815 1 1193
2 4816 1 1196
2 4817 1 1196
2 4818 1 1199
2 4819 1 1199
2 4820 1 1204
2 4821 1 1204
2 4822 1 1205
2 4823 1 1205
2 4824 1 1212
2 4825 1 1212
2 4826 1 1215
2 4827 1 1215
2 4828 1 1218
2 4829 1 1218
2 4830 1 1219
2 4831 1 1219
2 4832 1 1219
2 4833 1 1227
2 4834 1 1227
2 4835 1 1231
2 4836 1 1231
2 4837 1 1234
2 4838 1 1234
2 4839 1 1240
2 4840 1 1240
2 4841 1 1243
2 4842 1 1243
2 4843 1 1246
2 4844 1 1246
2 4845 1 1247
2 4846 1 1247
2 4847 1 1247
2 4848 1 1253
2 4849 1 1253
2 4850 1 1257
2 4851 1 1257
2 4852 1 1260
2 4853 1 1260
2 4854 1 1261
2 4855 1 1261
2 4856 1 1267
2 4857 1 1267
2 4858 1 1270
2 4859 1 1270
2 4860 1 1276
2 4861 1 1276
2 4862 1 1280
2 4863 1 1280
2 4864 1 1282
2 4865 1 1282
2 4866 1 1285
2 4867 1 1285
2 4868 1 1288
2 4869 1 1288
2 4870 1 1295
2 4871 1 1295
2 4872 1 1299
2 4873 1 1299
2 4874 1 1300
2 4875 1 1300
2 4876 1 1301
2 4877 1 1301
2 4878 1 1302
2 4879 1 1302
2 4880 1 1309
2 4881 1 1309
2 4882 1 1312
2 4883 1 1312
2 4884 1 1318
2 4885 1 1318
2 4886 1 1324
2 4887 1 1324
2 4888 1 1327
2 4889 1 1327
2 4890 1 1330
2 4891 1 1330
2 4892 1 1331
2 4893 1 1331
2 4894 1 1331
2 4895 1 1337
2 4896 1 1337
2 4897 1 1341
2 4898 1 1341
2 4899 1 1344
2 4900 1 1344
2 4901 1 1345
2 4902 1 1345
2 4903 1 1351
2 4904 1 1351
2 4905 1 1354
2 4906 1 1354
2 4907 1 1360
2 4908 1 1360
2 4909 1 1364
2 4910 1 1364
2 4911 1 1366
2 4912 1 1366
2 4913 1 1369
2 4914 1 1369
2 4915 1 1372
2 4916 1 1372
2 4917 1 1379
2 4918 1 1379
2 4919 1 1383
2 4920 1 1383
2 4921 1 1384
2 4922 1 1384
2 4923 1 1385
2 4924 1 1385
2 4925 1 1386
2 4926 1 1386
2 4927 1 1393
2 4928 1 1393
2 4929 1 1396
2 4930 1 1396
2 4931 1 1402
2 4932 1 1402
2 4933 1 1408
2 4934 1 1408
2 4935 1 1411
2 4936 1 1411
2 4937 1 1414
2 4938 1 1414
2 4939 1 1415
2 4940 1 1415
2 4941 1 1415
2 4942 1 1421
2 4943 1 1421
2 4944 1 1425
2 4945 1 1425
2 4946 1 1428
2 4947 1 1428
2 4948 1 1429
2 4949 1 1429
2 4950 1 1435
2 4951 1 1435
2 4952 1 1438
2 4953 1 1438
2 4954 1 1444
2 4955 1 1444
2 4956 1 1448
2 4957 1 1448
2 4958 1 1450
2 4959 1 1450
2 4960 1 1453
2 4961 1 1453
2 4962 1 1456
2 4963 1 1456
2 4964 1 1463
2 4965 1 1463
2 4966 1 1467
2 4967 1 1467
2 4968 1 1468
2 4969 1 1468
2 4970 1 1469
2 4971 1 1469
2 4972 1 1470
2 4973 1 1470
2 4974 1 1477
2 4975 1 1477
2 4976 1 1480
2 4977 1 1480
2 4978 1 1486
2 4979 1 1486
2 4980 1 1492
2 4981 1 1492
2 4982 1 1495
2 4983 1 1495
2 4984 1 1498
2 4985 1 1498
2 4986 1 1499
2 4987 1 1499
2 4988 1 1499
2 4989 1 1505
2 4990 1 1505
2 4991 1 1509
2 4992 1 1509
2 4993 1 1512
2 4994 1 1512
2 4995 1 1513
2 4996 1 1513
2 4997 1 1519
2 4998 1 1519
2 4999 1 1522
2 5000 1 1522
2 5001 1 1528
2 5002 1 1528
2 5003 1 1532
2 5004 1 1532
2 5005 1 1534
2 5006 1 1534
2 5007 1 1537
2 5008 1 1537
2 5009 1 1540
2 5010 1 1540
2 5011 1 1547
2 5012 1 1547
2 5013 1 1551
2 5014 1 1551
2 5015 1 1552
2 5016 1 1552
2 5017 1 1553
2 5018 1 1553
2 5019 1 1554
2 5020 1 1554
2 5021 1 1561
2 5022 1 1561
2 5023 1 1564
2 5024 1 1564
2 5025 1 1570
2 5026 1 1570
2 5027 1 1576
2 5028 1 1576
2 5029 1 1579
2 5030 1 1579
2 5031 1 1582
2 5032 1 1582
2 5033 1 1583
2 5034 1 1583
2 5035 1 1583
2 5036 1 1589
2 5037 1 1589
2 5038 1 1593
2 5039 1 1593
2 5040 1 1596
2 5041 1 1596
2 5042 1 1597
2 5043 1 1597
2 5044 1 1603
2 5045 1 1603
2 5046 1 1606
2 5047 1 1606
2 5048 1 1612
2 5049 1 1612
2 5050 1 1616
2 5051 1 1616
2 5052 1 1618
2 5053 1 1618
2 5054 1 1621
2 5055 1 1621
2 5056 1 1624
2 5057 1 1624
2 5058 1 1631
2 5059 1 1631
2 5060 1 1635
2 5061 1 1635
2 5062 1 1636
2 5063 1 1636
2 5064 1 1637
2 5065 1 1637
2 5066 1 1638
2 5067 1 1638
2 5068 1 1645
2 5069 1 1645
2 5070 1 1648
2 5071 1 1648
2 5072 1 1654
2 5073 1 1654
2 5074 1 1660
2 5075 1 1660
2 5076 1 1663
2 5077 1 1663
2 5078 1 1666
2 5079 1 1666
2 5080 1 1667
2 5081 1 1667
2 5082 1 1667
2 5083 1 1673
2 5084 1 1673
2 5085 1 1677
2 5086 1 1677
2 5087 1 1680
2 5088 1 1680
2 5089 1 1681
2 5090 1 1681
2 5091 1 1687
2 5092 1 1687
2 5093 1 1690
2 5094 1 1690
2 5095 1 1696
2 5096 1 1696
2 5097 1 1700
2 5098 1 1700
2 5099 1 1702
2 5100 1 1702
2 5101 1 1705
2 5102 1 1705
2 5103 1 1708
2 5104 1 1708
2 5105 1 1715
2 5106 1 1715
2 5107 1 1719
2 5108 1 1719
2 5109 1 1720
2 5110 1 1720
2 5111 1 1721
2 5112 1 1721
2 5113 1 1722
2 5114 1 1722
2 5115 1 1729
2 5116 1 1729
2 5117 1 1732
2 5118 1 1732
2 5119 1 1738
2 5120 1 1738
2 5121 1 1744
2 5122 1 1744
2 5123 1 1747
2 5124 1 1747
2 5125 1 1750
2 5126 1 1750
2 5127 1 1751
2 5128 1 1751
2 5129 1 1751
2 5130 1 1759
2 5131 1 1759
2 5132 1 1763
2 5133 1 1763
2 5134 1 1767
2 5135 1 1767
2 5136 1 1772
2 5137 1 1772
2 5138 1 1773
2 5139 1 1773
2 5140 1 1776
2 5141 1 1776
2 5142 1 1778
2 5143 1 1778
2 5144 1 1779
2 5145 1 1779
2 5146 1 1784
2 5147 1 1784
2 5148 1 1787
2 5149 1 1787
2 5150 1 1793
2 5151 1 1793
2 5152 1 1798
2 5153 1 1798
2 5154 1 1799
2 5155 1 1799
2 5156 1 1802
2 5157 1 1802
2 5158 1 1804
2 5159 1 1804
2 5160 1 1820
2 5161 1 1820
2 5162 1 1823
2 5163 1 1823
2 5164 1 1829
2 5165 1 1829
2 5166 1 1829
2 5167 1 1830
2 5168 1 1830
2 5169 1 1830
2 5170 1 1830
2 5171 1 1830
2 5172 1 1832
2 5173 1 1832
2 5174 1 1833
2 5175 1 1833
2 5176 1 1834
2 5177 1 1834
2 5178 1 1841
2 5179 1 1841
2 5180 1 1842
2 5181 1 1842
2 5182 1 1849
2 5183 1 1849
2 5184 1 1849
2 5185 1 1855
2 5186 1 1855
2 5187 1 1856
2 5188 1 1856
2 5189 1 1857
2 5190 1 1857
2 5191 1 1859
2 5192 1 1859
2 5193 1 1861
2 5194 1 1861
2 5195 1 1862
2 5196 1 1862
2 5197 1 1873
2 5198 1 1873
2 5199 1 1875
2 5200 1 1875
2 5201 1 1877
2 5202 1 1877
2 5203 1 1880
2 5204 1 1880
2 5205 1 1880
2 5206 1 1880
2 5207 1 1885
2 5208 1 1885
2 5209 1 1886
2 5210 1 1886
2 5211 1 1890
2 5212 1 1890
2 5213 1 1899
2 5214 1 1899
2 5215 1 1902
2 5216 1 1902
2 5217 1 1903
2 5218 1 1903
2 5219 1 1906
2 5220 1 1906
2 5221 1 1906
2 5222 1 1908
2 5223 1 1908
2 5224 1 1910
2 5225 1 1910
2 5226 1 1912
2 5227 1 1912
2 5228 1 1919
2 5229 1 1919
2 5230 1 1920
2 5231 1 1920
2 5232 1 1926
2 5233 1 1926
2 5234 1 1929
2 5235 1 1929
2 5236 1 1930
2 5237 1 1930
2 5238 1 1935
2 5239 1 1935
2 5240 1 1939
2 5241 1 1939
2 5242 1 1939
2 5243 1 1939
2 5244 1 1943
2 5245 1 1943
2 5246 1 1946
2 5247 1 1946
2 5248 1 1947
2 5249 1 1947
2 5250 1 1950
2 5251 1 1950
2 5252 1 1950
2 5253 1 1953
2 5254 1 1953
2 5255 1 1957
2 5256 1 1957
2 5257 1 1958
2 5258 1 1958
2 5259 1 1960
2 5260 1 1960
2 5261 1 1962
2 5262 1 1962
2 5263 1 1964
2 5264 1 1964
2 5265 1 1967
2 5266 1 1967
2 5267 1 1967
2 5268 1 1967
2 5269 1 1969
2 5270 1 1969
2 5271 1 1971
2 5272 1 1971
2 5273 1 1975
2 5274 1 1975
2 5275 1 1984
2 5276 1 1984
2 5277 1 1985
2 5278 1 1985
2 5279 1 1991
2 5280 1 1991
2 5281 1 1994
2 5282 1 1994
2 5283 1 1995
2 5284 1 1995
2 5285 1 1998
2 5286 1 1998
2 5287 1 2000
2 5288 1 2000
2 5289 1 2002
2 5290 1 2002
2 5291 1 2004
2 5292 1 2004
2 5293 1 2006
2 5294 1 2006
2 5295 1 2009
2 5296 1 2009
2 5297 1 2009
2 5298 1 2009
2 5299 1 2014
2 5300 1 2014
2 5301 1 2015
2 5302 1 2015
2 5303 1 2019
2 5304 1 2019
2 5305 1 2028
2 5306 1 2028
2 5307 1 2031
2 5308 1 2031
2 5309 1 2032
2 5310 1 2032
2 5311 1 2035
2 5312 1 2035
2 5313 1 2035
2 5314 1 2037
2 5315 1 2037
2 5316 1 2039
2 5317 1 2039
2 5318 1 2041
2 5319 1 2041
2 5320 1 2048
2 5321 1 2048
2 5322 1 2049
2 5323 1 2049
2 5324 1 2055
2 5325 1 2055
2 5326 1 2058
2 5327 1 2058
2 5328 1 2059
2 5329 1 2059
2 5330 1 2064
2 5331 1 2064
2 5332 1 2068
2 5333 1 2068
2 5334 1 2068
2 5335 1 2068
2 5336 1 2072
2 5337 1 2072
2 5338 1 2075
2 5339 1 2075
2 5340 1 2076
2 5341 1 2076
2 5342 1 2079
2 5343 1 2079
2 5344 1 2079
2 5345 1 2082
2 5346 1 2082
2 5347 1 2086
2 5348 1 2086
2 5349 1 2087
2 5350 1 2087
2 5351 1 2089
2 5352 1 2089
2 5353 1 2091
2 5354 1 2091
2 5355 1 2093
2 5356 1 2093
2 5357 1 2096
2 5358 1 2096
2 5359 1 2096
2 5360 1 2096
2 5361 1 2098
2 5362 1 2098
2 5363 1 2100
2 5364 1 2100
2 5365 1 2104
2 5366 1 2104
2 5367 1 2113
2 5368 1 2113
2 5369 1 2114
2 5370 1 2114
2 5371 1 2120
2 5372 1 2120
2 5373 1 2123
2 5374 1 2123
2 5375 1 2124
2 5376 1 2124
2 5377 1 2127
2 5378 1 2127
2 5379 1 2127
2 5380 1 2127
2 5381 1 2131
2 5382 1 2131
2 5383 1 2134
2 5384 1 2134
2 5385 1 2135
2 5386 1 2135
2 5387 1 2138
2 5388 1 2138
2 5389 1 2138
2 5390 1 2138
2 5391 1 2142
2 5392 1 2142
2 5393 1 2144
2 5394 1 2144
2 5395 1 2153
2 5396 1 2153
2 5397 1 2156
2 5398 1 2156
2 5399 1 2157
2 5400 1 2157
2 5401 1 2160
2 5402 1 2160
2 5403 1 2160
2 5404 1 2160
2 5405 1 2162
2 5406 1 2162
2 5407 1 2164
2 5408 1 2164
2 5409 1 2168
2 5410 1 2168
2 5411 1 2177
2 5412 1 2177
2 5413 1 2178
2 5414 1 2178
2 5415 1 2184
2 5416 1 2184
2 5417 1 2187
2 5418 1 2187
2 5419 1 2188
2 5420 1 2188
2 5421 1 2191
2 5422 1 2191
2 5423 1 2191
2 5424 1 2193
2 5425 1 2193
2 5426 1 2195
2 5427 1 2195
2 5428 1 2197
2 5429 1 2197
2 5430 1 2199
2 5431 1 2199
2 5432 1 2202
2 5433 1 2202
2 5434 1 2202
2 5435 1 2202
2 5436 1 2206
2 5437 1 2206
2 5438 1 2208
2 5439 1 2208
2 5440 1 2217
2 5441 1 2217
2 5442 1 2220
2 5443 1 2220
2 5444 1 2221
2 5445 1 2221
2 5446 1 2224
2 5447 1 2224
2 5448 1 2224
2 5449 1 2224
2 5450 1 2226
2 5451 1 2226
2 5452 1 2228
2 5453 1 2228
2 5454 1 2232
2 5455 1 2232
2 5456 1 2241
2 5457 1 2241
2 5458 1 2242
2 5459 1 2242
2 5460 1 2248
2 5461 1 2248
2 5462 1 2251
2 5463 1 2251
2 5464 1 2252
2 5465 1 2252
2 5466 1 2255
2 5467 1 2255
2 5468 1 2255
2 5469 1 2255
2 5470 1 2259
2 5471 1 2259
2 5472 1 2262
2 5473 1 2262
2 5474 1 2263
2 5475 1 2263
2 5476 1 2266
2 5477 1 2266
2 5478 1 2266
2 5479 1 2266
2 5480 1 2270
2 5481 1 2270
2 5482 1 2272
2 5483 1 2272
2 5484 1 2281
2 5485 1 2281
2 5486 1 2284
2 5487 1 2284
2 5488 1 2285
2 5489 1 2285
2 5490 1 2288
2 5491 1 2288
2 5492 1 2288
2 5493 1 2288
2 5494 1 2290
2 5495 1 2290
2 5496 1 2292
2 5497 1 2292
2 5498 1 2296
2 5499 1 2296
2 5500 1 2305
2 5501 1 2305
2 5502 1 2306
2 5503 1 2306
2 5504 1 2312
2 5505 1 2312
2 5506 1 2315
2 5507 1 2315
2 5508 1 2316
2 5509 1 2316
2 5510 1 2319
2 5511 1 2319
2 5512 1 2319
2 5513 1 2319
2 5514 1 2323
2 5515 1 2323
2 5516 1 2326
2 5517 1 2326
2 5518 1 2327
2 5519 1 2327
2 5520 1 2330
2 5521 1 2330
2 5522 1 2330
2 5523 1 2332
2 5524 1 2332
2 5525 1 2334
2 5526 1 2334
2 5527 1 2336
2 5528 1 2336
2 5529 1 2345
2 5530 1 2345
2 5531 1 2347
2 5532 1 2347
2 5533 1 2349
2 5534 1 2349
2 5535 1 2352
2 5536 1 2352
2 5537 1 2352
2 5538 1 2352
2 5539 1 2354
2 5540 1 2354
2 5541 1 2356
2 5542 1 2356
2 5543 1 2360
2 5544 1 2360
2 5545 1 2369
2 5546 1 2369
2 5547 1 2370
2 5548 1 2370
2 5549 1 2376
2 5550 1 2376
2 5551 1 2379
2 5552 1 2379
2 5553 1 2380
2 5554 1 2380
2 5555 1 2383
2 5556 1 2383
2 5557 1 2383
2 5558 1 2383
2 5559 1 2387
2 5560 1 2387
2 5561 1 2390
2 5562 1 2390
2 5563 1 2391
2 5564 1 2391
2 5565 1 2394
2 5566 1 2394
2 5567 1 2394
2 5568 1 2394
2 5569 1 2398
2 5570 1 2398
2 5571 1 2400
2 5572 1 2400
2 5573 1 2409
2 5574 1 2409
2 5575 1 2412
2 5576 1 2412
2 5577 1 2413
2 5578 1 2413
2 5579 1 2416
2 5580 1 2416
2 5581 1 2416
2 5582 1 2416
2 5583 1 2418
2 5584 1 2418
2 5585 1 2420
2 5586 1 2420
2 5587 1 2424
2 5588 1 2424
2 5589 1 2433
2 5590 1 2433
2 5591 1 2434
2 5592 1 2434
2 5593 1 2440
2 5594 1 2440
2 5595 1 2443
2 5596 1 2443
2 5597 1 2444
2 5598 1 2444
2 5599 1 2447
2 5600 1 2447
2 5601 1 2447
2 5602 1 2447
2 5603 1 2451
2 5604 1 2451
2 5605 1 2454
2 5606 1 2454
2 5607 1 2455
2 5608 1 2455
2 5609 1 2458
2 5610 1 2458
2 5611 1 2458
2 5612 1 2460
2 5613 1 2460
2 5614 1 2462
2 5615 1 2462
2 5616 1 2464
2 5617 1 2464
2 5618 1 2473
2 5619 1 2473
2 5620 1 2475
2 5621 1 2475
2 5622 1 2477
2 5623 1 2477
2 5624 1 2480
2 5625 1 2480
2 5626 1 2480
2 5627 1 2480
2 5628 1 2482
2 5629 1 2482
2 5630 1 2484
2 5631 1 2484
2 5632 1 2488
2 5633 1 2488
2 5634 1 2497
2 5635 1 2497
2 5636 1 2498
2 5637 1 2498
2 5638 1 2504
2 5639 1 2504
2 5640 1 2507
2 5641 1 2507
2 5642 1 2508
2 5643 1 2508
2 5644 1 2511
2 5645 1 2511
2 5646 1 2511
2 5647 1 2511
2 5648 1 2515
2 5649 1 2515
2 5650 1 2518
2 5651 1 2518
2 5652 1 2519
2 5653 1 2519
2 5654 1 2522
2 5655 1 2522
2 5656 1 2522
2 5657 1 2522
2 5658 1 2526
2 5659 1 2526
2 5660 1 2528
2 5661 1 2528
2 5662 1 2537
2 5663 1 2537
2 5664 1 2540
2 5665 1 2540
2 5666 1 2541
2 5667 1 2541
2 5668 1 2544
2 5669 1 2544
2 5670 1 2544
2 5671 1 2544
2 5672 1 2546
2 5673 1 2546
2 5674 1 2548
2 5675 1 2548
2 5676 1 2552
2 5677 1 2552
2 5678 1 2561
2 5679 1 2561
2 5680 1 2562
2 5681 1 2562
2 5682 1 2568
2 5683 1 2568
2 5684 1 2571
2 5685 1 2571
2 5686 1 2572
2 5687 1 2572
2 5688 1 2575
2 5689 1 2575
2 5690 1 2575
2 5691 1 2575
2 5692 1 2579
2 5693 1 2579
2 5694 1 2582
2 5695 1 2582
2 5696 1 2583
2 5697 1 2583
2 5698 1 2586
2 5699 1 2586
2 5700 1 2586
2 5701 1 2588
2 5702 1 2588
2 5703 1 2590
2 5704 1 2590
2 5705 1 2592
2 5706 1 2592
2 5707 1 2601
2 5708 1 2601
2 5709 1 2603
2 5710 1 2603
2 5711 1 2605
2 5712 1 2605
2 5713 1 2608
2 5714 1 2608
2 5715 1 2608
2 5716 1 2608
2 5717 1 2610
2 5718 1 2610
2 5719 1 2612
2 5720 1 2612
2 5721 1 2616
2 5722 1 2616
2 5723 1 2625
2 5724 1 2625
2 5725 1 2626
2 5726 1 2626
2 5727 1 2632
2 5728 1 2632
2 5729 1 2635
2 5730 1 2635
2 5731 1 2636
2 5732 1 2636
2 5733 1 2639
2 5734 1 2639
2 5735 1 2639
2 5736 1 2639
2 5737 1 2643
2 5738 1 2643
2 5739 1 2646
2 5740 1 2646
2 5741 1 2647
2 5742 1 2647
2 5743 1 2650
2 5744 1 2650
2 5745 1 2650
2 5746 1 2650
2 5747 1 2654
2 5748 1 2654
2 5749 1 2656
2 5750 1 2656
2 5751 1 2665
2 5752 1 2665
2 5753 1 2668
2 5754 1 2668
2 5755 1 2669
2 5756 1 2669
2 5757 1 2672
2 5758 1 2672
2 5759 1 2672
2 5760 1 2672
2 5761 1 2674
2 5762 1 2674
2 5763 1 2676
2 5764 1 2676
2 5765 1 2678
2 5766 1 2678
2 5767 1 2685
2 5768 1 2685
2 5769 1 2686
2 5770 1 2686
2 5771 1 2689
2 5772 1 2689
2 5773 1 2690
2 5774 1 2690
2 5775 1 2693
2 5776 1 2693
2 5777 1 2693
2 5778 1 2693
2 5779 1 2704
2 5780 1 2704
2 5781 1 2707
2 5782 1 2707
2 5783 1 2710
2 5784 1 2710
2 5785 1 2711
2 5786 1 2711
2 5787 1 2714
2 5788 1 2714
2 5789 1 2714
2 5790 1 2716
2 5791 1 2716
2 5792 1 2718
2 5793 1 2718
2 5794 1 2720
2 5795 1 2720
2 5796 1 2733
2 5797 1 2733
2 5798 1 2735
2 5799 1 2735
2 5800 1 2737
2 5801 1 2737
2 5802 1 2740
2 5803 1 2740
2 5804 1 2741
2 5805 1 2741
2 5806 1 2743
2 5807 1 2743
2 5808 1 2746
2 5809 1 2746
2 5810 1 2746
2 5811 1 2746
2 5812 1 2748
2 5813 1 2748
2 5814 1 2750
2 5815 1 2750
2 5816 1 2753
2 5817 1 2753
2 5818 1 2754
2 5819 1 2754
2 5820 1 2757
2 5821 1 2757
2 5822 1 2757
2 5823 1 2768
2 5824 1 2768
2 5825 1 2771
2 5826 1 2771
2 5827 1 2774
2 5828 1 2774
2 5829 1 2775
2 5830 1 2775
2 5831 1 2779
2 5832 1 2779
2 5833 1 2780
2 5834 1 2780
2 5835 1 2797
2 5836 1 2797
2 5837 1 2808
2 5838 1 2808
2 5839 1 2811
2 5840 1 2811
2 5841 1 2813
2 5842 1 2813
2 5843 1 2815
2 5844 1 2815
2 5845 1 2817
2 5846 1 2817
2 5847 1 2818
2 5848 1 2818
2 5849 1 2819
2 5850 1 2819
2 5851 1 2819
2 5852 1 2822
2 5853 1 2822
2 5854 1 2823
2 5855 1 2823
2 5856 1 2826
2 5857 1 2826
2 5858 1 2829
2 5859 1 2829
2 5860 1 2831
2 5861 1 2831
2 5862 1 2834
2 5863 1 2834
2 5864 1 2837
2 5865 1 2837
2 5866 1 2839
2 5867 1 2839
2 5868 1 2842
2 5869 1 2842
2 5870 1 2845
2 5871 1 2845
2 5872 1 2847
2 5873 1 2847
2 5874 1 2850
2 5875 1 2850
2 5876 1 2853
2 5877 1 2853
2 5878 1 2855
2 5879 1 2855
2 5880 1 2858
2 5881 1 2858
2 5882 1 2861
2 5883 1 2861
2 5884 1 2863
2 5885 1 2863
2 5886 1 2866
2 5887 1 2866
2 5888 1 2869
2 5889 1 2869
2 5890 1 2871
2 5891 1 2871
2 5892 1 2874
2 5893 1 2874
2 5894 1 2877
2 5895 1 2877
2 5896 1 2879
2 5897 1 2879
2 5898 1 2882
2 5899 1 2882
2 5900 1 2885
2 5901 1 2885
2 5902 1 2887
2 5903 1 2887
2 5904 1 2890
2 5905 1 2890
2 5906 1 2893
2 5907 1 2893
2 5908 1 2895
2 5909 1 2895
2 5910 1 2898
2 5911 1 2898
2 5912 1 2901
2 5913 1 2901
2 5914 1 2903
2 5915 1 2903
2 5916 1 2906
2 5917 1 2906
2 5918 1 2909
2 5919 1 2909
2 5920 1 2911
2 5921 1 2911
2 5922 1 2914
2 5923 1 2914
2 5924 1 2917
2 5925 1 2917
2 5926 1 2919
2 5927 1 2919
2 5928 1 2920
2 5929 1 2920
2 5930 1 2926
2 5931 1 2926
2 5932 1 2929
2 5933 1 2929
2 5934 1 2929
2 5935 1 2930
2 5936 1 2930
2 5937 1 2936
2 5938 1 2936
2 5939 1 2939
2 5940 1 2939
2 5941 1 2939
2 5942 1 2941
2 5943 1 2941
2 5944 1 2941
2 5945 1 2941
2 5946 1 2942
2 5947 1 2942
2 5948 1 2948
2 5949 1 2948
2 5950 1 2951
2 5951 1 2951
2 5952 1 2951
2 5953 1 2953
2 5954 1 2953
2 5955 1 2953
2 5956 1 2953
2 5957 1 2954
2 5958 1 2954
2 5959 1 2960
2 5960 1 2960
2 5961 1 2963
2 5962 1 2963
2 5963 1 2963
2 5964 1 2963
2 5965 1 2965
2 5966 1 2965
2 5967 1 2965
2 5968 1 2966
2 5969 1 2966
2 5970 1 2972
2 5971 1 2972
2 5972 1 2975
2 5973 1 2975
2 5974 1 2975
2 5975 1 2975
2 5976 1 2977
2 5977 1 2977
2 5978 1 2977
2 5979 1 2977
2 5980 1 2978
2 5981 1 2978
2 5982 1 2984
2 5983 1 2984
2 5984 1 2987
2 5985 1 2987
2 5986 1 2987
2 5987 1 2987
2 5988 1 2989
2 5989 1 2989
2 5990 1 2989
2 5991 1 2989
2 5992 1 2990
2 5993 1 2990
2 5994 1 2996
2 5995 1 2996
2 5996 1 2999
2 5997 1 2999
2 5998 1 2999
2 5999 1 3001
2 6000 1 3001
2 6001 1 3001
2 6002 1 3001
2 6003 1 3002
2 6004 1 3002
2 6005 1 3008
2 6006 1 3008
2 6007 1 3011
2 6008 1 3011
2 6009 1 3011
2 6010 1 3011
2 6011 1 3013
2 6012 1 3013
2 6013 1 3013
2 6014 1 3014
2 6015 1 3014
2 6016 1 3020
2 6017 1 3020
2 6018 1 3023
2 6019 1 3023
2 6020 1 3023
2 6021 1 3023
2 6022 1 3024
2 6023 1 3024
2 6024 1 3026
2 6025 1 3026
2 6026 1 3026
2 6027 1 3026
2 6028 1 3027
2 6029 1 3027
2 6030 1 3033
2 6031 1 3033
2 6032 1 3036
2 6033 1 3036
2 6034 1 3036
2 6035 1 3036
2 6036 1 3038
2 6037 1 3038
2 6038 1 3038
2 6039 1 3038
2 6040 1 3039
2 6041 1 3039
2 6042 1 3045
2 6043 1 3045
2 6044 1 3048
2 6045 1 3048
2 6046 1 3048
2 6047 1 3048
2 6048 1 3050
2 6049 1 3050
2 6050 1 3050
2 6051 1 3050
2 6052 1 3051
2 6053 1 3051
2 6054 1 3057
2 6055 1 3057
2 6056 1 3060
2 6057 1 3060
2 6058 1 3060
2 6059 1 3062
2 6060 1 3062
2 6061 1 3062
2 6062 1 3062
2 6063 1 3063
2 6064 1 3063
2 6065 1 3069
2 6066 1 3069
2 6067 1 3072
2 6068 1 3072
2 6069 1 3072
2 6070 1 3075
2 6071 1 3075
2 6072 1 3081
2 6073 1 3081
2 6074 1 3085
2 6075 1 3085
2 6076 1 3088
2 6077 1 3088
2 6078 1 3091
2 6079 1 3091
2 6080 1 3096
2 6081 1 3096
2 6082 1 3098
2 6083 1 3098
2 6084 1 3098
2 6085 1 3100
2 6086 1 3100
2 6087 1 3101
2 6088 1 3101
2 6089 1 3104
2 6090 1 3104
2 6091 1 3105
2 6092 1 3105
2 6093 1 3108
2 6094 1 3108
2 6095 1 3111
2 6096 1 3111
2 6097 1 3118
2 6098 1 3118
2 6099 1 3121
2 6100 1 3121
2 6101 1 3123
2 6102 1 3123
2 6103 1 3126
2 6104 1 3126
2 6105 1 3129
2 6106 1 3129
2 6107 1 3133
2 6108 1 3133
2 6109 1 3134
2 6110 1 3134
2 6111 1 3137
2 6112 1 3137
2 6113 1 3138
2 6114 1 3138
2 6115 1 3141
2 6116 1 3141
2 6117 1 3142
2 6118 1 3142
2 6119 1 3144
2 6120 1 3144
2 6121 1 3144
2 6122 1 3144
2 6123 1 3147
2 6124 1 3147
2 6125 1 3147
2 6126 1 3149
2 6127 1 3149
2 6128 1 3154
2 6129 1 3154
2 6130 1 3155
2 6131 1 3155
2 6132 1 3158
2 6133 1 3158
2 6134 1 3160
2 6135 1 3160
2 6136 1 3162
2 6137 1 3162
2 6138 1 3163
2 6139 1 3163
2 6140 1 3167
2 6141 1 3167
2 6142 1 3170
2 6143 1 3170
2 6144 1 3174
2 6145 1 3174
2 6146 1 3175
2 6147 1 3175
2 6148 1 3178
2 6149 1 3178
2 6150 1 3179
2 6151 1 3179
2 6152 1 3182
2 6153 1 3182
2 6154 1 3185
2 6155 1 3185
2 6156 1 3189
2 6157 1 3189
2 6158 1 3192
2 6159 1 3192
2 6160 1 3193
2 6161 1 3193
2 6162 1 3196
2 6163 1 3196
2 6164 1 3197
2 6165 1 3197
2 6166 1 3200
2 6167 1 3200
2 6168 1 3201
2 6169 1 3201
2 6170 1 3204
2 6171 1 3204
2 6172 1 3207
2 6173 1 3207
2 6174 1 3209
2 6175 1 3209
2 6176 1 3210
2 6177 1 3210
2 6178 1 3216
2 6179 1 3216
2 6180 1 3219
2 6181 1 3219
2 6182 1 3219
2 6183 1 3220
2 6184 1 3220
2 6185 1 3221
2 6186 1 3221
2 6187 1 3221
2 6188 1 3222
2 6189 1 3222
2 6190 1 3225
2 6191 1 3225
2 6192 1 3232
2 6193 1 3232
2 6194 1 3234
2 6195 1 3234
2 6196 1 3235
2 6197 1 3235
2 6198 1 3236
2 6199 1 3236
2 6200 1 3245
2 6201 1 3245
2 6202 1 3245
2 6203 1 3246
2 6204 1 3246
2 6205 1 3253
2 6206 1 3253
2 6207 1 3254
2 6208 1 3254
2 6209 1 3255
2 6210 1 3255
2 6211 1 3255
2 6212 1 3256
2 6213 1 3256
2 6214 1 3263
2 6215 1 3263
2 6216 1 3263
2 6217 1 3264
2 6218 1 3264
2 6219 1 3269
2 6220 1 3269
2 6221 1 3270
2 6222 1 3270
2 6223 1 3276
2 6224 1 3276
2 6225 1 3281
2 6226 1 3281
2 6227 1 3282
2 6228 1 3282
2 6229 1 3285
2 6230 1 3285
2 6231 1 3285
2 6232 1 3286
2 6233 1 3286
2 6234 1 3291
2 6235 1 3291
2 6236 1 3292
2 6237 1 3292
2 6238 1 3295
2 6239 1 3295
2 6240 1 3301
2 6241 1 3301
2 6242 1 3302
2 6243 1 3302
2 6244 1 3305
2 6245 1 3305
2 6246 1 3306
2 6247 1 3306
2 6248 1 3309
2 6249 1 3309
2 6250 1 3309
2 6251 1 3310
2 6252 1 3310
2 6253 1 3315
2 6254 1 3315
2 6255 1 3346
2 6256 1 3346
2 6257 1 3350
2 6258 1 3350
0 50 5 5 1 49
0 51 5 6 1 3449
0 52 5 6 1 3454
0 53 5 6 1 3460
0 54 5 6 1 3466
0 55 5 5 1 3472
0 56 5 6 1 3479
0 57 5 6 1 3486
0 58 5 5 1 3492
0 59 5 6 1 3499
0 60 5 6 1 3505
0 61 5 5 1 3511
0 62 5 6 1 3518
0 63 5 6 1 3525
0 64 5 5 1 3531
0 65 5 6 1 3538
0 66 5 6 1 3544
0 67 5 5 1 3550
0 68 5 6 1 3557
0 69 5 7 1 3564
0 70 5 6 1 3570
0 71 5 7 1 3577
0 72 5 7 1 3583
0 73 5 6 1 3589
0 74 5 7 1 3596
0 75 5 7 1 3603
0 76 5 6 1 3609
0 77 5 7 1 3616
0 78 5 7 1 3622
0 79 5 6 1 3628
0 80 5 7 1 3635
0 81 5 7 1 3642
0 82 5 5 1 3648
0 83 5 6 1 3655
0 84 5 6 1 3661
0 85 5 5 1 3667
0 86 5 6 1 3674
0 87 5 6 1 3681
0 88 5 5 1 3687
0 89 5 6 1 3694
0 90 5 6 1 3700
0 91 5 5 1 3706
0 92 5 6 1 3713
0 93 5 5 1 3720
0 94 5 6 1 3727
0 95 5 6 1 3734
0 96 5 5 1 3742
0 97 5 3 1 3750
0 98 5 4 1 3757
0 99 7 1 2 3743 4045
0 100 5 1 1 99
0 101 7 1 2 4037 3751
0 102 7 1 2 3758 101
0 103 5 2 1 102
0 104 7 2 2 100 4049
0 105 7 2 2 4031 4051
0 106 5 1 1 4053
0 107 7 1 2 3752 4054
0 108 5 1 1 107
0 109 7 2 2 4042 3759
0 110 5 1 1 4055
0 111 7 2 2 4038 4056
0 112 5 2 1 4057
0 113 7 1 2 3735 4058
0 114 5 1 1 113
0 115 7 2 2 108 114
0 116 5 2 1 4061
0 117 7 1 2 3753 4050
0 118 7 1 2 106 117
0 119 5 1 1 118
0 120 7 2 2 4059 119
0 121 5 1 1 4065
0 122 7 1 2 4032 121
0 123 5 2 1 122
0 124 7 1 2 3736 4066
0 125 5 1 1 124
0 126 7 2 2 4067 125
0 127 5 1 1 4069
0 128 7 2 2 4025 4070
0 129 5 2 1 4071
0 130 7 1 2 4052 4068
0 131 5 1 1 130
0 132 7 2 2 3754 4046
0 133 5 2 1 4075
0 134 7 2 2 3744 4076
0 135 5 1 1 4079
0 136 7 1 2 4033 4080
0 137 5 1 1 136
0 138 7 2 2 131 137
0 139 5 1 1 4081
0 140 7 1 2 4073 4082
0 141 5 2 1 140
0 142 7 2 2 4062 4083
0 143 5 1 1 4085
0 144 7 1 2 4026 143
0 145 5 2 1 144
0 146 7 1 2 3728 4086
0 147 5 1 1 146
0 148 7 2 2 4087 147
0 149 5 1 1 4089
0 150 7 2 2 4020 4090
0 151 5 2 1 4091
0 152 7 1 2 127 4088
0 153 5 1 1 152
0 154 7 1 2 4063 4072
0 155 5 1 1 154
0 156 7 2 2 153 155
0 157 5 1 1 4095
0 158 7 1 2 4093 157
0 159 5 2 1 158
0 160 7 1 2 4064 4074
0 161 5 1 1 160
0 162 7 1 2 139 161
0 163 5 1 1 162
0 164 7 3 2 4084 163
0 165 5 1 1 4099
0 166 7 1 2 4094 4100
0 167 5 1 1 166
0 168 7 1 2 4096 167
0 169 5 1 1 168
0 170 7 3 2 4097 169
0 171 5 1 1 4102
0 172 7 2 2 4098 165
0 173 5 1 1 4105
0 174 7 1 2 4021 173
0 175 5 2 1 174
0 176 7 1 2 3721 4106
0 177 5 1 1 176
0 178 7 2 2 4107 177
0 179 5 1 1 4109
0 180 7 2 2 4014 4110
0 181 5 2 1 4111
0 182 7 1 2 149 4108
0 183 5 1 1 182
0 184 7 1 2 4092 4101
0 185 5 1 1 184
0 186 7 2 2 183 185
0 187 5 1 1 4115
0 188 7 1 2 4113 187
0 189 5 2 1 188
0 190 7 2 2 171 4117
0 191 5 1 1 4119
0 192 7 1 2 4015 191
0 193 5 2 1 192
0 194 7 1 2 3714 4120
0 195 5 1 1 194
0 196 7 2 2 4121 195
0 197 5 1 1 4123
0 198 7 2 2 4009 4124
0 199 5 2 1 4125
0 200 7 1 2 179 4122
0 201 5 1 1 200
0 202 7 1 2 4103 4112
0 203 5 1 1 202
0 204 7 2 2 201 203
0 205 5 1 1 4129
0 206 7 1 2 4127 205
0 207 5 2 1 206
0 208 7 1 2 4104 4114
0 209 5 1 1 208
0 210 7 1 2 4116 209
0 211 5 1 1 210
0 212 7 3 2 4118 211
0 213 5 1 1 4133
0 214 7 1 2 4128 4134
0 215 5 1 1 214
0 216 7 1 2 4130 215
0 217 5 1 1 216
0 218 7 3 2 4131 217
0 219 5 1 1 4136
0 220 7 2 2 4132 213
0 221 5 1 1 4139
0 222 7 1 2 4010 221
0 223 5 2 1 222
0 224 7 1 2 3707 4140
0 225 5 1 1 224
0 226 7 2 2 4141 225
0 227 5 1 1 4143
0 228 7 2 2 4003 4144
0 229 5 2 1 4145
0 230 7 1 2 197 4142
0 231 5 1 1 230
0 232 7 1 2 4126 4135
0 233 5 1 1 232
0 234 7 2 2 231 233
0 235 5 1 1 4149
0 236 7 1 2 4147 235
0 237 5 2 1 236
0 238 7 2 2 219 4151
0 239 5 1 1 4153
0 240 7 1 2 4004 239
0 241 5 2 1 240
0 242 7 1 2 3701 4154
0 243 5 1 1 242
0 244 7 2 2 4155 243
0 245 5 1 1 4157
0 246 7 2 2 3997 4158
0 247 5 2 1 4159
0 248 7 1 2 227 4156
0 249 5 1 1 248
0 250 7 1 2 4137 4146
0 251 5 1 1 250
0 252 7 2 2 249 251
0 253 5 1 1 4163
0 254 7 1 2 4161 253
0 255 5 2 1 254
0 256 7 1 2 4138 4148
0 257 5 1 1 256
0 258 7 1 2 4150 257
0 259 5 1 1 258
0 260 7 3 2 4152 259
0 261 5 1 1 4167
0 262 7 1 2 4162 4168
0 263 5 1 1 262
0 264 7 1 2 4164 263
0 265 5 1 1 264
0 266 7 3 2 4165 265
0 267 5 1 1 4170
0 268 7 2 2 4166 261
0 269 5 1 1 4173
0 270 7 1 2 3998 269
0 271 5 2 1 270
0 272 7 1 2 3695 4174
0 273 5 1 1 272
0 274 7 2 2 4175 273
0 275 5 1 1 4177
0 276 7 2 2 3992 4178
0 277 5 2 1 4179
0 278 7 1 2 245 4176
0 279 5 1 1 278
0 280 7 1 2 4160 4169
0 281 5 1 1 280
0 282 7 2 2 279 281
0 283 5 1 1 4183
0 284 7 1 2 4181 283
0 285 5 2 1 284
0 286 7 2 2 267 4185
0 287 5 1 1 4187
0 288 7 1 2 3993 287
0 289 5 2 1 288
0 290 7 1 2 3688 4188
0 291 5 1 1 290
0 292 7 2 2 4189 291
0 293 5 1 1 4191
0 294 7 2 2 3986 4192
0 295 5 2 1 4193
0 296 7 1 2 275 4190
0 297 5 1 1 296
0 298 7 1 2 4171 4180
0 299 5 1 1 298
0 300 7 2 2 297 299
0 301 5 1 1 4197
0 302 7 1 2 4195 301
0 303 5 2 1 302
0 304 7 1 2 4172 4182
0 305 5 1 1 304
0 306 7 1 2 4184 305
0 307 5 1 1 306
0 308 7 3 2 4186 307
0 309 5 1 1 4201
0 310 7 1 2 4196 4202
0 311 5 1 1 310
0 312 7 1 2 4198 311
0 313 5 1 1 312
0 314 7 3 2 4199 313
0 315 5 1 1 4204
0 316 7 2 2 4200 309
0 317 5 1 1 4207
0 318 7 1 2 3987 317
0 319 5 2 1 318
0 320 7 1 2 3682 4208
0 321 5 1 1 320
0 322 7 2 2 4209 321
0 323 5 1 1 4211
0 324 7 2 2 3980 4212
0 325 5 2 1 4213
0 326 7 1 2 293 4210
0 327 5 1 1 326
0 328 7 1 2 4194 4203
0 329 5 1 1 328
0 330 7 2 2 327 329
0 331 5 1 1 4217
0 332 7 1 2 4215 331
0 333 5 2 1 332
0 334 7 2 2 315 4219
0 335 5 1 1 4221
0 336 7 1 2 3981 335
0 337 5 2 1 336
0 338 7 1 2 3675 4222
0 339 5 1 1 338
0 340 7 2 2 4223 339
0 341 5 1 1 4225
0 342 7 2 2 3975 4226
0 343 5 2 1 4227
0 344 7 1 2 323 4224
0 345 5 1 1 344
0 346 7 1 2 4205 4214
0 347 5 1 1 346
0 348 7 2 2 345 347
0 349 5 1 1 4231
0 350 7 1 2 4229 349
0 351 5 2 1 350
0 352 7 1 2 4206 4216
0 353 5 1 1 352
0 354 7 1 2 4218 353
0 355 5 1 1 354
0 356 7 3 2 4220 355
0 357 5 1 1 4235
0 358 7 1 2 4230 4236
0 359 5 1 1 358
0 360 7 1 2 4232 359
0 361 5 1 1 360
0 362 7 3 2 4233 361
0 363 5 1 1 4238
0 364 7 2 2 4234 357
0 365 5 1 1 4241
0 366 7 1 2 3976 365
0 367 5 2 1 366
0 368 7 1 2 3668 4242
0 369 5 1 1 368
0 370 7 2 2 4243 369
0 371 5 1 1 4245
0 372 7 2 2 3969 4246
0 373 5 2 1 4247
0 374 7 1 2 341 4244
0 375 5 1 1 374
0 376 7 1 2 4228 4237
0 377 5 1 1 376
0 378 7 2 2 375 377
0 379 5 1 1 4251
0 380 7 1 2 4249 379
0 381 5 2 1 380
0 382 7 2 2 363 4253
0 383 5 1 1 4255
0 384 7 1 2 3970 383
0 385 5 2 1 384
0 386 7 1 2 3662 4256
0 387 5 1 1 386
0 388 7 2 2 4257 387
0 389 5 1 1 4259
0 390 7 2 2 3963 4260
0 391 5 2 1 4261
0 392 7 1 2 371 4258
0 393 5 1 1 392
0 394 7 1 2 4239 4248
0 395 5 1 1 394
0 396 7 2 2 393 395
0 397 5 1 1 4265
0 398 7 1 2 4263 397
0 399 5 2 1 398
0 400 7 1 2 4240 4250
0 401 5 1 1 400
0 402 7 1 2 4252 401
0 403 5 1 1 402
0 404 7 3 2 4254 403
0 405 5 1 1 4269
0 406 7 1 2 4264 4270
0 407 5 1 1 406
0 408 7 1 2 4266 407
0 409 5 1 1 408
0 410 7 3 2 4267 409
0 411 5 1 1 4272
0 412 7 2 2 4268 405
0 413 5 1 1 4275
0 414 7 1 2 3964 413
0 415 5 2 1 414
0 416 7 1 2 3656 4276
0 417 5 1 1 416
0 418 7 2 2 4277 417
0 419 5 1 1 4279
0 420 7 2 2 3958 4280
0 421 5 2 1 4281
0 422 7 1 2 389 4278
0 423 5 1 1 422
0 424 7 1 2 4262 4271
0 425 5 1 1 424
0 426 7 2 2 423 425
0 427 5 1 1 4285
0 428 7 1 2 4283 427
0 429 5 2 1 428
0 430 7 2 2 411 4287
0 431 5 1 1 4289
0 432 7 1 2 3959 431
0 433 5 2 1 432
0 434 7 1 2 3649 4290
0 435 5 1 1 434
0 436 7 2 2 4291 435
0 437 5 1 1 4293
0 438 7 2 2 3951 4294
0 439 5 2 1 4295
0 440 7 1 2 419 4292
0 441 5 1 1 440
0 442 7 1 2 4273 4282
0 443 5 1 1 442
0 444 7 2 2 441 443
0 445 5 1 1 4299
0 446 7 1 2 4297 445
0 447 5 2 1 446
0 448 7 1 2 4274 4284
0 449 5 1 1 448
0 450 7 1 2 4286 449
0 451 5 1 1 450
0 452 7 3 2 4288 451
0 453 5 1 1 4303
0 454 7 1 2 4298 4304
0 455 5 1 1 454
0 456 7 1 2 4300 455
0 457 5 1 1 456
0 458 7 3 2 4301 457
0 459 5 1 1 4306
0 460 7 2 2 4302 453
0 461 5 1 1 4309
0 462 7 1 2 3952 461
0 463 5 2 1 462
0 464 7 1 2 3643 4310
0 465 5 1 1 464
0 466 7 2 2 4311 465
0 467 5 1 1 4313
0 468 7 2 2 3944 4314
0 469 5 2 1 4315
0 470 7 1 2 437 4312
0 471 5 1 1 470
0 472 7 1 2 4296 4305
0 473 5 1 1 472
0 474 7 2 2 471 473
0 475 5 1 1 4319
0 476 7 1 2 4317 475
0 477 5 2 1 476
0 478 7 2 2 459 4321
0 479 5 1 1 4323
0 480 7 1 2 3945 479
0 481 5 2 1 480
0 482 7 1 2 3636 4324
0 483 5 1 1 482
0 484 7 2 2 4325 483
0 485 5 1 1 4327
0 486 7 2 2 3938 4328
0 487 5 2 1 4329
0 488 7 1 2 467 4326
0 489 5 1 1 488
0 490 7 1 2 4307 4316
0 491 5 1 1 490
0 492 7 2 2 489 491
0 493 5 1 1 4333
0 494 7 1 2 4331 493
0 495 5 2 1 494
0 496 7 1 2 4308 4318
0 497 5 1 1 496
0 498 7 1 2 4320 497
0 499 5 1 1 498
0 500 7 3 2 4322 499
0 501 5 1 1 4337
0 502 7 1 2 4332 4338
0 503 5 1 1 502
0 504 7 1 2 4334 503
0 505 5 1 1 504
0 506 7 3 2 4335 505
0 507 5 1 1 4340
0 508 7 2 2 4336 501
0 509 5 1 1 4343
0 510 7 1 2 3939 509
0 511 5 2 1 510
0 512 7 1 2 3629 4344
0 513 5 1 1 512
0 514 7 2 2 4345 513
0 515 5 1 1 4347
0 516 7 2 2 3931 4348
0 517 5 2 1 4349
0 518 7 1 2 485 4346
0 519 5 1 1 518
0 520 7 1 2 4330 4339
0 521 5 1 1 520
0 522 7 2 2 519 521
0 523 5 1 1 4353
0 524 7 1 2 4351 523
0 525 5 2 1 524
0 526 7 2 2 507 4355
0 527 5 1 1 4357
0 528 7 1 2 3932 527
0 529 5 2 1 528
0 530 7 1 2 3623 4358
0 531 5 1 1 530
0 532 7 2 2 4359 531
0 533 5 1 1 4361
0 534 7 2 2 3924 4362
0 535 5 2 1 4363
0 536 7 1 2 515 4360
0 537 5 1 1 536
0 538 7 1 2 4341 4350
0 539 5 1 1 538
0 540 7 2 2 537 539
0 541 5 1 1 4367
0 542 7 1 2 4365 541
0 543 5 2 1 542
0 544 7 1 2 4342 4352
0 545 5 1 1 544
0 546 7 1 2 4354 545
0 547 5 1 1 546
0 548 7 3 2 4356 547
0 549 5 1 1 4371
0 550 7 1 2 4366 4372
0 551 5 1 1 550
0 552 7 1 2 4368 551
0 553 5 1 1 552
0 554 7 3 2 4369 553
0 555 5 1 1 4374
0 556 7 2 2 4370 549
0 557 5 1 1 4377
0 558 7 1 2 3925 557
0 559 5 2 1 558
0 560 7 1 2 3617 4378
0 561 5 1 1 560
0 562 7 2 2 4379 561
0 563 5 1 1 4381
0 564 7 2 2 3918 4382
0 565 5 2 1 4383
0 566 7 1 2 533 4380
0 567 5 1 1 566
0 568 7 1 2 4364 4373
0 569 5 1 1 568
0 570 7 2 2 567 569
0 571 5 1 1 4387
0 572 7 1 2 4385 571
0 573 5 2 1 572
0 574 7 2 2 555 4389
0 575 5 1 1 4391
0 576 7 1 2 3919 575
0 577 5 2 1 576
0 578 7 1 2 3610 4392
0 579 5 1 1 578
0 580 7 2 2 4393 579
0 581 5 1 1 4395
0 582 7 2 2 3911 4396
0 583 5 2 1 4397
0 584 7 1 2 563 4394
0 585 5 1 1 584
0 586 7 1 2 4375 4384
0 587 5 1 1 586
0 588 7 2 2 585 587
0 589 5 1 1 4401
0 590 7 1 2 4399 589
0 591 5 2 1 590
0 592 7 1 2 4376 4386
0 593 5 1 1 592
0 594 7 1 2 4388 593
0 595 5 1 1 594
0 596 7 3 2 4390 595
0 597 5 1 1 4405
0 598 7 1 2 4400 4406
0 599 5 1 1 598
0 600 7 1 2 4402 599
0 601 5 1 1 600
0 602 7 3 2 4403 601
0 603 5 1 1 4408
0 604 7 2 2 4404 597
0 605 5 1 1 4411
0 606 7 1 2 3912 605
0 607 5 2 1 606
0 608 7 1 2 3604 4412
0 609 5 1 1 608
0 610 7 2 2 4413 609
0 611 5 1 1 4415
0 612 7 2 2 3904 4416
0 613 5 2 1 4417
0 614 7 1 2 581 4414
0 615 5 1 1 614
0 616 7 1 2 4398 4407
0 617 5 1 1 616
0 618 7 2 2 615 617
0 619 5 1 1 4421
0 620 7 1 2 4419 619
0 621 5 2 1 620
0 622 7 2 2 603 4423
0 623 5 1 1 4425
0 624 7 1 2 3905 623
0 625 5 2 1 624
0 626 7 1 2 3597 4426
0 627 5 1 1 626
0 628 7 2 2 4427 627
0 629 5 1 1 4429
0 630 7 2 2 3898 4430
0 631 5 2 1 4431
0 632 7 1 2 611 4428
0 633 5 1 1 632
0 634 7 1 2 4409 4418
0 635 5 1 1 634
0 636 7 2 2 633 635
0 637 5 1 1 4435
0 638 7 1 2 4433 637
0 639 5 2 1 638
0 640 7 1 2 4410 4420
0 641 5 1 1 640
0 642 7 1 2 4422 641
0 643 5 1 1 642
0 644 7 3 2 4424 643
0 645 5 1 1 4439
0 646 7 1 2 4434 4440
0 647 5 1 1 646
0 648 7 1 2 4436 647
0 649 5 1 1 648
0 650 7 3 2 4437 649
0 651 5 1 1 4442
0 652 7 2 2 4438 645
0 653 5 1 1 4445
0 654 7 1 2 3899 653
0 655 5 2 1 654
0 656 7 1 2 3590 4446
0 657 5 1 1 656
0 658 7 2 2 4447 657
0 659 5 1 1 4449
0 660 7 2 2 3891 4450
0 661 5 2 1 4451
0 662 7 1 2 629 4448
0 663 5 1 1 662
0 664 7 1 2 4432 4441
0 665 5 1 1 664
0 666 7 2 2 663 665
0 667 5 1 1 4455
0 668 7 1 2 4453 667
0 669 5 2 1 668
0 670 7 2 2 651 4457
0 671 5 1 1 4459
0 672 7 1 2 3892 671
0 673 5 2 1 672
0 674 7 1 2 3584 4460
0 675 5 1 1 674
0 676 7 2 2 4461 675
0 677 5 1 1 4463
0 678 7 2 2 3884 4464
0 679 5 2 1 4465
0 680 7 1 2 659 4462
0 681 5 1 1 680
0 682 7 1 2 4443 4452
0 683 5 1 1 682
0 684 7 2 2 681 683
0 685 5 1 1 4469
0 686 7 1 2 4467 685
0 687 5 2 1 686
0 688 7 1 2 4444 4454
0 689 5 1 1 688
0 690 7 1 2 4456 689
0 691 5 1 1 690
0 692 7 3 2 4458 691
0 693 5 1 1 4473
0 694 7 1 2 4468 4474
0 695 5 1 1 694
0 696 7 1 2 4470 695
0 697 5 1 1 696
0 698 7 3 2 4471 697
0 699 5 1 1 4476
0 700 7 2 2 4472 693
0 701 5 1 1 4479
0 702 7 1 2 3885 701
0 703 5 2 1 702
0 704 7 1 2 3578 4480
0 705 5 1 1 704
0 706 7 2 2 4481 705
0 707 5 1 1 4483
0 708 7 2 2 3878 4484
0 709 5 2 1 4485
0 710 7 1 2 677 4482
0 711 5 1 1 710
0 712 7 1 2 4466 4475
0 713 5 1 1 712
0 714 7 2 2 711 713
0 715 5 1 1 4489
0 716 7 1 2 4487 715
0 717 5 2 1 716
0 718 7 2 2 699 4491
0 719 5 1 1 4493
0 720 7 1 2 3879 719
0 721 5 2 1 720
0 722 7 1 2 3571 4494
0 723 5 1 1 722
0 724 7 2 2 4495 723
0 725 5 1 1 4497
0 726 7 2 2 3871 4498
0 727 5 2 1 4499
0 728 7 1 2 707 4496
0 729 5 1 1 728
0 730 7 1 2 4477 4486
0 731 5 1 1 730
0 732 7 2 2 729 731
0 733 5 1 1 4503
0 734 7 1 2 4501 733
0 735 5 2 1 734
0 736 7 1 2 4478 4488
0 737 5 1 1 736
0 738 7 1 2 4490 737
0 739 5 1 1 738
0 740 7 3 2 4492 739
0 741 5 1 1 4507
0 742 7 1 2 4502 4508
0 743 5 1 1 742
0 744 7 1 2 4504 743
0 745 5 1 1 744
0 746 7 3 2 4505 745
0 747 5 1 1 4510
0 748 7 2 2 4506 741
0 749 5 1 1 4513
0 750 7 1 2 3872 749
0 751 5 2 1 750
0 752 7 1 2 3565 4514
0 753 5 1 1 752
0 754 7 2 2 4515 753
0 755 5 1 1 4517
0 756 7 2 2 3865 4518
0 757 5 2 1 4519
0 758 7 1 2 725 4516
0 759 5 1 1 758
0 760 7 1 2 4500 4509
0 761 5 1 1 760
0 762 7 2 2 759 761
0 763 5 1 1 4523
0 764 7 1 2 4521 763
0 765 5 2 1 764
0 766 7 2 2 747 4525
0 767 5 1 1 4527
0 768 7 1 2 3866 767
0 769 5 2 1 768
0 770 7 1 2 3558 4528
0 771 5 1 1 770
0 772 7 2 2 4529 771
0 773 5 1 1 4531
0 774 7 2 2 3860 4532
0 775 5 2 1 4533
0 776 7 1 2 755 4530
0 777 5 1 1 776
0 778 7 1 2 4511 4520
0 779 5 1 1 778
0 780 7 2 2 777 779
0 781 5 1 1 4537
0 782 7 1 2 4535 781
0 783 5 2 1 782
0 784 7 1 2 4512 4522
0 785 5 1 1 784
0 786 7 1 2 4524 785
0 787 5 1 1 786
0 788 7 3 2 4526 787
0 789 5 1 1 4541
0 790 7 1 2 4536 4542
0 791 5 1 1 790
0 792 7 1 2 4538 791
0 793 5 1 1 792
0 794 7 3 2 4539 793
0 795 5 1 1 4544
0 796 7 2 2 4540 789
0 797 5 1 1 4547
0 798 7 1 2 3861 797
0 799 5 2 1 798
0 800 7 1 2 3551 4548
0 801 5 1 1 800
0 802 7 2 2 4549 801
0 803 5 1 1 4551
0 804 7 2 2 3854 4552
0 805 5 2 1 4553
0 806 7 1 2 773 4550
0 807 5 1 1 806
0 808 7 1 2 4534 4543
0 809 5 1 1 808
0 810 7 2 2 807 809
0 811 5 1 1 4557
0 812 7 1 2 4555 811
0 813 5 2 1 812
0 814 7 2 2 795 4559
0 815 5 1 1 4561
0 816 7 1 2 3855 815
0 817 5 2 1 816
0 818 7 1 2 3545 4562
0 819 5 1 1 818
0 820 7 2 2 4563 819
0 821 5 1 1 4565
0 822 7 2 2 3848 4566
0 823 5 2 1 4567
0 824 7 1 2 803 4564
0 825 5 1 1 824
0 826 7 1 2 4545 4554
0 827 5 1 1 826
0 828 7 2 2 825 827
0 829 5 1 1 4571
0 830 7 1 2 4569 829
0 831 5 2 1 830
0 832 7 1 2 4546 4556
0 833 5 1 1 832
0 834 7 1 2 4558 833
0 835 5 1 1 834
0 836 7 3 2 4560 835
0 837 5 1 1 4575
0 838 7 1 2 4570 4576
0 839 5 1 1 838
0 840 7 1 2 4572 839
0 841 5 1 1 840
0 842 7 3 2 4573 841
0 843 5 1 1 4578
0 844 7 2 2 4574 837
0 845 5 1 1 4581
0 846 7 1 2 3849 845
0 847 5 2 1 846
0 848 7 1 2 3539 4582
0 849 5 1 1 848
0 850 7 2 2 4583 849
0 851 5 1 1 4585
0 852 7 2 2 3843 4586
0 853 5 2 1 4587
0 854 7 1 2 821 4584
0 855 5 1 1 854
0 856 7 1 2 4568 4577
0 857 5 1 1 856
0 858 7 2 2 855 857
0 859 5 1 1 4591
0 860 7 1 2 4589 859
0 861 5 2 1 860
0 862 7 2 2 843 4593
0 863 5 1 1 4595
0 864 7 1 2 3844 863
0 865 5 2 1 864
0 866 7 1 2 3532 4596
0 867 5 1 1 866
0 868 7 2 2 4597 867
0 869 5 1 1 4599
0 870 7 2 2 3837 4600
0 871 5 2 1 4601
0 872 7 1 2 851 4598
0 873 5 1 1 872
0 874 7 1 2 4579 4588
0 875 5 1 1 874
0 876 7 2 2 873 875
0 877 5 1 1 4605
0 878 7 1 2 4603 877
0 879 5 2 1 878
0 880 7 1 2 4580 4590
0 881 5 1 1 880
0 882 7 1 2 4592 881
0 883 5 1 1 882
0 884 7 3 2 4594 883
0 885 5 1 1 4609
0 886 7 1 2 4604 4610
0 887 5 1 1 886
0 888 7 1 2 4606 887
0 889 5 1 1 888
0 890 7 3 2 4607 889
0 891 5 1 1 4612
0 892 7 2 2 4608 885
0 893 5 1 1 4615
0 894 7 1 2 3838 893
0 895 5 2 1 894
0 896 7 1 2 3526 4616
0 897 5 1 1 896
0 898 7 2 2 4617 897
0 899 5 1 1 4619
0 900 7 2 2 3831 4620
0 901 5 2 1 4621
0 902 7 1 2 869 4618
0 903 5 1 1 902
0 904 7 1 2 4602 4611
0 905 5 1 1 904
0 906 7 2 2 903 905
0 907 5 1 1 4625
0 908 7 1 2 4623 907
0 909 5 2 1 908
0 910 7 2 2 891 4627
0 911 5 1 1 4629
0 912 7 1 2 3832 911
0 913 5 2 1 912
0 914 7 1 2 3519 4630
0 915 5 1 1 914
0 916 7 2 2 4631 915
0 917 5 1 1 4633
0 918 7 2 2 3826 4634
0 919 5 2 1 4635
0 920 7 1 2 899 4632
0 921 5 1 1 920
0 922 7 1 2 4613 4622
0 923 5 1 1 922
0 924 7 2 2 921 923
0 925 5 1 1 4639
0 926 7 1 2 4637 925
0 927 5 2 1 926
0 928 7 1 2 4614 4624
0 929 5 1 1 928
0 930 7 1 2 4626 929
0 931 5 1 1 930
0 932 7 3 2 4628 931
0 933 5 1 1 4643
0 934 7 1 2 4638 4644
0 935 5 1 1 934
0 936 7 1 2 4640 935
0 937 5 1 1 936
0 938 7 3 2 4641 937
0 939 5 1 1 4646
0 940 7 2 2 4642 933
0 941 5 1 1 4649
0 942 7 1 2 3827 941
0 943 5 2 1 942
0 944 7 1 2 3512 4650
0 945 5 1 1 944
0 946 7 2 2 4651 945
0 947 5 1 1 4653
0 948 7 2 2 3820 4654
0 949 5 2 1 4655
0 950 7 1 2 917 4652
0 951 5 1 1 950
0 952 7 1 2 4636 4645
0 953 5 1 1 952
0 954 7 2 2 951 953
0 955 5 1 1 4659
0 956 7 1 2 4657 955
0 957 5 2 1 956
0 958 7 2 2 939 4661
0 959 5 1 1 4663
0 960 7 1 2 3821 959
0 961 5 2 1 960
0 962 7 1 2 3506 4664
0 963 5 1 1 962
0 964 7 2 2 4665 963
0 965 5 1 1 4667
0 966 7 2 2 3814 4668
0 967 5 2 1 4669
0 968 7 1 2 947 4666
0 969 5 1 1 968
0 970 7 1 2 4647 4656
0 971 5 1 1 970
0 972 7 2 2 969 971
0 973 5 1 1 4673
0 974 7 1 2 4671 973
0 975 5 2 1 974
0 976 7 1 2 4648 4658
0 977 5 1 1 976
0 978 7 1 2 4660 977
0 979 5 1 1 978
0 980 7 3 2 4662 979
0 981 5 1 1 4677
0 982 7 1 2 4672 4678
0 983 5 1 1 982
0 984 7 1 2 4674 983
0 985 5 1 1 984
0 986 7 3 2 4675 985
0 987 5 1 1 4680
0 988 7 2 2 4676 981
0 989 5 1 1 4683
0 990 7 1 2 3815 989
0 991 5 2 1 990
0 992 7 1 2 3500 4684
0 993 5 1 1 992
0 994 7 2 2 4685 993
0 995 5 1 1 4687
0 996 7 2 2 3809 4688
0 997 5 2 1 4689
0 998 7 1 2 965 4686
0 999 5 1 1 998
0 1000 7 1 2 4670 4679
0 1001 5 1 1 1000
0 1002 7 2 2 999 1001
0 1003 5 1 1 4693
0 1004 7 1 2 4691 1003
0 1005 5 2 1 1004
0 1006 7 2 2 987 4695
0 1007 5 1 1 4697
0 1008 7 1 2 3810 1007
0 1009 5 2 1 1008
0 1010 7 1 2 3493 4698
0 1011 5 1 1 1010
0 1012 7 2 2 4699 1011
0 1013 5 1 1 4701
0 1014 7 2 2 3803 4702
0 1015 5 2 1 4703
0 1016 7 1 2 995 4700
0 1017 5 1 1 1016
0 1018 7 1 2 4681 4690
0 1019 5 1 1 1018
0 1020 7 2 2 1017 1019
0 1021 5 1 1 4707
0 1022 7 1 2 4705 1021
0 1023 5 2 1 1022
0 1024 7 1 2 4682 4692
0 1025 5 1 1 1024
0 1026 7 1 2 4694 1025
0 1027 5 1 1 1026
0 1028 7 3 2 4696 1027
0 1029 5 1 1 4711
0 1030 7 1 2 4706 4712
0 1031 5 1 1 1030
0 1032 7 1 2 4708 1031
0 1033 5 1 1 1032
0 1034 7 3 2 4709 1033
0 1035 5 1 1 4714
0 1036 7 2 2 4710 1029
0 1037 5 1 1 4717
0 1038 7 1 2 3804 1037
0 1039 5 2 1 1038
0 1040 7 1 2 3487 4718
0 1041 5 1 1 1040
0 1042 7 2 2 4719 1041
0 1043 5 1 1 4721
0 1044 7 2 2 3797 4722
0 1045 5 2 1 4723
0 1046 7 1 2 1013 4720
0 1047 5 1 1 1046
0 1048 7 1 2 4704 4713
0 1049 5 1 1 1048
0 1050 7 2 2 1047 1049
0 1051 5 1 1 4727
0 1052 7 1 2 4725 1051
0 1053 5 2 1 1052
0 1054 7 2 2 1035 4729
0 1055 5 1 1 4731
0 1056 7 1 2 3798 1055
0 1057 5 2 1 1056
0 1058 7 1 2 3480 4732
0 1059 5 1 1 1058
0 1060 7 2 2 4733 1059
0 1061 5 1 1 4735
0 1062 7 2 2 3792 4736
0 1063 5 2 1 4737
0 1064 7 1 2 1043 4734
0 1065 5 1 1 1064
0 1066 7 1 2 4715 4724
0 1067 5 1 1 1066
0 1068 7 2 2 1065 1067
0 1069 5 1 1 4741
0 1070 7 1 2 4739 1069
0 1071 5 2 1 1070
0 1072 7 1 2 4716 4726
0 1073 5 1 1 1072
0 1074 7 1 2 4728 1073
0 1075 5 1 1 1074
0 1076 7 3 2 4730 1075
0 1077 5 1 1 4745
0 1078 7 1 2 4740 4746
0 1079 5 1 1 1078
0 1080 7 1 2 4742 1079
0 1081 5 1 1 1080
0 1082 7 3 2 4743 1081
0 1083 5 1 1 4748
0 1084 7 2 2 4744 1077
0 1085 5 1 1 4751
0 1086 7 1 2 3793 1085
0 1087 5 2 1 1086
0 1088 7 1 2 3473 4752
0 1089 5 1 1 1088
0 1090 7 2 2 4753 1089
0 1091 5 1 1 4755
0 1092 7 2 2 3786 4756
0 1093 5 2 1 4757
0 1094 7 1 2 1061 4754
0 1095 5 1 1 1094
0 1096 7 1 2 4738 4747
0 1097 5 1 1 1096
0 1098 7 2 2 1095 1097
0 1099 5 1 1 4761
0 1100 7 1 2 4759 1099
0 1101 5 2 1 1100
0 1102 7 2 2 1083 4763
0 1103 5 1 1 4765
0 1104 7 1 2 3787 1103
0 1105 5 2 1 1104
0 1106 7 1 2 3467 4766
0 1107 5 1 1 1106
0 1108 7 2 2 4767 1107
0 1109 5 1 1 4769
0 1110 7 2 2 3780 4770
0 1111 5 2 1 4771
0 1112 7 1 2 1091 4768
0 1113 5 1 1 1112
0 1114 7 1 2 4749 4758
0 1115 5 1 1 1114
0 1116 7 2 2 1113 1115
0 1117 5 1 1 4775
0 1118 7 1 2 4773 1117
0 1119 5 2 1 1118
0 1120 7 1 2 4750 4760
0 1121 5 1 1 1120
0 1122 7 1 2 4762 1121
0 1123 5 1 1 1122
0 1124 7 3 2 4764 1123
0 1125 5 1 1 4779
0 1126 7 2 2 4777 1125
0 1127 5 1 1 4782
0 1128 7 1 2 3781 1127
0 1129 5 2 1 1128
0 1130 7 1 2 3461 4783
0 1131 5 1 1 1130
0 1132 7 3 2 4784 1131
0 1133 5 2 1 4786
0 1134 7 1 2 3774 4787
0 1135 5 2 1 1134
0 1136 7 1 2 1109 4785
0 1137 5 1 1 1136
0 1138 7 1 2 4772 4780
0 1139 5 1 1 1138
0 1140 7 2 2 1137 1139
0 1141 5 1 1 4793
0 1142 7 1 2 4791 1141
0 1143 5 2 1 1142
0 1144 7 1 2 4774 4781
0 1145 5 1 1 1144
0 1146 7 1 2 4776 1145
0 1147 5 1 1 1146
0 1148 7 2 2 4778 1147
0 1149 5 1 1 4797
0 1150 7 1 2 4792 4798
0 1151 5 1 1 1150
0 1152 7 1 2 4794 1151
0 1153 5 1 1 1152
0 1154 7 2 2 4795 1153
0 1155 5 1 1 4799
0 1156 7 2 2 4796 1149
0 1157 5 1 1 4801
0 1158 7 1 2 3455 4802
0 1159 5 2 1 1158
0 1160 7 2 2 4788 4803
0 1161 5 1 1 4805
0 1162 7 1 2 3775 1157
0 1163 5 3 1 1162
0 1164 7 1 2 4789 4807
0 1165 5 1 1 1164
0 1166 7 1 2 3763 3450
0 1167 7 1 2 1165 1166
0 1168 7 1 2 1161 1167
0 1169 5 1 1 1168
0 1170 7 2 2 3446 3768
0 1171 5 1 1 4810
0 1172 7 1 2 4808 4811
0 1173 7 1 2 4806 1172
0 1174 5 1 1 1173
0 1175 7 1 2 1169 1174
0 1176 5 1 1 1175
0 1177 7 1 2 1155 1176
0 1178 5 1 1 1177
0 1179 7 1 2 3447 4790
0 1180 5 1 1 1179
0 1181 7 1 2 3769 4800
0 1182 5 1 1 1181
0 1183 7 1 2 1180 1182
0 1184 5 1 1 1183
0 1185 7 1 2 4809 1171
0 1186 7 1 2 4804 1185
0 1187 7 1 2 1184 1186
0 1188 5 1 1 1187
0 1189 7 2 2 3745 110
0 1190 5 1 1 4812
0 1191 7 1 2 4039 4077
0 1192 5 1 1 1191
0 1193 7 2 2 1190 1192
0 1194 5 1 1 4814
0 1195 7 1 2 3737 4815
0 1196 5 2 1 1195
0 1197 7 1 2 4078 4813
0 1198 5 1 1 1197
0 1199 7 2 2 4060 1198
0 1200 5 1 1 4818
0 1201 7 1 2 4816 4819
0 1202 5 1 1 1201
0 1203 7 1 2 3738 1200
0 1204 5 2 1 1203
0 1205 7 2 2 1202 4820
0 1206 5 1 1 4822
0 1207 7 1 2 4027 4823
0 1208 5 1 1 1207
0 1209 7 1 2 4034 1194
0 1210 5 1 1 1209
0 1211 7 1 2 4817 1210
0 1212 7 2 2 4821 1211
0 1213 5 1 1 4824
0 1214 7 1 2 3729 4825
0 1215 5 2 1 1214
0 1216 7 1 2 3730 1206
0 1217 7 1 2 4826 1216
0 1218 5 2 1 1217
0 1219 7 3 2 1208 4828
0 1220 5 1 1 4830
0 1221 7 1 2 3722 1220
0 1222 5 1 1 1221
0 1223 7 1 2 4028 1213
0 1224 5 1 1 1223
0 1225 7 1 2 4827 1224
0 1226 7 1 2 4829 1225
0 1227 5 2 1 1226
0 1228 7 1 2 4831 4833
0 1229 5 1 1 1228
0 1230 7 1 2 3723 1229
0 1231 5 2 1 1230
0 1232 7 1 2 4832 4835
0 1233 5 1 1 1232
0 1234 7 2 2 1222 1233
0 1235 5 1 1 4837
0 1236 7 1 2 4016 4838
0 1237 5 1 1 1236
0 1238 7 1 2 4022 4834
0 1239 5 1 1 1238
0 1240 7 2 2 4836 1239
0 1241 5 1 1 4839
0 1242 7 1 2 3715 4840
0 1243 5 2 1 1242
0 1244 7 1 2 3716 1235
0 1245 7 1 2 4841 1244
0 1246 5 2 1 1245
0 1247 7 3 2 1237 4843
0 1248 5 1 1 4845
0 1249 7 1 2 4017 1241
0 1250 5 1 1 1249
0 1251 7 1 2 4842 1250
0 1252 7 1 2 4844 1251
0 1253 5 2 1 1252
0 1254 7 1 2 4846 4848
0 1255 5 1 1 1254
0 1256 7 1 2 3708 1255
0 1257 5 2 1 1256
0 1258 7 1 2 4011 4849
0 1259 5 1 1 1258
0 1260 7 2 2 4850 1259
0 1261 5 2 1 4852
0 1262 7 1 2 3709 1248
0 1263 5 1 1 1262
0 1264 7 1 2 4847 4851
0 1265 5 1 1 1264
0 1266 7 1 2 1263 1265
0 1267 5 2 1 1266
0 1268 7 1 2 4854 4856
0 1269 5 1 1 1268
0 1270 7 2 2 3702 1269
0 1271 5 1 1 4858
0 1272 7 1 2 4855 4859
0 1273 5 1 1 1272
0 1274 7 1 2 4005 4853
0 1275 5 1 1 1274
0 1276 7 2 2 1273 1275
0 1277 5 1 1 4860
0 1278 7 1 2 4006 4857
0 1279 5 1 1 1278
0 1280 7 2 2 1271 1279
0 1281 5 1 1 4862
0 1282 7 2 2 3696 1281
0 1283 5 1 1 4864
0 1284 7 1 2 4861 4865
0 1285 5 2 1 1284
0 1286 7 1 2 3999 4863
0 1287 5 1 1 1286
0 1288 7 2 2 1283 1287
0 1289 5 1 1 4868
0 1290 7 1 2 4866 1289
0 1291 5 1 1 1290
0 1292 7 1 2 3994 1291
0 1293 5 1 1 1292
0 1294 7 1 2 4000 1277
0 1295 5 2 1 1294
0 1296 7 1 2 4869 4870
0 1297 5 1 1 1296
0 1298 7 1 2 3689 1297
0 1299 5 2 1 1298
0 1300 7 2 2 1293 4872
0 1301 5 2 1 4874
0 1302 7 2 2 4867 4871
0 1303 5 1 1 4878
0 1304 7 1 2 3690 1303
0 1305 5 1 1 1304
0 1306 7 1 2 4873 4879
0 1307 5 1 1 1306
0 1308 7 1 2 1305 1307
0 1309 5 2 1 1308
0 1310 7 1 2 4876 4880
0 1311 5 1 1 1310
0 1312 7 2 2 3683 1311
0 1313 5 1 1 4882
0 1314 7 1 2 4877 4883
0 1315 5 1 1 1314
0 1316 7 1 2 3988 4875
0 1317 5 1 1 1316
0 1318 7 2 2 1315 1317
0 1319 5 1 1 4884
0 1320 7 1 2 3982 1319
0 1321 5 1 1 1320
0 1322 7 1 2 3989 4881
0 1323 5 1 1 1322
0 1324 7 2 2 1313 1323
0 1325 5 1 1 4886
0 1326 7 1 2 3676 4887
0 1327 5 2 1 1326
0 1328 7 1 2 3677 4885
0 1329 7 1 2 4888 1328
0 1330 5 2 1 1329
0 1331 7 3 2 1321 4890
0 1332 5 1 1 4892
0 1333 7 1 2 3983 1325
0 1334 5 1 1 1333
0 1335 7 1 2 4889 1334
0 1336 7 1 2 4891 1335
0 1337 5 2 1 1336
0 1338 7 1 2 4893 4895
0 1339 5 1 1 1338
0 1340 7 1 2 3669 1339
0 1341 5 2 1 1340
0 1342 7 1 2 3977 4896
0 1343 5 1 1 1342
0 1344 7 2 2 4897 1343
0 1345 5 2 1 4899
0 1346 7 1 2 3670 1332
0 1347 5 1 1 1346
0 1348 7 1 2 4894 4898
0 1349 5 1 1 1348
0 1350 7 1 2 1347 1349
0 1351 5 2 1 1350
0 1352 7 1 2 4901 4903
0 1353 5 1 1 1352
0 1354 7 2 2 3663 1353
0 1355 5 1 1 4905
0 1356 7 1 2 4902 4906
0 1357 5 1 1 1356
0 1358 7 1 2 3971 4900
0 1359 5 1 1 1358
0 1360 7 2 2 1357 1359
0 1361 5 1 1 4907
0 1362 7 1 2 3972 4904
0 1363 5 1 1 1362
0 1364 7 2 2 1355 1363
0 1365 5 1 1 4909
0 1366 7 2 2 3657 1365
0 1367 5 1 1 4911
0 1368 7 1 2 4908 4912
0 1369 5 2 1 1368
0 1370 7 1 2 3965 4910
0 1371 5 1 1 1370
0 1372 7 2 2 1367 1371
0 1373 5 1 1 4915
0 1374 7 1 2 4913 1373
0 1375 5 1 1 1374
0 1376 7 1 2 3960 1375
0 1377 5 1 1 1376
0 1378 7 1 2 3966 1361
0 1379 5 2 1 1378
0 1380 7 1 2 4916 4917
0 1381 5 1 1 1380
0 1382 7 1 2 3650 1381
0 1383 5 2 1 1382
0 1384 7 2 2 1377 4919
0 1385 5 2 1 4921
0 1386 7 2 2 4914 4918
0 1387 5 1 1 4925
0 1388 7 1 2 3651 1387
0 1389 5 1 1 1388
0 1390 7 1 2 4920 4926
0 1391 5 1 1 1390
0 1392 7 1 2 1389 1391
0 1393 5 2 1 1392
0 1394 7 1 2 4923 4927
0 1395 5 1 1 1394
0 1396 7 2 2 3644 1395
0 1397 5 1 1 4929
0 1398 7 1 2 4924 4930
0 1399 5 1 1 1398
0 1400 7 1 2 3953 4922
0 1401 5 1 1 1400
0 1402 7 2 2 1399 1401
0 1403 5 1 1 4931
0 1404 7 1 2 3946 1403
0 1405 5 1 1 1404
0 1406 7 1 2 3954 4928
0 1407 5 1 1 1406
0 1408 7 2 2 1397 1407
0 1409 5 1 1 4933
0 1410 7 1 2 3637 4934
0 1411 5 2 1 1410
0 1412 7 1 2 3638 4932
0 1413 7 1 2 4935 1412
0 1414 5 2 1 1413
0 1415 7 3 2 1405 4937
0 1416 5 1 1 4939
0 1417 7 1 2 3947 1409
0 1418 5 1 1 1417
0 1419 7 1 2 4936 1418
0 1420 7 1 2 4938 1419
0 1421 5 2 1 1420
0 1422 7 1 2 4940 4942
0 1423 5 1 1 1422
0 1424 7 1 2 3630 1423
0 1425 5 2 1 1424
0 1426 7 1 2 3940 4943
0 1427 5 1 1 1426
0 1428 7 2 2 4944 1427
0 1429 5 2 1 4946
0 1430 7 1 2 3631 1416
0 1431 5 1 1 1430
0 1432 7 1 2 4941 4945
0 1433 5 1 1 1432
0 1434 7 1 2 1431 1433
0 1435 5 2 1 1434
0 1436 7 1 2 4948 4950
0 1437 5 1 1 1436
0 1438 7 2 2 3624 1437
0 1439 5 1 1 4952
0 1440 7 1 2 4949 4953
0 1441 5 1 1 1440
0 1442 7 1 2 3933 4947
0 1443 5 1 1 1442
0 1444 7 2 2 1441 1443
0 1445 5 1 1 4954
0 1446 7 1 2 3934 4951
0 1447 5 1 1 1446
0 1448 7 2 2 1439 1447
0 1449 5 1 1 4956
0 1450 7 2 2 3618 1449
0 1451 5 1 1 4958
0 1452 7 1 2 4955 4959
0 1453 5 2 1 1452
0 1454 7 1 2 3926 4957
0 1455 5 1 1 1454
0 1456 7 2 2 1451 1455
0 1457 5 1 1 4962
0 1458 7 1 2 4960 1457
0 1459 5 1 1 1458
0 1460 7 1 2 3920 1459
0 1461 5 1 1 1460
0 1462 7 1 2 3927 1445
0 1463 5 2 1 1462
0 1464 7 1 2 4963 4964
0 1465 5 1 1 1464
0 1466 7 1 2 3611 1465
0 1467 5 2 1 1466
0 1468 7 2 2 1461 4966
0 1469 5 2 1 4968
0 1470 7 2 2 4961 4965
0 1471 5 1 1 4972
0 1472 7 1 2 3612 1471
0 1473 5 1 1 1472
0 1474 7 1 2 4967 4973
0 1475 5 1 1 1474
0 1476 7 1 2 1473 1475
0 1477 5 2 1 1476
0 1478 7 1 2 4970 4974
0 1479 5 1 1 1478
0 1480 7 2 2 3605 1479
0 1481 5 1 1 4976
0 1482 7 1 2 4971 4977
0 1483 5 1 1 1482
0 1484 7 1 2 3913 4969
0 1485 5 1 1 1484
0 1486 7 2 2 1483 1485
0 1487 5 1 1 4978
0 1488 7 1 2 3906 1487
0 1489 5 1 1 1488
0 1490 7 1 2 3914 4975
0 1491 5 1 1 1490
0 1492 7 2 2 1481 1491
0 1493 5 1 1 4980
0 1494 7 1 2 3598 4981
0 1495 5 2 1 1494
0 1496 7 1 2 3599 4979
0 1497 7 1 2 4982 1496
0 1498 5 2 1 1497
0 1499 7 3 2 1489 4984
0 1500 5 1 1 4986
0 1501 7 1 2 3907 1493
0 1502 5 1 1 1501
0 1503 7 1 2 4983 1502
0 1504 7 1 2 4985 1503
0 1505 5 2 1 1504
0 1506 7 1 2 4987 4989
0 1507 5 1 1 1506
0 1508 7 1 2 3591 1507
0 1509 5 2 1 1508
0 1510 7 1 2 3900 4990
0 1511 5 1 1 1510
0 1512 7 2 2 4991 1511
0 1513 5 2 1 4993
0 1514 7 1 2 3592 1500
0 1515 5 1 1 1514
0 1516 7 1 2 4988 4992
0 1517 5 1 1 1516
0 1518 7 1 2 1515 1517
0 1519 5 2 1 1518
0 1520 7 1 2 4995 4997
0 1521 5 1 1 1520
0 1522 7 2 2 3585 1521
0 1523 5 1 1 4999
0 1524 7 1 2 4996 5000
0 1525 5 1 1 1524
0 1526 7 1 2 3893 4994
0 1527 5 1 1 1526
0 1528 7 2 2 1525 1527
0 1529 5 1 1 5001
0 1530 7 1 2 3894 4998
0 1531 5 1 1 1530
0 1532 7 2 2 1523 1531
0 1533 5 1 1 5003
0 1534 7 2 2 3579 1533
0 1535 5 1 1 5005
0 1536 7 1 2 5002 5006
0 1537 5 2 1 1536
0 1538 7 1 2 3886 5004
0 1539 5 1 1 1538
0 1540 7 2 2 1535 1539
0 1541 5 1 1 5009
0 1542 7 1 2 5007 1541
0 1543 5 1 1 1542
0 1544 7 1 2 3880 1543
0 1545 5 1 1 1544
0 1546 7 1 2 3887 1529
0 1547 5 2 1 1546
0 1548 7 1 2 5010 5011
0 1549 5 1 1 1548
0 1550 7 1 2 3572 1549
0 1551 5 2 1 1550
0 1552 7 2 2 1545 5013
0 1553 5 2 1 5015
0 1554 7 2 2 5008 5012
0 1555 5 1 1 5019
0 1556 7 1 2 3573 1555
0 1557 5 1 1 1556
0 1558 7 1 2 5014 5020
0 1559 5 1 1 1558
0 1560 7 1 2 1557 1559
0 1561 5 2 1 1560
0 1562 7 1 2 5017 5021
0 1563 5 1 1 1562
0 1564 7 2 2 3566 1563
0 1565 5 1 1 5023
0 1566 7 1 2 5018 5024
0 1567 5 1 1 1566
0 1568 7 1 2 3873 5016
0 1569 5 1 1 1568
0 1570 7 2 2 1567 1569
0 1571 5 1 1 5025
0 1572 7 1 2 3867 1571
0 1573 5 1 1 1572
0 1574 7 1 2 3874 5022
0 1575 5 1 1 1574
0 1576 7 2 2 1565 1575
0 1577 5 1 1 5027
0 1578 7 1 2 3559 5028
0 1579 5 2 1 1578
0 1580 7 1 2 3560 5026
0 1581 7 1 2 5029 1580
0 1582 5 2 1 1581
0 1583 7 3 2 1573 5031
0 1584 5 1 1 5033
0 1585 7 1 2 3868 1577
0 1586 5 1 1 1585
0 1587 7 1 2 5030 1586
0 1588 7 1 2 5032 1587
0 1589 5 2 1 1588
0 1590 7 1 2 5034 5036
0 1591 5 1 1 1590
0 1592 7 1 2 3552 1591
0 1593 5 2 1 1592
0 1594 7 1 2 3862 5037
0 1595 5 1 1 1594
0 1596 7 2 2 5038 1595
0 1597 5 2 1 5040
0 1598 7 1 2 3553 1584
0 1599 5 1 1 1598
0 1600 7 1 2 5035 5039
0 1601 5 1 1 1600
0 1602 7 1 2 1599 1601
0 1603 5 2 1 1602
0 1604 7 1 2 5042 5044
0 1605 5 1 1 1604
0 1606 7 2 2 3546 1605
0 1607 5 1 1 5046
0 1608 7 1 2 5043 5047
0 1609 5 1 1 1608
0 1610 7 1 2 3856 5041
0 1611 5 1 1 1610
0 1612 7 2 2 1609 1611
0 1613 5 1 1 5048
0 1614 7 1 2 3857 5045
0 1615 5 1 1 1614
0 1616 7 2 2 1607 1615
0 1617 5 1 1 5050
0 1618 7 2 2 3540 1617
0 1619 5 1 1 5052
0 1620 7 1 2 5049 5053
0 1621 5 2 1 1620
0 1622 7 1 2 3850 5051
0 1623 5 1 1 1622
0 1624 7 2 2 1619 1623
0 1625 5 1 1 5056
0 1626 7 1 2 5054 1625
0 1627 5 1 1 1626
0 1628 7 1 2 3845 1627
0 1629 5 1 1 1628
0 1630 7 1 2 3851 1613
0 1631 5 2 1 1630
0 1632 7 1 2 5057 5058
0 1633 5 1 1 1632
0 1634 7 1 2 3533 1633
0 1635 5 2 1 1634
0 1636 7 2 2 1629 5060
0 1637 5 2 1 5062
0 1638 7 2 2 5055 5059
0 1639 5 1 1 5066
0 1640 7 1 2 3534 1639
0 1641 5 1 1 1640
0 1642 7 1 2 5061 5067
0 1643 5 1 1 1642
0 1644 7 1 2 1641 1643
0 1645 5 2 1 1644
0 1646 7 1 2 5064 5068
0 1647 5 1 1 1646
0 1648 7 2 2 3527 1647
0 1649 5 1 1 5070
0 1650 7 1 2 5065 5071
0 1651 5 1 1 1650
0 1652 7 1 2 3839 5063
0 1653 5 1 1 1652
0 1654 7 2 2 1651 1653
0 1655 5 1 1 5072
0 1656 7 1 2 3833 1655
0 1657 5 1 1 1656
0 1658 7 1 2 3840 5069
0 1659 5 1 1 1658
0 1660 7 2 2 1649 1659
0 1661 5 1 1 5074
0 1662 7 1 2 3520 5075
0 1663 5 2 1 1662
0 1664 7 1 2 3521 5073
0 1665 7 1 2 5076 1664
0 1666 5 2 1 1665
0 1667 7 3 2 1657 5078
0 1668 5 1 1 5080
0 1669 7 1 2 3834 1661
0 1670 5 1 1 1669
0 1671 7 1 2 5077 1670
0 1672 7 1 2 5079 1671
0 1673 5 2 1 1672
0 1674 7 1 2 5081 5083
0 1675 5 1 1 1674
0 1676 7 1 2 3513 1675
0 1677 5 2 1 1676
0 1678 7 1 2 3828 5084
0 1679 5 1 1 1678
0 1680 7 2 2 5085 1679
0 1681 5 2 1 5087
0 1682 7 1 2 3514 1668
0 1683 5 1 1 1682
0 1684 7 1 2 5082 5086
0 1685 5 1 1 1684
0 1686 7 1 2 1683 1685
0 1687 5 2 1 1686
0 1688 7 1 2 5089 5091
0 1689 5 1 1 1688
0 1690 7 2 2 3507 1689
0 1691 5 1 1 5093
0 1692 7 1 2 5090 5094
0 1693 5 1 1 1692
0 1694 7 1 2 3822 5088
0 1695 5 1 1 1694
0 1696 7 2 2 1693 1695
0 1697 5 1 1 5095
0 1698 7 1 2 3823 5092
0 1699 5 1 1 1698
0 1700 7 2 2 1691 1699
0 1701 5 1 1 5097
0 1702 7 2 2 3501 1701
0 1703 5 1 1 5099
0 1704 7 1 2 5096 5100
0 1705 5 2 1 1704
0 1706 7 1 2 3816 5098
0 1707 5 1 1 1706
0 1708 7 2 2 1703 1707
0 1709 5 1 1 5103
0 1710 7 1 2 5101 1709
0 1711 5 1 1 1710
0 1712 7 1 2 3811 1711
0 1713 5 1 1 1712
0 1714 7 1 2 3817 1697
0 1715 5 2 1 1714
0 1716 7 1 2 5104 5105
0 1717 5 1 1 1716
0 1718 7 1 2 3494 1717
0 1719 5 2 1 1718
0 1720 7 2 2 1713 5107
0 1721 5 2 1 5109
0 1722 7 2 2 5102 5106
0 1723 5 1 1 5113
0 1724 7 1 2 3495 1723
0 1725 5 1 1 1724
0 1726 7 1 2 5108 5114
0 1727 5 1 1 1726
0 1728 7 1 2 1725 1727
0 1729 5 2 1 1728
0 1730 7 1 2 5111 5115
0 1731 5 1 1 1730
0 1732 7 2 2 3488 1731
0 1733 5 1 1 5117
0 1734 7 1 2 5112 5118
0 1735 5 1 1 1734
0 1736 7 1 2 3805 5110
0 1737 5 1 1 1736
0 1738 7 2 2 1735 1737
0 1739 5 1 1 5119
0 1740 7 1 2 3799 1739
0 1741 5 1 1 1740
0 1742 7 1 2 3806 5116
0 1743 5 1 1 1742
0 1744 7 2 2 1733 1743
0 1745 5 1 1 5121
0 1746 7 1 2 3481 5122
0 1747 5 2 1 1746
0 1748 7 1 2 3482 5120
0 1749 7 1 2 5123 1748
0 1750 5 2 1 1749
0 1751 7 3 2 1741 5125
0 1752 5 1 1 5127
0 1753 7 1 2 3474 1752
0 1754 5 1 1 1753
0 1755 7 1 2 3800 1745
0 1756 5 1 1 1755
0 1757 7 1 2 5124 1756
0 1758 7 1 2 5126 1757
0 1759 5 2 1 1758
0 1760 7 1 2 5128 5130
0 1761 5 1 1 1760
0 1762 7 1 2 3475 1761
0 1763 5 2 1 1762
0 1764 7 1 2 5129 5132
0 1765 5 1 1 1764
0 1766 7 1 2 1754 1765
0 1767 5 2 1 1766
0 1768 7 1 2 3788 5134
0 1769 5 1 1 1768
0 1770 7 1 2 3794 5131
0 1771 5 1 1 1770
0 1772 7 2 2 5133 1771
0 1773 5 2 1 5136
0 1774 7 1 2 5135 5138
0 1775 5 1 1 1774
0 1776 7 2 2 3468 1775
0 1777 5 1 1 5140
0 1778 7 2 2 1769 1777
0 1779 5 2 1 5142
0 1780 7 1 2 5139 5141
0 1781 5 1 1 1780
0 1782 7 1 2 3789 5137
0 1783 5 1 1 1782
0 1784 7 2 2 1781 1783
0 1785 7 1 2 5144 5146
0 1786 5 1 1 1785
0 1787 7 2 2 3462 1786
0 1788 5 1 1 5148
0 1789 7 1 2 5145 5149
0 1790 5 1 1 1789
0 1791 7 1 2 3782 5143
0 1792 5 1 1 1791
0 1793 7 2 2 1790 1792
0 1794 7 1 2 3776 5150
0 1795 5 1 1 1794
0 1796 7 1 2 3783 5147
0 1797 5 1 1 1796
0 1798 7 2 2 1788 1797
0 1799 5 2 1 5152
0 1800 7 1 2 5151 5154
0 1801 5 1 1 1800
0 1802 7 2 2 3456 1801
0 1803 5 1 1 5156
0 1804 7 2 2 1795 1803
0 1805 5 1 1 5158
0 1806 7 1 2 5155 5157
0 1807 5 1 1 1806
0 1808 7 1 2 3777 5153
0 1809 5 1 1 1808
0 1810 7 1 2 3770 1809
0 1811 7 1 2 1807 1810
0 1812 5 1 1 1811
0 1813 7 1 2 1805 1812
0 1814 5 1 1 1813
0 1815 7 1 2 3771 5159
0 1816 5 1 1 1815
0 1817 7 1 2 3764 1816
0 1818 7 1 2 1814 1817
0 1819 5 1 1 1818
0 1820 7 2 2 3746 3755
0 1821 5 1 1 5160
0 1822 7 1 2 3760 1821
0 1823 5 2 1 1822
0 1824 7 1 2 4035 5162
0 1825 5 1 1 1824
0 1826 7 1 2 135 5163
0 1827 5 1 1 1826
0 1828 7 1 2 3739 1827
0 1829 5 3 1 1828
0 1830 7 5 2 1825 5164
0 1831 5 1 1 5167
0 1832 7 2 2 3761 5161
0 1833 5 2 1 5172
0 1834 7 2 2 3740 3747
0 1835 5 1 1 5176
0 1836 7 1 2 4043 1835
0 1837 5 1 1 1836
0 1838 7 1 2 4047 5177
0 1839 5 1 1 1838
0 1840 7 1 2 1837 1839
0 1841 7 2 2 5174 1840
0 1842 5 2 1 5178
0 1843 7 1 2 4029 5180
0 1844 5 1 1 1843
0 1845 7 1 2 4040 5175
0 1846 5 1 1 1845
0 1847 7 1 2 3748 5173
0 1848 5 1 1 1847
0 1849 7 3 2 1846 1848
0 1850 5 1 1 5182
0 1851 7 1 2 5168 5183
0 1852 5 1 1 1851
0 1853 7 1 2 5181 1852
0 1854 5 1 1 1853
0 1855 7 2 2 3731 1854
0 1856 5 2 1 5185
0 1857 7 2 2 1844 5187
0 1858 5 1 1 5189
0 1859 7 2 2 3724 5190
0 1860 7 1 2 5169 5191
0 1861 5 2 1 1860
0 1862 7 2 2 3732 5170
0 1863 5 1 1 5195
0 1864 7 1 2 5179 5196
0 1865 5 1 1 1864
0 1866 7 1 2 5165 1865
0 1867 5 1 1 1866
0 1868 7 1 2 1850 1867
0 1869 5 1 1 1868
0 1870 7 1 2 5166 5184
0 1871 7 1 2 1863 1870
0 1872 5 1 1 1871
0 1873 7 2 2 1869 1872
0 1874 7 1 2 5193 5197
0 1875 5 2 1 1874
0 1876 7 1 2 3725 5199
0 1877 5 2 1 1876
0 1878 7 1 2 4023 5198
0 1879 5 1 1 1878
0 1880 7 4 2 5201 1879
0 1881 5 1 1 5203
0 1882 7 1 2 1858 5202
0 1883 5 1 1 1882
0 1884 7 1 2 5192 5200
0 1885 5 2 1 1884
0 1886 7 2 2 1883 5207
0 1887 5 1 1 5209
0 1888 7 1 2 3717 5204
0 1889 7 1 2 5210 1888
0 1890 5 2 1 1889
0 1891 7 1 2 5171 5188
0 1892 5 1 1 1891
0 1893 7 1 2 1831 5186
0 1894 5 1 1 1893
0 1895 7 1 2 1892 1894
0 1896 7 1 2 5208 1895
0 1897 5 1 1 1896
0 1898 7 1 2 5194 1897
0 1899 5 2 1 1898
0 1900 7 1 2 5211 5213
0 1901 5 1 1 1900
0 1902 7 2 2 3718 1901
0 1903 5 2 1 5215
0 1904 7 1 2 4018 5214
0 1905 5 1 1 1904
0 1906 7 3 2 5217 1905
0 1907 5 1 1 5219
0 1908 7 2 2 3710 5220
0 1909 7 1 2 5205 5222
0 1910 5 2 1 1909
0 1911 7 1 2 5206 5216
0 1912 5 2 1 1911
0 1913 7 1 2 1881 5218
0 1914 5 1 1 1913
0 1915 7 1 2 5226 1914
0 1916 5 1 1 1915
0 1917 7 1 2 1887 5227
0 1918 5 1 1 1917
0 1919 7 2 2 5212 1918
0 1920 5 2 1 5228
0 1921 7 1 2 5223 5229
0 1922 5 1 1 1921
0 1923 7 1 2 1916 1922
0 1924 5 1 1 1923
0 1925 7 1 2 5224 1924
0 1926 5 2 1 1925
0 1927 7 1 2 5225 5230
0 1928 5 1 1 1927
0 1929 7 2 2 3711 1928
0 1930 5 2 1 5234
0 1931 7 1 2 5221 5236
0 1932 5 1 1 1931
0 1933 7 1 2 1907 5235
0 1934 5 1 1 1933
0 1935 7 2 2 1932 1934
0 1936 5 1 1 5238
0 1937 7 1 2 4012 5231
0 1938 5 1 1 1937
0 1939 7 4 2 5237 1938
0 1940 5 1 1 5240
0 1941 7 1 2 3703 5241
0 1942 7 1 2 1936 1941
0 1943 5 2 1 1942
0 1944 7 1 2 5232 5244
0 1945 5 1 1 1944
0 1946 7 2 2 3704 1945
0 1947 5 2 1 5246
0 1948 7 1 2 4007 5233
0 1949 5 1 1 1948
0 1950 7 3 2 5248 1949
0 1951 5 1 1 5250
0 1952 7 1 2 5242 5247
0 1953 5 2 1 1952
0 1954 7 1 2 5239 5253
0 1955 5 1 1 1954
0 1956 7 1 2 5245 1955
0 1957 5 2 1 1956
0 1958 7 2 2 3697 5251
0 1959 7 1 2 5243 5257
0 1960 5 2 1 1959
0 1961 7 1 2 5255 5259
0 1962 5 2 1 1961
0 1963 7 1 2 3698 5261
0 1964 5 2 1 1963
0 1965 7 1 2 4001 5256
0 1966 5 1 1 1965
0 1967 7 4 2 5263 1966
0 1968 5 1 1 5265
0 1969 7 2 2 3691 5266
0 1970 7 1 2 5252 5269
0 1971 5 2 1 1970
0 1972 7 1 2 1951 5264
0 1973 5 1 1 1972
0 1974 7 1 2 5258 5262
0 1975 5 2 1 1974
0 1976 7 1 2 1973 5273
0 1977 5 1 1 1976
0 1978 7 1 2 1940 5249
0 1979 5 1 1 1978
0 1980 7 1 2 5254 1979
0 1981 5 1 1 1980
0 1982 7 1 2 5274 1981
0 1983 5 1 1 1982
0 1984 7 2 2 5260 1983
0 1985 5 2 1 5275
0 1986 7 1 2 5270 5276
0 1987 5 1 1 1986
0 1988 7 1 2 1977 1987
0 1989 5 1 1 1988
0 1990 7 1 2 5271 1989
0 1991 5 2 1 1990
0 1992 7 1 2 5272 5277
0 1993 5 1 1 1992
0 1994 7 2 2 3692 1993
0 1995 5 2 1 5281
0 1996 7 1 2 3995 5278
0 1997 5 1 1 1996
0 1998 7 2 2 5283 1997
0 1999 5 1 1 5285
0 2000 7 2 2 3684 5286
0 2001 7 1 2 5267 5287
0 2002 5 2 1 2001
0 2003 7 1 2 5279 5289
0 2004 5 2 1 2003
0 2005 7 1 2 3685 5291
0 2006 5 2 1 2005
0 2007 7 1 2 3990 5280
0 2008 5 1 1 2007
0 2009 7 4 2 5293 2008
0 2010 5 1 1 5295
0 2011 7 1 2 1999 5294
0 2012 5 1 1 2011
0 2013 7 1 2 5288 5292
0 2014 5 2 1 2013
0 2015 7 2 2 2012 5299
0 2016 5 1 1 5301
0 2017 7 1 2 3678 5296
0 2018 7 1 2 5302 2017
0 2019 5 2 1 2018
0 2020 7 1 2 5268 5284
0 2021 5 1 1 2020
0 2022 7 1 2 1968 5282
0 2023 5 1 1 2022
0 2024 7 1 2 2021 2023
0 2025 7 1 2 5300 2024
0 2026 5 1 1 2025
0 2027 7 1 2 5290 2026
0 2028 5 2 1 2027
0 2029 7 1 2 5303 5305
0 2030 5 1 1 2029
0 2031 7 2 2 3679 2030
0 2032 5 2 1 5307
0 2033 7 1 2 3984 5306
0 2034 5 1 1 2033
0 2035 7 3 2 5309 2034
0 2036 5 1 1 5311
0 2037 7 2 2 3671 5312
0 2038 7 1 2 5297 5314
0 2039 5 2 1 2038
0 2040 7 1 2 5298 5308
0 2041 5 2 1 2040
0 2042 7 1 2 2010 5310
0 2043 5 1 1 2042
0 2044 7 1 2 5318 2043
0 2045 5 1 1 2044
0 2046 7 1 2 2016 5319
0 2047 5 1 1 2046
0 2048 7 2 2 5304 2047
0 2049 5 2 1 5320
0 2050 7 1 2 5315 5321
0 2051 5 1 1 2050
0 2052 7 1 2 2045 2051
0 2053 5 1 1 2052
0 2054 7 1 2 5316 2053
0 2055 5 2 1 2054
0 2056 7 1 2 5317 5322
0 2057 5 1 1 2056
0 2058 7 2 2 3672 2057
0 2059 5 2 1 5326
0 2060 7 1 2 5313 5328
0 2061 5 1 1 2060
0 2062 7 1 2 2036 5327
0 2063 5 1 1 2062
0 2064 7 2 2 2061 2063
0 2065 5 1 1 5330
0 2066 7 1 2 3978 5323
0 2067 5 1 1 2066
0 2068 7 4 2 5329 2067
0 2069 5 1 1 5332
0 2070 7 1 2 3664 5333
0 2071 7 1 2 2065 2070
0 2072 5 2 1 2071
0 2073 7 1 2 5324 5336
0 2074 5 1 1 2073
0 2075 7 2 2 3665 2074
0 2076 5 2 1 5338
0 2077 7 1 2 3973 5325
0 2078 5 1 1 2077
0 2079 7 3 2 5340 2078
0 2080 5 1 1 5342
0 2081 7 1 2 5334 5339
0 2082 5 2 1 2081
0 2083 7 1 2 5331 5345
0 2084 5 1 1 2083
0 2085 7 1 2 5337 2084
0 2086 5 2 1 2085
0 2087 7 2 2 3658 5343
0 2088 7 1 2 5335 5349
0 2089 5 2 1 2088
0 2090 7 1 2 5347 5351
0 2091 5 2 1 2090
0 2092 7 1 2 3659 5353
0 2093 5 2 1 2092
0 2094 7 1 2 3967 5348
0 2095 5 1 1 2094
0 2096 7 4 2 5355 2095
0 2097 5 1 1 5357
0 2098 7 2 2 3652 5358
0 2099 7 1 2 5344 5361
0 2100 5 2 1 2099
0 2101 7 1 2 2080 5356
0 2102 5 1 1 2101
0 2103 7 1 2 5350 5354
0 2104 5 2 1 2103
0 2105 7 1 2 2102 5365
0 2106 5 1 1 2105
0 2107 7 1 2 2069 5341
0 2108 5 1 1 2107
0 2109 7 1 2 5346 2108
0 2110 5 1 1 2109
0 2111 7 1 2 5366 2110
0 2112 5 1 1 2111
0 2113 7 2 2 5352 2112
0 2114 5 2 1 5367
0 2115 7 1 2 5362 5368
0 2116 5 1 1 2115
0 2117 7 1 2 2106 2116
0 2118 5 1 1 2117
0 2119 7 1 2 5363 2118
0 2120 5 2 1 2119
0 2121 7 1 2 5364 5369
0 2122 5 1 1 2121
0 2123 7 2 2 3653 2122
0 2124 5 2 1 5373
0 2125 7 1 2 3961 5370
0 2126 5 1 1 2125
0 2127 7 4 2 5375 2126
0 2128 5 1 1 5377
0 2129 7 1 2 3645 5359
0 2130 7 1 2 5378 2129
0 2131 5 2 1 2130
0 2132 7 1 2 5371 5381
0 2133 5 1 1 2132
0 2134 7 2 2 3646 2133
0 2135 5 2 1 5383
0 2136 7 1 2 3955 5372
0 2137 5 1 1 2136
0 2138 7 4 2 5385 2137
0 2139 5 1 1 5387
0 2140 7 1 2 3639 5379
0 2141 7 1 2 5388 2140
0 2142 5 2 1 2141
0 2143 7 1 2 5380 5384
0 2144 5 2 1 2143
0 2145 7 1 2 5360 5376
0 2146 5 1 1 2145
0 2147 7 1 2 2097 5374
0 2148 5 1 1 2147
0 2149 7 1 2 2146 2148
0 2150 7 1 2 5393 2149
0 2151 5 1 1 2150
0 2152 7 1 2 5382 2151
0 2153 5 2 1 2152
0 2154 7 1 2 5391 5395
0 2155 5 1 1 2154
0 2156 7 2 2 3640 2155
0 2157 5 2 1 5397
0 2158 7 1 2 3948 5396
0 2159 5 1 1 2158
0 2160 7 4 2 5399 2159
0 2161 5 1 1 5401
0 2162 7 2 2 3632 5402
0 2163 7 1 2 5389 5405
0 2164 5 2 1 2163
0 2165 7 1 2 2139 5400
0 2166 5 1 1 2165
0 2167 7 1 2 5390 5398
0 2168 5 2 1 2167
0 2169 7 1 2 2166 5409
0 2170 5 1 1 2169
0 2171 7 1 2 2128 5386
0 2172 5 1 1 2171
0 2173 7 1 2 5394 2172
0 2174 5 1 1 2173
0 2175 7 1 2 5410 2174
0 2176 5 1 1 2175
0 2177 7 2 2 5392 2176
0 2178 5 2 1 5411
0 2179 7 1 2 5406 5412
0 2180 5 1 1 2179
0 2181 7 1 2 2170 2180
0 2182 5 1 1 2181
0 2183 7 1 2 5407 2182
0 2184 5 2 1 2183
0 2185 7 1 2 5408 5413
0 2186 5 1 1 2185
0 2187 7 2 2 3633 2186
0 2188 5 2 1 5417
0 2189 7 1 2 3941 5414
0 2190 5 1 1 2189
0 2191 7 3 2 5419 2190
0 2192 5 1 1 5421
0 2193 7 2 2 3625 5422
0 2194 7 1 2 5403 5424
0 2195 5 2 1 2194
0 2196 7 1 2 5415 5426
0 2197 5 2 1 2196
0 2198 7 1 2 3626 5428
0 2199 5 2 1 2198
0 2200 7 1 2 3935 5416
0 2201 5 1 1 2200
0 2202 7 4 2 5430 2201
0 2203 5 1 1 5432
0 2204 7 1 2 3619 5423
0 2205 7 1 2 5433 2204
0 2206 5 2 1 2205
0 2207 7 1 2 5425 5429
0 2208 5 2 1 2207
0 2209 7 1 2 5404 5420
0 2210 5 1 1 2209
0 2211 7 1 2 2161 5418
0 2212 5 1 1 2211
0 2213 7 1 2 2210 2212
0 2214 7 1 2 5438 2213
0 2215 5 1 1 2214
0 2216 7 1 2 5427 2215
0 2217 5 2 1 2216
0 2218 7 1 2 5436 5440
0 2219 5 1 1 2218
0 2220 7 2 2 3620 2219
0 2221 5 2 1 5442
0 2222 7 1 2 3928 5441
0 2223 5 1 1 2222
0 2224 7 4 2 5444 2223
0 2225 5 1 1 5446
0 2226 7 2 2 3613 5447
0 2227 7 1 2 5434 5450
0 2228 5 2 1 2227
0 2229 7 1 2 2203 5445
0 2230 5 1 1 2229
0 2231 7 1 2 5435 5443
0 2232 5 2 1 2231
0 2233 7 1 2 2230 5454
0 2234 5 1 1 2233
0 2235 7 1 2 2192 5431
0 2236 5 1 1 2235
0 2237 7 1 2 5439 2236
0 2238 5 1 1 2237
0 2239 7 1 2 5455 2238
0 2240 5 1 1 2239
0 2241 7 2 2 5437 2240
0 2242 5 2 1 5456
0 2243 7 1 2 5451 5457
0 2244 5 1 1 2243
0 2245 7 1 2 2234 2244
0 2246 5 1 1 2245
0 2247 7 1 2 5452 2246
0 2248 5 2 1 2247
0 2249 7 1 2 5453 5458
0 2250 5 1 1 2249
0 2251 7 2 2 3614 2250
0 2252 5 2 1 5462
0 2253 7 1 2 3921 5459
0 2254 5 1 1 2253
0 2255 7 4 2 5464 2254
0 2256 5 1 1 5466
0 2257 7 1 2 3606 5448
0 2258 7 1 2 5467 2257
0 2259 5 2 1 2258
0 2260 7 1 2 5460 5470
0 2261 5 1 1 2260
0 2262 7 2 2 3607 2261
0 2263 5 2 1 5472
0 2264 7 1 2 3915 5461
0 2265 5 1 1 2264
0 2266 7 4 2 5474 2265
0 2267 5 1 1 5476
0 2268 7 1 2 3600 5468
0 2269 7 1 2 5477 2268
0 2270 5 2 1 2269
0 2271 7 1 2 5469 5473
0 2272 5 2 1 2271
0 2273 7 1 2 5449 5465
0 2274 5 1 1 2273
0 2275 7 1 2 2225 5463
0 2276 5 1 1 2275
0 2277 7 1 2 2274 2276
0 2278 7 1 2 5482 2277
0 2279 5 1 1 2278
0 2280 7 1 2 5471 2279
0 2281 5 2 1 2280
0 2282 7 1 2 5480 5484
0 2283 5 1 1 2282
0 2284 7 2 2 3601 2283
0 2285 5 2 1 5486
0 2286 7 1 2 3908 5485
0 2287 5 1 1 2286
0 2288 7 4 2 5488 2287
0 2289 5 1 1 5490
0 2290 7 2 2 3593 5491
0 2291 7 1 2 5478 5494
0 2292 5 2 1 2291
0 2293 7 1 2 2267 5489
0 2294 5 1 1 2293
0 2295 7 1 2 5479 5487
0 2296 5 2 1 2295
0 2297 7 1 2 2294 5498
0 2298 5 1 1 2297
0 2299 7 1 2 2256 5475
0 2300 5 1 1 2299
0 2301 7 1 2 5483 2300
0 2302 5 1 1 2301
0 2303 7 1 2 5499 2302
0 2304 5 1 1 2303
0 2305 7 2 2 5481 2304
0 2306 5 2 1 5500
0 2307 7 1 2 5495 5501
0 2308 5 1 1 2307
0 2309 7 1 2 2298 2308
0 2310 5 1 1 2309
0 2311 7 1 2 5496 2310
0 2312 5 2 1 2311
0 2313 7 1 2 5497 5502
0 2314 5 1 1 2313
0 2315 7 2 2 3594 2314
0 2316 5 2 1 5506
0 2317 7 1 2 3901 5503
0 2318 5 1 1 2317
0 2319 7 4 2 5508 2318
0 2320 5 1 1 5510
0 2321 7 1 2 3586 5492
0 2322 7 1 2 5511 2321
0 2323 5 2 1 2322
0 2324 7 1 2 5504 5514
0 2325 5 1 1 2324
0 2326 7 2 2 3587 2325
0 2327 5 2 1 5516
0 2328 7 1 2 3895 5505
0 2329 5 1 1 2328
0 2330 7 3 2 5518 2329
0 2331 5 1 1 5520
0 2332 7 2 2 3580 5521
0 2333 7 1 2 5512 5523
0 2334 5 2 1 2333
0 2335 7 1 2 5513 5517
0 2336 5 2 1 2335
0 2337 7 1 2 5493 5509
0 2338 5 1 1 2337
0 2339 7 1 2 2289 5507
0 2340 5 1 1 2339
0 2341 7 1 2 2338 2340
0 2342 7 1 2 5527 2341
0 2343 5 1 1 2342
0 2344 7 1 2 5515 2343
0 2345 5 2 1 2344
0 2346 7 1 2 5525 5529
0 2347 5 2 1 2346
0 2348 7 1 2 3581 5531
0 2349 5 2 1 2348
0 2350 7 1 2 3888 5530
0 2351 5 1 1 2350
0 2352 7 4 2 5533 2351
0 2353 5 1 1 5535
0 2354 7 2 2 3574 5536
0 2355 7 1 2 5522 5539
0 2356 5 2 1 2355
0 2357 7 1 2 2331 5534
0 2358 5 1 1 2357
0 2359 7 1 2 5524 5532
0 2360 5 2 1 2359
0 2361 7 1 2 2358 5543
0 2362 5 1 1 2361
0 2363 7 1 2 2320 5519
0 2364 5 1 1 2363
0 2365 7 1 2 5528 2364
0 2366 5 1 1 2365
0 2367 7 1 2 5544 2366
0 2368 5 1 1 2367
0 2369 7 2 2 5526 2368
0 2370 5 2 1 5545
0 2371 7 1 2 5540 5546
0 2372 5 1 1 2371
0 2373 7 1 2 2362 2372
0 2374 5 1 1 2373
0 2375 7 1 2 5541 2374
0 2376 5 2 1 2375
0 2377 7 1 2 5542 5547
0 2378 5 1 1 2377
0 2379 7 2 2 3575 2378
0 2380 5 2 1 5551
0 2381 7 1 2 3881 5548
0 2382 5 1 1 2381
0 2383 7 4 2 5553 2382
0 2384 5 1 1 5555
0 2385 7 1 2 3567 5537
0 2386 7 1 2 5556 2385
0 2387 5 2 1 2386
0 2388 7 1 2 5549 5559
0 2389 5 1 1 2388
0 2390 7 2 2 3568 2389
0 2391 5 2 1 5561
0 2392 7 1 2 3875 5550
0 2393 5 1 1 2392
0 2394 7 4 2 5563 2393
0 2395 5 1 1 5565
0 2396 7 1 2 3561 5557
0 2397 7 1 2 5566 2396
0 2398 5 2 1 2397
0 2399 7 1 2 5558 5562
0 2400 5 2 1 2399
0 2401 7 1 2 5538 5554
0 2402 5 1 1 2401
0 2403 7 1 2 2353 5552
0 2404 5 1 1 2403
0 2405 7 1 2 2402 2404
0 2406 7 1 2 5571 2405
0 2407 5 1 1 2406
0 2408 7 1 2 5560 2407
0 2409 5 2 1 2408
0 2410 7 1 2 5569 5573
0 2411 5 1 1 2410
0 2412 7 2 2 3562 2411
0 2413 5 2 1 5575
0 2414 7 1 2 3869 5574
0 2415 5 1 1 2414
0 2416 7 4 2 5577 2415
0 2417 5 1 1 5579
0 2418 7 2 2 3554 5580
0 2419 7 1 2 5567 5583
0 2420 5 2 1 2419
0 2421 7 1 2 2395 5578
0 2422 5 1 1 2421
0 2423 7 1 2 5568 5576
0 2424 5 2 1 2423
0 2425 7 1 2 2422 5587
0 2426 5 1 1 2425
0 2427 7 1 2 2384 5564
0 2428 5 1 1 2427
0 2429 7 1 2 5572 2428
0 2430 5 1 1 2429
0 2431 7 1 2 5588 2430
0 2432 5 1 1 2431
0 2433 7 2 2 5570 2432
0 2434 5 2 1 5589
0 2435 7 1 2 5584 5590
0 2436 5 1 1 2435
0 2437 7 1 2 2426 2436
0 2438 5 1 1 2437
0 2439 7 1 2 5585 2438
0 2440 5 2 1 2439
0 2441 7 1 2 5586 5591
0 2442 5 1 1 2441
0 2443 7 2 2 3555 2442
0 2444 5 2 1 5595
0 2445 7 1 2 3863 5592
0 2446 5 1 1 2445
0 2447 7 4 2 5597 2446
0 2448 5 1 1 5599
0 2449 7 1 2 3547 5581
0 2450 7 1 2 5600 2449
0 2451 5 2 1 2450
0 2452 7 1 2 5593 5603
0 2453 5 1 1 2452
0 2454 7 2 2 3548 2453
0 2455 5 2 1 5605
0 2456 7 1 2 3858 5594
0 2457 5 1 1 2456
0 2458 7 3 2 5607 2457
0 2459 5 1 1 5609
0 2460 7 2 2 3541 5610
0 2461 7 1 2 5601 5612
0 2462 5 2 1 2461
0 2463 7 1 2 5602 5606
0 2464 5 2 1 2463
0 2465 7 1 2 5582 5598
0 2466 5 1 1 2465
0 2467 7 1 2 2417 5596
0 2468 5 1 1 2467
0 2469 7 1 2 2466 2468
0 2470 7 1 2 5616 2469
0 2471 5 1 1 2470
0 2472 7 1 2 5604 2471
0 2473 5 2 1 2472
0 2474 7 1 2 5614 5618
0 2475 5 2 1 2474
0 2476 7 1 2 3542 5620
0 2477 5 2 1 2476
0 2478 7 1 2 3852 5619
0 2479 5 1 1 2478
0 2480 7 4 2 5622 2479
0 2481 5 1 1 5624
0 2482 7 2 2 3535 5625
0 2483 7 1 2 5611 5628
0 2484 5 2 1 2483
0 2485 7 1 2 2459 5623
0 2486 5 1 1 2485
0 2487 7 1 2 5613 5621
0 2488 5 2 1 2487
0 2489 7 1 2 2486 5632
0 2490 5 1 1 2489
0 2491 7 1 2 2448 5608
0 2492 5 1 1 2491
0 2493 7 1 2 5617 2492
0 2494 5 1 1 2493
0 2495 7 1 2 5633 2494
0 2496 5 1 1 2495
0 2497 7 2 2 5615 2496
0 2498 5 2 1 5634
0 2499 7 1 2 5629 5635
0 2500 5 1 1 2499
0 2501 7 1 2 2490 2500
0 2502 5 1 1 2501
0 2503 7 1 2 5630 2502
0 2504 5 2 1 2503
0 2505 7 1 2 5631 5636
0 2506 5 1 1 2505
0 2507 7 2 2 3536 2506
0 2508 5 2 1 5640
0 2509 7 1 2 3846 5637
0 2510 5 1 1 2509
0 2511 7 4 2 5642 2510
0 2512 5 1 1 5644
0 2513 7 1 2 3528 5626
0 2514 7 1 2 5645 2513
0 2515 5 2 1 2514
0 2516 7 1 2 5638 5648
0 2517 5 1 1 2516
0 2518 7 2 2 3529 2517
0 2519 5 2 1 5650
0 2520 7 1 2 3841 5639
0 2521 5 1 1 2520
0 2522 7 4 2 5652 2521
0 2523 5 1 1 5654
0 2524 7 1 2 3522 5646
0 2525 7 1 2 5655 2524
0 2526 5 2 1 2525
0 2527 7 1 2 5647 5651
0 2528 5 2 1 2527
0 2529 7 1 2 5627 5643
0 2530 5 1 1 2529
0 2531 7 1 2 2481 5641
0 2532 5 1 1 2531
0 2533 7 1 2 2530 2532
0 2534 7 1 2 5660 2533
0 2535 5 1 1 2534
0 2536 7 1 2 5649 2535
0 2537 5 2 1 2536
0 2538 7 1 2 5658 5662
0 2539 5 1 1 2538
0 2540 7 2 2 3523 2539
0 2541 5 2 1 5664
0 2542 7 1 2 3835 5663
0 2543 5 1 1 2542
0 2544 7 4 2 5666 2543
0 2545 5 1 1 5668
0 2546 7 2 2 3515 5669
0 2547 7 1 2 5656 5672
0 2548 5 2 1 2547
0 2549 7 1 2 2523 5667
0 2550 5 1 1 2549
0 2551 7 1 2 5657 5665
0 2552 5 2 1 2551
0 2553 7 1 2 2550 5676
0 2554 5 1 1 2553
0 2555 7 1 2 2512 5653
0 2556 5 1 1 2555
0 2557 7 1 2 5661 2556
0 2558 5 1 1 2557
0 2559 7 1 2 5677 2558
0 2560 5 1 1 2559
0 2561 7 2 2 5659 2560
0 2562 5 2 1 5678
0 2563 7 1 2 5673 5679
0 2564 5 1 1 2563
0 2565 7 1 2 2554 2564
0 2566 5 1 1 2565
0 2567 7 1 2 5674 2566
0 2568 5 2 1 2567
0 2569 7 1 2 5675 5680
0 2570 5 1 1 2569
0 2571 7 2 2 3516 2570
0 2572 5 2 1 5684
0 2573 7 1 2 3829 5681
0 2574 5 1 1 2573
0 2575 7 4 2 5686 2574
0 2576 5 1 1 5688
0 2577 7 1 2 3508 5670
0 2578 7 1 2 5689 2577
0 2579 5 2 1 2578
0 2580 7 1 2 5682 5692
0 2581 5 1 1 2580
0 2582 7 2 2 3509 2581
0 2583 5 2 1 5694
0 2584 7 1 2 3824 5683
0 2585 5 1 1 2584
0 2586 7 3 2 5696 2585
0 2587 5 1 1 5698
0 2588 7 2 2 3502 5699
0 2589 7 1 2 5690 5701
0 2590 5 2 1 2589
0 2591 7 1 2 5691 5695
0 2592 5 2 1 2591
0 2593 7 1 2 5671 5687
0 2594 5 1 1 2593
0 2595 7 1 2 2545 5685
0 2596 5 1 1 2595
0 2597 7 1 2 2594 2596
0 2598 7 1 2 5705 2597
0 2599 5 1 1 2598
0 2600 7 1 2 5693 2599
0 2601 5 2 1 2600
0 2602 7 1 2 5703 5707
0 2603 5 2 1 2602
0 2604 7 1 2 3503 5709
0 2605 5 2 1 2604
0 2606 7 1 2 3818 5708
0 2607 5 1 1 2606
0 2608 7 4 2 5711 2607
0 2609 5 1 1 5713
0 2610 7 2 2 3496 5714
0 2611 7 1 2 5700 5717
0 2612 5 2 1 2611
0 2613 7 1 2 2587 5712
0 2614 5 1 1 2613
0 2615 7 1 2 5702 5710
0 2616 5 2 1 2615
0 2617 7 1 2 2614 5721
0 2618 5 1 1 2617
0 2619 7 1 2 2576 5697
0 2620 5 1 1 2619
0 2621 7 1 2 5706 2620
0 2622 5 1 1 2621
0 2623 7 1 2 5722 2622
0 2624 5 1 1 2623
0 2625 7 2 2 5704 2624
0 2626 5 2 1 5723
0 2627 7 1 2 5718 5724
0 2628 5 1 1 2627
0 2629 7 1 2 2618 2628
0 2630 5 1 1 2629
0 2631 7 1 2 5719 2630
0 2632 5 2 1 2631
0 2633 7 1 2 5720 5725
0 2634 5 1 1 2633
0 2635 7 2 2 3497 2634
0 2636 5 2 1 5729
0 2637 7 1 2 3812 5726
0 2638 5 1 1 2637
0 2639 7 4 2 5731 2638
0 2640 5 1 1 5733
0 2641 7 1 2 3489 5715
0 2642 7 1 2 5734 2641
0 2643 5 2 1 2642
0 2644 7 1 2 5727 5737
0 2645 5 1 1 2644
0 2646 7 2 2 3490 2645
0 2647 5 2 1 5739
0 2648 7 1 2 3807 5728
0 2649 5 1 1 2648
0 2650 7 4 2 5741 2649
0 2651 5 1 1 5743
0 2652 7 1 2 3483 5735
0 2653 7 1 2 5744 2652
0 2654 5 2 1 2653
0 2655 7 1 2 5736 5740
0 2656 5 2 1 2655
0 2657 7 1 2 5716 5732
0 2658 5 1 1 2657
0 2659 7 1 2 2609 5730
0 2660 5 1 1 2659
0 2661 7 1 2 2658 2660
0 2662 7 1 2 5749 2661
0 2663 5 1 1 2662
0 2664 7 1 2 5738 2663
0 2665 5 2 1 2664
0 2666 7 1 2 5747 5751
0 2667 5 1 1 2666
0 2668 7 2 2 3484 2667
0 2669 5 2 1 5753
0 2670 7 1 2 3801 5752
0 2671 5 1 1 2670
0 2672 7 4 2 5755 2671
0 2673 5 1 1 5757
0 2674 7 2 2 3476 5758
0 2675 7 1 2 5745 5761
0 2676 5 2 1 2675
0 2677 7 1 2 5746 5754
0 2678 5 2 1 2677
0 2679 7 1 2 2640 5742
0 2680 5 1 1 2679
0 2681 7 1 2 5750 2680
0 2682 5 1 1 2681
0 2683 7 1 2 5765 2682
0 2684 5 1 1 2683
0 2685 7 2 2 5748 2684
0 2686 5 2 1 5767
0 2687 7 1 2 5763 5769
0 2688 5 1 1 2687
0 2689 7 2 2 3477 2688
0 2690 5 2 1 5771
0 2691 7 1 2 3795 5770
0 2692 5 1 1 2691
0 2693 7 4 2 5773 2692
0 2694 5 1 1 5775
0 2695 7 1 2 2651 5756
0 2696 5 1 1 2695
0 2697 7 1 2 5766 2696
0 2698 5 1 1 2697
0 2699 7 1 2 5762 5768
0 2700 5 1 1 2699
0 2701 7 1 2 2698 2700
0 2702 5 1 1 2701
0 2703 7 1 2 5764 2702
0 2704 5 2 1 2703
0 2705 7 1 2 3469 5759
0 2706 7 1 2 5776 2705
0 2707 5 2 1 2706
0 2708 7 1 2 5779 5781
0 2709 5 1 1 2708
0 2710 7 2 2 3470 2709
0 2711 5 2 1 5783
0 2712 7 1 2 3790 5780
0 2713 5 1 1 2712
0 2714 7 3 2 5785 2713
0 2715 5 1 1 5787
0 2716 7 2 2 3463 5788
0 2717 7 1 2 5777 5790
0 2718 5 2 1 2717
0 2719 7 1 2 5778 5784
0 2720 5 2 1 2719
0 2721 7 1 2 2694 5786
0 2722 5 1 1 2721
0 2723 7 1 2 5794 2722
0 2724 5 1 1 2723
0 2725 7 1 2 5760 5774
0 2726 5 1 1 2725
0 2727 7 1 2 2673 5772
0 2728 5 1 1 2727
0 2729 7 1 2 2726 2728
0 2730 7 1 2 5795 2729
0 2731 5 1 1 2730
0 2732 7 1 2 5782 2731
0 2733 5 2 1 2732
0 2734 7 1 2 5792 5796
0 2735 5 2 1 2734
0 2736 7 1 2 5791 5798
0 2737 5 2 1 2736
0 2738 7 1 2 2724 5800
0 2739 5 1 1 2738
0 2740 7 2 2 5793 2739
0 2741 5 2 1 5802
0 2742 7 1 2 3464 5799
0 2743 5 2 1 2742
0 2744 7 1 2 3784 5797
0 2745 5 1 1 2744
0 2746 7 4 2 5806 2745
0 2747 5 1 1 5808
0 2748 7 2 2 3457 5809
0 2749 7 1 2 5789 5812
0 2750 5 2 1 2749
0 2751 7 1 2 5804 5814
0 2752 5 1 1 2751
0 2753 7 2 2 3458 2752
0 2754 5 2 1 5816
0 2755 7 1 2 3778 5805
0 2756 5 1 1 2755
0 2757 7 3 2 5818 2756
0 2758 5 1 1 5820
0 2759 7 1 2 2715 5807
0 2760 5 1 1 2759
0 2761 7 1 2 5801 2760
0 2762 5 1 1 2761
0 2763 7 1 2 5803 5813
0 2764 5 1 1 2763
0 2765 7 1 2 2762 2764
0 2766 5 1 1 2765
0 2767 7 1 2 5815 2766
0 2768 5 2 1 2767
0 2769 7 1 2 3451 5810
0 2770 7 1 2 5821 2769
0 2771 5 2 1 2770
0 2772 7 1 2 5823 5825
0 2773 5 1 1 2772
0 2774 7 2 2 3452 2773
0 2775 5 2 1 5827
0 2776 7 1 2 2758 5829
0 2777 5 1 1 2776
0 2778 7 1 2 5822 5828
0 2779 5 2 1 2778
0 2780 7 2 2 2777 5831
0 2781 5 1 1 5833
0 2782 7 1 2 5811 5819
0 2783 5 1 1 2782
0 2784 7 1 2 2747 5817
0 2785 5 1 1 2784
0 2786 7 1 2 2783 2785
0 2787 7 1 2 5832 2786
0 2788 5 1 1 2787
0 2789 7 1 2 5826 2788
0 2790 5 1 1 2789
0 2791 7 1 2 3765 2790
0 2792 5 1 1 2791
0 2793 7 1 2 2781 2792
0 2794 5 1 1 2793
0 2795 7 1 2 3772 5824
0 2796 5 1 1 2795
0 2797 7 2 2 5830 2796
0 2798 5 1 1 5835
0 2799 7 1 2 5834 2798
0 2800 5 1 1 2799
0 2801 7 1 2 3766 5836
0 2802 5 1 1 2801
0 2803 7 1 2 2800 2802
0 2804 7 1 2 2794 2803
0 2805 5 1 1 2804
0 2806 7 1 2 1819 2805
0 2807 7 1 2 1188 2806
0 2808 7 2 2 1178 2807
0 2809 5 1 1 5837
0 2810 7 1 2 3779 3870
0 2811 5 2 1 2810
0 2812 7 1 2 3459 3563
0 2813 5 2 1 2812
0 2814 7 1 2 3773 3864
0 2815 5 2 1 2814
0 2816 7 1 2 3453 3556
0 2817 5 2 1 2816
0 2818 7 2 2 3448 3549
0 2819 5 3 1 5847
0 2820 7 1 2 5845 5849
0 2821 5 1 1 2820
0 2822 7 2 2 5843 2821
0 2823 5 2 1 5852
0 2824 7 1 2 5841 5854
0 2825 5 1 1 2824
0 2826 7 2 2 5839 2825
0 2827 5 1 1 5856
0 2828 7 1 2 3785 2827
0 2829 5 2 1 2828
0 2830 7 1 2 3465 5857
0 2831 5 2 1 2830
0 2832 7 1 2 3876 5860
0 2833 5 1 1 2832
0 2834 7 2 2 5858 2833
0 2835 5 1 1 5862
0 2836 7 1 2 3791 2835
0 2837 5 2 1 2836
0 2838 7 1 2 3471 5863
0 2839 5 2 1 2838
0 2840 7 1 2 3882 5866
0 2841 5 1 1 2840
0 2842 7 2 2 5864 2841
0 2843 5 1 1 5868
0 2844 7 1 2 3796 2843
0 2845 5 2 1 2844
0 2846 7 1 2 3478 5869
0 2847 5 2 1 2846
0 2848 7 1 2 3889 5872
0 2849 5 1 1 2848
0 2850 7 2 2 5870 2849
0 2851 5 1 1 5874
0 2852 7 1 2 3802 2851
0 2853 5 2 1 2852
0 2854 7 1 2 3485 5875
0 2855 5 2 1 2854
0 2856 7 1 2 3896 5878
0 2857 5 1 1 2856
0 2858 7 2 2 5876 2857
0 2859 5 1 1 5880
0 2860 7 1 2 3808 2859
0 2861 5 2 1 2860
0 2862 7 1 2 3491 5881
0 2863 5 2 1 2862
0 2864 7 1 2 3902 5884
0 2865 5 1 1 2864
0 2866 7 2 2 5882 2865
0 2867 5 1 1 5886
0 2868 7 1 2 3813 2867
0 2869 5 2 1 2868
0 2870 7 1 2 3498 5887
0 2871 5 2 1 2870
0 2872 7 1 2 3909 5890
0 2873 5 1 1 2872
0 2874 7 2 2 5888 2873
0 2875 5 1 1 5892
0 2876 7 1 2 3819 2875
0 2877 5 2 1 2876
0 2878 7 1 2 3504 5893
0 2879 5 2 1 2878
0 2880 7 1 2 3916 5896
0 2881 5 1 1 2880
0 2882 7 2 2 5894 2881
0 2883 5 1 1 5898
0 2884 7 1 2 3825 2883
0 2885 5 2 1 2884
0 2886 7 1 2 3510 5899
0 2887 5 2 1 2886
0 2888 7 1 2 3922 5902
0 2889 5 1 1 2888
0 2890 7 2 2 5900 2889
0 2891 5 1 1 5904
0 2892 7 1 2 3830 2891
0 2893 5 2 1 2892
0 2894 7 1 2 3517 5905
0 2895 5 2 1 2894
0 2896 7 1 2 3929 5908
0 2897 5 1 1 2896
0 2898 7 2 2 5906 2897
0 2899 5 1 1 5910
0 2900 7 1 2 3836 2899
0 2901 5 2 1 2900
0 2902 7 1 2 3524 5911
0 2903 5 2 1 2902
0 2904 7 1 2 3936 5914
0 2905 5 1 1 2904
0 2906 7 2 2 5912 2905
0 2907 5 1 1 5916
0 2908 7 1 2 3842 2907
0 2909 5 2 1 2908
0 2910 7 1 2 3530 5917
0 2911 5 2 1 2910
0 2912 7 1 2 3942 5920
0 2913 5 1 1 2912
0 2914 7 2 2 5918 2913
0 2915 5 1 1 5922
0 2916 7 1 2 3847 2915
0 2917 5 2 1 2916
0 2918 7 1 2 3537 5923
0 2919 5 2 1 2918
0 2920 7 2 2 5924 5926
0 2921 5 1 1 5928
0 2922 7 1 2 3641 5929
0 2923 5 1 1 2922
0 2924 7 1 2 3949 2921
0 2925 5 1 1 2924
0 2926 7 2 2 2923 2925
0 2927 5 1 1 5930
0 2928 7 1 2 3749 2927
0 2929 5 3 1 2928
0 2930 7 2 2 5919 5921
0 2931 5 1 1 5935
0 2932 7 1 2 3634 5936
0 2933 5 1 1 2932
0 2934 7 1 2 3943 2931
0 2935 5 1 1 2934
0 2936 7 2 2 2933 2935
0 2937 5 1 1 5937
0 2938 7 1 2 3741 2937
0 2939 5 3 1 2938
0 2940 7 1 2 4036 5938
0 2941 5 4 1 2940
0 2942 7 2 2 5913 5915
0 2943 5 1 1 5946
0 2944 7 1 2 3627 5947
0 2945 5 1 1 2944
0 2946 7 1 2 3937 2943
0 2947 5 1 1 2946
0 2948 7 2 2 2945 2947
0 2949 5 1 1 5948
0 2950 7 1 2 3733 2949
0 2951 5 3 1 2950
0 2952 7 1 2 4030 5949
0 2953 5 4 1 2952
0 2954 7 2 2 5907 5909
0 2955 5 1 1 5957
0 2956 7 1 2 3621 5958
0 2957 5 1 1 2956
0 2958 7 1 2 3930 2955
0 2959 5 1 1 2958
0 2960 7 2 2 2957 2959
0 2961 5 1 1 5959
0 2962 7 1 2 3726 2961
0 2963 5 4 1 2962
0 2964 7 1 2 4024 5960
0 2965 5 3 1 2964
0 2966 7 2 2 5901 5903
0 2967 5 1 1 5968
0 2968 7 1 2 3615 5969
0 2969 5 1 1 2968
0 2970 7 1 2 3923 2967
0 2971 5 1 1 2970
0 2972 7 2 2 2969 2971
0 2973 5 1 1 5970
0 2974 7 1 2 3719 2973
0 2975 5 4 1 2974
0 2976 7 1 2 4019 5971
0 2977 5 4 1 2976
0 2978 7 2 2 5895 5897
0 2979 5 1 1 5980
0 2980 7 1 2 3608 5981
0 2981 5 1 1 2980
0 2982 7 1 2 3917 2979
0 2983 5 1 1 2982
0 2984 7 2 2 2981 2983
0 2985 5 1 1 5982
0 2986 7 1 2 3712 2985
0 2987 5 4 1 2986
0 2988 7 1 2 4013 5983
0 2989 5 4 1 2988
0 2990 7 2 2 5889 5891
0 2991 5 1 1 5992
0 2992 7 1 2 3602 5993
0 2993 5 1 1 2992
0 2994 7 1 2 3910 2991
0 2995 5 1 1 2994
0 2996 7 2 2 2993 2995
0 2997 5 1 1 5994
0 2998 7 1 2 3705 2997
0 2999 5 3 1 2998
0 3000 7 1 2 4008 5995
0 3001 5 4 1 3000
0 3002 7 2 2 5883 5885
0 3003 5 1 1 6003
0 3004 7 1 2 3595 6004
0 3005 5 1 1 3004
0 3006 7 1 2 3903 3003
0 3007 5 1 1 3006
0 3008 7 2 2 3005 3007
0 3009 5 1 1 6005
0 3010 7 1 2 3699 3009
0 3011 5 4 1 3010
0 3012 7 1 2 4002 6006
0 3013 5 3 1 3012
0 3014 7 2 2 5877 5879
0 3015 5 1 1 6014
0 3016 7 1 2 3588 6015
0 3017 5 1 1 3016
0 3018 7 1 2 3897 3015
0 3019 5 1 1 3018
0 3020 7 2 2 3017 3019
0 3021 5 1 1 6016
0 3022 7 1 2 3996 6017
0 3023 5 4 1 3022
0 3024 7 2 2 6011 6018
0 3025 7 1 2 3693 3021
0 3026 5 4 1 3025
0 3027 7 2 2 5871 5873
0 3028 5 1 1 6028
0 3029 7 1 2 3582 6029
0 3030 5 1 1 3029
0 3031 7 1 2 3890 3028
0 3032 5 1 1 3031
0 3033 7 2 2 3030 3032
0 3034 5 1 1 6030
0 3035 7 1 2 3686 3034
0 3036 5 4 1 3035
0 3037 7 1 2 3991 6031
0 3038 5 4 1 3037
0 3039 7 2 2 5865 5867
0 3040 5 1 1 6040
0 3041 7 1 2 3576 6041
0 3042 5 1 1 3041
0 3043 7 1 2 3883 3040
0 3044 5 1 1 3043
0 3045 7 2 2 3042 3044
0 3046 5 1 1 6042
0 3047 7 1 2 3680 3046
0 3048 5 4 1 3047
0 3049 7 1 2 3985 6043
0 3050 5 4 1 3049
0 3051 7 2 2 5859 5861
0 3052 5 1 1 6052
0 3053 7 1 2 3569 6053
0 3054 5 1 1 3053
0 3055 7 1 2 3877 3052
0 3056 5 1 1 3055
0 3057 7 2 2 3054 3056
0 3058 5 1 1 6054
0 3059 7 1 2 3673 3058
0 3060 5 3 1 3059
0 3061 7 1 2 3979 6055
0 3062 5 4 1 3061
0 3063 7 2 2 5840 5842
0 3064 5 1 1 6063
0 3065 7 1 2 5853 3064
0 3066 5 1 1 3065
0 3067 7 1 2 5855 6064
0 3068 5 1 1 3067
0 3069 7 2 2 3066 3068
0 3070 5 1 1 6065
0 3071 7 1 2 3974 3070
0 3072 5 3 1 3071
0 3073 7 1 2 3666 6066
0 3074 5 1 1 3073
0 3075 7 2 2 5844 5846
0 3076 5 1 1 6070
0 3077 7 1 2 5848 3076
0 3078 5 1 1 3077
0 3079 7 1 2 5850 6071
0 3080 5 1 1 3079
0 3081 7 2 2 3078 3080
0 3082 5 1 1 6072
0 3083 7 1 2 3660 6073
0 3084 5 1 1 3083
0 3085 7 2 2 3074 3084
0 3086 5 1 1 6074
0 3087 7 1 2 6067 3086
0 3088 5 2 1 3087
0 3089 7 1 2 3767 3859
0 3090 5 1 1 3089
0 3091 7 2 2 5851 3090
0 3092 5 1 1 6078
0 3093 7 1 2 3962 6079
0 3094 5 1 1 3093
0 3095 7 1 2 3968 3082
0 3096 5 2 1 3095
0 3097 7 1 2 3094 6080
0 3098 7 3 2 6068 3097
0 3099 5 1 1 6082
0 3100 7 2 2 6076 3099
0 3101 5 2 1 6085
0 3102 7 1 2 6059 6087
0 3103 5 1 1 3102
0 3104 7 2 2 6056 3103
0 3105 5 2 1 6089
0 3106 7 1 2 6048 6091
0 3107 5 1 1 3106
0 3108 7 2 2 6044 3107
0 3109 5 1 1 6093
0 3110 7 1 2 6036 3109
0 3111 5 2 1 3110
0 3112 7 1 2 6032 6095
0 3113 7 1 2 6024 3112
0 3114 5 1 1 3113
0 3115 7 1 2 6022 3114
0 3116 5 1 1 3115
0 3117 7 1 2 6007 3116
0 3118 5 2 1 3117
0 3119 7 1 2 5999 6097
0 3120 5 1 1 3119
0 3121 7 2 2 5996 3120
0 3122 5 1 1 6099
0 3123 7 2 2 5988 3122
0 3124 5 1 1 6101
0 3125 7 1 2 5984 3124
0 3126 5 2 1 3125
0 3127 7 1 2 5976 6103
0 3128 5 1 1 3127
0 3129 7 2 2 5972 3128
0 3130 5 1 1 6105
0 3131 7 1 2 5965 3130
0 3132 5 1 1 3131
0 3133 7 2 2 5961 3132
0 3134 5 2 1 6107
0 3135 7 1 2 5953 6109
0 3136 5 1 1 3135
0 3137 7 2 2 5950 3136
0 3138 5 2 1 6111
0 3139 7 1 2 5942 6113
0 3140 5 1 1 3139
0 3141 7 2 2 5939 3140
0 3142 5 2 1 6115
0 3143 7 1 2 4041 5931
0 3144 5 4 1 3143
0 3145 7 1 2 6117 6119
0 3146 5 1 1 3145
0 3147 7 3 2 5932 3146
0 3148 5 1 1 6123
0 3149 7 2 2 3654 3092
0 3150 5 1 1 6126
0 3151 7 1 2 6081 6127
0 3152 7 1 2 6069 3151
0 3153 5 1 1 3152
0 3154 7 2 2 6077 3153
0 3155 5 2 1 6128
0 3156 7 1 2 6060 6130
0 3157 5 1 1 3156
0 3158 7 2 2 6057 3157
0 3159 5 1 1 6132
0 3160 7 2 2 6049 3159
0 3161 5 1 1 6134
0 3162 7 2 2 6045 3161
0 3163 5 2 1 6136
0 3164 7 1 2 6037 6138
0 3165 5 1 1 3164
0 3166 7 1 2 6033 3165
0 3167 5 2 1 3166
0 3168 7 1 2 6019 6140
0 3169 5 1 1 3168
0 3170 7 2 2 6025 3169
0 3171 5 1 1 6142
0 3172 7 1 2 6012 3171
0 3173 5 1 1 3172
0 3174 7 2 2 6008 3173
0 3175 5 2 1 6144
0 3176 7 1 2 6000 6146
0 3177 5 1 1 3176
0 3178 7 2 2 5997 3177
0 3179 5 2 1 6148
0 3180 7 1 2 5989 6150
0 3181 5 1 1 3180
0 3182 7 2 2 5985 3181
0 3183 7 1 2 5973 6152
0 3184 5 1 1 3183
0 3185 7 2 2 5966 5977
0 3186 7 1 2 3184 6154
0 3187 5 1 1 3186
0 3188 7 1 2 5962 3187
0 3189 5 2 1 3188
0 3190 7 1 2 5954 6156
0 3191 5 1 1 3190
0 3192 7 2 2 5951 3191
0 3193 5 2 1 6158
0 3194 7 1 2 5943 6160
0 3195 5 1 1 3194
0 3196 7 2 2 5940 3195
0 3197 5 2 1 6162
0 3198 7 1 2 6120 6164
0 3199 5 1 1 3198
0 3200 7 2 2 5933 3199
0 3201 5 2 1 6166
0 3202 7 1 2 3950 5927
0 3203 5 1 1 3202
0 3204 7 2 2 5925 3203
0 3205 5 1 1 6170
0 3206 7 1 2 3853 3205
0 3207 5 2 1 3206
0 3208 7 1 2 3543 6171
0 3209 5 2 1 3208
0 3210 7 2 2 6172 6174
0 3211 5 1 1 6176
0 3212 7 1 2 3647 6177
0 3213 5 1 1 3212
0 3214 7 1 2 3956 3211
0 3215 5 1 1 3214
0 3216 7 2 2 3213 3215
0 3217 5 1 1 6178
0 3218 7 1 2 3756 3217
0 3219 5 3 1 3218
0 3220 7 2 2 4044 6179
0 3221 5 3 1 6183
0 3222 7 2 2 6180 6185
0 3223 5 1 1 6188
0 3224 7 1 2 6168 6189
0 3225 5 2 1 3224
0 3226 7 1 2 3148 6190
0 3227 5 1 1 3226
0 3228 7 1 2 6181 6124
0 3229 5 1 1 3228
0 3230 7 1 2 3957 6175
0 3231 5 1 1 3230
0 3232 7 2 2 6173 3231
0 3233 5 1 1 6192
0 3234 7 2 2 3762 3233
0 3235 5 2 1 6194
0 3236 7 2 2 6186 6196
0 3237 7 1 2 3229 6198
0 3238 7 1 2 3227 3237
0 3239 5 1 1 3238
0 3240 7 1 2 6125 6195
0 3241 7 1 2 6184 3240
0 3242 5 1 1 3241
0 3243 7 1 2 3239 3242
0 3244 5 1 1 3243
0 3245 7 3 2 5934 6121
0 3246 5 2 1 6200
0 3247 7 1 2 6116 6203
0 3248 5 1 1 3247
0 3249 7 1 2 6118 6201
0 3250 5 1 1 3249
0 3251 7 1 2 3248 3250
0 3252 5 1 1 3251
0 3253 7 2 2 4048 6193
0 3254 5 2 1 6205
0 3255 7 3 2 5941 5944
0 3256 5 2 1 6209
0 3257 7 1 2 6112 6212
0 3258 5 1 1 3257
0 3259 7 1 2 6114 6210
0 3260 5 1 1 3259
0 3261 7 1 2 3258 3260
0 3262 5 1 1 3261
0 3263 7 3 2 5952 5955
0 3264 5 2 1 6214
0 3265 7 1 2 6110 6217
0 3266 5 1 1 3265
0 3267 7 1 2 6108 6215
0 3268 5 1 1 3267
0 3269 7 2 2 5963 5967
0 3270 5 2 1 6219
0 3271 7 1 2 6106 6220
0 3272 5 1 1 3271
0 3273 7 1 2 5978 6221
0 3274 5 1 1 3273
0 3275 7 1 2 5974 5979
0 3276 5 2 1 3275
0 3277 7 1 2 6104 6223
0 3278 5 1 1 3277
0 3279 7 1 2 5986 6102
0 3280 5 1 1 3279
0 3281 7 2 2 5987 5990
0 3282 5 2 1 6225
0 3283 7 1 2 6100 6227
0 3284 5 1 1 3283
0 3285 7 3 2 5998 6001
0 3286 5 2 1 6229
0 3287 7 1 2 6009 6232
0 3288 5 1 1 3287
0 3289 7 1 2 6098 6230
0 3290 5 1 1 3289
0 3291 7 2 2 6010 6013
0 3292 5 2 1 6234
0 3293 7 1 2 6026 6236
0 3294 5 1 1 3293
0 3295 7 2 2 6020 6027
0 3296 5 1 1 6238
0 3297 7 1 2 6096 6239
0 3298 5 1 1 3297
0 3299 7 1 2 6034 3298
0 3300 5 1 1 3299
0 3301 7 2 2 6035 6038
0 3302 5 2 1 6240
0 3303 7 1 2 6094 6242
0 3304 5 1 1 3303
0 3305 7 2 2 6046 6050
0 3306 5 2 1 6244
0 3307 7 1 2 6090 6245
0 3308 5 1 1 3307
0 3309 7 3 2 6058 6061
0 3310 5 2 1 6248
0 3311 7 1 2 6088 6249
0 3312 5 1 1 3311
0 3313 7 1 2 6075 3150
0 3314 7 1 2 6083 3313
0 3315 5 2 1 3314
0 3316 7 1 2 6086 6251
0 3317 5 1 1 3316
0 3318 7 1 2 6253 3317
0 3319 7 1 2 3312 3318
0 3320 5 1 1 3319
0 3321 7 1 2 6092 6246
0 3322 5 1 1 3321
0 3323 7 1 2 3320 3322
0 3324 7 1 2 3308 3323
0 3325 5 1 1 3324
0 3326 7 1 2 3304 3325
0 3327 7 1 2 3300 3326
0 3328 7 1 2 3294 3327
0 3329 7 1 2 3290 3328
0 3330 7 1 2 3288 3329
0 3331 7 1 2 3284 3330
0 3332 7 1 2 3280 3331
0 3333 5 1 1 3332
0 3334 7 1 2 3278 3333
0 3335 7 1 2 3274 3334
0 3336 7 1 2 3272 3335
0 3337 7 1 2 3268 3336
0 3338 7 1 2 3266 3337
0 3339 7 1 2 3262 3338
0 3340 7 1 2 6207 3339
0 3341 7 1 2 3252 3340
0 3342 7 1 2 3244 3341
0 3343 5 1 1 3342
0 3344 7 1 2 6169 6187
0 3345 5 1 1 3344
0 3346 7 2 2 6182 3345
0 3347 5 1 1 6255
0 3348 7 1 2 6206 3347
0 3349 5 1 1 3348
0 3350 7 2 2 6208 6256
0 3351 5 1 1 6257
0 3352 7 1 2 3349 3351
0 3353 5 1 1 3352
0 3354 7 1 2 6167 3223
0 3355 5 1 1 3354
0 3356 7 1 2 6161 6211
0 3357 5 1 1 3356
0 3358 7 1 2 6159 6213
0 3359 5 1 1 3358
0 3360 7 1 2 5964 6218
0 3361 5 1 1 3360
0 3362 7 1 2 6157 6216
0 3363 5 1 1 3362
0 3364 7 1 2 5975 6222
0 3365 5 1 1 3364
0 3366 7 1 2 6153 6224
0 3367 5 1 1 3366
0 3368 7 1 2 6149 6226
0 3369 5 1 1 3368
0 3370 7 1 2 6151 6228
0 3371 5 1 1 3370
0 3372 7 1 2 6147 6233
0 3373 5 1 1 3372
0 3374 7 1 2 6145 6231
0 3375 5 1 1 3374
0 3376 7 1 2 6021 6237
0 3377 5 1 1 3376
0 3378 7 1 2 6143 6235
0 3379 5 1 1 3378
0 3380 7 1 2 6141 3296
0 3381 5 1 1 3380
0 3382 7 1 2 6137 6241
0 3383 5 1 1 3382
0 3384 7 1 2 6047 6135
0 3385 5 1 1 3384
0 3386 7 1 2 6133 6247
0 3387 5 1 1 3386
0 3388 7 1 2 6129 6250
0 3389 5 1 1 3388
0 3390 7 1 2 6131 6252
0 3391 5 1 1 3390
0 3392 7 1 2 6254 3391
0 3393 7 1 2 3389 3392
0 3394 5 1 1 3393
0 3395 7 1 2 3387 3394
0 3396 7 1 2 3385 3395
0 3397 5 1 1 3396
0 3398 7 1 2 6139 6243
0 3399 5 1 1 3398
0 3400 7 1 2 3397 3399
0 3401 7 1 2 3383 3400
0 3402 7 1 2 3381 3401
0 3403 7 1 2 3379 3402
0 3404 7 1 2 3377 3403
0 3405 7 1 2 3375 3404
0 3406 7 1 2 3373 3405
0 3407 7 1 2 3371 3406
0 3408 7 1 2 3369 3407
0 3409 5 1 1 3408
0 3410 7 1 2 3367 3409
0 3411 7 1 2 3365 3410
0 3412 7 1 2 3363 3411
0 3413 7 1 2 3361 3412
0 3414 7 1 2 3359 3413
0 3415 7 1 2 3357 3414
0 3416 7 1 2 6197 3415
0 3417 7 1 2 6204 6163
0 3418 5 1 1 3417
0 3419 7 1 2 6202 6165
0 3420 5 1 1 3419
0 3421 7 1 2 3418 3420
0 3422 7 1 2 3416 3421
0 3423 7 1 2 6191 3422
0 3424 7 1 2 3355 3423
0 3425 7 1 2 3353 3424
0 3426 5 1 1 3425
0 3427 7 1 2 3343 3426
0 3428 5 1 1 3427
0 3429 7 1 2 2809 3428
0 3430 5 1 1 3429
0 3431 7 1 2 6062 6084
0 3432 7 1 2 6051 3431
0 3433 7 1 2 6039 3432
0 3434 7 1 2 6023 3433
0 3435 7 1 2 6002 3434
0 3436 7 1 2 5991 3435
0 3437 7 1 2 6155 3436
0 3438 7 1 2 5956 3437
0 3439 7 1 2 5945 3438
0 3440 7 1 2 6122 3439
0 3441 7 1 2 6199 3440
0 3442 7 1 2 6258 3441
0 3443 7 1 2 5838 3442
0 3444 5 1 1 3443
0 3445 7 1 2 3430 3444
3 9999 5 0 1 3445
