1 0 0 1 0
1 1 0 2 0
2 26 1 1
2 27 1 1
1 2 0 2 0
2 350 1 2
2 351 1 2
1 3 0 2 0
2 352 1 3
2 353 1 3
1 4 0 4 0
2 354 1 4
2 355 1 4
2 356 1 4
2 357 1 4
1 5 0 8 0
2 358 1 5
2 359 1 5
2 360 1 5
2 361 1 5
2 362 1 5
2 363 1 5
2 364 1 5
2 365 1 5
1 6 0 8 0
2 366 1 6
2 367 1 6
2 368 1 6
2 369 1 6
2 370 1 6
2 371 1 6
2 372 1 6
2 373 1 6
1 7 0 6 0
2 374 1 7
2 375 1 7
2 376 1 7
2 377 1 7
2 378 1 7
2 379 1 7
1 8 0 2 0
2 380 1 8
2 381 1 8
1 9 0 2 0
2 382 1 9
2 383 1 9
1 10 0 2 0
2 384 1 10
2 385 1 10
1 11 0 2 0
2 386 1 11
2 387 1 11
1 12 0 2 0
2 388 1 12
2 389 1 12
1 13 0 2 0
2 390 1 13
2 391 1 13
1 14 0 2 0
2 392 1 14
2 393 1 14
1 15 0 2 0
2 394 1 15
2 395 1 15
1 16 0 2 0
2 396 1 16
2 397 1 16
1 17 0 0 0
1 18 0 0 0
1 19 0 0 0
1 20 0 0 0
1 21 0 2 0
2 398 1 21
2 399 1 21
1 22 0 2 0
2 400 1 22
2 401 1 22
1 23 0 2 0
2 402 1 23
2 403 1 23
1 24 0 2 0
2 404 1 24
2 405 1 24
1 25 0 4 0
2 406 1 25
2 407 1 25
2 408 1 25
2 409 1 25
2 410 1 31
2 411 1 31
2 412 1 31
2 413 1 31
2 414 1 31
2 415 1 32
2 416 1 32
2 417 1 32
2 418 1 32
2 419 1 32
2 420 1 32
2 421 1 33
2 422 1 33
2 423 1 33
2 424 1 33
2 425 1 33
2 426 1 33
2 427 1 34
2 428 1 34
2 429 1 34
2 430 1 34
2 431 1 34
2 432 1 48
2 433 1 48
2 434 1 48
2 435 1 49
2 436 1 49
2 437 1 49
2 438 1 50
2 439 1 50
2 440 1 51
2 441 1 51
2 442 1 51
2 443 1 51
2 444 1 51
2 445 1 52
2 446 1 52
2 447 1 53
2 448 1 53
2 449 1 60
2 450 1 60
2 451 1 62
2 452 1 62
2 453 1 62
2 454 1 63
2 455 1 63
2 456 1 65
2 457 1 65
2 458 1 68
2 459 1 68
2 460 1 73
2 461 1 73
2 462 1 75
2 463 1 75
2 464 1 77
2 465 1 77
2 466 1 85
2 467 1 85
2 468 1 85
2 469 1 85
2 470 1 85
2 471 1 86
2 472 1 86
2 473 1 86
2 474 1 88
2 475 1 88
2 476 1 88
2 477 1 92
2 478 1 92
2 479 1 92
2 480 1 92
2 481 1 95
2 482 1 95
2 483 1 96
2 484 1 96
2 485 1 101
2 486 1 101
2 487 1 103
2 488 1 103
2 489 1 105
2 490 1 105
2 491 1 105
2 492 1 105
2 493 1 105
2 494 1 105
2 495 1 113
2 496 1 113
2 497 1 113
2 498 1 113
2 499 1 113
2 500 1 113
2 501 1 114
2 502 1 114
2 503 1 114
2 504 1 119
2 505 1 119
2 506 1 121
2 507 1 121
2 508 1 130
2 509 1 130
2 510 1 131
2 511 1 131
2 512 1 131
2 513 1 131
2 514 1 132
2 515 1 132
2 516 1 133
2 517 1 133
2 518 1 133
2 519 1 133
2 520 1 134
2 521 1 134
2 522 1 134
2 523 1 134
2 524 1 145
2 525 1 145
2 526 1 149
2 527 1 149
2 528 1 157
2 529 1 157
2 530 1 157
2 531 1 158
2 532 1 158
2 533 1 170
2 534 1 170
2 535 1 170
2 536 1 171
2 537 1 171
2 538 1 171
2 539 1 171
2 540 1 172
2 541 1 172
2 542 1 172
2 543 1 173
2 544 1 173
2 545 1 173
2 546 1 173
2 547 1 174
2 548 1 174
2 549 1 174
2 550 1 205
2 551 1 205
2 552 1 224
2 553 1 224
2 554 1 228
2 555 1 228
2 556 1 232
2 557 1 232
2 558 1 243
2 559 1 243
2 560 1 244
2 561 1 244
2 562 1 253
2 563 1 253
2 564 1 255
2 565 1 255
2 566 1 265
2 567 1 265
2 568 1 300
2 569 1 300
2 570 1 300
0 28 5 1 1 26
0 29 5 1 1 350
0 30 5 1 1 352
0 31 5 5 1 354
0 32 5 6 1 358
0 33 5 6 1 366
0 34 5 5 1 374
0 35 5 1 1 380
0 36 5 1 1 382
0 37 5 1 1 384
0 38 5 1 1 386
0 39 5 1 1 388
0 40 5 1 1 390
0 41 5 1 1 392
0 42 5 1 1 394
0 43 5 1 1 396
0 44 5 1 1 398
0 45 5 1 1 400
0 46 5 1 1 402
0 47 5 1 1 404
0 48 5 3 1 406
0 49 7 3 2 39 399
0 50 5 2 1 435
0 51 7 5 2 389 44
0 52 5 2 1 440
0 53 7 2 2 438 445
0 54 7 1 2 381 397
0 55 5 1 1 54
0 56 7 1 2 35 43
0 57 5 1 1 56
0 58 7 1 2 0 57
0 59 5 1 1 58
0 60 7 2 2 55 59
0 61 5 1 1 449
0 62 7 3 2 353 387
0 63 5 2 1 451
0 64 7 1 2 351 385
0 65 5 2 1 64
0 66 7 1 2 27 383
0 67 5 1 1 66
0 68 7 2 2 456 67
0 69 7 1 2 454 458
0 70 7 1 2 450 69
0 71 5 1 1 70
0 72 7 1 2 30 38
0 73 5 2 1 72
0 74 7 1 2 29 37
0 75 5 2 1 74
0 76 7 1 2 28 36
0 77 5 2 1 76
0 78 7 1 2 462 464
0 79 5 1 1 78
0 80 7 1 2 455 457
0 81 7 1 2 79 80
0 82 5 1 1 81
0 83 7 1 2 460 82
0 84 7 1 2 71 83
0 85 5 5 1 84
0 86 7 3 2 410 415
0 87 7 1 2 421 427
0 88 7 3 2 432 87
0 89 7 1 2 471 474
0 90 7 1 2 466 89
0 91 5 1 1 90
0 92 7 4 2 355 452
0 93 5 1 1 477
0 94 7 1 2 367 375
0 95 7 2 2 407 94
0 96 7 2 2 359 481
0 97 7 1 2 478 483
0 98 5 1 1 97
0 99 7 1 2 91 98
0 100 5 1 1 99
0 101 7 2 2 395 47
0 102 5 1 1 485
0 103 7 2 2 42 405
0 104 5 1 1 487
0 105 7 6 2 102 104
0 106 7 1 2 100 489
0 107 5 1 1 106
0 108 7 1 2 408 486
0 109 5 1 1 108
0 110 7 1 2 433 488
0 111 5 1 1 110
0 112 7 1 2 109 111
0 113 5 6 1 112
0 114 7 3 2 422 376
0 115 5 1 1 501
0 116 7 1 2 472 502
0 117 7 1 2 467 116
0 118 5 1 1 117
0 119 7 2 2 368 428
0 120 5 1 1 504
0 121 7 2 2 360 505
0 122 7 1 2 479 506
0 123 5 1 1 122
0 124 7 1 2 118 123
0 125 5 1 1 124
0 126 7 1 2 495 125
0 127 5 1 1 126
0 128 7 1 2 107 127
0 129 5 1 1 128
0 130 7 2 2 41 403
0 131 5 4 1 508
0 132 7 2 2 393 46
0 133 5 4 1 514
0 134 7 4 2 510 516
0 135 5 1 1 520
0 136 7 1 2 129 521
0 137 5 1 1 136
0 138 7 1 2 429 517
0 139 5 1 1 138
0 140 7 1 2 377 511
0 141 5 1 1 140
0 142 7 1 2 139 141
0 143 7 1 2 496 142
0 144 5 1 1 143
0 145 7 2 2 378 409
0 146 5 1 1 524
0 147 7 1 2 512 146
0 148 5 1 1 147
0 149 7 2 2 430 434
0 150 5 1 1 526
0 151 7 1 2 518 150
0 152 5 1 1 151
0 153 7 1 2 490 152
0 154 7 1 2 148 153
0 155 5 1 1 154
0 156 7 1 2 144 155
0 157 5 3 1 156
0 158 7 2 2 361 423
0 159 7 1 2 480 531
0 160 5 1 1 159
0 161 7 1 2 369 473
0 162 7 1 2 468 161
0 163 5 1 1 162
0 164 7 1 2 160 163
0 165 5 1 1 164
0 166 7 1 2 528 165
0 167 5 1 1 166
0 168 7 1 2 137 167
0 169 5 1 1 168
0 170 7 3 2 391 45
0 171 5 4 1 533
0 172 7 3 2 40 401
0 173 5 4 1 540
0 174 7 3 2 536 543
0 175 5 1 1 547
0 176 7 1 2 169 548
0 177 5 1 1 176
0 178 7 1 2 482 534
0 179 5 1 1 178
0 180 7 1 2 475 541
0 181 5 1 1 180
0 182 7 1 2 179 181
0 183 5 1 1 182
0 184 7 1 2 491 183
0 185 5 1 1 184
0 186 7 1 2 120 544
0 187 5 1 1 186
0 188 7 1 2 115 537
0 189 5 1 1 188
0 190 7 1 2 187 189
0 191 7 1 2 497 190
0 192 5 1 1 191
0 193 7 1 2 185 192
0 194 5 1 1 193
0 195 7 1 2 522 194
0 196 5 1 1 195
0 197 7 1 2 424 538
0 198 5 1 1 197
0 199 7 1 2 370 545
0 200 5 1 1 199
0 201 7 1 2 198 200
0 202 7 1 2 529 201
0 203 5 1 1 202
0 204 7 1 2 196 203
0 205 5 2 1 204
0 206 7 1 2 416 93
0 207 5 1 1 206
0 208 7 1 2 411 469
0 209 5 1 1 208
0 210 7 1 2 362 209
0 211 5 1 1 210
0 212 7 1 2 207 211
0 213 7 1 2 550 212
0 214 5 1 1 213
0 215 7 1 2 177 214
0 216 5 1 1 215
0 217 7 1 2 447 216
0 218 5 1 1 217
0 219 7 1 2 412 441
0 220 5 1 1 219
0 221 7 1 2 356 448
0 222 5 1 1 221
0 223 7 1 2 220 222
0 224 5 2 1 223
0 225 7 1 2 363 175
0 226 5 1 1 225
0 227 7 1 2 417 539
0 228 5 2 1 227
0 229 7 1 2 226 554
0 230 7 1 2 552 229
0 231 5 1 1 230
0 232 7 2 2 413 436
0 233 7 1 2 364 535
0 234 7 1 2 556 233
0 235 5 1 1 234
0 236 7 1 2 231 235
0 237 5 1 1 236
0 238 7 1 2 379 498
0 239 5 1 1 238
0 240 7 1 2 492 527
0 241 5 1 1 240
0 242 7 1 2 239 241
0 243 5 2 1 242
0 244 7 2 2 425 509
0 245 5 1 1 560
0 246 7 1 2 558 561
0 247 5 1 1 246
0 248 7 1 2 431 499
0 249 5 1 1 248
0 250 7 1 2 493 525
0 251 5 1 1 250
0 252 7 1 2 249 251
0 253 5 2 1 252
0 254 7 1 2 426 519
0 255 5 2 1 254
0 256 7 1 2 371 135
0 257 5 1 1 256
0 258 7 1 2 564 257
0 259 7 1 2 562 258
0 260 5 1 1 259
0 261 7 1 2 247 260
0 262 5 1 1 261
0 263 7 1 2 237 262
0 264 5 1 1 263
0 265 7 2 2 418 542
0 266 5 1 1 566
0 267 7 1 2 553 567
0 268 5 1 1 267
0 269 7 1 2 546 555
0 270 5 1 1 269
0 271 7 1 2 557 266
0 272 7 1 2 270 271
0 273 5 1 1 272
0 274 7 1 2 268 273
0 275 5 1 1 274
0 276 7 1 2 372 515
0 277 7 1 2 563 276
0 278 5 1 1 277
0 279 7 1 2 513 565
0 280 5 1 1 279
0 281 7 1 2 245 280
0 282 7 1 2 559 281
0 283 5 1 1 282
0 284 7 1 2 278 283
0 285 5 1 1 284
0 286 7 1 2 275 285
0 287 5 1 1 286
0 288 7 1 2 264 287
0 289 5 1 1 288
0 290 7 1 2 465 61
0 291 5 1 1 290
0 292 7 1 2 459 291
0 293 5 1 1 292
0 294 7 1 2 461 463
0 295 7 1 2 293 294
0 296 7 1 2 289 295
0 297 5 1 1 296
0 298 7 1 2 442 532
0 299 5 1 1 298
0 300 7 3 2 419 437
0 301 7 1 2 373 568
0 302 5 1 1 301
0 303 7 1 2 299 302
0 304 5 1 1 303
0 305 7 1 2 530 304
0 306 5 1 1 305
0 307 7 1 2 443 484
0 308 5 1 1 307
0 309 7 1 2 476 569
0 310 5 1 1 309
0 311 7 1 2 308 310
0 312 5 1 1 311
0 313 7 1 2 494 312
0 314 5 1 1 313
0 315 7 1 2 503 570
0 316 5 1 1 315
0 317 7 1 2 444 507
0 318 5 1 1 317
0 319 7 1 2 316 318
0 320 5 1 1 319
0 321 7 1 2 500 320
0 322 5 1 1 321
0 323 7 1 2 314 322
0 324 5 1 1 323
0 325 7 1 2 523 324
0 326 5 1 1 325
0 327 7 1 2 306 326
0 328 5 1 1 327
0 329 7 1 2 549 328
0 330 5 1 1 329
0 331 7 1 2 420 446
0 332 5 1 1 331
0 333 7 1 2 365 439
0 334 5 1 1 333
0 335 7 1 2 332 334
0 336 7 1 2 551 335
0 337 5 1 1 336
0 338 7 1 2 330 337
0 339 5 1 1 338
0 340 7 1 2 357 470
0 341 5 1 1 340
0 342 7 1 2 414 453
0 343 5 1 1 342
0 344 7 1 2 341 343
0 345 5 1 1 344
0 346 7 1 2 339 345
0 347 5 1 1 346
0 348 7 1 2 297 347
0 349 7 1 2 218 348
3 799 5 0 1 349
