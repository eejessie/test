1 0 0 8 0
2 32 1 0
2 1937 1 0
2 1938 1 0
2 1939 1 0
2 1940 1 0
2 1941 1 0
2 1942 1 0
2 1943 1 0
1 1 0 8 0
2 1944 1 1
2 1945 1 1
2 1946 1 1
2 1947 1 1
2 1948 1 1
2 1949 1 1
2 1950 1 1
2 1951 1 1
1 2 0 8 0
2 1952 1 2
2 1953 1 2
2 1954 1 2
2 1955 1 2
2 1956 1 2
2 1957 1 2
2 1958 1 2
2 1959 1 2
1 3 0 9 0
2 1960 1 3
2 1961 1 3
2 1962 1 3
2 1963 1 3
2 1964 1 3
2 1965 1 3
2 1966 1 3
2 1967 1 3
2 1968 1 3
1 4 0 8 0
2 1969 1 4
2 1970 1 4
2 1971 1 4
2 1972 1 4
2 1973 1 4
2 1974 1 4
2 1975 1 4
2 1976 1 4
1 5 0 9 0
2 1977 1 5
2 1978 1 5
2 1979 1 5
2 1980 1 5
2 1981 1 5
2 1982 1 5
2 1983 1 5
2 1984 1 5
2 1985 1 5
1 6 0 8 0
2 1986 1 6
2 1987 1 6
2 1988 1 6
2 1989 1 6
2 1990 1 6
2 1991 1 6
2 1992 1 6
2 1993 1 6
1 7 0 8 0
2 1994 1 7
2 1995 1 7
2 1996 1 7
2 1997 1 7
2 1998 1 7
2 1999 1 7
2 2000 1 7
2 2001 1 7
1 8 0 8 0
2 2002 1 8
2 2003 1 8
2 2004 1 8
2 2005 1 8
2 2006 1 8
2 2007 1 8
2 2008 1 8
2 2009 1 8
1 9 0 8 0
2 2010 1 9
2 2011 1 9
2 2012 1 9
2 2013 1 9
2 2014 1 9
2 2015 1 9
2 2016 1 9
2 2017 1 9
1 10 0 9 0
2 2018 1 10
2 2019 1 10
2 2020 1 10
2 2021 1 10
2 2022 1 10
2 2023 1 10
2 2024 1 10
2 2025 1 10
2 2026 1 10
1 11 0 8 0
2 2027 1 11
2 2028 1 11
2 2029 1 11
2 2030 1 11
2 2031 1 11
2 2032 1 11
2 2033 1 11
2 2034 1 11
1 12 0 8 0
2 2035 1 12
2 2036 1 12
2 2037 1 12
2 2038 1 12
2 2039 1 12
2 2040 1 12
2 2041 1 12
2 2042 1 12
1 13 0 8 0
2 2043 1 13
2 2044 1 13
2 2045 1 13
2 2046 1 13
2 2047 1 13
2 2048 1 13
2 2049 1 13
2 2050 1 13
1 14 0 8 0
2 2051 1 14
2 2052 1 14
2 2053 1 14
2 2054 1 14
2 2055 1 14
2 2056 1 14
2 2057 1 14
2 2058 1 14
1 15 0 8 0
2 2059 1 15
2 2060 1 15
2 2061 1 15
2 2062 1 15
2 2063 1 15
2 2064 1 15
2 2065 1 15
2 2066 1 15
1 16 0 2 0
2 2067 1 16
2 2068 1 16
1 17 0 2 0
2 2069 1 17
2 2070 1 17
1 18 0 2 0
2 2071 1 18
2 2072 1 18
1 19 0 2 0
2 2073 1 19
2 2074 1 19
1 20 0 2 0
2 2075 1 20
2 2076 1 20
1 21 0 2 0
2 2077 1 21
2 2078 1 21
1 22 0 2 0
2 2079 1 22
2 2080 1 22
1 23 0 2 0
2 2081 1 23
2 2082 1 23
1 24 0 2 0
2 2083 1 24
2 2084 1 24
1 25 0 2 0
2 2085 1 25
2 2086 1 25
1 26 0 2 0
2 2087 1 26
2 2088 1 26
1 27 0 2 0
2 2089 1 27
2 2090 1 27
1 28 0 2 0
2 2091 1 28
2 2092 1 28
1 29 0 2 0
2 2093 1 29
2 2094 1 29
1 30 0 2 0
2 2095 1 30
2 2096 1 30
1 31 0 2 0
2 2097 1 31
2 2098 1 31
2 2099 1 33
2 2100 1 33
2 2101 1 33
2 2102 1 49
2 2103 1 49
2 2104 1 51
2 2105 1 51
2 2106 1 52
2 2107 1 52
2 2108 1 53
2 2109 1 53
2 2110 1 55
2 2111 1 55
2 2112 1 58
2 2113 1 58
2 2114 1 61
2 2115 1 61
2 2116 1 64
2 2117 1 64
2 2118 1 65
2 2119 1 65
2 2120 1 67
2 2121 1 67
2 2122 1 69
2 2123 1 69
2 2124 1 75
2 2125 1 75
2 2126 1 78
2 2127 1 78
2 2128 1 78
2 2129 1 82
2 2130 1 82
2 2131 1 83
2 2132 1 83
2 2133 1 85
2 2134 1 85
2 2135 1 88
2 2136 1 88
2 2137 1 89
2 2138 1 89
2 2139 1 93
2 2140 1 93
2 2141 1 96
2 2142 1 96
2 2143 1 97
2 2144 1 97
2 2145 1 101
2 2146 1 101
2 2147 1 104
2 2148 1 104
2 2149 1 105
2 2150 1 105
2 2151 1 109
2 2152 1 109
2 2153 1 112
2 2154 1 112
2 2155 1 113
2 2156 1 113
2 2157 1 115
2 2158 1 115
2 2159 1 118
2 2160 1 118
2 2161 1 119
2 2162 1 119
2 2163 1 123
2 2164 1 123
2 2165 1 126
2 2166 1 126
2 2167 1 127
2 2168 1 127
2 2169 1 131
2 2170 1 131
2 2171 1 134
2 2172 1 134
2 2173 1 135
2 2174 1 135
2 2175 1 139
2 2176 1 139
2 2177 1 142
2 2178 1 142
2 2179 1 143
2 2180 1 143
2 2181 1 147
2 2182 1 147
2 2183 1 150
2 2184 1 150
2 2185 1 151
2 2186 1 151
2 2187 1 155
2 2188 1 155
2 2189 1 158
2 2190 1 158
2 2191 1 159
2 2192 1 159
2 2193 1 163
2 2194 1 163
2 2195 1 166
2 2196 1 166
2 2197 1 167
2 2198 1 167
2 2199 1 171
2 2200 1 171
2 2201 1 174
2 2202 1 174
2 2203 1 175
2 2204 1 175
2 2205 1 177
2 2206 1 177
2 2207 1 179
2 2208 1 179
2 2209 1 181
2 2210 1 181
2 2211 1 182
2 2212 1 182
2 2213 1 183
2 2214 1 183
2 2215 1 184
2 2216 1 184
2 2217 1 186
2 2218 1 186
2 2219 1 187
2 2220 1 187
2 2221 1 191
2 2222 1 191
2 2223 1 194
2 2224 1 194
2 2225 1 195
2 2226 1 195
2 2227 1 199
2 2228 1 199
2 2229 1 202
2 2230 1 202
2 2231 1 203
2 2232 1 203
2 2233 1 207
2 2234 1 207
2 2235 1 210
2 2236 1 210
2 2237 1 211
2 2238 1 211
2 2239 1 215
2 2240 1 215
2 2241 1 218
2 2242 1 218
2 2243 1 219
2 2244 1 219
2 2245 1 223
2 2246 1 223
2 2247 1 226
2 2248 1 226
2 2249 1 227
2 2250 1 227
2 2251 1 231
2 2252 1 231
2 2253 1 234
2 2254 1 234
2 2255 1 235
2 2256 1 235
2 2257 1 239
2 2258 1 239
2 2259 1 242
2 2260 1 242
2 2261 1 243
2 2262 1 243
2 2263 1 245
2 2264 1 245
2 2265 1 248
2 2266 1 248
2 2267 1 251
2 2268 1 251
2 2269 1 255
2 2270 1 255
2 2271 1 258
2 2272 1 258
2 2273 1 259
2 2274 1 259
2 2275 1 263
2 2276 1 263
2 2277 1 266
2 2278 1 266
2 2279 1 267
2 2280 1 267
2 2281 1 269
2 2282 1 269
2 2283 1 272
2 2284 1 272
2 2285 1 273
2 2286 1 273
2 2287 1 275
2 2288 1 275
2 2289 1 281
2 2290 1 281
2 2291 1 284
2 2292 1 284
2 2293 1 287
2 2294 1 287
2 2295 1 290
2 2296 1 290
2 2297 1 293
2 2298 1 293
2 2299 1 297
2 2300 1 297
2 2301 1 300
2 2302 1 300
2 2303 1 301
2 2304 1 301
2 2305 1 305
2 2306 1 305
2 2307 1 308
2 2308 1 308
2 2309 1 309
2 2310 1 309
2 2311 1 311
2 2312 1 311
2 2313 1 314
2 2314 1 314
2 2315 1 317
2 2316 1 317
2 2317 1 321
2 2318 1 321
2 2319 1 324
2 2320 1 324
2 2321 1 325
2 2322 1 325
2 2323 1 329
2 2324 1 329
2 2325 1 332
2 2326 1 332
2 2327 1 333
2 2328 1 333
2 2329 1 337
2 2330 1 337
2 2331 1 340
2 2332 1 340
2 2333 1 341
2 2334 1 341
2 2335 1 345
2 2336 1 345
2 2337 1 348
2 2338 1 348
2 2339 1 349
2 2340 1 349
2 2341 1 353
2 2342 1 353
2 2343 1 356
2 2344 1 356
2 2345 1 357
2 2346 1 357
2 2347 1 359
2 2348 1 359
2 2349 1 362
2 2350 1 362
2 2351 1 363
2 2352 1 363
2 2353 1 367
2 2354 1 367
2 2355 1 370
2 2356 1 370
2 2357 1 371
2 2358 1 371
2 2359 1 373
2 2360 1 373
2 2361 1 375
2 2362 1 375
2 2363 1 378
2 2364 1 378
2 2365 1 379
2 2366 1 379
2 2367 1 381
2 2368 1 381
2 2369 1 383
2 2370 1 383
2 2371 1 385
2 2372 1 385
2 2373 1 387
2 2374 1 387
2 2375 1 388
2 2376 1 388
2 2377 1 389
2 2378 1 389
2 2379 1 390
2 2380 1 390
2 2381 1 391
2 2382 1 391
2 2383 1 392
2 2384 1 392
2 2385 1 393
2 2386 1 393
2 2387 1 394
2 2388 1 394
2 2389 1 396
2 2390 1 396
2 2391 1 399
2 2392 1 399
2 2393 1 403
2 2394 1 403
2 2395 1 406
2 2396 1 406
2 2397 1 409
2 2398 1 409
2 2399 1 413
2 2400 1 413
2 2401 1 416
2 2402 1 416
2 2403 1 417
2 2404 1 417
2 2405 1 420
2 2406 1 420
2 2407 1 421
2 2408 1 421
2 2409 1 425
2 2410 1 425
2 2411 1 428
2 2412 1 428
2 2413 1 429
2 2414 1 429
2 2415 1 433
2 2416 1 433
2 2417 1 436
2 2418 1 436
2 2419 1 437
2 2420 1 437
2 2421 1 441
2 2422 1 441
2 2423 1 444
2 2424 1 444
2 2425 1 447
2 2426 1 447
2 2427 1 451
2 2428 1 451
2 2429 1 454
2 2430 1 454
2 2431 1 457
2 2432 1 457
2 2433 1 461
2 2434 1 461
2 2435 1 464
2 2436 1 464
2 2437 1 465
2 2438 1 465
2 2439 1 467
2 2440 1 467
2 2441 1 470
2 2442 1 470
2 2443 1 471
2 2444 1 471
2 2445 1 475
2 2446 1 475
2 2447 1 478
2 2448 1 478
2 2449 1 479
2 2450 1 479
2 2451 1 483
2 2452 1 483
2 2453 1 486
2 2454 1 486
2 2455 1 487
2 2456 1 487
2 2457 1 491
2 2458 1 491
2 2459 1 494
2 2460 1 494
2 2461 1 495
2 2462 1 495
2 2463 1 499
2 2464 1 499
2 2465 1 502
2 2466 1 502
2 2467 1 503
2 2468 1 503
2 2469 1 507
2 2470 1 507
2 2471 1 510
2 2472 1 510
2 2473 1 511
2 2474 1 511
2 2475 1 513
2 2476 1 513
2 2477 1 519
2 2478 1 519
2 2479 1 522
2 2480 1 522
2 2481 1 525
2 2482 1 525
2 2483 1 528
2 2484 1 528
2 2485 1 531
2 2486 1 531
2 2487 1 535
2 2488 1 535
2 2489 1 538
2 2490 1 538
2 2491 1 539
2 2492 1 539
2 2493 1 543
2 2494 1 543
2 2495 1 546
2 2496 1 546
2 2497 1 547
2 2498 1 547
2 2499 1 551
2 2500 1 551
2 2501 1 554
2 2502 1 554
2 2503 1 555
2 2504 1 555
2 2505 1 559
2 2506 1 559
2 2507 1 562
2 2508 1 562
2 2509 1 563
2 2510 1 563
2 2511 1 567
2 2512 1 567
2 2513 1 570
2 2514 1 570
2 2515 1 571
2 2516 1 571
2 2517 1 575
2 2518 1 575
2 2519 1 578
2 2520 1 578
2 2521 1 579
2 2522 1 579
2 2523 1 583
2 2524 1 583
2 2525 1 586
2 2526 1 586
2 2527 1 587
2 2528 1 587
2 2529 1 589
2 2530 1 589
2 2531 1 592
2 2532 1 592
2 2533 1 595
2 2534 1 595
2 2535 1 599
2 2536 1 599
2 2537 1 602
2 2538 1 602
2 2539 1 603
2 2540 1 603
2 2541 1 607
2 2542 1 607
2 2543 1 610
2 2544 1 610
2 2545 1 611
2 2546 1 611
2 2547 1 615
2 2548 1 615
2 2549 1 618
2 2550 1 618
2 2551 1 619
2 2552 1 619
2 2553 1 623
2 2554 1 623
2 2555 1 626
2 2556 1 626
2 2557 1 627
2 2558 1 627
2 2559 1 633
2 2560 1 633
2 2561 1 636
2 2562 1 636
2 2563 1 637
2 2564 1 637
2 2565 1 641
2 2566 1 641
2 2567 1 644
2 2568 1 644
2 2569 1 645
2 2570 1 645
2 2571 1 649
2 2572 1 649
2 2573 1 652
2 2574 1 652
2 2575 1 653
2 2576 1 653
2 2577 1 657
2 2578 1 657
2 2579 1 660
2 2580 1 660
2 2581 1 661
2 2582 1 661
2 2583 1 663
2 2584 1 663
2 2585 1 666
2 2586 1 666
2 2587 1 669
2 2588 1 669
2 2589 1 673
2 2590 1 673
2 2591 1 676
2 2592 1 676
2 2593 1 677
2 2594 1 677
2 2595 1 681
2 2596 1 681
2 2597 1 684
2 2598 1 684
2 2599 1 687
2 2600 1 687
2 2601 1 689
2 2602 1 689
2 2603 1 691
2 2604 1 691
2 2605 1 693
2 2606 1 693
2 2607 1 695
2 2608 1 695
2 2609 1 697
2 2610 1 697
2 2611 1 699
2 2612 1 699
2 2613 1 700
2 2614 1 700
2 2615 1 701
2 2616 1 701
2 2617 1 701
2 2618 1 704
2 2619 1 704
2 2620 1 707
2 2621 1 707
2 2622 1 715
2 2623 1 715
2 2624 1 718
2 2625 1 718
2 2626 1 719
2 2627 1 719
2 2628 1 723
2 2629 1 723
2 2630 1 726
2 2631 1 726
2 2632 1 729
2 2633 1 729
2 2634 1 731
2 2635 1 731
2 2636 1 733
2 2637 1 733
2 2638 1 735
2 2639 1 735
2 2640 1 736
2 2641 1 736
2 2642 1 738
2 2643 1 738
2 2644 1 739
2 2645 1 739
2 2646 1 743
2 2647 1 743
2 2648 1 746
2 2649 1 746
2 2650 1 747
2 2651 1 747
2 2652 1 751
2 2653 1 751
2 2654 1 754
2 2655 1 754
2 2656 1 755
2 2657 1 755
2 2658 1 759
2 2659 1 759
2 2660 1 762
2 2661 1 762
2 2662 1 763
2 2663 1 763
2 2664 1 767
2 2665 1 767
2 2666 1 770
2 2667 1 770
2 2668 1 771
2 2669 1 771
2 2670 1 775
2 2671 1 775
2 2672 1 778
2 2673 1 778
2 2674 1 779
2 2675 1 779
2 2676 1 783
2 2677 1 783
2 2678 1 786
2 2679 1 786
2 2680 1 787
2 2681 1 787
2 2682 1 791
2 2683 1 791
2 2684 1 794
2 2685 1 794
2 2686 1 795
2 2687 1 795
2 2688 1 799
2 2689 1 799
2 2690 1 802
2 2691 1 802
2 2692 1 803
2 2693 1 803
2 2694 1 807
2 2695 1 807
2 2696 1 810
2 2697 1 810
2 2698 1 811
2 2699 1 811
2 2700 1 815
2 2701 1 815
2 2702 1 818
2 2703 1 818
2 2704 1 819
2 2705 1 819
2 2706 1 823
2 2707 1 823
2 2708 1 826
2 2709 1 826
2 2710 1 827
2 2711 1 827
2 2712 1 831
2 2713 1 831
2 2714 1 834
2 2715 1 834
2 2716 1 835
2 2717 1 835
2 2718 1 835
2 2719 1 835
2 2720 1 836
2 2721 1 836
2 2722 1 836
2 2723 1 839
2 2724 1 839
2 2725 1 839
2 2726 1 839
2 2727 1 840
2 2728 1 840
2 2729 1 840
2 2730 1 842
2 2731 1 842
2 2732 1 842
2 2733 1 844
2 2734 1 844
2 2735 1 844
2 2736 1 847
2 2737 1 847
2 2738 1 847
2 2739 1 847
2 2740 1 848
2 2741 1 848
2 2742 1 848
2 2743 1 850
2 2744 1 850
2 2745 1 850
2 2746 1 852
2 2747 1 852
2 2748 1 852
2 2749 1 855
2 2750 1 855
2 2751 1 855
2 2752 1 855
2 2753 1 856
2 2754 1 856
2 2755 1 856
2 2756 1 858
2 2757 1 858
2 2758 1 858
2 2759 1 860
2 2760 1 860
2 2761 1 860
2 2762 1 863
2 2763 1 863
2 2764 1 863
2 2765 1 863
2 2766 1 864
2 2767 1 864
2 2768 1 864
2 2769 1 866
2 2770 1 866
2 2771 1 866
2 2772 1 868
2 2773 1 868
2 2774 1 868
2 2775 1 871
2 2776 1 871
2 2777 1 871
2 2778 1 871
2 2779 1 872
2 2780 1 872
2 2781 1 872
2 2782 1 874
2 2783 1 874
2 2784 1 874
2 2785 1 876
2 2786 1 876
2 2787 1 876
2 2788 1 879
2 2789 1 879
2 2790 1 879
2 2791 1 879
2 2792 1 880
2 2793 1 880
2 2794 1 880
2 2795 1 882
2 2796 1 882
2 2797 1 882
2 2798 1 884
2 2799 1 884
2 2800 1 884
2 2801 1 887
2 2802 1 887
2 2803 1 887
2 2804 1 887
2 2805 1 888
2 2806 1 888
2 2807 1 888
2 2808 1 890
2 2809 1 890
2 2810 1 890
2 2811 1 892
2 2812 1 892
2 2813 1 892
2 2814 1 895
2 2815 1 895
2 2816 1 895
2 2817 1 895
2 2818 1 896
2 2819 1 896
2 2820 1 896
2 2821 1 898
2 2822 1 898
2 2823 1 898
2 2824 1 900
2 2825 1 900
2 2826 1 900
2 2827 1 903
2 2828 1 903
2 2829 1 904
2 2830 1 904
2 2831 1 904
2 2832 1 906
2 2833 1 906
2 2834 1 906
2 2835 1 908
2 2836 1 908
2 2837 1 908
2 2838 1 911
2 2839 1 911
2 2840 1 911
2 2841 1 911
2 2842 1 912
2 2843 1 912
2 2844 1 912
2 2845 1 914
2 2846 1 914
2 2847 1 914
2 2848 1 916
2 2849 1 916
2 2850 1 916
2 2851 1 919
2 2852 1 919
2 2853 1 919
2 2854 1 919
2 2855 1 920
2 2856 1 920
2 2857 1 920
2 2858 1 922
2 2859 1 922
2 2860 1 922
2 2861 1 924
2 2862 1 924
2 2863 1 924
2 2864 1 927
2 2865 1 927
2 2866 1 927
2 2867 1 927
2 2868 1 928
2 2869 1 928
2 2870 1 928
2 2871 1 930
2 2872 1 930
2 2873 1 930
2 2874 1 932
2 2875 1 932
2 2876 1 932
2 2877 1 933
2 2878 1 933
2 2879 1 933
2 2880 1 935
2 2881 1 935
2 2882 1 936
2 2883 1 936
2 2884 1 936
2 2885 1 936
2 2886 1 936
2 2887 1 939
2 2888 1 939
2 2889 1 940
2 2890 1 940
2 2891 1 943
2 2892 1 943
2 2893 1 944
2 2894 1 944
2 2895 1 947
2 2896 1 947
2 2897 1 948
2 2898 1 948
2 2899 1 951
2 2900 1 951
2 2901 1 952
2 2902 1 952
2 2903 1 955
2 2904 1 955
2 2905 1 956
2 2906 1 956
2 2907 1 959
2 2908 1 959
2 2909 1 960
2 2910 1 960
2 2911 1 963
2 2912 1 963
2 2913 1 964
2 2914 1 964
2 2915 1 967
2 2916 1 967
2 2917 1 968
2 2918 1 968
2 2919 1 971
2 2920 1 971
2 2921 1 972
2 2922 1 972
2 2923 1 975
2 2924 1 975
2 2925 1 976
2 2926 1 976
2 2927 1 979
2 2928 1 979
2 2929 1 980
2 2930 1 980
2 2931 1 983
2 2932 1 983
2 2933 1 984
2 2934 1 984
2 2935 1 987
2 2936 1 987
2 2937 1 987
2 2938 1 987
2 2939 1 988
2 2940 1 988
2 2941 1 988
2 2942 1 990
2 2943 1 990
2 2944 1 990
2 2945 1 992
2 2946 1 992
2 2947 1 992
2 2948 1 993
2 2949 1 993
2 2950 1 993
2 2951 1 994
2 2952 1 994
2 2953 1 999
2 2954 1 999
2 2955 1 999
2 2956 1 1000
2 2957 1 1000
2 2958 1 1002
2 2959 1 1002
2 2960 1 1002
2 2961 1 1004
2 2962 1 1004
2 2963 1 1004
2 2964 1 1005
2 2965 1 1005
2 2966 1 1005
2 2967 1 1006
2 2968 1 1006
2 2969 1 1009
2 2970 1 1009
2 2971 1 1009
2 2972 1 1009
2 2973 1 1010
2 2974 1 1010
2 2975 1 1010
2 2976 1 1012
2 2977 1 1012
2 2978 1 1012
2 2979 1 1014
2 2980 1 1014
2 2981 1 1014
2 2982 1 1017
2 2983 1 1017
2 2984 1 1018
2 2985 1 1018
2 2986 1 1021
2 2987 1 1021
2 2988 1 1022
2 2989 1 1022
2 2990 1 1024
2 2991 1 1024
2 2992 1 1026
2 2993 1 1026
2 2994 1 1027
2 2995 1 1027
2 2996 1 1030
2 2997 1 1030
2 2998 1 1031
2 2999 1 1031
2 3000 1 1031
2 3001 1 1032
2 3002 1 1032
2 3003 1 1037
2 3004 1 1037
2 3005 1 1037
2 3006 1 1038
2 3007 1 1038
2 3008 1 1039
2 3009 1 1039
2 3010 1 1039
2 3011 1 1040
2 3012 1 1040
2 3013 1 1045
2 3014 1 1045
2 3015 1 1045
2 3016 1 1046
2 3017 1 1046
2 3018 1 1048
2 3019 1 1048
2 3020 1 1049
2 3021 1 1049
2 3022 1 1049
2 3023 1 1050
2 3024 1 1050
2 3025 1 1055
2 3026 1 1055
2 3027 1 1055
2 3028 1 1056
2 3029 1 1056
2 3030 1 1058
2 3031 1 1058
2 3032 1 1059
2 3033 1 1059
2 3034 1 1059
2 3035 1 1060
2 3036 1 1060
2 3037 1 1065
2 3038 1 1065
2 3039 1 1065
2 3040 1 1066
2 3041 1 1066
2 3042 1 1068
2 3043 1 1068
2 3044 1 1069
2 3045 1 1069
2 3046 1 1069
2 3047 1 1070
2 3048 1 1070
2 3049 1 1075
2 3050 1 1075
2 3051 1 1075
2 3052 1 1076
2 3053 1 1076
2 3054 1 1078
2 3055 1 1078
2 3056 1 1079
2 3057 1 1079
2 3058 1 1079
2 3059 1 1080
2 3060 1 1080
2 3061 1 1085
2 3062 1 1085
2 3063 1 1085
2 3064 1 1086
2 3065 1 1086
2 3066 1 1088
2 3067 1 1088
2 3068 1 1089
2 3069 1 1089
2 3070 1 1089
2 3071 1 1090
2 3072 1 1090
2 3073 1 1095
2 3074 1 1095
2 3075 1 1095
2 3076 1 1096
2 3077 1 1096
2 3078 1 1098
2 3079 1 1098
2 3080 1 1099
2 3081 1 1099
2 3082 1 1099
2 3083 1 1100
2 3084 1 1100
2 3085 1 1105
2 3086 1 1105
2 3087 1 1105
2 3088 1 1106
2 3089 1 1106
2 3090 1 1108
2 3091 1 1108
2 3092 1 1109
2 3093 1 1109
2 3094 1 1109
2 3095 1 1110
2 3096 1 1110
2 3097 1 1115
2 3098 1 1115
2 3099 1 1115
2 3100 1 1116
2 3101 1 1116
2 3102 1 1118
2 3103 1 1118
2 3104 1 1119
2 3105 1 1119
2 3106 1 1119
2 3107 1 1120
2 3108 1 1120
2 3109 1 1125
2 3110 1 1125
2 3111 1 1125
2 3112 1 1126
2 3113 1 1126
2 3114 1 1128
2 3115 1 1128
2 3116 1 1129
2 3117 1 1129
2 3118 1 1129
2 3119 1 1130
2 3120 1 1130
2 3121 1 1135
2 3122 1 1135
2 3123 1 1135
2 3124 1 1136
2 3125 1 1136
2 3126 1 1138
2 3127 1 1138
2 3128 1 1139
2 3129 1 1139
2 3130 1 1139
2 3131 1 1140
2 3132 1 1140
2 3133 1 1145
2 3134 1 1145
2 3135 1 1145
2 3136 1 1146
2 3137 1 1146
2 3138 1 1148
2 3139 1 1148
2 3140 1 1149
2 3141 1 1149
2 3142 1 1149
2 3143 1 1150
2 3144 1 1150
2 3145 1 1155
2 3146 1 1155
2 3147 1 1158
2 3148 1 1158
2 3149 1 1160
2 3150 1 1160
2 3151 1 1160
2 3152 1 1161
2 3153 1 1161
2 3154 1 1161
2 3155 1 1162
2 3156 1 1162
2 3157 1 1163
2 3158 1 1163
2 3159 1 1164
2 3160 1 1164
2 3161 1 1167
2 3162 1 1167
2 3163 1 1170
2 3164 1 1170
2 3165 1 1171
2 3166 1 1171
2 3167 1 1175
2 3168 1 1175
2 3169 1 1178
2 3170 1 1178
2 3171 1 1179
2 3172 1 1179
2 3173 1 1183
2 3174 1 1183
2 3175 1 1186
2 3176 1 1186
2 3177 1 1187
2 3178 1 1187
2 3179 1 1191
2 3180 1 1191
2 3181 1 1194
2 3182 1 1194
2 3183 1 1195
2 3184 1 1195
2 3185 1 1199
2 3186 1 1199
2 3187 1 1202
2 3188 1 1202
2 3189 1 1203
2 3190 1 1203
2 3191 1 1207
2 3192 1 1207
2 3193 1 1210
2 3194 1 1210
2 3195 1 1211
2 3196 1 1211
2 3197 1 1215
2 3198 1 1215
2 3199 1 1218
2 3200 1 1218
2 3201 1 1219
2 3202 1 1219
2 3203 1 1223
2 3204 1 1223
2 3205 1 1226
2 3206 1 1226
2 3207 1 1227
2 3208 1 1227
2 3209 1 1231
2 3210 1 1231
2 3211 1 1234
2 3212 1 1234
2 3213 1 1235
2 3214 1 1235
2 3215 1 1239
2 3216 1 1239
2 3217 1 1242
2 3218 1 1242
2 3219 1 1243
2 3220 1 1243
2 3221 1 1247
2 3222 1 1247
2 3223 1 1250
2 3224 1 1250
2 3225 1 1251
2 3226 1 1251
2 3227 1 1255
2 3228 1 1255
2 3229 1 1258
2 3230 1 1258
2 3231 1 1259
2 3232 1 1259
2 3233 1 1263
2 3234 1 1263
2 3235 1 1266
2 3236 1 1266
2 3237 1 1267
2 3238 1 1267
2 3239 1 1271
2 3240 1 1271
2 3241 1 1272
2 3242 1 1272
2 3243 1 1277
2 3244 1 1277
2 3245 1 1280
2 3246 1 1280
2 3247 1 1283
2 3248 1 1283
2 3249 1 1289
2 3250 1 1289
2 3251 1 1295
2 3252 1 1295
2 3253 1 1301
2 3254 1 1301
2 3255 1 1309
2 3256 1 1309
2 3257 1 1317
2 3258 1 1317
2 3259 1 1325
2 3260 1 1325
2 3261 1 1333
2 3262 1 1333
2 3263 1 1341
2 3264 1 1341
2 3265 1 1345
2 3266 1 1345
2 3267 1 1353
2 3268 1 1353
2 3269 1 1361
2 3270 1 1361
2 3271 1 1363
2 3272 1 1363
2 3273 1 1380
2 3274 1 1380
2 3275 1 1388
2 3276 1 1388
2 3277 1 1425
2 3278 1 1425
2 3279 1 1441
2 3280 1 1441
2 3281 1 1464
2 3282 1 1464
2 3283 1 1465
2 3284 1 1465
2 3285 1 1468
2 3286 1 1468
2 3287 1 1469
2 3288 1 1469
2 3289 1 1472
2 3290 1 1472
2 3291 1 1473
2 3292 1 1473
2 3293 1 1476
2 3294 1 1476
2 3295 1 1477
2 3296 1 1477
2 3297 1 1480
2 3298 1 1480
2 3299 1 1481
2 3300 1 1481
2 3301 1 1484
2 3302 1 1484
2 3303 1 1485
2 3304 1 1485
2 3305 1 1488
2 3306 1 1488
2 3307 1 1489
2 3308 1 1489
2 3309 1 1492
2 3310 1 1492
2 3311 1 1493
2 3312 1 1493
2 3313 1 1496
2 3314 1 1496
2 3315 1 1497
2 3316 1 1497
2 3317 1 1500
2 3318 1 1500
2 3319 1 1501
2 3320 1 1501
2 3321 1 1504
2 3322 1 1504
2 3323 1 1505
2 3324 1 1505
2 3325 1 1510
2 3326 1 1510
2 3327 1 1510
2 3328 1 1511
2 3329 1 1511
2 3330 1 1516
2 3331 1 1516
2 3332 1 1516
2 3333 1 1517
2 3334 1 1517
2 3335 1 1519
2 3336 1 1519
2 3337 1 1524
2 3338 1 1524
2 3339 1 1524
2 3340 1 1525
2 3341 1 1525
2 3342 1 1530
2 3343 1 1530
2 3344 1 1530
2 3345 1 1531
2 3346 1 1531
2 3347 1 1533
2 3348 1 1533
2 3349 1 1538
2 3350 1 1538
2 3351 1 1538
2 3352 1 1539
2 3353 1 1539
2 3354 1 1541
2 3355 1 1541
2 3356 1 1546
2 3357 1 1546
2 3358 1 1546
2 3359 1 1547
2 3360 1 1547
2 3361 1 1549
2 3362 1 1549
2 3363 1 1554
2 3364 1 1554
2 3365 1 1554
2 3366 1 1555
2 3367 1 1555
2 3368 1 1557
2 3369 1 1557
2 3370 1 1562
2 3371 1 1562
2 3372 1 1562
2 3373 1 1563
2 3374 1 1563
2 3375 1 1565
2 3376 1 1565
2 3377 1 1570
2 3378 1 1570
2 3379 1 1570
2 3380 1 1571
2 3381 1 1571
2 3382 1 1573
2 3383 1 1573
2 3384 1 1578
2 3385 1 1578
2 3386 1 1578
2 3387 1 1579
2 3388 1 1579
2 3389 1 1581
2 3390 1 1581
2 3391 1 1586
2 3392 1 1586
2 3393 1 1586
2 3394 1 1587
2 3395 1 1587
2 3396 1 1589
2 3397 1 1589
2 3398 1 1594
2 3399 1 1594
2 3400 1 1594
2 3401 1 1597
2 3402 1 1597
2 3403 1 1598
2 3404 1 1598
2 3405 1 1599
2 3406 1 1599
2 3407 1 1602
2 3408 1 1602
2 3409 1 1605
2 3410 1 1605
2 3411 1 1606
2 3412 1 1606
2 3413 1 1610
2 3414 1 1610
2 3415 1 1613
2 3416 1 1613
2 3417 1 1614
2 3418 1 1614
2 3419 1 1618
2 3420 1 1618
2 3421 1 1621
2 3422 1 1621
2 3423 1 1622
2 3424 1 1622
2 3425 1 1626
2 3426 1 1626
2 3427 1 1629
2 3428 1 1629
2 3429 1 1630
2 3430 1 1630
2 3431 1 1634
2 3432 1 1634
2 3433 1 1637
2 3434 1 1637
2 3435 1 1638
2 3436 1 1638
2 3437 1 1642
2 3438 1 1642
2 3439 1 1645
2 3440 1 1645
2 3441 1 1646
2 3442 1 1646
2 3443 1 1650
2 3444 1 1650
2 3445 1 1653
2 3446 1 1653
2 3447 1 1654
2 3448 1 1654
2 3449 1 1658
2 3450 1 1658
2 3451 1 1661
2 3452 1 1661
2 3453 1 1662
2 3454 1 1662
2 3455 1 1666
2 3456 1 1666
2 3457 1 1669
2 3458 1 1669
2 3459 1 1670
2 3460 1 1670
2 3461 1 1674
2 3462 1 1674
2 3463 1 1677
2 3464 1 1677
2 3465 1 1678
2 3466 1 1678
2 3467 1 1682
2 3468 1 1682
2 3469 1 1683
2 3470 1 1683
2 3471 1 1688
2 3472 1 1688
2 3473 1 1688
2 3474 1 1689
2 3475 1 1689
2 3476 1 1691
2 3477 1 1691
2 3478 1 1694
2 3479 1 1694
2 3480 1 1697
2 3481 1 1697
2 3482 1 1700
2 3483 1 1700
2 3484 1 1708
2 3485 1 1708
2 3486 1 1716
2 3487 1 1716
2 3488 1 1724
2 3489 1 1724
2 3490 1 1732
2 3491 1 1732
2 3492 1 1740
2 3493 1 1740
2 3494 1 1748
2 3495 1 1748
2 3496 1 1756
2 3497 1 1756
2 3498 1 1760
2 3499 1 1760
2 3500 1 1768
2 3501 1 1768
2 3502 1 1778
2 3503 1 1778
2 3504 1 1795
2 3505 1 1795
2 3506 1 1803
2 3507 1 1803
2 3508 1 1842
2 3509 1 1842
2 3510 1 1846
2 3511 1 1846
2 3512 1 1850
2 3513 1 1850
2 3514 1 1851
2 3515 1 1851
2 3516 1 1856
2 3517 1 1856
2 3518 1 1856
2 3519 1 1857
2 3520 1 1857
2 3521 1 1859
2 3522 1 1859
2 3523 1 1862
2 3524 1 1862
2 3525 1 1865
2 3526 1 1865
2 3527 1 1871
2 3528 1 1871
2 3529 1 1875
2 3530 1 1875
2 3531 1 1875
2 3532 1 1876
2 3533 1 1876
2 3534 1 1881
2 3535 1 1881
2 3536 1 1884
2 3537 1 1884
2 3538 1 1887
2 3539 1 1887
2 3540 1 1890
2 3541 1 1890
2 3542 1 1893
2 3543 1 1893
2 3544 1 1902
2 3545 1 1902
2 3546 1 1905
2 3547 1 1905
2 3548 1 1906
2 3549 1 1906
2 3550 1 1912
2 3551 1 1912
2 3552 1 1915
2 3553 1 1915
2 3554 1 1918
2 3555 1 1918
0 33 5 3 1 2067
0 34 5 1 1 2069
0 35 5 1 1 2071
0 36 5 1 1 2073
0 37 5 1 1 2075
0 38 5 1 1 2077
0 39 5 1 1 2079
0 40 5 1 1 2081
0 41 5 1 1 2083
0 42 5 1 1 2085
0 43 5 1 1 2087
0 44 5 1 1 2089
0 45 5 1 1 2091
0 46 5 1 1 2093
0 47 5 1 1 2095
0 48 5 1 1 2097
0 49 7 2 2 1994 2059
0 50 5 1 1 2102
0 51 7 2 2 1986 2051
0 52 5 2 1 2104
0 53 7 2 2 1977 2060
0 54 5 1 1 2108
0 55 7 2 2 1995 2043
0 56 5 1 1 2110
0 57 7 1 2 2109 2111
0 58 5 2 1 57
0 59 7 1 2 54 56
0 60 5 1 1 59
0 61 7 2 2 60 2112
0 62 5 1 1 2114
0 63 7 1 2 2105 2115
0 64 5 2 1 63
0 65 7 2 2 2113 2116
0 66 5 1 1 2118
0 67 7 2 2 1987 2061
0 68 5 1 1 2120
0 69 7 2 2 1996 2052
0 70 5 1 1 2122
0 71 7 1 2 68 2123
0 72 5 1 1 71
0 73 7 1 2 2121 70
0 74 5 1 1 73
0 75 7 2 2 72 74
0 76 5 1 1 2124
0 77 7 1 2 66 76
0 78 5 3 1 77
0 79 7 1 2 2106 2126
0 80 5 1 1 79
0 81 7 1 2 2103 80
0 82 5 2 1 81
0 83 7 2 2 1969 2062
0 84 5 1 1 2131
0 85 7 2 2 1997 2035
0 86 5 1 1 2133
0 87 7 1 2 2132 2134
0 88 5 2 1 87
0 89 7 2 2 1988 2044
0 90 5 1 1 2137
0 91 7 1 2 84 86
0 92 5 1 1 91
0 93 7 2 2 2135 92
0 94 5 1 1 2139
0 95 7 1 2 2138 2140
0 96 5 2 1 95
0 97 7 2 2 2136 2141
0 98 5 1 1 2143
0 99 7 1 2 2107 62
0 100 5 1 1 99
0 101 7 2 2 2117 100
0 102 5 1 1 2145
0 103 7 1 2 98 2146
0 104 5 2 1 103
0 105 7 2 2 1978 2053
0 106 5 1 1 2149
0 107 7 1 2 90 94
0 108 5 1 1 107
0 109 7 2 2 2142 108
0 110 5 1 1 2151
0 111 7 1 2 2150 2152
0 112 5 2 1 111
0 113 7 2 2 1960 2063
0 114 5 1 1 2155
0 115 7 2 2 1998 2027
0 116 5 1 1 2157
0 117 7 1 2 2156 2158
0 118 5 2 1 117
0 119 7 2 2 1989 2036
0 120 5 1 1 2161
0 121 7 1 2 114 116
0 122 5 1 1 121
0 123 7 2 2 2159 122
0 124 5 1 1 2163
0 125 7 1 2 2162 2164
0 126 5 2 1 125
0 127 7 2 2 2160 2165
0 128 5 1 1 2167
0 129 7 1 2 106 110
0 130 5 1 1 129
0 131 7 2 2 2153 130
0 132 5 1 1 2169
0 133 7 1 2 128 2170
0 134 5 2 1 133
0 135 7 2 2 2154 2171
0 136 5 1 1 2173
0 137 7 1 2 2144 102
0 138 5 1 1 137
0 139 7 2 2 2147 138
0 140 5 1 1 2175
0 141 7 1 2 136 2176
0 142 5 2 1 141
0 143 7 2 2 2148 2177
0 144 5 1 1 2179
0 145 7 1 2 2119 2125
0 146 5 1 1 145
0 147 7 2 2 2127 146
0 148 5 1 1 2181
0 149 7 1 2 144 2182
0 150 5 2 1 149
0 151 7 2 2 1970 2054
0 152 5 1 1 2185
0 153 7 1 2 120 124
0 154 5 1 1 153
0 155 7 2 2 2166 154
0 156 5 1 1 2187
0 157 7 1 2 2186 2188
0 158 5 2 1 157
0 159 7 2 2 1979 2045
0 160 5 1 1 2191
0 161 7 1 2 152 156
0 162 5 1 1 161
0 163 7 2 2 2189 162
0 164 5 1 1 2193
0 165 7 1 2 2192 2194
0 166 5 2 1 165
0 167 7 2 2 2190 2195
0 168 5 1 1 2197
0 169 7 1 2 2168 132
0 170 5 1 1 169
0 171 7 2 2 2172 170
0 172 5 1 1 2199
0 173 7 1 2 168 2200
0 174 5 2 1 173
0 175 7 2 2 1952 2064
0 176 5 1 1 2203
0 177 7 2 2 1999 2002
0 178 5 1 1 2205
0 179 7 2 2 1990 2010
0 180 5 1 1 2207
0 181 7 2 2 2206 2208
0 182 5 2 1 2209
0 183 7 2 2 2018 2210
0 184 5 2 1 2213
0 185 7 1 2 2204 2214
0 186 5 2 1 185
0 187 7 2 2 2000 2019
0 188 5 1 1 2219
0 189 7 1 2 176 2215
0 190 5 1 1 189
0 191 7 2 2 2217 190
0 192 5 1 1 2221
0 193 7 1 2 2220 2222
0 194 5 2 1 193
0 195 7 2 2 2218 2223
0 196 5 1 1 2225
0 197 7 1 2 160 164
0 198 5 1 1 197
0 199 7 2 2 2196 198
0 200 5 1 1 2227
0 201 7 1 2 196 2228
0 202 5 2 1 201
0 203 7 2 2 1980 2037
0 204 5 1 1 2231
0 205 7 1 2 188 192
0 206 5 1 1 205
0 207 7 2 2 2224 206
0 208 5 1 1 2233
0 209 7 1 2 2232 2234
0 210 5 2 1 209
0 211 7 2 2 1991 2028
0 212 5 1 1 2237
0 213 7 1 2 204 208
0 214 5 1 1 213
0 215 7 2 2 2235 214
0 216 5 1 1 2239
0 217 7 1 2 2238 2240
0 218 5 2 1 217
0 219 7 2 2 2236 2241
0 220 5 1 1 2243
0 221 7 1 2 2226 200
0 222 5 1 1 221
0 223 7 2 2 2229 222
0 224 5 1 1 2245
0 225 7 1 2 220 2246
0 226 5 2 1 225
0 227 7 2 2 2230 2247
0 228 5 1 1 2249
0 229 7 1 2 2198 172
0 230 5 1 1 229
0 231 7 2 2 2201 230
0 232 5 1 1 2251
0 233 7 1 2 228 2252
0 234 5 2 1 233
0 235 7 2 2 2202 2253
0 236 5 1 1 2255
0 237 7 1 2 2174 140
0 238 5 1 1 237
0 239 7 2 2 2178 238
0 240 5 1 1 2257
0 241 7 1 2 236 2258
0 242 5 2 1 241
0 243 7 2 2 1961 2055
0 244 5 1 1 2261
0 245 7 2 2 1971 2046
0 246 5 1 1 2263
0 247 7 1 2 2262 2264
0 248 5 2 1 247
0 249 7 1 2 212 216
0 250 5 1 1 249
0 251 7 2 2 2242 250
0 252 5 1 1 2267
0 253 7 1 2 244 246
0 254 5 1 1 253
0 255 7 2 2 2265 254
0 256 5 1 1 2269
0 257 7 1 2 2268 2270
0 258 5 2 1 257
0 259 7 2 2 2266 2271
0 260 5 1 1 2273
0 261 7 1 2 2244 224
0 262 5 1 1 261
0 263 7 2 2 2248 262
0 264 5 1 1 2275
0 265 7 1 2 260 2276
0 266 5 2 1 265
0 267 7 2 2 1981 2029
0 268 5 1 1 2279
0 269 7 2 2 1953 2056
0 270 5 1 1 2281
0 271 7 1 2 2280 2282
0 272 5 2 1 271
0 273 7 2 2 1944 2065
0 274 5 1 1 2285
0 275 7 2 2 1972 2038
0 276 5 1 1 2287
0 277 7 1 2 1992 2020
0 278 5 1 1 277
0 279 7 1 2 2211 278
0 280 5 1 1 279
0 281 7 2 2 2216 280
0 282 5 1 1 2289
0 283 7 1 2 2288 2290
0 284 5 2 1 283
0 285 7 1 2 276 282
0 286 5 1 1 285
0 287 7 2 2 2291 286
0 288 5 1 1 2293
0 289 7 1 2 2286 2294
0 290 5 2 1 289
0 291 7 1 2 274 288
0 292 5 1 1 291
0 293 7 2 2 2295 292
0 294 5 1 1 2297
0 295 7 1 2 268 270
0 296 5 1 1 295
0 297 7 2 2 2283 296
0 298 5 1 1 2299
0 299 7 1 2 2298 2300
0 300 5 2 1 299
0 301 7 2 2 2284 2301
0 302 5 1 1 2303
0 303 7 1 2 252 256
0 304 5 1 1 303
0 305 7 2 2 2272 304
0 306 5 1 1 2305
0 307 7 1 2 302 2306
0 308 5 2 1 307
0 309 7 2 2 2001 2011
0 310 5 1 1 2309
0 311 7 2 2 1962 2047
0 312 5 1 1 2311
0 313 7 1 2 2310 2312
0 314 5 2 1 313
0 315 7 1 2 294 298
0 316 5 1 1 315
0 317 7 2 2 2302 316
0 318 5 1 1 2315
0 319 7 1 2 310 312
0 320 5 1 1 319
0 321 7 2 2 2313 320
0 322 5 1 1 2317
0 323 7 1 2 2316 2318
0 324 5 2 1 323
0 325 7 2 2 2314 2319
0 326 5 1 1 2321
0 327 7 1 2 2304 306
0 328 5 1 1 327
0 329 7 2 2 2307 328
0 330 5 1 1 2323
0 331 7 1 2 326 2324
0 332 5 2 1 331
0 333 7 2 2 2308 2325
0 334 5 1 1 2327
0 335 7 1 2 2274 264
0 336 5 1 1 335
0 337 7 2 2 2277 336
0 338 5 1 1 2329
0 339 7 1 2 334 2330
0 340 5 2 1 339
0 341 7 2 2 2278 2331
0 342 5 1 1 2333
0 343 7 1 2 2250 232
0 344 5 1 1 343
0 345 7 2 2 2254 344
0 346 5 1 1 2335
0 347 7 1 2 342 2336
0 348 5 2 1 347
0 349 7 2 2 2292 2296
0 350 5 1 1 2339
0 351 7 1 2 2322 330
0 352 5 1 1 351
0 353 7 2 2 2326 352
0 354 5 1 1 2341
0 355 7 1 2 350 2342
0 356 5 2 1 355
0 357 7 2 2 1982 2021
0 358 5 1 1 2345
0 359 7 2 2 1973 2030
0 360 5 1 1 2347
0 361 7 1 2 2346 2348
0 362 5 2 1 361
0 363 7 2 2 1945 2057
0 364 5 1 1 2351
0 365 7 1 2 358 360
0 366 5 1 1 365
0 367 7 2 2 2349 366
0 368 5 1 1 2353
0 369 7 1 2 2352 2354
0 370 5 2 1 369
0 371 7 2 2 2350 2355
0 372 5 1 1 2357
0 373 7 2 2 1954 2048
0 374 5 1 1 2359
0 375 7 2 2 32 2066
0 376 5 1 1 2361
0 377 7 1 2 2360 2362
0 378 5 2 1 377
0 379 7 2 2 1963 2039
0 380 5 1 1 2365
0 381 7 2 2 1974 2012
0 382 5 1 1 2367
0 383 7 2 2 1937 2031
0 384 5 1 1 2369
0 385 7 2 2 1955 2013
0 386 5 1 1 2371
0 387 7 2 2 2370 2372
0 388 5 2 1 2373
0 389 7 2 2 1964 2374
0 390 5 2 1 2377
0 391 7 2 2 2368 2378
0 392 5 2 1 2381
0 393 7 2 2 1983 2382
0 394 5 2 1 2385
0 395 7 1 2 2366 2386
0 396 5 2 1 395
0 397 7 1 2 380 2387
0 398 5 1 1 397
0 399 7 2 2 2389 398
0 400 5 1 1 2391
0 401 7 1 2 178 180
0 402 5 1 1 401
0 403 7 2 2 2212 402
0 404 5 1 1 2393
0 405 7 1 2 2392 2394
0 406 5 2 1 405
0 407 7 1 2 400 404
0 408 5 1 1 407
0 409 7 2 2 2395 408
0 410 5 1 1 2397
0 411 7 1 2 374 376
0 412 5 1 1 411
0 413 7 2 2 2363 412
0 414 5 1 1 2399
0 415 7 1 2 2398 2400
0 416 5 2 1 415
0 417 7 2 2 2364 2401
0 418 5 1 1 2403
0 419 7 1 2 372 418
0 420 5 2 1 419
0 421 7 2 2 2390 2396
0 422 5 1 1 2407
0 423 7 1 2 2358 2404
0 424 5 1 1 423
0 425 7 2 2 2405 424
0 426 5 1 1 2409
0 427 7 1 2 422 2410
0 428 5 2 1 427
0 429 7 2 2 2406 2411
0 430 5 1 1 2413
0 431 7 1 2 2340 354
0 432 5 1 1 431
0 433 7 2 2 2343 432
0 434 5 1 1 2415
0 435 7 1 2 430 2416
0 436 5 2 1 435
0 437 7 2 2 2344 2417
0 438 5 1 1 2419
0 439 7 1 2 2328 338
0 440 5 1 1 439
0 441 7 2 2 2332 440
0 442 5 1 1 2421
0 443 7 1 2 438 2422
0 444 5 2 1 443
0 445 7 1 2 318 322
0 446 5 1 1 445
0 447 7 2 2 2320 446
0 448 5 1 1 2425
0 449 7 1 2 2408 426
0 450 5 1 1 449
0 451 7 2 2 2412 450
0 452 5 1 1 2427
0 453 7 1 2 2426 2428
0 454 5 2 1 453
0 455 7 1 2 364 368
0 456 5 1 1 455
0 457 7 2 2 2356 456
0 458 5 1 1 2431
0 459 7 1 2 410 414
0 460 5 1 1 459
0 461 7 2 2 2402 460
0 462 5 1 1 2433
0 463 7 1 2 2432 2434
0 464 5 2 1 463
0 465 7 2 2 1965 2032
0 466 5 1 1 2437
0 467 7 2 2 1956 2040
0 468 5 1 1 2439
0 469 7 1 2 2438 2440
0 470 5 2 1 469
0 471 7 2 2 1946 2049
0 472 5 1 1 2443
0 473 7 1 2 466 468
0 474 5 1 1 473
0 475 7 2 2 2441 474
0 476 5 1 1 2445
0 477 7 1 2 2444 2446
0 478 5 2 1 477
0 479 7 2 2 2442 2447
0 480 5 1 1 2449
0 481 7 1 2 458 462
0 482 5 1 1 481
0 483 7 2 2 2435 482
0 484 5 1 1 2451
0 485 7 1 2 480 2452
0 486 5 2 1 485
0 487 7 2 2 2436 2453
0 488 5 1 1 2455
0 489 7 1 2 448 452
0 490 5 1 1 489
0 491 7 2 2 2429 490
0 492 5 1 1 2457
0 493 7 1 2 488 2458
0 494 5 2 1 493
0 495 7 2 2 2430 2459
0 496 5 1 1 2461
0 497 7 1 2 2414 434
0 498 5 1 1 497
0 499 7 2 2 2418 498
0 500 5 1 1 2463
0 501 7 1 2 496 2464
0 502 5 2 1 501
0 503 7 2 2 1938 2058
0 504 5 1 1 2467
0 505 7 1 2 472 476
0 506 5 1 1 505
0 507 7 2 2 2448 506
0 508 5 1 1 2469
0 509 7 1 2 2468 2470
0 510 5 2 1 509
0 511 7 2 2 1993 2003
0 512 5 1 1 2473
0 513 7 2 2 1975 2022
0 514 5 1 1 2475
0 515 7 1 2 1984 2014
0 516 5 1 1 515
0 517 7 1 2 2383 516
0 518 5 1 1 517
0 519 7 2 2 2388 518
0 520 5 1 1 2477
0 521 7 1 2 2476 2478
0 522 5 2 1 521
0 523 7 1 2 514 520
0 524 5 1 1 523
0 525 7 2 2 2479 524
0 526 5 1 1 2481
0 527 7 1 2 2474 2482
0 528 5 2 1 527
0 529 7 1 2 512 526
0 530 5 1 1 529
0 531 7 2 2 2483 530
0 532 5 1 1 2485
0 533 7 1 2 504 508
0 534 5 1 1 533
0 535 7 2 2 2471 534
0 536 5 1 1 2487
0 537 7 1 2 2486 2488
0 538 5 2 1 537
0 539 7 2 2 2472 2489
0 540 5 1 1 2491
0 541 7 1 2 2450 484
0 542 5 1 1 541
0 543 7 2 2 2454 542
0 544 5 1 1 2493
0 545 7 1 2 540 2494
0 546 5 2 1 545
0 547 7 2 2 2480 2484
0 548 5 1 1 2497
0 549 7 1 2 2492 544
0 550 5 1 1 549
0 551 7 2 2 2495 550
0 552 5 1 1 2499
0 553 7 1 2 548 2500
0 554 5 2 1 553
0 555 7 2 2 2496 2501
0 556 5 1 1 2503
0 557 7 1 2 2456 492
0 558 5 1 1 557
0 559 7 2 2 2460 558
0 560 5 1 1 2505
0 561 7 1 2 556 2506
0 562 5 2 1 561
0 563 7 2 2 1966 2023
0 564 5 1 1 2509
0 565 7 1 2 382 2379
0 566 5 1 1 565
0 567 7 2 2 2384 566
0 568 5 1 1 2511
0 569 7 1 2 2510 2512
0 570 5 2 1 569
0 571 7 2 2 1985 2004
0 572 5 1 1 2515
0 573 7 1 2 564 568
0 574 5 1 1 573
0 575 7 2 2 2513 574
0 576 5 1 1 2517
0 577 7 1 2 2516 2518
0 578 5 2 1 577
0 579 7 2 2 2514 2519
0 580 5 1 1 2521
0 581 7 1 2 532 536
0 582 5 1 1 581
0 583 7 2 2 2490 582
0 584 5 1 1 2523
0 585 7 1 2 580 2524
0 586 5 2 1 585
0 587 7 2 2 1957 2033
0 588 5 1 1 2527
0 589 7 2 2 1939 2050
0 590 5 1 1 2529
0 591 7 1 2 2528 2530
0 592 5 2 1 591
0 593 7 1 2 572 576
0 594 5 1 1 593
0 595 7 2 2 2520 594
0 596 5 1 1 2533
0 597 7 1 2 588 590
0 598 5 1 1 597
0 599 7 2 2 2531 598
0 600 5 1 1 2535
0 601 7 1 2 2534 2536
0 602 5 2 1 601
0 603 7 2 2 2532 2537
0 604 5 1 1 2539
0 605 7 1 2 2522 584
0 606 5 1 1 605
0 607 7 2 2 2525 606
0 608 5 1 1 2541
0 609 7 1 2 604 2542
0 610 5 2 1 609
0 611 7 2 2 2526 2543
0 612 5 1 1 2545
0 613 7 1 2 2498 552
0 614 5 1 1 613
0 615 7 2 2 2502 614
0 616 5 1 1 2547
0 617 7 1 2 612 2548
0 618 5 2 1 617
0 619 7 2 2 1947 2041
0 620 5 1 1 2551
0 621 7 1 2 596 600
0 622 5 1 1 621
0 623 7 2 2 2538 622
0 624 5 1 1 2553
0 625 7 1 2 2552 2554
0 626 5 2 1 625
0 627 7 2 2 1958 2024
0 628 5 1 1 2557
0 629 7 1 2 1967 2015
0 630 5 1 1 629
0 631 7 1 2 2375 630
0 632 5 1 1 631
0 633 7 2 2 2380 632
0 634 5 1 1 2559
0 635 7 1 2 2558 2560
0 636 5 2 1 635
0 637 7 2 2 1976 2005
0 638 5 1 1 2563
0 639 7 1 2 628 634
0 640 5 1 1 639
0 641 7 2 2 2561 640
0 642 5 1 1 2565
0 643 7 1 2 2564 2566
0 644 5 2 1 643
0 645 7 2 2 2562 2567
0 646 5 1 1 2569
0 647 7 1 2 620 624
0 648 5 1 1 647
0 649 7 2 2 2555 648
0 650 5 1 1 2571
0 651 7 1 2 646 2572
0 652 5 2 1 651
0 653 7 2 2 2556 2573
0 654 5 1 1 2575
0 655 7 1 2 2540 608
0 656 5 1 1 655
0 657 7 2 2 2544 656
0 658 5 1 1 2577
0 659 7 1 2 654 2578
0 660 5 2 1 659
0 661 7 2 2 1940 2042
0 662 5 1 1 2581
0 663 7 2 2 1948 2034
0 664 5 1 1 2583
0 665 7 1 2 2582 2584
0 666 5 2 1 665
0 667 7 1 2 638 642
0 668 5 1 1 667
0 669 7 2 2 2568 668
0 670 5 1 1 2587
0 671 7 1 2 662 664
0 672 5 1 1 671
0 673 7 2 2 2585 672
0 674 5 1 1 2589
0 675 7 1 2 2588 2590
0 676 5 2 1 675
0 677 7 2 2 2586 2591
0 678 5 1 1 2593
0 679 7 1 2 2570 650
0 680 5 1 1 679
0 681 7 2 2 2574 680
0 682 5 1 1 2595
0 683 7 1 2 678 2596
0 684 5 2 1 683
0 685 7 1 2 670 674
0 686 5 1 1 685
0 687 7 2 2 2592 686
0 688 5 1 1 2599
0 689 7 2 2 1949 2025
0 690 5 1 1 2601
0 691 7 2 2 1968 2006
0 692 5 1 1 2603
0 693 7 2 2 2602 2604
0 694 5 1 1 2605
0 695 7 2 2 1950 2016
0 696 5 1 1 2607
0 697 7 2 2 1941 2026
0 698 5 1 1 2609
0 699 7 2 2 2608 2610
0 700 5 2 1 2611
0 701 7 3 2 694 2613
0 702 5 1 1 2615
0 703 7 1 2 2600 702
0 704 5 2 1 703
0 705 7 1 2 384 386
0 706 5 1 1 705
0 707 7 2 2 2376 706
0 708 5 1 1 2620
0 709 7 1 2 690 692
0 710 5 1 1 709
0 711 7 1 2 2616 710
0 712 5 1 1 711
0 713 7 1 2 2606 2612
0 714 5 1 1 713
0 715 7 2 2 712 714
0 716 5 1 1 2622
0 717 7 1 2 2621 716
0 718 5 2 1 717
0 719 7 2 2 1959 2007
0 720 5 1 1 2626
0 721 7 1 2 696 698
0 722 5 1 1 721
0 723 7 2 2 2614 722
0 724 5 1 1 2628
0 725 7 1 2 2627 2629
0 726 5 2 1 725
0 727 7 1 2 720 724
0 728 5 1 1 727
0 729 7 2 2 2630 728
0 730 5 1 1 2632
0 731 7 2 2 1942 2017
0 732 5 1 1 2634
0 733 7 2 2 1951 2008
0 734 5 1 1 2636
0 735 7 2 2 2635 2637
0 736 5 2 1 2638
0 737 7 1 2 2633 2639
0 738 5 2 1 737
0 739 7 2 2 2631 2642
0 740 5 1 1 2644
0 741 7 1 2 708 2623
0 742 5 1 1 741
0 743 7 2 2 2624 742
0 744 5 1 1 2646
0 745 7 1 2 740 2647
0 746 5 2 1 745
0 747 7 2 2 2625 2648
0 748 5 1 1 2650
0 749 7 1 2 688 2617
0 750 5 1 1 749
0 751 7 2 2 2618 750
0 752 5 1 1 2652
0 753 7 1 2 748 2653
0 754 5 2 1 753
0 755 7 2 2 2619 2654
0 756 5 1 1 2656
0 757 7 1 2 2594 682
0 758 5 1 1 757
0 759 7 2 2 2597 758
0 760 5 1 1 2658
0 761 7 1 2 756 2659
0 762 5 2 1 761
0 763 7 2 2 2598 2660
0 764 5 1 1 2662
0 765 7 1 2 2576 658
0 766 5 1 1 765
0 767 7 2 2 2579 766
0 768 5 1 1 2664
0 769 7 1 2 764 2665
0 770 5 2 1 769
0 771 7 2 2 2580 2666
0 772 5 1 1 2668
0 773 7 1 2 2546 616
0 774 5 1 1 773
0 775 7 2 2 2549 774
0 776 5 1 1 2670
0 777 7 1 2 772 2671
0 778 5 2 1 777
0 779 7 2 2 2550 2672
0 780 5 1 1 2674
0 781 7 1 2 2504 560
0 782 5 1 1 781
0 783 7 2 2 2507 782
0 784 5 1 1 2676
0 785 7 1 2 780 2677
0 786 5 2 1 785
0 787 7 2 2 2508 2678
0 788 5 1 1 2680
0 789 7 1 2 2462 500
0 790 5 1 1 789
0 791 7 2 2 2465 790
0 792 5 1 1 2682
0 793 7 1 2 788 2683
0 794 5 2 1 793
0 795 7 2 2 2466 2684
0 796 5 1 1 2686
0 797 7 1 2 2420 442
0 798 5 1 1 797
0 799 7 2 2 2423 798
0 800 5 1 1 2688
0 801 7 1 2 796 2689
0 802 5 2 1 801
0 803 7 2 2 2424 2690
0 804 5 1 1 2692
0 805 7 1 2 2334 346
0 806 5 1 1 805
0 807 7 2 2 2337 806
0 808 5 1 1 2694
0 809 7 1 2 804 2695
0 810 5 2 1 809
0 811 7 2 2 2338 2696
0 812 5 1 1 2698
0 813 7 1 2 2256 240
0 814 5 1 1 813
0 815 7 2 2 2259 814
0 816 5 1 1 2700
0 817 7 1 2 812 2701
0 818 5 2 1 817
0 819 7 2 2 2260 2702
0 820 5 1 1 2704
0 821 7 1 2 2180 148
0 822 5 1 1 821
0 823 7 2 2 2183 822
0 824 5 1 1 2706
0 825 7 1 2 820 2707
0 826 5 2 1 825
0 827 7 2 2 2184 2708
0 828 5 1 1 2710
0 829 7 1 2 2128 50
0 830 5 1 1 829
0 831 7 2 2 2129 830
0 832 5 1 1 2712
0 833 7 1 2 828 2713
0 834 5 2 1 833
0 835 7 4 2 2130 2714
0 836 5 3 1 2716
0 837 7 1 2 2699 816
0 838 5 1 1 837
0 839 7 4 2 2703 838
0 840 5 3 1 2723
0 841 7 1 2 45 2724
0 842 5 3 1 841
0 843 7 1 2 2092 2727
0 844 5 3 1 843
0 845 7 1 2 2693 808
0 846 5 1 1 845
0 847 7 4 2 2697 846
0 848 5 3 1 2736
0 849 7 1 2 44 2737
0 850 5 3 1 849
0 851 7 1 2 2090 2740
0 852 5 3 1 851
0 853 7 1 2 2687 800
0 854 5 1 1 853
0 855 7 4 2 2691 854
0 856 5 3 1 2749
0 857 7 1 2 43 2750
0 858 5 3 1 857
0 859 7 1 2 2088 2753
0 860 5 3 1 859
0 861 7 1 2 2681 792
0 862 5 1 1 861
0 863 7 4 2 2685 862
0 864 5 3 1 2762
0 865 7 1 2 42 2763
0 866 5 3 1 865
0 867 7 1 2 2086 2766
0 868 5 3 1 867
0 869 7 1 2 2675 784
0 870 5 1 1 869
0 871 7 4 2 2679 870
0 872 5 3 1 2775
0 873 7 1 2 41 2776
0 874 5 3 1 873
0 875 7 1 2 2084 2779
0 876 5 3 1 875
0 877 7 1 2 2669 776
0 878 5 1 1 877
0 879 7 4 2 2673 878
0 880 5 3 1 2788
0 881 7 1 2 40 2789
0 882 5 3 1 881
0 883 7 1 2 2082 2792
0 884 5 3 1 883
0 885 7 1 2 2663 768
0 886 5 1 1 885
0 887 7 4 2 2667 886
0 888 5 3 1 2801
0 889 7 1 2 39 2802
0 890 5 3 1 889
0 891 7 1 2 2080 2805
0 892 5 3 1 891
0 893 7 1 2 2657 760
0 894 5 1 1 893
0 895 7 4 2 2661 894
0 896 5 3 1 2814
0 897 7 1 2 38 2815
0 898 5 3 1 897
0 899 7 1 2 2078 2818
0 900 5 3 1 899
0 901 7 1 2 2651 752
0 902 5 1 1 901
0 903 7 2 2 2655 902
0 904 5 3 1 2827
0 905 7 1 2 37 2828
0 906 5 3 1 905
0 907 7 1 2 2076 2829
0 908 5 3 1 907
0 909 7 1 2 2645 744
0 910 5 1 1 909
0 911 7 4 2 2649 910
0 912 5 3 1 2838
0 913 7 1 2 36 2839
0 914 5 3 1 913
0 915 7 1 2 2074 2842
0 916 5 3 1 915
0 917 7 1 2 730 2640
0 918 5 1 1 917
0 919 7 4 2 2643 918
0 920 5 3 1 2851
0 921 7 1 2 35 2852
0 922 5 3 1 921
0 923 7 1 2 2072 2855
0 924 5 3 1 923
0 925 7 1 2 732 734
0 926 5 1 1 925
0 927 7 4 2 2641 926
0 928 5 3 1 2864
0 929 7 1 2 34 2865
0 930 5 3 1 929
0 931 7 1 2 2070 2868
0 932 5 3 1 931
0 933 7 3 2 1943 2009
0 934 5 1 1 2877
0 935 7 2 2 2068 934
0 936 5 5 1 2880
0 937 7 1 2 2874 2882
0 938 5 1 1 937
0 939 7 2 2 2871 938
0 940 5 2 1 2887
0 941 7 1 2 2861 2889
0 942 5 1 1 941
0 943 7 2 2 2858 942
0 944 5 2 1 2891
0 945 7 1 2 2848 2893
0 946 5 1 1 945
0 947 7 2 2 2845 946
0 948 5 2 1 2895
0 949 7 1 2 2835 2897
0 950 5 1 1 949
0 951 7 2 2 2832 950
0 952 5 2 1 2899
0 953 7 1 2 2824 2901
0 954 5 1 1 953
0 955 7 2 2 2821 954
0 956 5 2 1 2903
0 957 7 1 2 2811 2905
0 958 5 1 1 957
0 959 7 2 2 2808 958
0 960 5 2 1 2907
0 961 7 1 2 2798 2909
0 962 5 1 1 961
0 963 7 2 2 2795 962
0 964 5 2 1 2911
0 965 7 1 2 2785 2913
0 966 5 1 1 965
0 967 7 2 2 2782 966
0 968 5 2 1 2915
0 969 7 1 2 2772 2917
0 970 5 1 1 969
0 971 7 2 2 2769 970
0 972 5 2 1 2919
0 973 7 1 2 2759 2921
0 974 5 1 1 973
0 975 7 2 2 2756 974
0 976 5 2 1 2923
0 977 7 1 2 2746 2925
0 978 5 1 1 977
0 979 7 2 2 2743 978
0 980 5 2 1 2927
0 981 7 1 2 2733 2929
0 982 5 1 1 981
0 983 7 2 2 2730 982
0 984 5 2 1 2931
0 985 7 1 2 2705 824
0 986 5 1 1 985
0 987 7 4 2 2709 986
0 988 5 3 1 2935
0 989 7 1 2 46 2936
0 990 5 3 1 989
0 991 7 1 2 2094 2939
0 992 5 3 1 991
0 993 7 3 2 2942 2945
0 994 5 2 1 2948
0 995 7 1 2 2932 2951
0 996 5 1 1 995
0 997 7 1 2 2933 2949
0 998 5 1 1 997
0 999 7 3 2 996 998
0 1000 5 2 1 2953
0 1001 7 1 2 48 2720
0 1002 5 3 1 1001
0 1003 7 1 2 2098 2717
0 1004 5 3 1 1003
0 1005 7 3 2 2958 2961
0 1006 5 2 1 2964
0 1007 7 1 2 2711 832
0 1008 5 1 1 1007
0 1009 7 4 2 2715 1008
0 1010 5 3 1 2969
0 1011 7 1 2 47 2970
0 1012 5 3 1 1011
0 1013 7 1 2 2096 2973
0 1014 5 3 1 1013
0 1015 7 1 2 2946 2934
0 1016 5 1 1 1015
0 1017 7 2 2 2943 1016
0 1018 5 2 1 2982
0 1019 7 1 2 2979 2984
0 1020 5 1 1 1019
0 1021 7 2 2 2976 1020
0 1022 5 2 1 2986
0 1023 7 1 2 2967 2988
0 1024 5 2 1 1023
0 1025 7 1 2 2965 2987
0 1026 5 2 1 1025
0 1027 7 2 2 2990 2992
0 1028 5 1 1 2994
0 1029 7 1 2 2954 1028
0 1030 5 2 1 1029
0 1031 7 3 2 2734 2731
0 1032 5 2 1 2998
0 1033 7 1 2 3001 2928
0 1034 5 1 1 1033
0 1035 7 1 2 2999 2930
0 1036 5 1 1 1035
0 1037 7 3 2 1034 1036
0 1038 5 2 1 3003
0 1039 7 3 2 2980 2977
0 1040 5 2 1 3008
0 1041 7 1 2 3011 2983
0 1042 5 1 1 1041
0 1043 7 1 2 3009 2985
0 1044 5 1 1 1043
0 1045 7 3 2 1042 1044
0 1046 5 2 1 3013
0 1047 7 1 2 3004 3014
0 1048 5 2 1 1047
0 1049 7 3 2 2744 2747
0 1050 5 2 1 3020
0 1051 7 1 2 2924 3023
0 1052 5 1 1 1051
0 1053 7 1 2 2926 3021
0 1054 5 1 1 1053
0 1055 7 3 2 1052 1054
0 1056 5 2 1 3025
0 1057 7 1 2 2955 3026
0 1058 5 2 1 1057
0 1059 7 3 2 2757 2760
0 1060 5 2 1 3032
0 1061 7 1 2 2920 3035
0 1062 5 1 1 1061
0 1063 7 1 2 2922 3033
0 1064 5 1 1 1063
0 1065 7 3 2 1062 1064
0 1066 5 2 1 3037
0 1067 7 1 2 3005 3038
0 1068 5 2 1 1067
0 1069 7 3 2 2770 2773
0 1070 5 2 1 3044
0 1071 7 1 2 2916 3047
0 1072 5 1 1 1071
0 1073 7 1 2 2918 3045
0 1074 5 1 1 1073
0 1075 7 3 2 1072 1074
0 1076 5 2 1 3049
0 1077 7 1 2 3027 3050
0 1078 5 2 1 1077
0 1079 7 3 2 2783 2786
0 1080 5 2 1 3056
0 1081 7 1 2 2912 3059
0 1082 5 1 1 1081
0 1083 7 1 2 2914 3057
0 1084 5 1 1 1083
0 1085 7 3 2 1082 1084
0 1086 5 2 1 3061
0 1087 7 1 2 3039 3062
0 1088 5 2 1 1087
0 1089 7 3 2 2796 2799
0 1090 5 2 1 3068
0 1091 7 1 2 2908 3071
0 1092 5 1 1 1091
0 1093 7 1 2 2910 3069
0 1094 5 1 1 1093
0 1095 7 3 2 1092 1094
0 1096 5 2 1 3073
0 1097 7 1 2 3051 3074
0 1098 5 2 1 1097
0 1099 7 3 2 2809 2812
0 1100 5 2 1 3080
0 1101 7 1 2 2904 3083
0 1102 5 1 1 1101
0 1103 7 1 2 2906 3081
0 1104 5 1 1 1103
0 1105 7 3 2 1102 1104
0 1106 5 2 1 3085
0 1107 7 1 2 3063 3086
0 1108 5 2 1 1107
0 1109 7 3 2 2822 2825
0 1110 5 2 1 3092
0 1111 7 1 2 2900 3095
0 1112 5 1 1 1111
0 1113 7 1 2 2902 3093
0 1114 5 1 1 1113
0 1115 7 3 2 1112 1114
0 1116 5 2 1 3097
0 1117 7 1 2 3075 3098
0 1118 5 2 1 1117
0 1119 7 3 2 2833 2836
0 1120 5 2 1 3104
0 1121 7 1 2 2896 3107
0 1122 5 1 1 1121
0 1123 7 1 2 2898 3105
0 1124 5 1 1 1123
0 1125 7 3 2 1122 1124
0 1126 5 2 1 3109
0 1127 7 1 2 3087 3110
0 1128 5 2 1 1127
0 1129 7 3 2 2846 2849
0 1130 5 2 1 3116
0 1131 7 1 2 2892 3119
0 1132 5 1 1 1131
0 1133 7 1 2 2894 3117
0 1134 5 1 1 1133
0 1135 7 3 2 1132 1134
0 1136 5 2 1 3121
0 1137 7 1 2 3099 3122
0 1138 5 2 1 1137
0 1139 7 3 2 2859 2862
0 1140 5 2 1 3128
0 1141 7 1 2 2888 3131
0 1142 5 1 1 1141
0 1143 7 1 2 2890 3129
0 1144 5 1 1 1143
0 1145 7 3 2 1142 1144
0 1146 5 2 1 3133
0 1147 7 1 2 3111 3134
0 1148 5 2 1 1147
0 1149 7 3 2 2872 2875
0 1150 5 2 1 3140
0 1151 7 1 2 2881 3141
0 1152 5 1 1 1151
0 1153 7 1 2 2883 3143
0 1154 5 1 1 1153
0 1155 7 2 2 1152 1154
0 1156 5 1 1 3145
0 1157 7 1 2 3123 1156
0 1158 5 2 1 1157
0 1159 7 1 2 2099 2878
0 1160 5 3 1 1159
0 1161 7 3 2 2884 3149
0 1162 5 2 1 3152
0 1163 7 2 2 3135 3155
0 1164 5 2 1 3157
0 1165 7 1 2 3124 3146
0 1166 5 1 1 1165
0 1167 7 2 2 3147 1166
0 1168 5 1 1 3161
0 1169 7 1 2 3158 3162
0 1170 5 2 1 1169
0 1171 7 2 2 3148 3163
0 1172 5 1 1 3165
0 1173 7 1 2 3112 3136
0 1174 5 1 1 1173
0 1175 7 2 2 3138 1174
0 1176 5 1 1 3167
0 1177 7 1 2 1172 3168
0 1178 5 2 1 1177
0 1179 7 2 2 3139 3169
0 1180 5 1 1 3171
0 1181 7 1 2 3100 3125
0 1182 5 1 1 1181
0 1183 7 2 2 3126 1182
0 1184 5 1 1 3173
0 1185 7 1 2 1180 3174
0 1186 5 2 1 1185
0 1187 7 2 2 3127 3175
0 1188 5 1 1 3177
0 1189 7 1 2 3088 3113
0 1190 5 1 1 1189
0 1191 7 2 2 3114 1190
0 1192 5 1 1 3179
0 1193 7 1 2 1188 3180
0 1194 5 2 1 1193
0 1195 7 2 2 3115 3181
0 1196 5 1 1 3183
0 1197 7 1 2 3076 3101
0 1198 5 1 1 1197
0 1199 7 2 2 3102 1198
0 1200 5 1 1 3185
0 1201 7 1 2 1196 3186
0 1202 5 2 1 1201
0 1203 7 2 2 3103 3187
0 1204 5 1 1 3189
0 1205 7 1 2 3064 3089
0 1206 5 1 1 1205
0 1207 7 2 2 3090 1206
0 1208 5 1 1 3191
0 1209 7 1 2 1204 3192
0 1210 5 2 1 1209
0 1211 7 2 2 3091 3193
0 1212 5 1 1 3195
0 1213 7 1 2 3052 3077
0 1214 5 1 1 1213
0 1215 7 2 2 3078 1214
0 1216 5 1 1 3197
0 1217 7 1 2 1212 3198
0 1218 5 2 1 1217
0 1219 7 2 2 3079 3199
0 1220 5 1 1 3201
0 1221 7 1 2 3040 3065
0 1222 5 1 1 1221
0 1223 7 2 2 3066 1222
0 1224 5 1 1 3203
0 1225 7 1 2 1220 3204
0 1226 5 2 1 1225
0 1227 7 2 2 3067 3205
0 1228 5 1 1 3207
0 1229 7 1 2 3028 3053
0 1230 5 1 1 1229
0 1231 7 2 2 3054 1230
0 1232 5 1 1 3209
0 1233 7 1 2 1228 3210
0 1234 5 2 1 1233
0 1235 7 2 2 3055 3211
0 1236 5 1 1 3213
0 1237 7 1 2 3006 3041
0 1238 5 1 1 1237
0 1239 7 2 2 3042 1238
0 1240 5 1 1 3215
0 1241 7 1 2 1236 3216
0 1242 5 2 1 1241
0 1243 7 2 2 3043 3217
0 1244 5 1 1 3219
0 1245 7 1 2 2956 3029
0 1246 5 1 1 1245
0 1247 7 2 2 3030 1246
0 1248 5 1 1 3221
0 1249 7 1 2 1244 3222
0 1250 5 2 1 1249
0 1251 7 2 2 3031 3223
0 1252 5 1 1 3225
0 1253 7 1 2 3007 3016
0 1254 5 1 1 1253
0 1255 7 2 2 3018 1254
0 1256 5 1 1 3227
0 1257 7 1 2 1252 3228
0 1258 5 2 1 1257
0 1259 7 2 2 3019 3229
0 1260 5 1 1 3231
0 1261 7 1 2 2957 2995
0 1262 5 1 1 1261
0 1263 7 2 2 2996 1262
0 1264 5 1 1 3233
0 1265 7 1 2 1260 3234
0 1266 5 2 1 1265
0 1267 7 2 2 2997 3235
0 1268 5 1 1 3237
0 1269 7 1 2 2962 2989
0 1270 5 1 1 1269
0 1271 7 2 2 2959 1270
0 1272 5 2 1 3239
0 1273 7 1 2 3015 3241
0 1274 5 1 1 1273
0 1275 7 1 2 3017 3240
0 1276 5 1 1 1275
0 1277 7 2 2 1274 1276
0 1278 5 1 1 3243
0 1279 7 1 2 1268 1278
0 1280 5 2 1 1279
0 1281 7 1 2 3238 3244
0 1282 5 1 1 1281
0 1283 7 2 2 3245 1282
0 1284 5 1 1 3247
0 1285 7 1 2 2721 1284
0 1286 5 1 1 1285
0 1287 7 1 2 3226 1256
0 1288 5 1 1 1287
0 1289 7 2 2 3230 1288
0 1290 5 1 1 3249
0 1291 7 1 2 2937 1290
0 1292 5 1 1 1291
0 1293 7 1 2 3214 1240
0 1294 5 1 1 1293
0 1295 7 2 2 3218 1294
0 1296 5 1 1 3251
0 1297 7 1 2 2738 1296
0 1298 5 1 1 1297
0 1299 7 1 2 3208 1232
0 1300 5 1 1 1299
0 1301 7 2 2 3212 1300
0 1302 5 1 1 3253
0 1303 7 1 2 2754 3254
0 1304 5 1 1 1303
0 1305 7 1 2 2751 1302
0 1306 5 1 1 1305
0 1307 7 1 2 3202 1224
0 1308 5 1 1 1307
0 1309 7 2 2 3206 1308
0 1310 5 1 1 3255
0 1311 7 1 2 2767 3256
0 1312 5 1 1 1311
0 1313 7 1 2 2764 1310
0 1314 5 1 1 1313
0 1315 7 1 2 3196 1216
0 1316 5 1 1 1315
0 1317 7 2 2 3200 1316
0 1318 5 1 1 3257
0 1319 7 1 2 2780 3258
0 1320 5 1 1 1319
0 1321 7 1 2 2777 1318
0 1322 5 1 1 1321
0 1323 7 1 2 3190 1208
0 1324 5 1 1 1323
0 1325 7 2 2 3194 1324
0 1326 5 1 1 3259
0 1327 7 1 2 2793 3260
0 1328 5 1 1 1327
0 1329 7 1 2 2790 1326
0 1330 5 1 1 1329
0 1331 7 1 2 3184 1200
0 1332 5 1 1 1331
0 1333 7 2 2 3188 1332
0 1334 5 1 1 3261
0 1335 7 1 2 2806 3262
0 1336 5 1 1 1335
0 1337 7 1 2 2803 1334
0 1338 5 1 1 1337
0 1339 7 1 2 3172 1184
0 1340 5 1 1 1339
0 1341 7 2 2 3176 1340
0 1342 5 1 1 3263
0 1343 7 1 2 3166 1176
0 1344 5 1 1 1343
0 1345 7 2 2 3170 1344
0 1346 5 1 1 3265
0 1347 7 1 2 2843 3266
0 1348 5 1 1 1347
0 1349 7 1 2 2840 1346
0 1350 5 1 1 1349
0 1351 7 1 2 3159 1168
0 1352 5 1 1 1351
0 1353 7 2 2 3164 1352
0 1354 5 1 1 3267
0 1355 7 1 2 2856 3268
0 1356 5 1 1 1355
0 1357 7 1 2 2853 1354
0 1358 5 1 1 1357
0 1359 7 1 2 3137 3153
0 1360 5 1 1 1359
0 1361 7 2 2 2100 3144
0 1362 5 1 1 3269
0 1363 7 2 2 2885 1362
0 1364 5 1 1 3271
0 1365 7 1 2 2866 3272
0 1366 5 1 1 1365
0 1367 7 1 2 3160 1366
0 1368 7 1 2 1360 1367
0 1369 5 1 1 1368
0 1370 7 1 2 2869 1364
0 1371 5 1 1 1370
0 1372 7 1 2 1369 1371
0 1373 5 1 1 1372
0 1374 7 1 2 1358 1373
0 1375 5 1 1 1374
0 1376 7 1 2 1356 1375
0 1377 5 1 1 1376
0 1378 7 1 2 1350 1377
0 1379 5 1 1 1378
0 1380 7 2 2 1348 1379
0 1381 5 1 1 3273
0 1382 7 1 2 3264 1381
0 1383 5 1 1 1382
0 1384 7 1 2 1342 3274
0 1385 5 1 1 1384
0 1386 7 1 2 2830 1385
0 1387 5 1 1 1386
0 1388 7 2 2 1383 1387
0 1389 5 1 1 3275
0 1390 7 1 2 2816 3276
0 1391 5 1 1 1390
0 1392 7 1 2 3178 1192
0 1393 5 1 1 1392
0 1394 7 1 2 3182 1393
0 1395 7 1 2 1391 1394
0 1396 5 1 1 1395
0 1397 7 1 2 2819 1389
0 1398 5 1 1 1397
0 1399 7 1 2 1396 1398
0 1400 5 1 1 1399
0 1401 7 1 2 1338 1400
0 1402 5 1 1 1401
0 1403 7 1 2 1336 1402
0 1404 5 1 1 1403
0 1405 7 1 2 1330 1404
0 1406 5 1 1 1405
0 1407 7 1 2 1328 1406
0 1408 5 1 1 1407
0 1409 7 1 2 1322 1408
0 1410 5 1 1 1409
0 1411 7 1 2 1320 1410
0 1412 5 1 1 1411
0 1413 7 1 2 1314 1412
0 1414 5 1 1 1413
0 1415 7 1 2 1312 1414
0 1416 5 1 1 1415
0 1417 7 1 2 1306 1416
0 1418 5 1 1 1417
0 1419 7 1 2 1304 1418
0 1420 5 1 1 1419
0 1421 7 1 2 1298 1420
0 1422 5 1 1 1421
0 1423 7 1 2 3220 1248
0 1424 5 1 1 1423
0 1425 7 2 2 3224 1424
0 1426 5 1 1 3277
0 1427 7 1 2 2728 3278
0 1428 5 1 1 1427
0 1429 7 1 2 2741 3252
0 1430 5 1 1 1429
0 1431 7 1 2 1428 1430
0 1432 7 1 2 1422 1431
0 1433 5 1 1 1432
0 1434 7 1 2 2725 1426
0 1435 5 1 1 1434
0 1436 7 1 2 1433 1435
0 1437 7 1 2 1292 1436
0 1438 5 1 1 1437
0 1439 7 1 2 3232 1264
0 1440 5 1 1 1439
0 1441 7 2 2 3236 1440
0 1442 5 1 1 3279
0 1443 7 1 2 2974 3280
0 1444 5 1 1 1443
0 1445 7 1 2 2940 3250
0 1446 5 1 1 1445
0 1447 7 1 2 1444 1446
0 1448 7 1 2 1438 1447
0 1449 5 1 1 1448
0 1450 7 1 2 2971 1442
0 1451 5 1 1 1450
0 1452 7 1 2 1449 1451
0 1453 7 1 2 1286 1452
0 1454 5 1 1 1453
0 1455 7 1 2 2718 3248
0 1456 5 1 1 1455
0 1457 7 1 2 2991 3242
0 1458 7 1 2 3246 1457
0 1459 7 1 2 1456 1458
0 1460 7 1 2 1454 1459
0 1461 5 1 1 1460
0 1462 7 1 2 2873 3150
0 1463 5 1 1 1462
0 1464 7 2 2 2876 1463
0 1465 5 2 1 3281
0 1466 7 1 2 2860 3283
0 1467 5 1 1 1466
0 1468 7 2 2 2863 1467
0 1469 5 2 1 3285
0 1470 7 1 2 2847 3287
0 1471 5 1 1 1470
0 1472 7 2 2 2850 1471
0 1473 5 2 1 3289
0 1474 7 1 2 2834 3291
0 1475 5 1 1 1474
0 1476 7 2 2 2837 1475
0 1477 5 2 1 3293
0 1478 7 1 2 2823 3295
0 1479 5 1 1 1478
0 1480 7 2 2 2826 1479
0 1481 5 2 1 3297
0 1482 7 1 2 2810 3299
0 1483 5 1 1 1482
0 1484 7 2 2 2813 1483
0 1485 5 2 1 3301
0 1486 7 1 2 2797 3303
0 1487 5 1 1 1486
0 1488 7 2 2 2800 1487
0 1489 5 2 1 3305
0 1490 7 1 2 2784 3307
0 1491 5 1 1 1490
0 1492 7 2 2 2787 1491
0 1493 5 2 1 3309
0 1494 7 1 2 2771 3311
0 1495 5 1 1 1494
0 1496 7 2 2 2774 1495
0 1497 5 2 1 3313
0 1498 7 1 2 2758 3315
0 1499 5 1 1 1498
0 1500 7 2 2 2761 1499
0 1501 5 2 1 3317
0 1502 7 1 2 2745 3319
0 1503 5 1 1 1502
0 1504 7 2 2 2748 1503
0 1505 5 2 1 3321
0 1506 7 1 2 3000 3323
0 1507 5 1 1 1506
0 1508 7 1 2 3002 3322
0 1509 5 1 1 1508
0 1510 7 3 2 1507 1509
0 1511 5 2 1 3325
0 1512 7 1 2 3034 3316
0 1513 5 1 1 1512
0 1514 7 1 2 3036 3314
0 1515 5 1 1 1514
0 1516 7 3 2 1513 1515
0 1517 5 2 1 3330
0 1518 7 1 2 3326 3331
0 1519 5 2 1 1518
0 1520 7 1 2 3022 3320
0 1521 5 1 1 1520
0 1522 7 1 2 3024 3318
0 1523 5 1 1 1522
0 1524 7 3 2 1521 1523
0 1525 5 2 1 3337
0 1526 7 1 2 3046 3312
0 1527 5 1 1 1526
0 1528 7 1 2 3048 3310
0 1529 5 1 1 1528
0 1530 7 3 2 1527 1529
0 1531 5 2 1 3342
0 1532 7 1 2 3338 3343
0 1533 5 2 1 1532
0 1534 7 1 2 3058 3308
0 1535 5 1 1 1534
0 1536 7 1 2 3060 3306
0 1537 5 1 1 1536
0 1538 7 3 2 1535 1537
0 1539 5 2 1 3349
0 1540 7 1 2 3332 3350
0 1541 5 2 1 1540
0 1542 7 1 2 3070 3304
0 1543 5 1 1 1542
0 1544 7 1 2 3072 3302
0 1545 5 1 1 1544
0 1546 7 3 2 1543 1545
0 1547 5 2 1 3356
0 1548 7 1 2 3344 3357
0 1549 5 2 1 1548
0 1550 7 1 2 3082 3300
0 1551 5 1 1 1550
0 1552 7 1 2 3084 3298
0 1553 5 1 1 1552
0 1554 7 3 2 1551 1553
0 1555 5 2 1 3363
0 1556 7 1 2 3351 3364
0 1557 5 2 1 1556
0 1558 7 1 2 3094 3296
0 1559 5 1 1 1558
0 1560 7 1 2 3096 3294
0 1561 5 1 1 1560
0 1562 7 3 2 1559 1561
0 1563 5 2 1 3370
0 1564 7 1 2 3358 3371
0 1565 5 2 1 1564
0 1566 7 1 2 3106 3292
0 1567 5 1 1 1566
0 1568 7 1 2 3108 3290
0 1569 5 1 1 1568
0 1570 7 3 2 1567 1569
0 1571 5 2 1 3377
0 1572 7 1 2 3365 3378
0 1573 5 2 1 1572
0 1574 7 1 2 3118 3288
0 1575 5 1 1 1574
0 1576 7 1 2 3120 3286
0 1577 5 1 1 1576
0 1578 7 3 2 1575 1577
0 1579 5 2 1 3384
0 1580 7 1 2 3372 3385
0 1581 5 2 1 1580
0 1582 7 1 2 3130 3284
0 1583 5 1 1 1582
0 1584 7 1 2 3132 3282
0 1585 5 1 1 1584
0 1586 7 3 2 1583 1585
0 1587 5 2 1 3391
0 1588 7 1 2 3379 3392
0 1589 5 2 1 1588
0 1590 7 1 2 3142 3151
0 1591 5 1 1 1590
0 1592 7 1 2 2879 3270
0 1593 5 1 1 1592
0 1594 7 3 2 1591 1593
0 1595 5 1 1 3398
0 1596 7 1 2 3386 3399
0 1597 5 2 1 1596
0 1598 7 2 2 3156 3393
0 1599 5 2 1 3403
0 1600 7 1 2 3387 1595
0 1601 5 1 1 1600
0 1602 7 2 2 3401 1601
0 1603 5 1 1 3407
0 1604 7 1 2 3404 3408
0 1605 5 2 1 1604
0 1606 7 2 2 3402 3409
0 1607 5 1 1 3411
0 1608 7 1 2 3380 3394
0 1609 5 1 1 1608
0 1610 7 2 2 3396 1609
0 1611 5 1 1 3413
0 1612 7 1 2 1607 3414
0 1613 5 2 1 1612
0 1614 7 2 2 3397 3415
0 1615 5 1 1 3417
0 1616 7 1 2 3373 3388
0 1617 5 1 1 1616
0 1618 7 2 2 3389 1617
0 1619 5 1 1 3419
0 1620 7 1 2 1615 3420
0 1621 5 2 1 1620
0 1622 7 2 2 3390 3421
0 1623 5 1 1 3423
0 1624 7 1 2 3366 3381
0 1625 5 1 1 1624
0 1626 7 2 2 3382 1625
0 1627 5 1 1 3425
0 1628 7 1 2 1623 3426
0 1629 5 2 1 1628
0 1630 7 2 2 3383 3427
0 1631 5 1 1 3429
0 1632 7 1 2 3359 3374
0 1633 5 1 1 1632
0 1634 7 2 2 3375 1633
0 1635 5 1 1 3431
0 1636 7 1 2 1631 3432
0 1637 5 2 1 1636
0 1638 7 2 2 3376 3433
0 1639 5 1 1 3435
0 1640 7 1 2 3352 3367
0 1641 5 1 1 1640
0 1642 7 2 2 3368 1641
0 1643 5 1 1 3437
0 1644 7 1 2 1639 3438
0 1645 5 2 1 1644
0 1646 7 2 2 3369 3439
0 1647 5 1 1 3441
0 1648 7 1 2 3345 3360
0 1649 5 1 1 1648
0 1650 7 2 2 3361 1649
0 1651 5 1 1 3443
0 1652 7 1 2 1647 3444
0 1653 5 2 1 1652
0 1654 7 2 2 3362 3445
0 1655 5 1 1 3447
0 1656 7 1 2 3333 3353
0 1657 5 1 1 1656
0 1658 7 2 2 3354 1657
0 1659 5 1 1 3449
0 1660 7 1 2 1655 3450
0 1661 5 2 1 1660
0 1662 7 2 2 3355 3451
0 1663 5 1 1 3453
0 1664 7 1 2 3340 3346
0 1665 5 1 1 1664
0 1666 7 2 2 3347 1665
0 1667 5 1 1 3455
0 1668 7 1 2 1663 3456
0 1669 5 2 1 1668
0 1670 7 2 2 3348 3457
0 1671 5 1 1 3459
0 1672 7 1 2 3328 3334
0 1673 5 1 1 1672
0 1674 7 2 2 3335 1673
0 1675 5 1 1 3461
0 1676 7 1 2 1671 3462
0 1677 5 2 1 1676
0 1678 7 2 2 3336 3463
0 1679 5 1 1 3465
0 1680 7 1 2 2732 3324
0 1681 5 1 1 1680
0 1682 7 2 2 2735 1681
0 1683 5 2 1 3467
0 1684 7 1 2 2952 3468
0 1685 5 1 1 1684
0 1686 7 1 2 2950 3469
0 1687 5 1 1 1686
0 1688 7 3 2 1685 1687
0 1689 5 2 1 3471
0 1690 7 1 2 3472 3339
0 1691 5 2 1 1690
0 1692 7 1 2 3474 3341
0 1693 5 1 1 1692
0 1694 7 2 2 3476 1693
0 1695 5 1 1 3478
0 1696 7 1 2 1679 3479
0 1697 5 2 1 1696
0 1698 7 1 2 3466 1695
0 1699 5 1 1 1698
0 1700 7 2 2 3480 1699
0 1701 5 1 1 3482
0 1702 7 1 2 2729 3483
0 1703 5 1 1 1702
0 1704 7 1 2 2726 1701
0 1705 5 1 1 1704
0 1706 7 1 2 3460 1675
0 1707 5 1 1 1706
0 1708 7 2 2 3464 1707
0 1709 5 1 1 3484
0 1710 7 1 2 2742 3485
0 1711 5 1 1 1710
0 1712 7 1 2 2739 1709
0 1713 5 1 1 1712
0 1714 7 1 2 3454 1667
0 1715 5 1 1 1714
0 1716 7 2 2 3458 1715
0 1717 5 1 1 3486
0 1718 7 1 2 2755 3487
0 1719 5 1 1 1718
0 1720 7 1 2 2752 1717
0 1721 5 1 1 1720
0 1722 7 1 2 3448 1659
0 1723 5 1 1 1722
0 1724 7 2 2 3452 1723
0 1725 5 1 1 3488
0 1726 7 1 2 2768 3489
0 1727 5 1 1 1726
0 1728 7 1 2 2765 1725
0 1729 5 1 1 1728
0 1730 7 1 2 3442 1651
0 1731 5 1 1 1730
0 1732 7 2 2 3446 1731
0 1733 5 1 1 3490
0 1734 7 1 2 2781 3491
0 1735 5 1 1 1734
0 1736 7 1 2 2778 1733
0 1737 5 1 1 1736
0 1738 7 1 2 3436 1643
0 1739 5 1 1 1738
0 1740 7 2 2 3440 1739
0 1741 5 1 1 3492
0 1742 7 1 2 2794 3493
0 1743 5 1 1 1742
0 1744 7 1 2 2791 1741
0 1745 5 1 1 1744
0 1746 7 1 2 3430 1635
0 1747 5 1 1 1746
0 1748 7 2 2 3434 1747
0 1749 5 1 1 3494
0 1750 7 1 2 2807 3495
0 1751 5 1 1 1750
0 1752 7 1 2 2804 1749
0 1753 5 1 1 1752
0 1754 7 1 2 3418 1619
0 1755 5 1 1 1754
0 1756 7 2 2 3422 1755
0 1757 5 1 1 3496
0 1758 7 1 2 3412 1611
0 1759 5 1 1 1758
0 1760 7 2 2 3416 1759
0 1761 5 1 1 3498
0 1762 7 1 2 2844 3499
0 1763 5 1 1 1762
0 1764 7 1 2 2841 1761
0 1765 5 1 1 1764
0 1766 7 1 2 3405 1603
0 1767 5 1 1 1766
0 1768 7 2 2 3410 1767
0 1769 5 1 1 3500
0 1770 7 1 2 2857 3501
0 1771 5 1 1 1770
0 1772 7 1 2 2854 1769
0 1773 5 1 1 1772
0 1774 7 1 2 3154 3395
0 1775 5 1 1 1774
0 1776 7 1 2 2101 3400
0 1777 5 1 1 1776
0 1778 7 2 2 2886 1777
0 1779 5 1 1 3502
0 1780 7 1 2 2867 3503
0 1781 5 1 1 1780
0 1782 7 1 2 3406 1781
0 1783 7 1 2 1775 1782
0 1784 5 1 1 1783
0 1785 7 1 2 2870 1779
0 1786 5 1 1 1785
0 1787 7 1 2 1784 1786
0 1788 5 1 1 1787
0 1789 7 1 2 1773 1788
0 1790 5 1 1 1789
0 1791 7 1 2 1771 1790
0 1792 5 1 1 1791
0 1793 7 1 2 1765 1792
0 1794 5 1 1 1793
0 1795 7 2 2 1763 1794
0 1796 5 1 1 3504
0 1797 7 1 2 3497 1796
0 1798 5 1 1 1797
0 1799 7 1 2 1757 3505
0 1800 5 1 1 1799
0 1801 7 1 2 2831 1800
0 1802 5 1 1 1801
0 1803 7 2 2 1798 1802
0 1804 5 1 1 3506
0 1805 7 1 2 2817 3507
0 1806 5 1 1 1805
0 1807 7 1 2 3424 1627
0 1808 5 1 1 1807
0 1809 7 1 2 3428 1808
0 1810 7 1 2 1806 1809
0 1811 5 1 1 1810
0 1812 7 1 2 2820 1804
0 1813 5 1 1 1812
0 1814 7 1 2 1811 1813
0 1815 5 1 1 1814
0 1816 7 1 2 1753 1815
0 1817 5 1 1 1816
0 1818 7 1 2 1751 1817
0 1819 5 1 1 1818
0 1820 7 1 2 1745 1819
0 1821 5 1 1 1820
0 1822 7 1 2 1743 1821
0 1823 5 1 1 1822
0 1824 7 1 2 1737 1823
0 1825 5 1 1 1824
0 1826 7 1 2 1735 1825
0 1827 5 1 1 1826
0 1828 7 1 2 1729 1827
0 1829 5 1 1 1828
0 1830 7 1 2 1727 1829
0 1831 5 1 1 1830
0 1832 7 1 2 1721 1831
0 1833 5 1 1 1832
0 1834 7 1 2 1719 1833
0 1835 5 1 1 1834
0 1836 7 1 2 1713 1835
0 1837 5 1 1 1836
0 1838 7 1 2 1711 1837
0 1839 5 1 1 1838
0 1840 7 1 2 1705 1839
0 1841 5 1 1 1840
0 1842 7 2 2 1703 1841
0 1843 5 1 1 3508
0 1844 7 1 2 2938 3509
0 1845 5 1 1 1844
0 1846 7 2 2 3477 3481
0 1847 5 1 1 3510
0 1848 7 1 2 2944 3470
0 1849 5 1 1 1848
0 1850 7 2 2 2947 1849
0 1851 5 2 1 3512
0 1852 7 1 2 3012 3513
0 1853 5 1 1 1852
0 1854 7 1 2 3010 3514
0 1855 5 1 1 1854
0 1856 7 3 2 1853 1855
0 1857 5 2 1 3516
0 1858 7 1 2 3327 3517
0 1859 5 2 1 1858
0 1860 7 1 2 3329 3519
0 1861 5 1 1 1860
0 1862 7 2 2 3521 1861
0 1863 5 1 1 3523
0 1864 7 1 2 1847 3524
0 1865 5 2 1 1864
0 1866 7 1 2 3511 1863
0 1867 5 1 1 1866
0 1868 7 1 2 3525 1867
0 1869 7 1 2 1845 1868
0 1870 5 1 1 1869
0 1871 7 2 2 3522 3526
0 1872 5 1 1 3527
0 1873 7 1 2 2978 3515
0 1874 5 1 1 1873
0 1875 7 3 2 2981 1874
0 1876 5 2 1 3529
0 1877 7 1 2 2966 3532
0 1878 5 1 1 1877
0 1879 7 1 2 2968 3530
0 1880 5 1 1 1879
0 1881 7 2 2 1878 1880
0 1882 5 1 1 3534
0 1883 7 1 2 3473 3535
0 1884 5 2 1 1883
0 1885 7 1 2 3475 1882
0 1886 5 1 1 1885
0 1887 7 2 2 3536 1886
0 1888 5 1 1 3538
0 1889 7 1 2 1872 3539
0 1890 5 2 1 1889
0 1891 7 1 2 3528 1888
0 1892 5 1 1 1891
0 1893 7 2 2 3540 1892
0 1894 5 1 1 3542
0 1895 7 1 2 2975 3543
0 1896 5 1 1 1895
0 1897 7 1 2 2941 1843
0 1898 5 1 1 1897
0 1899 7 1 2 1896 1898
0 1900 7 1 2 1870 1899
0 1901 5 1 1 1900
0 1902 7 2 2 3537 3541
0 1903 5 1 1 3544
0 1904 7 1 2 2963 3531
0 1905 5 2 1 1904
0 1906 7 2 2 2960 3546
0 1907 5 1 1 3548
0 1908 7 1 2 3520 3549
0 1909 5 1 1 1908
0 1910 7 1 2 3518 1907
0 1911 5 1 1 1910
0 1912 7 2 2 1909 1911
0 1913 5 1 1 3550
0 1914 7 1 2 1903 3551
0 1915 5 2 1 1914
0 1916 7 1 2 3545 1913
0 1917 5 1 1 1916
0 1918 7 2 2 3552 1917
0 1919 5 1 1 3554
0 1920 7 1 2 2722 1919
0 1921 5 1 1 1920
0 1922 7 1 2 2972 1894
0 1923 5 1 1 1922
0 1924 7 1 2 1921 1923
0 1925 7 1 2 1901 1924
0 1926 5 1 1 1925
0 1927 7 1 2 2719 3555
0 1928 5 1 1 1927
0 1929 7 1 2 2993 3533
0 1930 5 1 1 1929
0 1931 7 1 2 3547 1930
0 1932 7 1 2 3553 1931
0 1933 7 1 2 1928 1932
0 1934 7 1 2 1926 1933
0 1935 5 1 1 1934
0 1936 7 1 2 1461 1935
3 4299 5 0 1 1936
